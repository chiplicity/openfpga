magic
tech EFS8A
magscale 1 2
timestamp 1604349425
<< locali >>
rect 175249 272375 175283 276625
rect 175341 262651 175375 269621
rect 175341 250343 175375 259965
rect 175341 243407 175375 243577
rect 154825 233615 154859 233785
rect 164393 233479 164427 233785
rect 255749 233547 255783 233649
rect 255749 233513 255933 233547
rect 156239 233309 156389 233343
rect 61261 232663 61295 232901
rect 247745 232799 247779 232969
rect 161173 231507 161207 232697
rect 248481 232595 248515 232901
rect 256485 232595 256519 233241
rect 59605 225251 59639 225421
rect 60893 225319 60927 225489
rect 60985 225387 61019 225489
rect 60985 225353 61077 225387
rect 56293 224707 56327 225013
rect 56385 224571 56419 224877
rect 58869 223687 58903 225013
rect 59329 224367 59363 225081
rect 61445 224979 61479 225217
rect 157769 225115 157803 226849
rect 60893 224435 60927 224877
rect 61537 224571 61571 224877
rect 157401 224707 157435 225081
rect 253725 224911 253759 225421
rect 61537 224537 61813 224571
rect 59329 224333 59513 224367
rect 59329 224027 59363 224265
rect 250321 224163 250355 224741
rect 252529 224707 252563 224809
rect 253725 224299 253759 224537
rect 253817 224163 253851 224265
rect 23817 181119 23851 181289
rect 58133 175475 58167 181221
rect 58869 180167 58903 181357
rect 60433 180031 60467 181017
rect 60893 180779 60927 181221
rect 251517 181187 251551 181357
rect 62825 180915 62859 181017
rect 62917 180167 62951 180881
rect 63377 180575 63411 180677
rect 156941 180507 156975 181085
rect 63929 179963 63963 180269
rect 153169 179963 153203 180201
rect 153353 180099 153387 180269
rect 157217 180235 157251 180881
rect 248849 180847 248883 181085
rect 159149 180167 159183 180745
rect 248757 180303 248791 180813
rect 249677 180235 249711 181017
rect 250413 180167 250447 180677
rect 154917 179895 154951 179997
rect 157493 179963 157527 180065
rect 251057 180031 251091 180745
rect 254277 180643 254311 181153
rect 155285 179827 155319 179929
rect 103765 175475 103799 175645
rect 200365 175475 200399 175781
rect 205149 175679 205183 175781
rect 152065 172959 152099 173061
rect 153077 172891 153111 173061
rect 151973 172211 152007 172857
rect 152341 172007 152375 172857
rect 153261 172143 153295 172721
rect 156757 172687 156791 172857
rect 161357 172687 161391 172857
rect 256025 171735 256059 172313
rect 173041 157183 173075 160345
rect 134033 154803 134067 154973
rect 228333 145419 228367 145929
rect 176261 144739 176295 145385
rect 228333 145283 228367 145385
rect 60985 138755 61019 139129
rect 61077 138823 61111 139061
rect 61169 138959 61203 139129
rect 61261 138687 61295 139673
rect 61353 138891 61387 138993
rect 61353 138857 61997 138891
rect 69909 138619 69943 139197
rect 70553 139027 70587 139537
rect 156849 139469 157677 139503
rect 156113 139027 156147 139401
rect 156849 138959 156883 139469
rect 244617 139435 244651 139673
rect 250045 139435 250079 139945
rect 250723 139877 250965 139911
rect 250413 139741 250965 139775
rect 250413 139299 250447 139741
rect 158965 138619 158999 139265
rect 252069 138619 252103 139605
rect 252253 138823 252287 139333
rect 253541 139163 253575 139401
rect 253633 138959 253667 139129
rect 59237 130595 59271 131173
rect 59237 130561 59697 130595
rect 60341 130459 60375 130969
rect 60709 130867 60743 131309
rect 60801 130391 60835 131377
rect 60893 130595 60927 130833
rect 64941 130391 64975 131377
rect 155745 131207 155779 131513
rect 157217 131479 157251 131513
rect 157217 131445 157527 131479
rect 155135 130833 155285 130867
rect 157401 130799 157435 131377
rect 157493 131275 157527 131445
rect 157493 131241 157769 131275
rect 157861 131071 157895 131649
rect 249401 131547 249435 131717
rect 245077 130799 245111 130969
rect 156055 130629 156147 130663
rect 64941 130357 65033 130391
rect 62365 130255 62399 130357
rect 156113 130323 156147 130629
rect 157033 130527 157067 130765
rect 63779 130289 63929 130323
rect 158321 130323 158355 130629
rect 246365 130595 246399 131445
rect 249861 130731 249895 131105
rect 250229 131003 250263 131377
rect 250597 130901 250689 130935
rect 250597 130663 250631 130901
rect 250781 130867 250815 131513
rect 251149 130663 251183 130833
rect 252161 130731 252195 131649
rect 228425 120531 228459 124713
rect 292825 110263 292859 112473
rect 228517 90883 228551 95745
rect 60157 87279 60191 87517
rect 60985 87211 61019 87449
rect 58961 86803 58995 87109
rect 155561 86735 155595 87517
rect 157435 87109 157527 87143
rect 156607 86497 156883 86531
rect 156849 86463 156883 86497
rect 157217 86463 157251 86973
rect 157493 86939 157527 87109
rect 250781 87007 250815 87517
rect 157401 86123 157435 86905
rect 251241 86735 251275 86905
rect 251241 86701 251517 86735
rect 86837 81839 86871 83845
rect 58685 78507 58719 78609
rect 60341 78235 60375 78337
rect 62089 78099 62123 78609
rect 62273 78235 62307 78473
rect 62181 78099 62215 78201
rect 89781 77691 89815 83913
rect 93645 81839 93679 83845
rect 94933 80751 94967 83845
rect 96681 81907 96715 83981
rect 109837 81907 109871 83845
rect 99717 81771 99751 81873
rect 99659 81737 99751 81771
rect 100177 81159 100211 81805
rect 111217 80139 111251 83845
rect 112505 81839 112539 83845
rect 115173 81635 115207 83845
rect 117933 81567 117967 83845
rect 120601 81499 120635 83913
rect 123269 81431 123303 83845
rect 124741 80139 124775 83913
rect 126029 81363 126063 83845
rect 128697 81295 128731 83845
rect 196961 81771 196995 81941
rect 156021 78711 156055 79425
rect 158413 78439 158447 79017
rect 249401 78575 249435 78745
rect 157401 78031 157435 78065
rect 157401 77997 157493 78031
rect 157309 77895 157343 77997
rect 157309 77861 157493 77895
rect 135781 58583 135815 58753
<< viali >>
rect 175249 276625 175283 276659
rect 175249 272341 175283 272375
rect 175341 269621 175375 269655
rect 175341 262617 175375 262651
rect 175341 259965 175375 259999
rect 175341 250309 175375 250343
rect 175341 243577 175375 243611
rect 175341 243373 175375 243407
rect 154825 233785 154859 233819
rect 154825 233581 154859 233615
rect 164393 233785 164427 233819
rect 255749 233649 255783 233683
rect 255933 233513 255967 233547
rect 164393 233445 164427 233479
rect 156205 233309 156239 233343
rect 156389 233309 156423 233343
rect 256485 233241 256519 233275
rect 247745 232969 247779 233003
rect 61261 232901 61295 232935
rect 247745 232765 247779 232799
rect 248481 232901 248515 232935
rect 61261 232629 61295 232663
rect 161173 232697 161207 232731
rect 248481 232561 248515 232595
rect 256485 232561 256519 232595
rect 161173 231473 161207 231507
rect 157769 226849 157803 226883
rect 60893 225489 60927 225523
rect 59605 225421 59639 225455
rect 60985 225489 61019 225523
rect 61077 225353 61111 225387
rect 60893 225285 60927 225319
rect 59605 225217 59639 225251
rect 61445 225217 61479 225251
rect 59329 225081 59363 225115
rect 56293 225013 56327 225047
rect 58869 225013 58903 225047
rect 56293 224673 56327 224707
rect 56385 224877 56419 224911
rect 56385 224537 56419 224571
rect 61445 224945 61479 224979
rect 157401 225081 157435 225115
rect 157769 225081 157803 225115
rect 253725 225421 253759 225455
rect 60893 224877 60927 224911
rect 61537 224877 61571 224911
rect 253725 224877 253759 224911
rect 252529 224809 252563 224843
rect 157401 224673 157435 224707
rect 250321 224741 250355 224775
rect 61813 224537 61847 224571
rect 60893 224401 60927 224435
rect 59513 224333 59547 224367
rect 59329 224265 59363 224299
rect 252529 224673 252563 224707
rect 253725 224537 253759 224571
rect 253725 224265 253759 224299
rect 253817 224265 253851 224299
rect 250321 224129 250355 224163
rect 253817 224129 253851 224163
rect 59329 223993 59363 224027
rect 58869 223653 58903 223687
rect 58869 181357 58903 181391
rect 23817 181289 23851 181323
rect 23817 181085 23851 181119
rect 58133 181221 58167 181255
rect 251517 181357 251551 181391
rect 60893 181221 60927 181255
rect 58869 180133 58903 180167
rect 60433 181017 60467 181051
rect 251517 181153 251551 181187
rect 254277 181153 254311 181187
rect 156941 181085 156975 181119
rect 62825 181017 62859 181051
rect 62825 180881 62859 180915
rect 62917 180881 62951 180915
rect 60893 180745 60927 180779
rect 63377 180677 63411 180711
rect 63377 180541 63411 180575
rect 248849 181085 248883 181119
rect 156941 180473 156975 180507
rect 157217 180881 157251 180915
rect 62917 180133 62951 180167
rect 63929 180269 63963 180303
rect 60433 179997 60467 180031
rect 153353 180269 153387 180303
rect 63929 179929 63963 179963
rect 153169 180201 153203 180235
rect 248757 180813 248791 180847
rect 248849 180813 248883 180847
rect 249677 181017 249711 181051
rect 157217 180201 157251 180235
rect 159149 180745 159183 180779
rect 248757 180269 248791 180303
rect 251057 180745 251091 180779
rect 249677 180201 249711 180235
rect 250413 180677 250447 180711
rect 159149 180133 159183 180167
rect 250413 180133 250447 180167
rect 153353 180065 153387 180099
rect 157493 180065 157527 180099
rect 153169 179929 153203 179963
rect 154917 179997 154951 180031
rect 254277 180609 254311 180643
rect 251057 179997 251091 180031
rect 154917 179861 154951 179895
rect 155285 179929 155319 179963
rect 157493 179929 157527 179963
rect 155285 179793 155319 179827
rect 200365 175781 200399 175815
rect 58133 175441 58167 175475
rect 103765 175645 103799 175679
rect 103765 175441 103799 175475
rect 205149 175781 205183 175815
rect 205149 175645 205183 175679
rect 200365 175441 200399 175475
rect 152065 173061 152099 173095
rect 152065 172925 152099 172959
rect 153077 173061 153111 173095
rect 151973 172857 152007 172891
rect 151973 172177 152007 172211
rect 152341 172857 152375 172891
rect 153077 172857 153111 172891
rect 156757 172857 156791 172891
rect 153261 172721 153295 172755
rect 156757 172653 156791 172687
rect 161357 172857 161391 172891
rect 161357 172653 161391 172687
rect 153261 172109 153295 172143
rect 256025 172313 256059 172347
rect 152341 171973 152375 172007
rect 256025 171701 256059 171735
rect 173041 160345 173075 160379
rect 173041 157149 173075 157183
rect 134033 154973 134067 155007
rect 134033 154769 134067 154803
rect 228333 145929 228367 145963
rect 176261 145385 176295 145419
rect 228333 145385 228367 145419
rect 228333 145249 228367 145283
rect 176261 144705 176295 144739
rect 250045 139945 250079 139979
rect 61261 139673 61295 139707
rect 60985 139129 61019 139163
rect 61169 139129 61203 139163
rect 61077 139061 61111 139095
rect 61169 138925 61203 138959
rect 61077 138789 61111 138823
rect 60985 138721 61019 138755
rect 244617 139673 244651 139707
rect 70553 139537 70587 139571
rect 69909 139197 69943 139231
rect 61353 138993 61387 139027
rect 61997 138857 62031 138891
rect 61261 138653 61295 138687
rect 157677 139469 157711 139503
rect 70553 138993 70587 139027
rect 156113 139401 156147 139435
rect 156113 138993 156147 139027
rect 244617 139401 244651 139435
rect 250689 139877 250723 139911
rect 250965 139877 250999 139911
rect 250045 139401 250079 139435
rect 250965 139741 250999 139775
rect 156849 138925 156883 138959
rect 158965 139265 158999 139299
rect 250413 139265 250447 139299
rect 252069 139605 252103 139639
rect 69909 138585 69943 138619
rect 158965 138585 158999 138619
rect 253541 139401 253575 139435
rect 252253 139333 252287 139367
rect 253541 139129 253575 139163
rect 253633 139129 253667 139163
rect 253633 138925 253667 138959
rect 252253 138789 252287 138823
rect 252069 138585 252103 138619
rect 249401 131717 249435 131751
rect 157861 131649 157895 131683
rect 155745 131513 155779 131547
rect 60801 131377 60835 131411
rect 60709 131309 60743 131343
rect 59237 131173 59271 131207
rect 60341 130969 60375 131003
rect 59697 130561 59731 130595
rect 60709 130833 60743 130867
rect 60341 130425 60375 130459
rect 64941 131377 64975 131411
rect 60893 130833 60927 130867
rect 60893 130561 60927 130595
rect 157217 131513 157251 131547
rect 155745 131173 155779 131207
rect 157401 131377 157435 131411
rect 155101 130833 155135 130867
rect 155285 130833 155319 130867
rect 157769 131241 157803 131275
rect 252161 131649 252195 131683
rect 249401 131513 249435 131547
rect 250781 131513 250815 131547
rect 157861 131037 157895 131071
rect 246365 131445 246399 131479
rect 157033 130765 157067 130799
rect 157401 130765 157435 130799
rect 245077 130969 245111 131003
rect 245077 130765 245111 130799
rect 156021 130629 156055 130663
rect 60801 130357 60835 130391
rect 62365 130357 62399 130391
rect 65033 130357 65067 130391
rect 157033 130493 157067 130527
rect 158321 130629 158355 130663
rect 63745 130289 63779 130323
rect 63929 130289 63963 130323
rect 156113 130289 156147 130323
rect 250229 131377 250263 131411
rect 249861 131105 249895 131139
rect 250229 130969 250263 131003
rect 249861 130697 249895 130731
rect 250689 130901 250723 130935
rect 250781 130833 250815 130867
rect 251149 130833 251183 130867
rect 250597 130629 250631 130663
rect 252161 130697 252195 130731
rect 251149 130629 251183 130663
rect 246365 130561 246399 130595
rect 158321 130289 158355 130323
rect 62365 130221 62399 130255
rect 228425 124713 228459 124747
rect 228425 120497 228459 120531
rect 292825 112473 292859 112507
rect 292825 110229 292859 110263
rect 228517 95745 228551 95779
rect 228517 90849 228551 90883
rect 60157 87517 60191 87551
rect 155561 87517 155595 87551
rect 60157 87245 60191 87279
rect 60985 87449 61019 87483
rect 60985 87177 61019 87211
rect 58961 87109 58995 87143
rect 58961 86769 58995 86803
rect 250781 87517 250815 87551
rect 157401 87109 157435 87143
rect 155561 86701 155595 86735
rect 157217 86973 157251 87007
rect 156573 86497 156607 86531
rect 156849 86429 156883 86463
rect 250781 86973 250815 87007
rect 157217 86429 157251 86463
rect 157401 86905 157435 86939
rect 157493 86905 157527 86939
rect 251241 86905 251275 86939
rect 251517 86701 251551 86735
rect 157401 86089 157435 86123
rect 96681 83981 96715 84015
rect 89781 83913 89815 83947
rect 86837 83845 86871 83879
rect 86837 81805 86871 81839
rect 58685 78609 58719 78643
rect 58685 78473 58719 78507
rect 62089 78609 62123 78643
rect 60341 78337 60375 78371
rect 60341 78201 60375 78235
rect 62273 78473 62307 78507
rect 62089 78065 62123 78099
rect 62181 78201 62215 78235
rect 62273 78201 62307 78235
rect 62181 78065 62215 78099
rect 93645 83845 93679 83879
rect 93645 81805 93679 81839
rect 94933 83845 94967 83879
rect 120601 83913 120635 83947
rect 109837 83845 109871 83879
rect 96681 81873 96715 81907
rect 99717 81873 99751 81907
rect 109837 81873 109871 81907
rect 111217 83845 111251 83879
rect 99625 81737 99659 81771
rect 100177 81805 100211 81839
rect 100177 81125 100211 81159
rect 94933 80717 94967 80751
rect 112505 83845 112539 83879
rect 112505 81805 112539 81839
rect 115173 83845 115207 83879
rect 115173 81601 115207 81635
rect 117933 83845 117967 83879
rect 117933 81533 117967 81567
rect 124741 83913 124775 83947
rect 120601 81465 120635 81499
rect 123269 83845 123303 83879
rect 123269 81397 123303 81431
rect 111217 80105 111251 80139
rect 126029 83845 126063 83879
rect 126029 81329 126063 81363
rect 128697 83845 128731 83879
rect 196961 81941 196995 81975
rect 196961 81737 196995 81771
rect 128697 81261 128731 81295
rect 124741 80105 124775 80139
rect 156021 79425 156055 79459
rect 156021 78677 156055 78711
rect 158413 79017 158447 79051
rect 249401 78745 249435 78779
rect 249401 78541 249435 78575
rect 158413 78405 158447 78439
rect 157401 78065 157435 78099
rect 157309 77997 157343 78031
rect 157493 77997 157527 78031
rect 157493 77861 157527 77895
rect 89781 77657 89815 77691
rect 135781 58753 135815 58787
rect 135781 58549 135815 58583
<< metal1 >>
rect 34658 299396 34664 299448
rect 34716 299436 34722 299448
rect 211942 299436 211948 299448
rect 34716 299408 211948 299436
rect 34716 299396 34722 299408
rect 211942 299396 211948 299408
rect 212000 299396 212006 299448
rect 248742 299396 248748 299448
rect 248800 299436 248806 299448
rect 267234 299436 267240 299448
rect 248800 299408 267240 299436
rect 248800 299396 248806 299408
rect 267234 299396 267240 299408
rect 267292 299396 267298 299448
rect 101726 299328 101732 299380
rect 101784 299368 101790 299380
rect 292534 299368 292540 299380
rect 101784 299340 292540 299368
rect 101784 299328 101790 299340
rect 292534 299328 292540 299340
rect 292592 299328 292598 299380
rect 34566 299260 34572 299312
rect 34624 299300 34630 299312
rect 285450 299300 285456 299312
rect 34624 299272 285456 299300
rect 34624 299260 34630 299272
rect 285450 299260 285456 299272
rect 285508 299260 285514 299312
rect 28218 298648 28224 298700
rect 28276 298688 28282 298700
rect 29138 298688 29144 298700
rect 28276 298660 29144 298688
rect 28276 298648 28282 298660
rect 29138 298648 29144 298660
rect 29196 298648 29202 298700
rect 138434 298648 138440 298700
rect 138492 298688 138498 298700
rect 139538 298688 139544 298700
rect 138492 298660 139544 298688
rect 138492 298648 138498 298660
rect 139538 298648 139544 298660
rect 139596 298648 139602 298700
rect 65018 295112 65024 295164
rect 65076 295152 65082 295164
rect 96206 295152 96212 295164
rect 65076 295124 96212 295152
rect 65076 295112 65082 295124
rect 96206 295112 96212 295124
rect 96264 295112 96270 295164
rect 139538 295112 139544 295164
rect 139596 295152 139602 295164
rect 203846 295152 203852 295164
rect 139596 295124 203852 295152
rect 139596 295112 139602 295124
rect 203846 295112 203852 295124
rect 203904 295112 203910 295164
rect 123530 294636 123536 294688
rect 123588 294676 123594 294688
rect 264750 294676 264756 294688
rect 123588 294648 264756 294676
rect 123588 294636 123594 294648
rect 264750 294636 264756 294648
rect 264808 294636 264814 294688
rect 13406 294568 13412 294620
rect 13464 294608 13470 294620
rect 190506 294608 190512 294620
rect 13464 294580 190512 294608
rect 13464 294568 13470 294580
rect 190506 294568 190512 294580
rect 190564 294568 190570 294620
rect 217186 294568 217192 294620
rect 217244 294608 217250 294620
rect 265854 294608 265860 294620
rect 217244 294580 265860 294608
rect 217244 294568 217250 294580
rect 265854 294568 265860 294580
rect 265912 294568 265918 294620
rect 110190 294500 110196 294552
rect 110248 294540 110254 294552
rect 292626 294540 292632 294552
rect 110248 294512 292632 294540
rect 110248 294500 110254 294512
rect 292626 294500 292632 294512
rect 292684 294500 292690 294552
rect 13222 286204 13228 286256
rect 13280 286244 13286 286256
rect 20214 286244 20220 286256
rect 13280 286216 20220 286244
rect 13280 286204 13286 286216
rect 20214 286204 20220 286216
rect 20272 286204 20278 286256
rect 175234 276656 175240 276668
rect 175195 276628 175240 276656
rect 175234 276616 175240 276628
rect 175292 276616 175298 276668
rect 79554 274440 79560 274492
rect 79612 274480 79618 274492
rect 114790 274480 114796 274492
rect 79612 274452 114796 274480
rect 79612 274440 79618 274452
rect 114790 274440 114796 274452
rect 114848 274440 114854 274492
rect 173394 274440 173400 274492
rect 173452 274480 173458 274492
rect 208814 274480 208820 274492
rect 173452 274452 208820 274480
rect 173452 274440 173458 274452
rect 208814 274440 208820 274452
rect 208872 274440 208878 274492
rect 218842 274440 218848 274492
rect 218900 274480 218906 274492
rect 225282 274480 225288 274492
rect 218900 274452 225288 274480
rect 218900 274440 218906 274452
rect 225282 274440 225288 274452
rect 225340 274440 225346 274492
rect 175234 272372 175240 272384
rect 175195 272344 175240 272372
rect 175234 272332 175240 272344
rect 175292 272332 175298 272384
rect 175234 269612 175240 269664
rect 175292 269652 175298 269664
rect 175329 269655 175387 269661
rect 175329 269652 175341 269655
rect 175292 269624 175341 269652
rect 175292 269612 175298 269624
rect 175329 269621 175341 269624
rect 175375 269621 175387 269655
rect 175329 269615 175387 269621
rect 265854 266824 265860 266876
rect 265912 266864 265918 266876
rect 300078 266864 300084 266876
rect 265912 266836 300084 266864
rect 265912 266824 265918 266836
rect 300078 266824 300084 266836
rect 300136 266824 300142 266876
rect 78910 264036 78916 264088
rect 78968 264076 78974 264088
rect 124450 264076 124456 264088
rect 78968 264048 124456 264076
rect 78968 264036 78974 264048
rect 124450 264036 124456 264048
rect 124508 264076 124514 264088
rect 125738 264076 125744 264088
rect 124508 264048 125744 264076
rect 124508 264036 124514 264048
rect 125738 264036 125744 264048
rect 125796 264036 125802 264088
rect 143034 264036 143040 264088
rect 143092 264076 143098 264088
rect 225190 264076 225196 264088
rect 143092 264048 225196 264076
rect 143092 264036 143098 264048
rect 225190 264036 225196 264048
rect 225248 264036 225254 264088
rect 198878 263968 198884 264020
rect 198936 264008 198942 264020
rect 233470 264008 233476 264020
rect 198936 263980 233476 264008
rect 198936 263968 198942 263980
rect 233470 263968 233476 263980
rect 233528 263968 233534 264020
rect 125738 263356 125744 263408
rect 125796 263396 125802 263408
rect 132730 263396 132736 263408
rect 125796 263368 132736 263396
rect 125796 263356 125802 263368
rect 132730 263356 132736 263368
rect 132788 263396 132794 263408
rect 139630 263396 139636 263408
rect 132788 263368 139636 263396
rect 132788 263356 132794 263368
rect 139630 263356 139636 263368
rect 139688 263356 139694 263408
rect 105038 262676 105044 262728
rect 105096 262716 105102 262728
rect 139630 262716 139636 262728
rect 105096 262688 139636 262716
rect 105096 262676 105102 262688
rect 139630 262676 139636 262688
rect 139688 262676 139694 262728
rect 47078 262608 47084 262660
rect 47136 262648 47142 262660
rect 131350 262648 131356 262660
rect 47136 262620 131356 262648
rect 47136 262608 47142 262620
rect 131350 262608 131356 262620
rect 131408 262608 131414 262660
rect 175326 262648 175332 262660
rect 175287 262620 175332 262648
rect 175326 262608 175332 262620
rect 175384 262608 175390 262660
rect 80106 261452 80112 261504
rect 80164 261492 80170 261504
rect 87190 261492 87196 261504
rect 80164 261464 87196 261492
rect 80164 261452 80170 261464
rect 87190 261452 87196 261464
rect 87248 261452 87254 261504
rect 173578 261452 173584 261504
rect 173636 261492 173642 261504
rect 181950 261492 181956 261504
rect 173636 261464 181956 261492
rect 173636 261452 173642 261464
rect 181950 261452 181956 261464
rect 182008 261452 182014 261504
rect 80198 261384 80204 261436
rect 80256 261424 80262 261436
rect 87282 261424 87288 261436
rect 80256 261396 87288 261424
rect 80256 261384 80262 261396
rect 87282 261384 87288 261396
rect 87340 261384 87346 261436
rect 173670 261384 173676 261436
rect 173728 261424 173734 261436
rect 181766 261424 181772 261436
rect 173728 261396 181772 261424
rect 173728 261384 173734 261396
rect 181766 261384 181772 261396
rect 181824 261384 181830 261436
rect 95378 260636 95384 260688
rect 95436 260676 95442 260688
rect 109546 260676 109552 260688
rect 95436 260648 109552 260676
rect 95436 260636 95442 260648
rect 109546 260636 109552 260648
rect 109604 260636 109610 260688
rect 189218 260636 189224 260688
rect 189276 260676 189282 260688
rect 203846 260676 203852 260688
rect 189276 260648 203852 260676
rect 189276 260636 189282 260648
rect 203846 260636 203852 260648
rect 203904 260636 203910 260688
rect 80106 260160 80112 260212
rect 80164 260200 80170 260212
rect 85166 260200 85172 260212
rect 80164 260172 85172 260200
rect 80164 260160 80170 260172
rect 85166 260160 85172 260172
rect 85224 260160 85230 260212
rect 80198 260092 80204 260144
rect 80256 260132 80262 260144
rect 85074 260132 85080 260144
rect 80256 260104 85080 260132
rect 80256 260092 80262 260104
rect 85074 260092 85080 260104
rect 85132 260092 85138 260144
rect 172842 260092 172848 260144
rect 172900 260132 172906 260144
rect 179006 260132 179012 260144
rect 172900 260104 179012 260132
rect 172900 260092 172906 260104
rect 179006 260092 179012 260104
rect 179064 260092 179070 260144
rect 173578 260024 173584 260076
rect 173636 260064 173642 260076
rect 179098 260064 179104 260076
rect 173636 260036 179104 260064
rect 173636 260024 173642 260036
rect 179098 260024 179104 260036
rect 179156 260024 179162 260076
rect 229974 260024 229980 260076
rect 230032 260064 230038 260076
rect 233470 260064 233476 260076
rect 230032 260036 233476 260064
rect 230032 260024 230038 260036
rect 233470 260024 233476 260036
rect 233528 260024 233534 260076
rect 175326 259996 175332 260008
rect 175287 259968 175332 259996
rect 175326 259956 175332 259968
rect 175384 259956 175390 260008
rect 173394 259344 173400 259396
rect 173452 259384 173458 259396
rect 175694 259384 175700 259396
rect 173452 259356 175700 259384
rect 173452 259344 173458 259356
rect 175694 259344 175700 259356
rect 175752 259344 175758 259396
rect 80198 258664 80204 258716
rect 80256 258704 80262 258716
rect 84430 258704 84436 258716
rect 80256 258676 84436 258704
rect 80256 258664 80262 258676
rect 84430 258664 84436 258676
rect 84488 258664 84494 258716
rect 173578 258664 173584 258716
rect 173636 258704 173642 258716
rect 178914 258704 178920 258716
rect 173636 258676 178920 258704
rect 173636 258664 173642 258676
rect 178914 258664 178920 258676
rect 178972 258664 178978 258716
rect 79830 258596 79836 258648
rect 79888 258636 79894 258648
rect 82406 258636 82412 258648
rect 79888 258608 82412 258636
rect 79888 258596 79894 258608
rect 82406 258596 82412 258608
rect 82464 258596 82470 258648
rect 88478 258528 88484 258580
rect 88536 258568 88542 258580
rect 129510 258568 129516 258580
rect 88536 258540 129516 258568
rect 88536 258528 88542 258540
rect 129510 258528 129516 258540
rect 129568 258528 129574 258580
rect 182318 258528 182324 258580
rect 182376 258568 182382 258580
rect 223534 258568 223540 258580
rect 182376 258540 223540 258568
rect 182376 258528 182382 258540
rect 223534 258528 223540 258540
rect 223592 258528 223598 258580
rect 173302 257984 173308 258036
rect 173360 258024 173366 258036
rect 175602 258024 175608 258036
rect 173360 257996 175608 258024
rect 173360 257984 173366 257996
rect 175602 257984 175608 257996
rect 175660 257984 175666 258036
rect 229422 257712 229428 257764
rect 229480 257752 229486 257764
rect 233562 257752 233568 257764
rect 229480 257724 233568 257752
rect 229480 257712 229486 257724
rect 233562 257712 233568 257724
rect 233620 257712 233626 257764
rect 80014 257644 80020 257696
rect 80072 257684 80078 257696
rect 82314 257684 82320 257696
rect 80072 257656 82320 257684
rect 80072 257644 80078 257656
rect 82314 257644 82320 257656
rect 82372 257644 82378 257696
rect 229514 257508 229520 257560
rect 229572 257548 229578 257560
rect 233470 257548 233476 257560
rect 229572 257520 233476 257548
rect 229572 257508 229578 257520
rect 233470 257508 233476 257520
rect 233528 257508 233534 257560
rect 173578 257304 173584 257356
rect 173636 257344 173642 257356
rect 175510 257344 175516 257356
rect 173636 257316 175516 257344
rect 173636 257304 173642 257316
rect 175510 257304 175516 257316
rect 175568 257304 175574 257356
rect 80198 257236 80204 257288
rect 80256 257276 80262 257288
rect 81670 257276 81676 257288
rect 80256 257248 81676 257276
rect 80256 257236 80262 257248
rect 81670 257236 81676 257248
rect 81728 257236 81734 257288
rect 131350 257236 131356 257288
rect 131408 257276 131414 257288
rect 132730 257276 132736 257288
rect 131408 257248 132736 257276
rect 131408 257236 131414 257248
rect 132730 257236 132736 257248
rect 132788 257276 132794 257288
rect 134202 257276 134208 257288
rect 132788 257248 134208 257276
rect 132788 257236 132794 257248
rect 134202 257236 134208 257248
rect 134260 257236 134266 257288
rect 229606 257236 229612 257288
rect 229664 257276 229670 257288
rect 233470 257276 233476 257288
rect 229664 257248 233476 257276
rect 229664 257236 229670 257248
rect 233470 257236 233476 257248
rect 233528 257236 233534 257288
rect 82406 257168 82412 257220
rect 82464 257208 82470 257220
rect 87190 257208 87196 257220
rect 82464 257180 87196 257208
rect 82464 257168 82470 257180
rect 87190 257168 87196 257180
rect 87248 257168 87254 257220
rect 131534 257168 131540 257220
rect 131592 257208 131598 257220
rect 140550 257208 140556 257220
rect 131592 257180 140556 257208
rect 131592 257168 131598 257180
rect 140550 257168 140556 257180
rect 140608 257168 140614 257220
rect 179006 257168 179012 257220
rect 179064 257208 179070 257220
rect 182318 257208 182324 257220
rect 179064 257180 182324 257208
rect 179064 257168 179070 257180
rect 182318 257168 182324 257180
rect 182376 257168 182382 257220
rect 226202 257168 226208 257220
rect 226260 257208 226266 257220
rect 234298 257208 234304 257220
rect 226260 257180 234304 257208
rect 226260 257168 226266 257180
rect 234298 257168 234304 257180
rect 234356 257168 234362 257220
rect 131350 257100 131356 257152
rect 131408 257140 131414 257152
rect 140274 257140 140280 257152
rect 131408 257112 140280 257140
rect 131408 257100 131414 257112
rect 140274 257100 140280 257112
rect 140332 257100 140338 257152
rect 179098 257100 179104 257152
rect 179156 257140 179162 257152
rect 182226 257140 182232 257152
rect 179156 257112 182232 257140
rect 179156 257100 179162 257112
rect 182226 257100 182232 257112
rect 182284 257100 182290 257152
rect 226294 257100 226300 257152
rect 226352 257140 226358 257152
rect 234666 257140 234672 257152
rect 226352 257112 234672 257140
rect 226352 257100 226358 257112
rect 234666 257100 234672 257112
rect 234724 257100 234730 257152
rect 131442 257032 131448 257084
rect 131500 257072 131506 257084
rect 140366 257072 140372 257084
rect 131500 257044 140372 257072
rect 131500 257032 131506 257044
rect 140366 257032 140372 257044
rect 140424 257032 140430 257084
rect 175694 257032 175700 257084
rect 175752 257072 175758 257084
rect 182042 257072 182048 257084
rect 175752 257044 182048 257072
rect 175752 257032 175758 257044
rect 182042 257032 182048 257044
rect 182100 257032 182106 257084
rect 225374 257032 225380 257084
rect 225432 257072 225438 257084
rect 234114 257072 234120 257084
rect 225432 257044 234120 257072
rect 225432 257032 225438 257044
rect 234114 257032 234120 257044
rect 234172 257032 234178 257084
rect 85166 256964 85172 257016
rect 85224 257004 85230 257016
rect 87282 257004 87288 257016
rect 85224 256976 87288 257004
rect 85224 256964 85230 256976
rect 87282 256964 87288 256976
rect 87340 256964 87346 257016
rect 85074 256760 85080 256812
rect 85132 256800 85138 256812
rect 87558 256800 87564 256812
rect 85132 256772 87564 256800
rect 85132 256760 85138 256772
rect 87558 256760 87564 256772
rect 87616 256760 87622 256812
rect 173118 256420 173124 256472
rect 173176 256460 173182 256472
rect 175786 256460 175792 256472
rect 173176 256432 175792 256460
rect 173176 256420 173182 256432
rect 175786 256420 175792 256432
rect 175844 256420 175850 256472
rect 173302 256080 173308 256132
rect 173360 256120 173366 256132
rect 175694 256120 175700 256132
rect 173360 256092 175700 256120
rect 173360 256080 173366 256092
rect 175694 256080 175700 256092
rect 175752 256080 175758 256132
rect 80106 255944 80112 255996
rect 80164 255984 80170 255996
rect 82130 255984 82136 255996
rect 80164 255956 82136 255984
rect 80164 255944 80170 255956
rect 82130 255944 82136 255956
rect 82188 255944 82194 255996
rect 80198 255876 80204 255928
rect 80256 255916 80262 255928
rect 81762 255916 81768 255928
rect 80256 255888 81768 255916
rect 80256 255876 80262 255888
rect 81762 255876 81768 255888
rect 81820 255876 81826 255928
rect 230158 255876 230164 255928
rect 230216 255916 230222 255928
rect 233470 255916 233476 255928
rect 230216 255888 233476 255916
rect 230216 255876 230222 255888
rect 233470 255876 233476 255888
rect 233528 255876 233534 255928
rect 82314 255808 82320 255860
rect 82372 255848 82378 255860
rect 87190 255848 87196 255860
rect 82372 255820 87196 255848
rect 82372 255808 82378 255820
rect 87190 255808 87196 255820
rect 87248 255808 87254 255860
rect 131534 255808 131540 255860
rect 131592 255848 131598 255860
rect 139814 255848 139820 255860
rect 131592 255820 139820 255848
rect 131592 255808 131598 255820
rect 139814 255808 139820 255820
rect 139872 255808 139878 255860
rect 175602 255808 175608 255860
rect 175660 255848 175666 255860
rect 181858 255848 181864 255860
rect 175660 255820 181864 255848
rect 175660 255808 175666 255820
rect 181858 255808 181864 255820
rect 181916 255808 181922 255860
rect 225558 255808 225564 255860
rect 225616 255848 225622 255860
rect 234758 255848 234764 255860
rect 225616 255820 234764 255848
rect 225616 255808 225622 255820
rect 234758 255808 234764 255820
rect 234816 255808 234822 255860
rect 81670 255740 81676 255792
rect 81728 255780 81734 255792
rect 87282 255780 87288 255792
rect 81728 255752 87288 255780
rect 81728 255740 81734 255752
rect 87282 255740 87288 255752
rect 87340 255740 87346 255792
rect 131626 255740 131632 255792
rect 131684 255780 131690 255792
rect 139630 255780 139636 255792
rect 131684 255752 139636 255780
rect 131684 255740 131690 255752
rect 139630 255740 139636 255752
rect 139688 255740 139694 255792
rect 175510 255740 175516 255792
rect 175568 255780 175574 255792
rect 182226 255780 182232 255792
rect 175568 255752 182232 255780
rect 175568 255740 175574 255752
rect 182226 255740 182232 255752
rect 182284 255740 182290 255792
rect 226386 255740 226392 255792
rect 226444 255780 226450 255792
rect 233838 255780 233844 255792
rect 226444 255752 233844 255780
rect 226444 255740 226450 255752
rect 233838 255740 233844 255752
rect 233896 255740 233902 255792
rect 84430 255672 84436 255724
rect 84488 255712 84494 255724
rect 87374 255712 87380 255724
rect 84488 255684 87380 255712
rect 84488 255672 84494 255684
rect 87374 255672 87380 255684
rect 87432 255672 87438 255724
rect 131442 255672 131448 255724
rect 131500 255712 131506 255724
rect 139906 255712 139912 255724
rect 131500 255684 139912 255712
rect 131500 255672 131506 255684
rect 139906 255672 139912 255684
rect 139964 255672 139970 255724
rect 178914 255672 178920 255724
rect 178972 255712 178978 255724
rect 182318 255712 182324 255724
rect 178972 255684 182324 255712
rect 178972 255672 178978 255684
rect 182318 255672 182324 255684
rect 182376 255672 182382 255724
rect 226294 255672 226300 255724
rect 226352 255712 226358 255724
rect 229974 255712 229980 255724
rect 226352 255684 229980 255712
rect 226352 255672 226358 255684
rect 229974 255672 229980 255684
rect 230032 255672 230038 255724
rect 131350 255604 131356 255656
rect 131408 255644 131414 255656
rect 140090 255644 140096 255656
rect 131408 255616 140096 255644
rect 131408 255604 131414 255616
rect 140090 255604 140096 255616
rect 140148 255604 140154 255656
rect 225926 255604 225932 255656
rect 225984 255644 225990 255656
rect 229422 255644 229428 255656
rect 225984 255616 229428 255644
rect 225984 255604 225990 255616
rect 229422 255604 229428 255616
rect 229480 255604 229486 255656
rect 80106 254584 80112 254636
rect 80164 254624 80170 254636
rect 80164 254596 85764 254624
rect 80164 254584 80170 254596
rect 80198 254448 80204 254500
rect 80256 254488 80262 254500
rect 84982 254488 84988 254500
rect 80256 254460 84988 254488
rect 80256 254448 80262 254460
rect 84982 254448 84988 254460
rect 85040 254448 85046 254500
rect 85736 254420 85764 254596
rect 173210 254516 173216 254568
rect 173268 254556 173274 254568
rect 173268 254528 178500 254556
rect 173268 254516 173274 254528
rect 173486 254448 173492 254500
rect 173544 254488 173550 254500
rect 173544 254460 178408 254488
rect 173544 254448 173550 254460
rect 87374 254420 87380 254432
rect 85736 254392 87380 254420
rect 87374 254380 87380 254392
rect 87432 254380 87438 254432
rect 131534 254380 131540 254432
rect 131592 254420 131598 254432
rect 139722 254420 139728 254432
rect 131592 254392 139728 254420
rect 131592 254380 131598 254392
rect 139722 254380 139728 254392
rect 139780 254380 139786 254432
rect 81762 254312 81768 254364
rect 81820 254352 81826 254364
rect 87282 254352 87288 254364
rect 81820 254324 87288 254352
rect 81820 254312 81826 254324
rect 87282 254312 87288 254324
rect 87340 254312 87346 254364
rect 131350 254312 131356 254364
rect 131408 254352 131414 254364
rect 139998 254352 140004 254364
rect 131408 254324 140004 254352
rect 131408 254312 131414 254324
rect 139998 254312 140004 254324
rect 140056 254312 140062 254364
rect 178380 254352 178408 254460
rect 178472 254420 178500 254528
rect 182042 254420 182048 254432
rect 178472 254392 182048 254420
rect 182042 254380 182048 254392
rect 182100 254380 182106 254432
rect 225926 254380 225932 254432
rect 225984 254420 225990 254432
rect 230158 254420 230164 254432
rect 225984 254392 230164 254420
rect 225984 254380 225990 254392
rect 230158 254380 230164 254392
rect 230216 254380 230222 254432
rect 182134 254352 182140 254364
rect 178380 254324 182140 254352
rect 182134 254312 182140 254324
rect 182192 254312 182198 254364
rect 131442 254244 131448 254296
rect 131500 254284 131506 254296
rect 139630 254284 139636 254296
rect 131500 254256 139636 254284
rect 131500 254244 131506 254256
rect 139630 254244 139636 254256
rect 139688 254244 139694 254296
rect 175786 254244 175792 254296
rect 175844 254284 175850 254296
rect 182226 254284 182232 254296
rect 175844 254256 182232 254284
rect 175844 254244 175850 254256
rect 182226 254244 182232 254256
rect 182284 254244 182290 254296
rect 82130 254176 82136 254228
rect 82188 254216 82194 254228
rect 87190 254216 87196 254228
rect 82188 254188 87196 254216
rect 82188 254176 82194 254188
rect 87190 254176 87196 254188
rect 87248 254176 87254 254228
rect 175694 254176 175700 254228
rect 175752 254216 175758 254228
rect 182318 254216 182324 254228
rect 175752 254188 182324 254216
rect 175752 254176 175758 254188
rect 182318 254176 182324 254188
rect 182376 254176 182382 254228
rect 226294 254108 226300 254160
rect 226352 254148 226358 254160
rect 229514 254148 229520 254160
rect 226352 254120 229520 254148
rect 226352 254108 226358 254120
rect 229514 254108 229520 254120
rect 229572 254108 229578 254160
rect 226294 253972 226300 254024
rect 226352 254012 226358 254024
rect 229606 254012 229612 254024
rect 226352 253984 229612 254012
rect 226352 253972 226358 253984
rect 229606 253972 229612 253984
rect 229664 253972 229670 254024
rect 84982 253768 84988 253820
rect 85040 253808 85046 253820
rect 87190 253808 87196 253820
rect 85040 253780 87196 253808
rect 85040 253768 85046 253780
rect 87190 253768 87196 253780
rect 87248 253768 87254 253820
rect 80106 253224 80112 253276
rect 80164 253264 80170 253276
rect 80164 253236 85764 253264
rect 80164 253224 80170 253236
rect 80198 253088 80204 253140
rect 80256 253128 80262 253140
rect 80256 253100 85672 253128
rect 80256 253088 80262 253100
rect 85644 252992 85672 253100
rect 85736 253060 85764 253236
rect 173210 253156 173216 253208
rect 173268 253196 173274 253208
rect 173268 253168 178500 253196
rect 173268 253156 173274 253168
rect 173486 253088 173492 253140
rect 173544 253128 173550 253140
rect 173544 253100 178408 253128
rect 173544 253088 173550 253100
rect 87190 253060 87196 253072
rect 85736 253032 87196 253060
rect 87190 253020 87196 253032
rect 87248 253020 87254 253072
rect 131442 253020 131448 253072
rect 131500 253060 131506 253072
rect 139814 253060 139820 253072
rect 131500 253032 139820 253060
rect 131500 253020 131506 253032
rect 139814 253020 139820 253032
rect 139872 253020 139878 253072
rect 87282 252992 87288 253004
rect 85644 252964 87288 252992
rect 87282 252952 87288 252964
rect 87340 252952 87346 253004
rect 131534 252952 131540 253004
rect 131592 252992 131598 253004
rect 139630 252992 139636 253004
rect 131592 252964 139636 252992
rect 131592 252952 131598 252964
rect 139630 252952 139636 252964
rect 139688 252952 139694 253004
rect 178380 252992 178408 253100
rect 178472 253060 178500 253168
rect 230618 253088 230624 253140
rect 230676 253128 230682 253140
rect 233654 253128 233660 253140
rect 230676 253100 233660 253128
rect 230676 253088 230682 253100
rect 233654 253088 233660 253100
rect 233712 253088 233718 253140
rect 182318 253060 182324 253072
rect 178472 253032 182324 253060
rect 182318 253020 182324 253032
rect 182376 253020 182382 253072
rect 226294 253020 226300 253072
rect 226352 253060 226358 253072
rect 233930 253060 233936 253072
rect 226352 253032 233936 253060
rect 226352 253020 226358 253032
rect 233930 253020 233936 253032
rect 233988 253020 233994 253072
rect 181398 252992 181404 253004
rect 178380 252964 181404 252992
rect 181398 252952 181404 252964
rect 181456 252952 181462 253004
rect 226386 252952 226392 253004
rect 226444 252992 226450 253004
rect 233562 252992 233568 253004
rect 226444 252964 233568 252992
rect 226444 252952 226450 252964
rect 233562 252952 233568 252964
rect 233620 252952 233626 253004
rect 131350 252884 131356 252936
rect 131408 252924 131414 252936
rect 139906 252924 139912 252936
rect 131408 252896 139912 252924
rect 131408 252884 131414 252896
rect 139906 252884 139912 252896
rect 139964 252884 139970 252936
rect 226294 252884 226300 252936
rect 226352 252924 226358 252936
rect 233746 252924 233752 252936
rect 226352 252896 233752 252924
rect 226352 252884 226358 252896
rect 233746 252884 233752 252896
rect 233804 252884 233810 252936
rect 225650 252816 225656 252868
rect 225708 252856 225714 252868
rect 233470 252856 233476 252868
rect 225708 252828 233476 252856
rect 225708 252816 225714 252828
rect 233470 252816 233476 252828
rect 233528 252816 233534 252868
rect 80198 252340 80204 252392
rect 80256 252380 80262 252392
rect 87190 252380 87196 252392
rect 80256 252352 87196 252380
rect 80256 252340 80262 252352
rect 87190 252340 87196 252352
rect 87248 252340 87254 252392
rect 131350 252340 131356 252392
rect 131408 252380 131414 252392
rect 140550 252380 140556 252392
rect 131408 252352 140556 252380
rect 131408 252340 131414 252352
rect 140550 252340 140556 252352
rect 140608 252340 140614 252392
rect 173578 252340 173584 252392
rect 173636 252380 173642 252392
rect 182318 252380 182324 252392
rect 173636 252352 182324 252380
rect 173636 252340 173642 252352
rect 182318 252340 182324 252352
rect 182376 252340 182382 252392
rect 80198 251728 80204 251780
rect 80256 251768 80262 251780
rect 80256 251740 85764 251768
rect 80256 251728 80262 251740
rect 85736 251632 85764 251740
rect 173486 251728 173492 251780
rect 173544 251768 173550 251780
rect 173544 251740 178316 251768
rect 173544 251728 173550 251740
rect 131350 251660 131356 251712
rect 131408 251700 131414 251712
rect 140182 251700 140188 251712
rect 131408 251672 140188 251700
rect 131408 251660 131414 251672
rect 140182 251660 140188 251672
rect 140240 251660 140246 251712
rect 178288 251700 178316 251740
rect 181766 251700 181772 251712
rect 178288 251672 181772 251700
rect 181766 251660 181772 251672
rect 181824 251660 181830 251712
rect 225374 251660 225380 251712
rect 225432 251700 225438 251712
rect 233562 251700 233568 251712
rect 225432 251672 233568 251700
rect 225432 251660 225438 251672
rect 233562 251660 233568 251672
rect 233620 251660 233626 251712
rect 87190 251632 87196 251644
rect 85736 251604 87196 251632
rect 87190 251592 87196 251604
rect 87248 251592 87254 251644
rect 226386 251592 226392 251644
rect 226444 251632 226450 251644
rect 233470 251632 233476 251644
rect 226444 251604 233476 251632
rect 226444 251592 226450 251604
rect 233470 251592 233476 251604
rect 233528 251592 233534 251644
rect 226294 251524 226300 251576
rect 226352 251564 226358 251576
rect 230618 251564 230624 251576
rect 226352 251536 230624 251564
rect 226352 251524 226358 251536
rect 230618 251524 230624 251536
rect 230676 251524 230682 251576
rect 80198 251048 80204 251100
rect 80256 251088 80262 251100
rect 87190 251088 87196 251100
rect 80256 251060 87196 251088
rect 80256 251048 80262 251060
rect 87190 251048 87196 251060
rect 87248 251048 87254 251100
rect 131350 251048 131356 251100
rect 131408 251088 131414 251100
rect 140642 251088 140648 251100
rect 131408 251060 140648 251088
rect 131408 251048 131414 251060
rect 140642 251048 140648 251060
rect 140700 251048 140706 251100
rect 173486 251048 173492 251100
rect 173544 251088 173550 251100
rect 182318 251088 182324 251100
rect 173544 251060 182324 251088
rect 173544 251048 173550 251060
rect 182318 251048 182324 251060
rect 182376 251048 182382 251100
rect 80106 250980 80112 251032
rect 80164 251020 80170 251032
rect 87282 251020 87288 251032
rect 80164 250992 87288 251020
rect 80164 250980 80170 250992
rect 87282 250980 87288 250992
rect 87340 250980 87346 251032
rect 131442 250980 131448 251032
rect 131500 251020 131506 251032
rect 140550 251020 140556 251032
rect 131500 250992 140556 251020
rect 131500 250980 131506 250992
rect 140550 250980 140556 250992
rect 140608 250980 140614 251032
rect 173578 250980 173584 251032
rect 173636 251020 173642 251032
rect 182226 251020 182232 251032
rect 173636 250992 182232 251020
rect 173636 250980 173642 250992
rect 182226 250980 182232 250992
rect 182284 250980 182290 251032
rect 175329 250343 175387 250349
rect 175329 250309 175341 250343
rect 175375 250340 175387 250343
rect 175418 250340 175424 250352
rect 175375 250312 175424 250340
rect 175375 250309 175387 250312
rect 175329 250303 175387 250309
rect 175418 250300 175424 250312
rect 175476 250300 175482 250352
rect 131350 250232 131356 250284
rect 131408 250272 131414 250284
rect 140550 250272 140556 250284
rect 131408 250244 140556 250272
rect 131408 250232 131414 250244
rect 140550 250232 140556 250244
rect 140608 250232 140614 250284
rect 226294 250232 226300 250284
rect 226352 250272 226358 250284
rect 233562 250272 233568 250284
rect 226352 250244 233568 250272
rect 226352 250232 226358 250244
rect 233562 250232 233568 250244
rect 233620 250232 233626 250284
rect 225926 250164 225932 250216
rect 225984 250204 225990 250216
rect 233470 250204 233476 250216
rect 225984 250176 233476 250204
rect 225984 250164 225990 250176
rect 233470 250164 233476 250176
rect 233528 250164 233534 250216
rect 80106 249620 80112 249672
rect 80164 249660 80170 249672
rect 87190 249660 87196 249672
rect 80164 249632 87196 249660
rect 80164 249620 80170 249632
rect 87190 249620 87196 249632
rect 87248 249620 87254 249672
rect 131810 249620 131816 249672
rect 131868 249660 131874 249672
rect 140458 249660 140464 249672
rect 131868 249632 140464 249660
rect 131868 249620 131874 249632
rect 140458 249620 140464 249632
rect 140516 249620 140522 249672
rect 173578 249620 173584 249672
rect 173636 249660 173642 249672
rect 182318 249660 182324 249672
rect 173636 249632 182324 249660
rect 173636 249620 173642 249632
rect 182318 249620 182324 249632
rect 182376 249620 182382 249672
rect 225558 249620 225564 249672
rect 225616 249660 225622 249672
rect 233562 249660 233568 249672
rect 225616 249632 233568 249660
rect 225616 249620 225622 249632
rect 233562 249620 233568 249632
rect 233620 249620 233626 249672
rect 80198 249552 80204 249604
rect 80256 249592 80262 249604
rect 87282 249592 87288 249604
rect 80256 249564 87288 249592
rect 80256 249552 80262 249564
rect 87282 249552 87288 249564
rect 87340 249552 87346 249604
rect 131350 249552 131356 249604
rect 131408 249592 131414 249604
rect 139998 249592 140004 249604
rect 131408 249564 140004 249592
rect 131408 249552 131414 249564
rect 139998 249552 140004 249564
rect 140056 249552 140062 249604
rect 173670 249552 173676 249604
rect 173728 249592 173734 249604
rect 182226 249592 182232 249604
rect 173728 249564 182232 249592
rect 173728 249552 173734 249564
rect 182226 249552 182232 249564
rect 182284 249552 182290 249604
rect 226294 249552 226300 249604
rect 226352 249592 226358 249604
rect 233470 249592 233476 249604
rect 226352 249564 233476 249592
rect 226352 249552 226358 249564
rect 233470 249552 233476 249564
rect 233528 249552 233534 249604
rect 131350 248940 131356 248992
rect 131408 248980 131414 248992
rect 131408 248952 137560 248980
rect 131408 248940 131414 248952
rect 79278 248872 79284 248924
rect 79336 248912 79342 248924
rect 87190 248912 87196 248924
rect 79336 248884 87196 248912
rect 79336 248872 79342 248884
rect 87190 248872 87196 248884
rect 87248 248872 87254 248924
rect 137532 248912 137560 248952
rect 140366 248912 140372 248924
rect 137532 248884 140372 248912
rect 140366 248872 140372 248884
rect 140424 248872 140430 248924
rect 173210 248872 173216 248924
rect 173268 248912 173274 248924
rect 181582 248912 181588 248924
rect 173268 248884 181588 248912
rect 173268 248872 173274 248884
rect 181582 248872 181588 248884
rect 181640 248872 181646 248924
rect 80198 248804 80204 248856
rect 80256 248844 80262 248856
rect 87374 248844 87380 248856
rect 80256 248816 87380 248844
rect 80256 248804 80262 248816
rect 87374 248804 87380 248816
rect 87432 248804 87438 248856
rect 173578 248804 173584 248856
rect 173636 248844 173642 248856
rect 182318 248844 182324 248856
rect 173636 248816 182324 248844
rect 173636 248804 173642 248816
rect 182318 248804 182324 248816
rect 182376 248804 182382 248856
rect 226294 248260 226300 248312
rect 226352 248300 226358 248312
rect 233562 248300 233568 248312
rect 226352 248272 233568 248300
rect 226352 248260 226358 248272
rect 233562 248260 233568 248272
rect 233620 248260 233626 248312
rect 131350 248192 131356 248244
rect 131408 248232 131414 248244
rect 140366 248232 140372 248244
rect 131408 248204 140372 248232
rect 131408 248192 131414 248204
rect 140366 248192 140372 248204
rect 140424 248192 140430 248244
rect 226386 248192 226392 248244
rect 226444 248232 226450 248244
rect 233470 248232 233476 248244
rect 226444 248204 233476 248232
rect 226444 248192 226450 248204
rect 233470 248192 233476 248204
rect 233528 248192 233534 248244
rect 85902 247716 85908 247768
rect 85960 247756 85966 247768
rect 88018 247756 88024 247768
rect 85960 247728 88024 247756
rect 85960 247716 85966 247728
rect 88018 247716 88024 247728
rect 88076 247716 88082 247768
rect 131810 247716 131816 247768
rect 131868 247756 131874 247768
rect 137054 247756 137060 247768
rect 131868 247728 137060 247756
rect 131868 247716 131874 247728
rect 137054 247716 137060 247728
rect 137112 247716 137118 247768
rect 132546 247648 132552 247700
rect 132604 247688 132610 247700
rect 137514 247688 137520 247700
rect 132604 247660 137520 247688
rect 132604 247648 132610 247660
rect 137514 247648 137520 247660
rect 137572 247648 137578 247700
rect 226294 247648 226300 247700
rect 226352 247688 226358 247700
rect 234390 247688 234396 247700
rect 226352 247660 234396 247688
rect 226352 247648 226358 247660
rect 234390 247648 234396 247660
rect 234448 247648 234454 247700
rect 86086 247580 86092 247632
rect 86144 247620 86150 247632
rect 87190 247620 87196 247632
rect 86144 247592 87196 247620
rect 86144 247580 86150 247592
rect 87190 247580 87196 247592
rect 87248 247580 87254 247632
rect 131442 247580 131448 247632
rect 131500 247620 131506 247632
rect 131500 247592 138204 247620
rect 131500 247580 131506 247592
rect 79278 247512 79284 247564
rect 79336 247552 79342 247564
rect 88386 247552 88392 247564
rect 79336 247524 88392 247552
rect 79336 247512 79342 247524
rect 88386 247512 88392 247524
rect 88444 247512 88450 247564
rect 138176 247552 138204 247592
rect 226386 247580 226392 247632
rect 226444 247620 226450 247632
rect 234482 247620 234488 247632
rect 226444 247592 234488 247620
rect 226444 247580 226450 247592
rect 234482 247580 234488 247592
rect 234540 247580 234546 247632
rect 140366 247552 140372 247564
rect 138176 247524 140372 247552
rect 140366 247512 140372 247524
rect 140424 247512 140430 247564
rect 173210 247512 173216 247564
rect 173268 247552 173274 247564
rect 181122 247552 181128 247564
rect 173268 247524 181128 247552
rect 173268 247512 173274 247524
rect 181122 247512 181128 247524
rect 181180 247512 181186 247564
rect 80198 247444 80204 247496
rect 80256 247484 80262 247496
rect 88294 247484 88300 247496
rect 80256 247456 88300 247484
rect 80256 247444 80262 247456
rect 88294 247444 88300 247456
rect 88352 247444 88358 247496
rect 173578 247444 173584 247496
rect 173636 247484 173642 247496
rect 181030 247484 181036 247496
rect 173636 247456 181036 247484
rect 173636 247444 173642 247456
rect 181030 247444 181036 247456
rect 181088 247444 181094 247496
rect 137514 247240 137520 247292
rect 137572 247280 137578 247292
rect 140642 247280 140648 247292
rect 137572 247252 140648 247280
rect 137572 247240 137578 247252
rect 140642 247240 140648 247252
rect 140700 247240 140706 247292
rect 80014 246356 80020 246408
rect 80072 246396 80078 246408
rect 87190 246396 87196 246408
rect 80072 246368 87196 246396
rect 80072 246356 80078 246368
rect 87190 246356 87196 246368
rect 87248 246356 87254 246408
rect 131442 246356 131448 246408
rect 131500 246396 131506 246408
rect 137238 246396 137244 246408
rect 131500 246368 137244 246396
rect 131500 246356 131506 246368
rect 137238 246356 137244 246368
rect 137296 246356 137302 246408
rect 173946 246356 173952 246408
rect 174004 246396 174010 246408
rect 182318 246396 182324 246408
rect 174004 246368 182324 246396
rect 174004 246356 174010 246368
rect 182318 246356 182324 246368
rect 182376 246356 182382 246408
rect 226294 246356 226300 246408
rect 226352 246396 226358 246408
rect 233654 246396 233660 246408
rect 226352 246368 233660 246396
rect 226352 246356 226358 246368
rect 233654 246356 233660 246368
rect 233712 246356 233718 246408
rect 132178 246288 132184 246340
rect 132236 246328 132242 246340
rect 140642 246328 140648 246340
rect 132236 246300 140648 246328
rect 132236 246288 132242 246300
rect 140642 246288 140648 246300
rect 140700 246288 140706 246340
rect 226386 246288 226392 246340
rect 226444 246328 226450 246340
rect 233562 246328 233568 246340
rect 226444 246300 233568 246328
rect 226444 246288 226450 246300
rect 233562 246288 233568 246300
rect 233620 246288 233626 246340
rect 131350 246220 131356 246272
rect 131408 246260 131414 246272
rect 140182 246260 140188 246272
rect 131408 246232 140188 246260
rect 131408 246220 131414 246232
rect 140182 246220 140188 246232
rect 140240 246220 140246 246272
rect 225650 246220 225656 246272
rect 225708 246260 225714 246272
rect 233470 246260 233476 246272
rect 225708 246232 233476 246260
rect 225708 246220 225714 246232
rect 233470 246220 233476 246232
rect 233528 246220 233534 246272
rect 79278 246152 79284 246204
rect 79336 246192 79342 246204
rect 86086 246192 86092 246204
rect 79336 246164 86092 246192
rect 79336 246152 79342 246164
rect 86086 246152 86092 246164
rect 86144 246152 86150 246204
rect 137054 246084 137060 246136
rect 137112 246124 137118 246136
rect 140550 246124 140556 246136
rect 137112 246096 140556 246124
rect 137112 246084 137118 246096
rect 140550 246084 140556 246096
rect 140608 246084 140614 246136
rect 173578 246084 173584 246136
rect 173636 246124 173642 246136
rect 180846 246124 180852 246136
rect 173636 246096 180852 246124
rect 173636 246084 173642 246096
rect 180846 246084 180852 246096
rect 180904 246084 180910 246136
rect 137238 245948 137244 246000
rect 137296 245988 137302 246000
rect 140366 245988 140372 246000
rect 137296 245960 140372 245988
rect 137296 245948 137302 245960
rect 140366 245948 140372 245960
rect 140424 245948 140430 246000
rect 80198 245880 80204 245932
rect 80256 245920 80262 245932
rect 85902 245920 85908 245932
rect 80256 245892 85908 245920
rect 80256 245880 80262 245892
rect 85902 245880 85908 245892
rect 85960 245880 85966 245932
rect 173486 245676 173492 245728
rect 173544 245716 173550 245728
rect 180938 245716 180944 245728
rect 173544 245688 180944 245716
rect 173544 245676 173550 245688
rect 180938 245676 180944 245688
rect 180996 245676 181002 245728
rect 225558 245200 225564 245252
rect 225616 245240 225622 245252
rect 227950 245240 227956 245252
rect 225616 245212 227956 245240
rect 225616 245200 225622 245212
rect 227950 245200 227956 245212
rect 228008 245200 228014 245252
rect 131810 244996 131816 245048
rect 131868 245036 131874 245048
rect 135950 245036 135956 245048
rect 131868 245008 135956 245036
rect 131868 244996 131874 245008
rect 135950 244996 135956 245008
rect 136008 244996 136014 245048
rect 131350 244928 131356 244980
rect 131408 244968 131414 244980
rect 135858 244968 135864 244980
rect 131408 244940 135864 244968
rect 131408 244928 131414 244940
rect 135858 244928 135864 244940
rect 135916 244928 135922 244980
rect 226202 244928 226208 244980
rect 226260 244968 226266 244980
rect 228042 244968 228048 244980
rect 226260 244940 228048 244968
rect 226260 244928 226266 244940
rect 228042 244928 228048 244940
rect 228100 244928 228106 244980
rect 131994 244860 132000 244912
rect 132052 244900 132058 244912
rect 139630 244900 139636 244912
rect 132052 244872 139636 244900
rect 132052 244860 132058 244872
rect 139630 244860 139636 244872
rect 139688 244860 139694 244912
rect 226386 244860 226392 244912
rect 226444 244900 226450 244912
rect 228134 244900 228140 244912
rect 226444 244872 228140 244900
rect 226444 244860 226450 244872
rect 228134 244860 228140 244872
rect 228192 244860 228198 244912
rect 131442 244792 131448 244844
rect 131500 244832 131506 244844
rect 139722 244832 139728 244844
rect 131500 244804 139728 244832
rect 131500 244792 131506 244804
rect 139722 244792 139728 244804
rect 139780 244792 139786 244844
rect 226294 244792 226300 244844
rect 226352 244832 226358 244844
rect 233470 244832 233476 244844
rect 226352 244804 233476 244832
rect 226352 244792 226358 244804
rect 233470 244792 233476 244804
rect 233528 244792 233534 244844
rect 80106 244724 80112 244776
rect 80164 244764 80170 244776
rect 87098 244764 87104 244776
rect 80164 244736 87104 244764
rect 80164 244724 80170 244736
rect 87098 244724 87104 244736
rect 87156 244724 87162 244776
rect 173578 244724 173584 244776
rect 173636 244764 173642 244776
rect 180754 244764 180760 244776
rect 173636 244736 180760 244764
rect 173636 244724 173642 244736
rect 180754 244724 180760 244736
rect 180812 244724 180818 244776
rect 80198 244656 80204 244708
rect 80256 244696 80262 244708
rect 87006 244696 87012 244708
rect 80256 244668 87012 244696
rect 80256 244656 80262 244668
rect 87006 244656 87012 244668
rect 87064 244656 87070 244708
rect 172842 244656 172848 244708
rect 172900 244696 172906 244708
rect 180662 244696 180668 244708
rect 172900 244668 180668 244696
rect 172900 244656 172906 244668
rect 180662 244656 180668 244668
rect 180720 244656 180726 244708
rect 131350 243636 131356 243688
rect 131408 243676 131414 243688
rect 136778 243676 136784 243688
rect 131408 243648 136784 243676
rect 131408 243636 131414 243648
rect 136778 243636 136784 243648
rect 136836 243636 136842 243688
rect 131442 243568 131448 243620
rect 131500 243608 131506 243620
rect 136686 243608 136692 243620
rect 131500 243580 136692 243608
rect 131500 243568 131506 243580
rect 136686 243568 136692 243580
rect 136744 243568 136750 243620
rect 175329 243611 175387 243617
rect 175329 243577 175341 243611
rect 175375 243608 175387 243611
rect 175418 243608 175424 243620
rect 175375 243580 175424 243608
rect 175375 243577 175387 243580
rect 175329 243571 175387 243577
rect 175418 243568 175424 243580
rect 175476 243568 175482 243620
rect 225742 243568 225748 243620
rect 225800 243608 225806 243620
rect 233654 243608 233660 243620
rect 225800 243580 233660 243608
rect 225800 243568 225806 243580
rect 233654 243568 233660 243580
rect 233712 243568 233718 243620
rect 79922 243500 79928 243552
rect 79980 243540 79986 243552
rect 87190 243540 87196 243552
rect 79980 243512 87196 243540
rect 79980 243500 79986 243512
rect 87190 243500 87196 243512
rect 87248 243500 87254 243552
rect 131534 243500 131540 243552
rect 131592 243540 131598 243552
rect 139354 243540 139360 243552
rect 131592 243512 139360 243540
rect 131592 243500 131598 243512
rect 139354 243500 139360 243512
rect 139412 243500 139418 243552
rect 173854 243500 173860 243552
rect 173912 243540 173918 243552
rect 181214 243540 181220 243552
rect 173912 243512 181220 243540
rect 173912 243500 173918 243512
rect 181214 243500 181220 243512
rect 181272 243500 181278 243552
rect 226202 243500 226208 243552
rect 226260 243540 226266 243552
rect 233838 243540 233844 243552
rect 226260 243512 233844 243540
rect 226260 243500 226266 243512
rect 233838 243500 233844 243512
rect 233896 243500 233902 243552
rect 80106 243432 80112 243484
rect 80164 243472 80170 243484
rect 87282 243472 87288 243484
rect 80164 243444 87288 243472
rect 80164 243432 80170 243444
rect 87282 243432 87288 243444
rect 87340 243432 87346 243484
rect 131626 243432 131632 243484
rect 131684 243472 131690 243484
rect 139538 243472 139544 243484
rect 131684 243444 139544 243472
rect 131684 243432 131690 243444
rect 139538 243432 139544 243444
rect 139596 243432 139602 243484
rect 173486 243432 173492 243484
rect 173544 243472 173550 243484
rect 182318 243472 182324 243484
rect 173544 243444 182324 243472
rect 173544 243432 173550 243444
rect 182318 243432 182324 243444
rect 182376 243432 182382 243484
rect 226294 243432 226300 243484
rect 226352 243472 226358 243484
rect 233746 243472 233752 243484
rect 226352 243444 233752 243472
rect 226352 243432 226358 243444
rect 233746 243432 233752 243444
rect 233804 243432 233810 243484
rect 80198 243364 80204 243416
rect 80256 243404 80262 243416
rect 86914 243404 86920 243416
rect 80256 243376 86920 243404
rect 80256 243364 80262 243376
rect 86914 243364 86920 243376
rect 86972 243364 86978 243416
rect 175326 243404 175332 243416
rect 175287 243376 175332 243404
rect 175326 243364 175332 243376
rect 175384 243364 175390 243416
rect 228042 243364 228048 243416
rect 228100 243404 228106 243416
rect 233470 243404 233476 243416
rect 228100 243376 233476 243404
rect 228100 243364 228106 243376
rect 233470 243364 233476 243376
rect 233528 243364 233534 243416
rect 227950 243296 227956 243348
rect 228008 243336 228014 243348
rect 233562 243336 233568 243348
rect 228008 243308 233568 243336
rect 228008 243296 228014 243308
rect 233562 243296 233568 243308
rect 233620 243296 233626 243348
rect 173578 243160 173584 243212
rect 173636 243200 173642 243212
rect 180846 243200 180852 243212
rect 173636 243172 180852 243200
rect 173636 243160 173642 243172
rect 180846 243160 180852 243172
rect 180904 243160 180910 243212
rect 80198 242752 80204 242804
rect 80256 242792 80262 242804
rect 86822 242792 86828 242804
rect 80256 242764 86828 242792
rect 80256 242752 80262 242764
rect 86822 242752 86828 242764
rect 86880 242752 86886 242804
rect 172842 242752 172848 242804
rect 172900 242792 172906 242804
rect 180938 242792 180944 242804
rect 172900 242764 180944 242792
rect 172900 242752 172906 242764
rect 180938 242752 180944 242764
rect 180996 242752 181002 242804
rect 79278 242208 79284 242260
rect 79336 242248 79342 242260
rect 87190 242248 87196 242260
rect 79336 242220 87196 242248
rect 79336 242208 79342 242220
rect 87190 242208 87196 242220
rect 87248 242208 87254 242260
rect 131350 242208 131356 242260
rect 131408 242248 131414 242260
rect 136134 242248 136140 242260
rect 131408 242220 136140 242248
rect 131408 242208 131414 242220
rect 136134 242208 136140 242220
rect 136192 242208 136198 242260
rect 173762 242208 173768 242260
rect 173820 242248 173826 242260
rect 182318 242248 182324 242260
rect 173820 242220 182324 242248
rect 173820 242208 173826 242220
rect 182318 242208 182324 242220
rect 182376 242208 182382 242260
rect 226018 242208 226024 242260
rect 226076 242248 226082 242260
rect 228686 242248 228692 242260
rect 226076 242220 228692 242248
rect 226076 242208 226082 242220
rect 228686 242208 228692 242220
rect 228744 242208 228750 242260
rect 131442 242140 131448 242192
rect 131500 242180 131506 242192
rect 136226 242180 136232 242192
rect 131500 242152 136232 242180
rect 131500 242140 131506 242152
rect 136226 242140 136232 242152
rect 136284 242140 136290 242192
rect 226294 242140 226300 242192
rect 226352 242180 226358 242192
rect 226352 242152 228732 242180
rect 226352 242140 226358 242152
rect 131534 242072 131540 242124
rect 131592 242112 131598 242124
rect 139446 242112 139452 242124
rect 131592 242084 139452 242112
rect 131592 242072 131598 242084
rect 139446 242072 139452 242084
rect 139504 242072 139510 242124
rect 226386 242072 226392 242124
rect 226444 242112 226450 242124
rect 228594 242112 228600 242124
rect 226444 242084 228600 242112
rect 226444 242072 226450 242084
rect 228594 242072 228600 242084
rect 228652 242072 228658 242124
rect 228704 242112 228732 242152
rect 233562 242112 233568 242124
rect 228704 242084 233568 242112
rect 233562 242072 233568 242084
rect 233620 242072 233626 242124
rect 79094 242004 79100 242056
rect 79152 242044 79158 242056
rect 87558 242044 87564 242056
rect 79152 242016 87564 242044
rect 79152 242004 79158 242016
rect 87558 242004 87564 242016
rect 87616 242004 87622 242056
rect 135858 242004 135864 242056
rect 135916 242044 135922 242056
rect 140550 242044 140556 242056
rect 135916 242016 140556 242044
rect 135916 242004 135922 242016
rect 140550 242004 140556 242016
rect 140608 242004 140614 242056
rect 173578 242004 173584 242056
rect 173636 242044 173642 242056
rect 182226 242044 182232 242056
rect 173636 242016 182232 242044
rect 173636 242004 173642 242016
rect 182226 242004 182232 242016
rect 182284 242004 182290 242056
rect 228134 242004 228140 242056
rect 228192 242044 228198 242056
rect 233470 242044 233476 242056
rect 228192 242016 233476 242044
rect 228192 242004 228198 242016
rect 233470 242004 233476 242016
rect 233528 242004 233534 242056
rect 264750 242004 264756 242056
rect 264808 242044 264814 242056
rect 300170 242044 300176 242056
rect 264808 242016 300176 242044
rect 264808 242004 264814 242016
rect 300170 242004 300176 242016
rect 300228 242004 300234 242056
rect 80198 241936 80204 241988
rect 80256 241976 80262 241988
rect 87650 241976 87656 241988
rect 80256 241948 87656 241976
rect 80256 241936 80262 241948
rect 87650 241936 87656 241948
rect 87708 241936 87714 241988
rect 135950 241936 135956 241988
rect 136008 241976 136014 241988
rect 140182 241976 140188 241988
rect 136008 241948 140188 241976
rect 136008 241936 136014 241948
rect 140182 241936 140188 241948
rect 140240 241936 140246 241988
rect 173670 241936 173676 241988
rect 173728 241976 173734 241988
rect 182042 241976 182048 241988
rect 173728 241948 182048 241976
rect 173728 241936 173734 241948
rect 182042 241936 182048 241948
rect 182100 241936 182106 241988
rect 178914 240712 178920 240764
rect 178972 240752 178978 240764
rect 181582 240752 181588 240764
rect 178972 240724 181588 240752
rect 178972 240712 178978 240724
rect 181582 240712 181588 240724
rect 181640 240712 181646 240764
rect 85074 240644 85080 240696
rect 85132 240684 85138 240696
rect 87374 240684 87380 240696
rect 85132 240656 87380 240684
rect 85132 240644 85138 240656
rect 87374 240644 87380 240656
rect 87432 240644 87438 240696
rect 131350 240644 131356 240696
rect 131408 240684 131414 240696
rect 139262 240684 139268 240696
rect 131408 240656 139268 240684
rect 131408 240644 131414 240656
rect 139262 240644 139268 240656
rect 139320 240644 139326 240696
rect 226018 240644 226024 240696
rect 226076 240684 226082 240696
rect 234114 240684 234120 240696
rect 226076 240656 234120 240684
rect 226076 240644 226082 240656
rect 234114 240644 234120 240656
rect 234172 240644 234178 240696
rect 109914 240440 109920 240492
rect 109972 240480 109978 240492
rect 141010 240480 141016 240492
rect 109972 240452 141016 240480
rect 109972 240440 109978 240452
rect 141010 240440 141016 240452
rect 141068 240440 141074 240492
rect 203110 239760 203116 239812
rect 203168 239800 203174 239812
rect 203846 239800 203852 239812
rect 203168 239772 203852 239800
rect 203168 239760 203174 239772
rect 203846 239760 203852 239772
rect 203904 239760 203910 239812
rect 80198 239216 80204 239268
rect 80256 239256 80262 239268
rect 87466 239256 87472 239268
rect 80256 239228 87472 239256
rect 80256 239216 80262 239228
rect 87466 239216 87472 239228
rect 87524 239216 87530 239268
rect 136778 239216 136784 239268
rect 136836 239256 136842 239268
rect 140550 239256 140556 239268
rect 136836 239228 140556 239256
rect 136836 239216 136842 239228
rect 140550 239216 140556 239228
rect 140608 239216 140614 239268
rect 173670 239216 173676 239268
rect 173728 239256 173734 239268
rect 182134 239256 182140 239268
rect 173728 239228 182140 239256
rect 173728 239216 173734 239228
rect 182134 239216 182140 239228
rect 182192 239216 182198 239268
rect 226570 239216 226576 239268
rect 226628 239256 226634 239268
rect 233470 239256 233476 239268
rect 226628 239228 233476 239256
rect 226628 239216 226634 239228
rect 233470 239216 233476 239228
rect 233528 239216 233534 239268
rect 136686 239148 136692 239200
rect 136744 239188 136750 239200
rect 140642 239188 140648 239200
rect 136744 239160 140648 239188
rect 136744 239148 136750 239160
rect 140642 239148 140648 239160
rect 140700 239148 140706 239200
rect 80198 237856 80204 237908
rect 80256 237896 80262 237908
rect 86546 237896 86552 237908
rect 80256 237868 86552 237896
rect 80256 237856 80262 237868
rect 86546 237856 86552 237868
rect 86604 237856 86610 237908
rect 228686 237856 228692 237908
rect 228744 237896 228750 237908
rect 233470 237896 233476 237908
rect 228744 237868 233476 237896
rect 228744 237856 228750 237868
rect 233470 237856 233476 237868
rect 233528 237856 233534 237908
rect 136226 237788 136232 237840
rect 136284 237828 136290 237840
rect 140550 237828 140556 237840
rect 136284 237800 140556 237828
rect 136284 237788 136290 237800
rect 140550 237788 140556 237800
rect 140608 237788 140614 237840
rect 228594 237788 228600 237840
rect 228652 237828 228658 237840
rect 233562 237828 233568 237840
rect 228652 237800 233568 237828
rect 228652 237788 228658 237800
rect 233562 237788 233568 237800
rect 233620 237788 233626 237840
rect 136134 237516 136140 237568
rect 136192 237556 136198 237568
rect 140274 237556 140280 237568
rect 136192 237528 140280 237556
rect 136192 237516 136198 237528
rect 140274 237516 140280 237528
rect 140332 237516 140338 237568
rect 173578 237380 173584 237432
rect 173636 237420 173642 237432
rect 180386 237420 180392 237432
rect 173636 237392 180392 237420
rect 173636 237380 173642 237392
rect 180386 237380 180392 237392
rect 180444 237380 180450 237432
rect 80198 237312 80204 237364
rect 80256 237352 80262 237364
rect 86454 237352 86460 237364
rect 80256 237324 86460 237352
rect 80256 237312 80262 237324
rect 86454 237312 86460 237324
rect 86512 237312 86518 237364
rect 173394 236904 173400 236956
rect 173452 236944 173458 236956
rect 180294 236944 180300 236956
rect 173452 236916 180300 236944
rect 173452 236904 173458 236916
rect 180294 236904 180300 236916
rect 180352 236904 180358 236956
rect 173578 236496 173584 236548
rect 173636 236536 173642 236548
rect 178914 236536 178920 236548
rect 173636 236508 178920 236536
rect 173636 236496 173642 236508
rect 178914 236496 178920 236508
rect 178972 236496 178978 236548
rect 80198 235272 80204 235324
rect 80256 235312 80262 235324
rect 85074 235312 85080 235324
rect 80256 235284 85080 235312
rect 80256 235272 80262 235284
rect 85074 235272 85080 235284
rect 85132 235272 85138 235324
rect 154813 233819 154871 233825
rect 154813 233785 154825 233819
rect 154859 233816 154871 233819
rect 164381 233819 164439 233825
rect 164381 233816 164393 233819
rect 154859 233788 164393 233816
rect 154859 233785 154871 233788
rect 154813 233779 154871 233785
rect 164381 233785 164393 233788
rect 164427 233785 164439 233819
rect 164381 233779 164439 233785
rect 151774 233708 151780 233760
rect 151832 233748 151838 233760
rect 163182 233748 163188 233760
rect 151832 233720 163188 233748
rect 151832 233708 151838 233720
rect 163182 233708 163188 233720
rect 163240 233708 163246 233760
rect 249110 233708 249116 233760
rect 249168 233748 249174 233760
rect 259230 233748 259236 233760
rect 249168 233720 259236 233748
rect 249168 233708 249174 233720
rect 259230 233708 259236 233720
rect 259288 233708 259294 233760
rect 60878 233640 60884 233692
rect 60936 233680 60942 233692
rect 60936 233652 66444 233680
rect 60936 233640 60942 233652
rect 60142 233572 60148 233624
rect 60200 233612 60206 233624
rect 66416 233612 66444 233652
rect 154902 233640 154908 233692
rect 154960 233680 154966 233692
rect 167874 233680 167880 233692
rect 154960 233652 167880 233680
rect 154960 233640 154966 233652
rect 167874 233640 167880 233652
rect 167932 233640 167938 233692
rect 249294 233640 249300 233692
rect 249352 233680 249358 233692
rect 255737 233683 255795 233689
rect 255737 233680 255749 233683
rect 249352 233652 255749 233680
rect 249352 233640 249358 233652
rect 255737 233649 255749 233652
rect 255783 233649 255795 233683
rect 259782 233680 259788 233692
rect 255737 233643 255795 233649
rect 255844 233652 259788 233680
rect 71642 233612 71648 233624
rect 60200 233584 66352 233612
rect 66416 233584 71648 233612
rect 60200 233572 60206 233584
rect 57934 233504 57940 233556
rect 57992 233544 57998 233556
rect 66214 233544 66220 233556
rect 57992 233516 66220 233544
rect 57992 233504 57998 233516
rect 66214 233504 66220 233516
rect 66272 233504 66278 233556
rect 60602 233436 60608 233488
rect 60660 233476 60666 233488
rect 66324 233476 66352 233584
rect 71642 233572 71648 233584
rect 71700 233572 71706 233624
rect 154626 233572 154632 233624
rect 154684 233612 154690 233624
rect 154813 233615 154871 233621
rect 154813 233612 154825 233615
rect 154684 233584 154825 233612
rect 154684 233572 154690 233584
rect 154813 233581 154825 233584
rect 154859 233581 154871 233615
rect 154813 233575 154871 233581
rect 247730 233572 247736 233624
rect 247788 233612 247794 233624
rect 255844 233612 255872 233652
rect 259782 233640 259788 233652
rect 259840 233640 259846 233692
rect 247788 233584 255872 233612
rect 247788 233572 247794 233584
rect 138158 233504 138164 233556
rect 138216 233544 138222 233556
rect 142850 233544 142856 233556
rect 138216 233516 142856 233544
rect 138216 233504 138222 233516
rect 142850 233504 142856 233516
rect 142908 233504 142914 233556
rect 153154 233504 153160 233556
rect 153212 233544 153218 233556
rect 153212 233516 156512 233544
rect 153212 233504 153218 233516
rect 72378 233476 72384 233488
rect 60660 233448 61200 233476
rect 66324 233448 72384 233476
rect 60660 233436 60666 233448
rect 61172 233340 61200 233448
rect 72378 233436 72384 233448
rect 72436 233436 72442 233488
rect 137974 233436 137980 233488
rect 138032 233476 138038 233488
rect 143954 233476 143960 233488
rect 138032 233448 143960 233476
rect 138032 233436 138038 233448
rect 143954 233436 143960 233448
rect 144012 233436 144018 233488
rect 61246 233368 61252 233420
rect 61304 233408 61310 233420
rect 74402 233408 74408 233420
rect 61304 233380 74408 233408
rect 61304 233368 61310 233380
rect 74402 233368 74408 233380
rect 74460 233368 74466 233420
rect 137882 233368 137888 233420
rect 137940 233408 137946 233420
rect 144598 233408 144604 233420
rect 137940 233380 144604 233408
rect 137940 233368 137946 233380
rect 144598 233368 144604 233380
rect 144656 233368 144662 233420
rect 153246 233368 153252 233420
rect 153304 233408 153310 233420
rect 156484 233408 156512 233516
rect 159502 233504 159508 233556
rect 159560 233544 159566 233556
rect 162078 233544 162084 233556
rect 159560 233516 162084 233544
rect 159560 233504 159566 233516
rect 162078 233504 162084 233516
rect 162136 233504 162142 233556
rect 248650 233504 248656 233556
rect 248708 233544 248714 233556
rect 255826 233544 255832 233556
rect 248708 233516 255832 233544
rect 248708 233504 248714 233516
rect 255826 233504 255832 233516
rect 255884 233504 255890 233556
rect 255921 233547 255979 233553
rect 255921 233513 255933 233547
rect 255967 233544 255979 233547
rect 261990 233544 261996 233556
rect 255967 233516 261996 233544
rect 255967 233513 255979 233516
rect 255921 233507 255979 233513
rect 261990 233504 261996 233516
rect 262048 233504 262054 233556
rect 164381 233479 164439 233485
rect 164381 233445 164393 233479
rect 164427 233476 164439 233479
rect 166678 233476 166684 233488
rect 164427 233448 166684 233476
rect 164427 233445 164439 233448
rect 164381 233439 164439 233445
rect 166678 233436 166684 233448
rect 166736 233436 166742 233488
rect 248926 233436 248932 233488
rect 248984 233476 248990 233488
rect 261438 233476 261444 233488
rect 248984 233448 261444 233476
rect 248984 233436 248990 233448
rect 261438 233436 261444 233448
rect 261496 233436 261502 233488
rect 164930 233408 164936 233420
rect 153304 233380 156328 233408
rect 156484 233380 164936 233408
rect 153304 233368 153310 233380
rect 61172 233312 65616 233340
rect 57658 233232 57664 233284
rect 57716 233272 57722 233284
rect 65478 233272 65484 233284
rect 57716 233244 65484 233272
rect 57716 233232 57722 233244
rect 65478 233232 65484 233244
rect 65536 233232 65542 233284
rect 65588 233272 65616 233312
rect 154534 233300 154540 233352
rect 154592 233340 154598 233352
rect 156098 233340 156104 233352
rect 154592 233312 156104 233340
rect 154592 233300 154598 233312
rect 156098 233300 156104 233312
rect 156156 233300 156162 233352
rect 156193 233343 156251 233349
rect 156193 233309 156205 233343
rect 156239 233309 156251 233343
rect 156193 233303 156251 233309
rect 73022 233272 73028 233284
rect 65588 233244 73028 233272
rect 73022 233232 73028 233244
rect 73080 233232 73086 233284
rect 138066 233232 138072 233284
rect 138124 233272 138130 233284
rect 143770 233272 143776 233284
rect 138124 233244 143776 233272
rect 138124 233232 138130 233244
rect 143770 233232 143776 233244
rect 143828 233232 143834 233284
rect 153706 233232 153712 233284
rect 153764 233272 153770 233284
rect 156208 233272 156236 233303
rect 153764 233244 156236 233272
rect 156300 233272 156328 233380
rect 164930 233368 164936 233380
rect 164988 233368 164994 233420
rect 249018 233368 249024 233420
rect 249076 233408 249082 233420
rect 255550 233408 255556 233420
rect 249076 233380 255556 233408
rect 249076 233368 249082 233380
rect 255550 233368 255556 233380
rect 255608 233368 255614 233420
rect 156377 233343 156435 233349
rect 156377 233309 156389 233343
rect 156423 233340 156435 233343
rect 166126 233340 166132 233352
rect 156423 233312 166132 233340
rect 156423 233309 156435 233312
rect 156377 233303 156435 233309
rect 166126 233300 166132 233312
rect 166184 233300 166190 233352
rect 165942 233272 165948 233284
rect 156300 233244 165948 233272
rect 153764 233232 153770 233244
rect 165942 233232 165948 233244
rect 166000 233232 166006 233284
rect 246994 233232 247000 233284
rect 247052 233272 247058 233284
rect 249570 233272 249576 233284
rect 247052 233244 249576 233272
rect 247052 233232 247058 233244
rect 249570 233232 249576 233244
rect 249628 233232 249634 233284
rect 256378 233272 256384 233284
rect 249680 233244 256384 233272
rect 61706 233164 61712 233216
rect 61764 233204 61770 233216
rect 62074 233204 62080 233216
rect 61764 233176 62080 233204
rect 61764 233164 61770 233176
rect 62074 233164 62080 233176
rect 62132 233164 62138 233216
rect 62258 233164 62264 233216
rect 62316 233204 62322 233216
rect 75782 233204 75788 233216
rect 62316 233176 75788 233204
rect 62316 233164 62322 233176
rect 75782 233164 75788 233176
rect 75840 233164 75846 233216
rect 137790 233164 137796 233216
rect 137848 233204 137854 233216
rect 145150 233204 145156 233216
rect 137848 233176 145156 233204
rect 137848 233164 137854 233176
rect 145150 233164 145156 233176
rect 145208 233164 145214 233216
rect 151590 233164 151596 233216
rect 151648 233204 151654 233216
rect 156190 233204 156196 233216
rect 151648 233176 156196 233204
rect 151648 233164 151654 233176
rect 156190 233164 156196 233176
rect 156248 233164 156254 233216
rect 168610 233204 168616 233216
rect 156392 233176 168616 233204
rect 53242 233096 53248 233148
rect 53300 233136 53306 233148
rect 62350 233136 62356 233148
rect 53300 233108 62356 233136
rect 53300 233096 53306 233108
rect 62350 233096 62356 233108
rect 62408 233096 62414 233148
rect 62442 233096 62448 233148
rect 62500 233136 62506 233148
rect 76426 233136 76432 233148
rect 62500 233108 76432 233136
rect 62500 233096 62506 233108
rect 76426 233096 76432 233108
rect 76484 233096 76490 233148
rect 155270 233096 155276 233148
rect 155328 233136 155334 233148
rect 156392 233136 156420 233176
rect 168610 233164 168616 233176
rect 168668 233164 168674 233216
rect 231814 233164 231820 233216
rect 231872 233204 231878 233216
rect 239174 233204 239180 233216
rect 231872 233176 239180 233204
rect 231872 233164 231878 233176
rect 239174 233164 239180 233176
rect 239232 233164 239238 233216
rect 245338 233164 245344 233216
rect 245396 233204 245402 233216
rect 249386 233204 249392 233216
rect 245396 233176 249392 233204
rect 245396 233164 245402 233176
rect 249386 233164 249392 233176
rect 249444 233164 249450 233216
rect 249478 233164 249484 233216
rect 249536 233204 249542 233216
rect 249680 233204 249708 233244
rect 256378 233232 256384 233244
rect 256436 233232 256442 233284
rect 256473 233275 256531 233281
rect 256473 233241 256485 233275
rect 256519 233272 256531 233275
rect 258954 233272 258960 233284
rect 256519 233244 258960 233272
rect 256519 233241 256531 233244
rect 256473 233235 256531 233241
rect 258954 233232 258960 233244
rect 259012 233232 259018 233284
rect 249536 233176 249708 233204
rect 249536 233164 249542 233176
rect 250306 233164 250312 233216
rect 250364 233204 250370 233216
rect 263094 233204 263100 233216
rect 250364 233176 263100 233204
rect 250364 233164 250370 233176
rect 263094 233164 263100 233176
rect 263152 233164 263158 233216
rect 167322 233136 167328 233148
rect 155328 233108 156420 233136
rect 156484 233108 167328 233136
rect 155328 233096 155334 233108
rect 38154 233028 38160 233080
rect 38212 233068 38218 233080
rect 49194 233068 49200 233080
rect 38212 233040 49200 233068
rect 38212 233028 38218 233040
rect 49194 233028 49200 233040
rect 49252 233028 49258 233080
rect 62074 233028 62080 233080
rect 62132 233068 62138 233080
rect 75046 233068 75052 233080
rect 62132 233040 75052 233068
rect 62132 233028 62138 233040
rect 75046 233028 75052 233040
rect 75104 233028 75110 233080
rect 137606 233028 137612 233080
rect 137664 233068 137670 233080
rect 145702 233068 145708 233080
rect 137664 233040 145708 233068
rect 137664 233028 137670 233040
rect 145702 233028 145708 233040
rect 145760 233028 145766 233080
rect 150486 233028 150492 233080
rect 150544 233068 150550 233080
rect 154810 233068 154816 233080
rect 150544 233040 154816 233068
rect 150544 233028 150550 233040
rect 154810 233028 154816 233040
rect 154868 233028 154874 233080
rect 156484 233068 156512 233108
rect 167322 233096 167328 233108
rect 167380 233096 167386 233148
rect 248466 233096 248472 233148
rect 248524 233136 248530 233148
rect 261070 233136 261076 233148
rect 248524 233108 261076 233136
rect 248524 233096 248530 233108
rect 261070 233096 261076 233108
rect 261128 233096 261134 233148
rect 161802 233068 161808 233080
rect 154920 233040 156512 233068
rect 156576 233040 161808 233068
rect 56002 232960 56008 233012
rect 56060 233000 56066 233012
rect 66030 233000 66036 233012
rect 56060 232972 66036 233000
rect 56060 232960 56066 232972
rect 66030 232960 66036 232972
rect 66088 232960 66094 233012
rect 154718 232960 154724 233012
rect 154776 233000 154782 233012
rect 154920 233000 154948 233040
rect 156576 233000 156604 233040
rect 161802 233028 161808 233040
rect 161860 233028 161866 233080
rect 231722 233028 231728 233080
rect 231780 233068 231786 233080
rect 239634 233068 239640 233080
rect 231780 233040 239640 233068
rect 231780 233028 231786 233040
rect 239634 233028 239640 233040
rect 239692 233028 239698 233080
rect 245798 233028 245804 233080
rect 245856 233068 245862 233080
rect 249662 233068 249668 233080
rect 245856 233040 249668 233068
rect 245856 233028 245862 233040
rect 249662 233028 249668 233040
rect 249720 233028 249726 233080
rect 249846 233028 249852 233080
rect 249904 233068 249910 233080
rect 262542 233068 262548 233080
rect 249904 233040 262548 233068
rect 249904 233028 249910 233040
rect 262542 233028 262548 233040
rect 262600 233028 262606 233080
rect 154776 232972 154948 233000
rect 155288 232972 156604 233000
rect 154776 232960 154782 232972
rect 61249 232935 61307 232941
rect 61249 232901 61261 232935
rect 61295 232932 61307 232935
rect 63638 232932 63644 232944
rect 61295 232904 63644 232932
rect 61295 232901 61307 232904
rect 61249 232895 61307 232901
rect 63638 232892 63644 232904
rect 63696 232892 63702 232944
rect 152786 232892 152792 232944
rect 152844 232932 152850 232944
rect 155178 232932 155184 232944
rect 152844 232904 155184 232932
rect 152844 232892 152850 232904
rect 155178 232892 155184 232904
rect 155236 232892 155242 232944
rect 56646 232824 56652 232876
rect 56704 232864 56710 232876
rect 66398 232864 66404 232876
rect 56704 232836 66404 232864
rect 56704 232824 56710 232836
rect 66398 232824 66404 232836
rect 66456 232824 66462 232876
rect 150578 232824 150584 232876
rect 150636 232864 150642 232876
rect 155288 232864 155316 232972
rect 242486 232960 242492 233012
rect 242544 233000 242550 233012
rect 247638 233000 247644 233012
rect 242544 232972 247644 233000
rect 242544 232960 242550 232972
rect 247638 232960 247644 232972
rect 247696 232960 247702 233012
rect 247733 233003 247791 233009
rect 247733 232969 247745 233003
rect 247779 233000 247791 233003
rect 258310 233000 258316 233012
rect 247779 232972 258316 233000
rect 247779 232969 247791 232972
rect 247733 232963 247791 232969
rect 258310 232960 258316 232972
rect 258368 232960 258374 233012
rect 158030 232892 158036 232944
rect 158088 232932 158094 232944
rect 161158 232932 161164 232944
rect 158088 232904 161164 232932
rect 158088 232892 158094 232904
rect 161158 232892 161164 232904
rect 161216 232892 161222 232944
rect 243590 232892 243596 232944
rect 243648 232932 243654 232944
rect 248282 232932 248288 232944
rect 243648 232904 248288 232932
rect 243648 232892 243654 232904
rect 248282 232892 248288 232904
rect 248340 232892 248346 232944
rect 248469 232935 248527 232941
rect 248469 232901 248481 232935
rect 248515 232932 248527 232935
rect 256930 232932 256936 232944
rect 248515 232904 256936 232932
rect 248515 232901 248527 232904
rect 248469 232895 248527 232901
rect 256930 232892 256936 232904
rect 256988 232892 256994 232944
rect 150636 232836 155316 232864
rect 150636 232824 150642 232836
rect 159778 232824 159784 232876
rect 159836 232864 159842 232876
rect 162630 232864 162636 232876
rect 159836 232836 162636 232864
rect 159836 232824 159842 232836
rect 162630 232824 162636 232836
rect 162688 232824 162694 232876
rect 244142 232824 244148 232876
rect 244200 232864 244206 232876
rect 247546 232864 247552 232876
rect 244200 232836 247552 232864
rect 244200 232824 244206 232836
rect 247546 232824 247552 232836
rect 247604 232824 247610 232876
rect 254170 232864 254176 232876
rect 248484 232836 254176 232864
rect 59314 232756 59320 232808
rect 59372 232796 59378 232808
rect 59372 232768 68376 232796
rect 59372 232756 59378 232768
rect 58026 232688 58032 232740
rect 58084 232728 58090 232740
rect 61338 232728 61344 232740
rect 58084 232700 61344 232728
rect 58084 232688 58090 232700
rect 61338 232688 61344 232700
rect 61396 232688 61402 232740
rect 61522 232688 61528 232740
rect 61580 232728 61586 232740
rect 68238 232728 68244 232740
rect 61580 232700 68244 232728
rect 61580 232688 61586 232700
rect 68238 232688 68244 232700
rect 68296 232688 68302 232740
rect 60786 232620 60792 232672
rect 60844 232660 60850 232672
rect 61249 232663 61307 232669
rect 61249 232660 61261 232663
rect 60844 232632 61261 232660
rect 60844 232620 60850 232632
rect 61249 232629 61261 232632
rect 61295 232629 61307 232663
rect 61249 232623 61307 232629
rect 61614 232620 61620 232672
rect 61672 232660 61678 232672
rect 67594 232660 67600 232672
rect 61672 232632 67600 232660
rect 61672 232620 61678 232632
rect 67594 232620 67600 232632
rect 67652 232620 67658 232672
rect 68348 232660 68376 232768
rect 149842 232756 149848 232808
rect 149900 232796 149906 232808
rect 151866 232796 151872 232808
rect 149900 232768 151872 232796
rect 149900 232756 149906 232768
rect 151866 232756 151872 232768
rect 151924 232756 151930 232808
rect 151958 232756 151964 232808
rect 152016 232796 152022 232808
rect 156282 232796 156288 232808
rect 152016 232768 156288 232796
rect 152016 232756 152022 232768
rect 156282 232756 156288 232768
rect 156340 232756 156346 232808
rect 156834 232756 156840 232808
rect 156892 232796 156898 232808
rect 160054 232796 160060 232808
rect 156892 232768 160060 232796
rect 156892 232756 156898 232768
rect 160054 232756 160060 232768
rect 160112 232756 160118 232808
rect 246718 232756 246724 232808
rect 246776 232796 246782 232808
rect 247733 232799 247791 232805
rect 247733 232796 247745 232799
rect 246776 232768 247745 232796
rect 246776 232756 246782 232768
rect 247733 232765 247745 232768
rect 247779 232765 247791 232799
rect 247733 232759 247791 232765
rect 248006 232756 248012 232808
rect 248064 232796 248070 232808
rect 248484 232796 248512 232836
rect 254170 232824 254176 232836
rect 254228 232824 254234 232876
rect 248064 232768 248512 232796
rect 248064 232756 248070 232768
rect 248558 232756 248564 232808
rect 248616 232796 248622 232808
rect 254722 232796 254728 232808
rect 248616 232768 254728 232796
rect 248616 232756 248622 232768
rect 254722 232756 254728 232768
rect 254780 232756 254786 232808
rect 153338 232688 153344 232740
rect 153396 232728 153402 232740
rect 158214 232728 158220 232740
rect 153396 232700 158220 232728
rect 153396 232688 153402 232700
rect 158214 232688 158220 232700
rect 158272 232688 158278 232740
rect 158582 232688 158588 232740
rect 158640 232728 158646 232740
rect 160974 232728 160980 232740
rect 158640 232700 160980 232728
rect 158640 232688 158646 232700
rect 160974 232688 160980 232700
rect 161032 232688 161038 232740
rect 161161 232731 161219 232737
rect 161161 232697 161173 232731
rect 161207 232728 161219 232731
rect 169070 232728 169076 232740
rect 161207 232700 169076 232728
rect 161207 232697 161219 232700
rect 161161 232691 161219 232697
rect 169070 232688 169076 232700
rect 169128 232688 169134 232740
rect 247178 232688 247184 232740
rect 247236 232728 247242 232740
rect 258678 232728 258684 232740
rect 247236 232700 258684 232728
rect 247236 232688 247242 232700
rect 258678 232688 258684 232700
rect 258736 232688 258742 232740
rect 70998 232660 71004 232672
rect 68348 232632 71004 232660
rect 70998 232620 71004 232632
rect 71056 232620 71062 232672
rect 153982 232620 153988 232672
rect 154040 232660 154046 232672
rect 154994 232660 155000 232672
rect 154040 232632 155000 232660
rect 154040 232620 154046 232632
rect 154994 232620 155000 232632
rect 155052 232620 155058 232672
rect 155086 232620 155092 232672
rect 155144 232660 155150 232672
rect 158306 232660 158312 232672
rect 155144 232632 158312 232660
rect 155144 232620 155150 232632
rect 158306 232620 158312 232632
rect 158364 232620 158370 232672
rect 159042 232620 159048 232672
rect 159100 232660 159106 232672
rect 161066 232660 161072 232672
rect 159100 232632 161072 232660
rect 159100 232620 159106 232632
rect 161066 232620 161072 232632
rect 161124 232620 161130 232672
rect 231630 232620 231636 232672
rect 231688 232660 231694 232672
rect 238530 232660 238536 232672
rect 231688 232632 238536 232660
rect 231688 232620 231694 232632
rect 238530 232620 238536 232632
rect 238588 232620 238594 232672
rect 244418 232620 244424 232672
rect 244476 232660 244482 232672
rect 247362 232660 247368 232672
rect 244476 232632 247368 232660
rect 244476 232620 244482 232632
rect 247362 232620 247368 232632
rect 247420 232620 247426 232672
rect 248098 232620 248104 232672
rect 248156 232660 248162 232672
rect 249938 232660 249944 232672
rect 248156 232632 249944 232660
rect 248156 232620 248162 232632
rect 249938 232620 249944 232632
rect 249996 232620 250002 232672
rect 252054 232620 252060 232672
rect 252112 232660 252118 232672
rect 257022 232660 257028 232672
rect 252112 232632 257028 232660
rect 252112 232620 252118 232632
rect 257022 232620 257028 232632
rect 257080 232620 257086 232672
rect 57290 232552 57296 232604
rect 57348 232592 57354 232604
rect 61430 232592 61436 232604
rect 57348 232564 61436 232592
rect 57348 232552 57354 232564
rect 61430 232552 61436 232564
rect 61488 232552 61494 232604
rect 61798 232552 61804 232604
rect 61856 232592 61862 232604
rect 63454 232592 63460 232604
rect 61856 232564 63460 232592
rect 61856 232552 61862 232564
rect 63454 232552 63460 232564
rect 63512 232552 63518 232604
rect 67962 232552 67968 232604
rect 68020 232592 68026 232604
rect 70262 232592 70268 232604
rect 68020 232564 70268 232592
rect 68020 232552 68026 232564
rect 70262 232552 70268 232564
rect 70320 232552 70326 232604
rect 157478 232552 157484 232604
rect 157536 232592 157542 232604
rect 159870 232592 159876 232604
rect 157536 232564 159876 232592
rect 157536 232552 157542 232564
rect 159870 232552 159876 232564
rect 159928 232552 159934 232604
rect 231538 232552 231544 232604
rect 231596 232592 231602 232604
rect 237978 232592 237984 232604
rect 231596 232564 237984 232592
rect 231596 232552 231602 232564
rect 237978 232552 237984 232564
rect 238036 232552 238042 232604
rect 245798 232552 245804 232604
rect 245856 232592 245862 232604
rect 248469 232595 248527 232601
rect 248469 232592 248481 232595
rect 245856 232564 248481 232592
rect 245856 232552 245862 232564
rect 248469 232561 248481 232564
rect 248515 232561 248527 232595
rect 248469 232555 248527 232561
rect 253066 232552 253072 232604
rect 253124 232592 253130 232604
rect 256473 232595 256531 232601
rect 256473 232592 256485 232595
rect 253124 232564 256485 232592
rect 253124 232552 253130 232564
rect 256473 232561 256485 232564
rect 256519 232561 256531 232595
rect 256473 232555 256531 232561
rect 62166 232484 62172 232536
rect 62224 232524 62230 232536
rect 66858 232524 66864 232536
rect 62224 232496 66864 232524
rect 62224 232484 62230 232496
rect 66858 232484 66864 232496
rect 66916 232484 66922 232536
rect 67870 232484 67876 232536
rect 67928 232524 67934 232536
rect 69618 232524 69624 232536
rect 67928 232496 69624 232524
rect 67928 232484 67934 232496
rect 69618 232484 69624 232496
rect 69676 232484 69682 232536
rect 151038 232484 151044 232536
rect 151096 232524 151102 232536
rect 153430 232524 153436 232536
rect 151096 232496 153436 232524
rect 151096 232484 151102 232496
rect 153430 232484 153436 232496
rect 153488 232484 153494 232536
rect 156374 232484 156380 232536
rect 156432 232524 156438 232536
rect 159134 232524 159140 232536
rect 156432 232496 159140 232524
rect 156432 232484 156438 232496
rect 159134 232484 159140 232496
rect 159192 232484 159198 232536
rect 231446 232484 231452 232536
rect 231504 232524 231510 232536
rect 237610 232524 237616 232536
rect 231504 232496 237616 232524
rect 231504 232484 231510 232496
rect 237610 232484 237616 232496
rect 237668 232484 237674 232536
rect 243038 232484 243044 232536
rect 243096 232524 243102 232536
rect 246994 232524 247000 232536
rect 243096 232496 247000 232524
rect 243096 232484 243102 232496
rect 246994 232484 247000 232496
rect 247052 232484 247058 232536
rect 248190 232484 248196 232536
rect 248248 232524 248254 232536
rect 260334 232524 260340 232536
rect 248248 232496 260340 232524
rect 248248 232484 248254 232496
rect 260334 232484 260340 232496
rect 260392 232484 260398 232536
rect 60050 232416 60056 232468
rect 60108 232456 60114 232468
rect 61154 232456 61160 232468
rect 60108 232428 61160 232456
rect 60108 232416 60114 232428
rect 61154 232416 61160 232428
rect 61212 232416 61218 232468
rect 61982 232416 61988 232468
rect 62040 232456 62046 232468
rect 68974 232456 68980 232468
rect 62040 232428 68980 232456
rect 62040 232416 62046 232428
rect 68974 232416 68980 232428
rect 69032 232416 69038 232468
rect 158398 232416 158404 232468
rect 158456 232456 158462 232468
rect 159686 232456 159692 232468
rect 158456 232428 159692 232456
rect 158456 232416 158462 232428
rect 159686 232416 159692 232428
rect 159744 232416 159750 232468
rect 162354 232416 162360 232468
rect 162412 232456 162418 232468
rect 163826 232456 163832 232468
rect 162412 232428 163832 232456
rect 162412 232416 162418 232428
rect 163826 232416 163832 232428
rect 163884 232416 163890 232468
rect 231354 232416 231360 232468
rect 231412 232456 231418 232468
rect 236874 232456 236880 232468
rect 231412 232428 236880 232456
rect 231412 232416 231418 232428
rect 236874 232416 236880 232428
rect 236932 232416 236938 232468
rect 241566 232416 241572 232468
rect 241624 232456 241630 232468
rect 245430 232456 245436 232468
rect 241624 232428 245436 232456
rect 241624 232416 241630 232428
rect 245430 232416 245436 232428
rect 245488 232416 245494 232468
rect 246442 232416 246448 232468
rect 246500 232456 246506 232468
rect 251410 232456 251416 232468
rect 246500 232428 251416 232456
rect 246500 232416 246506 232428
rect 251410 232416 251416 232428
rect 251468 232416 251474 232468
rect 256194 232416 256200 232468
rect 256252 232456 256258 232468
rect 257482 232456 257488 232468
rect 256252 232428 257488 232456
rect 256252 232416 256258 232428
rect 257482 232416 257488 232428
rect 257540 232416 257546 232468
rect 155730 231464 155736 231516
rect 155788 231504 155794 231516
rect 161161 231507 161219 231513
rect 161161 231504 161173 231507
rect 155788 231476 161173 231504
rect 155788 231464 155794 231476
rect 161161 231473 161173 231476
rect 161207 231473 161219 231507
rect 161161 231467 161219 231473
rect 126474 229628 126480 229680
rect 126532 229668 126538 229680
rect 159594 229668 159600 229680
rect 126532 229640 159600 229668
rect 126532 229628 126538 229640
rect 159594 229628 159600 229640
rect 159652 229628 159658 229680
rect 220498 229628 220504 229680
rect 220556 229668 220562 229680
rect 254722 229668 254728 229680
rect 220556 229640 254728 229668
rect 220556 229628 220562 229640
rect 254722 229628 254728 229640
rect 254780 229628 254786 229680
rect 137698 228200 137704 228252
rect 137756 228240 137762 228252
rect 146806 228240 146812 228252
rect 137756 228212 146812 228240
rect 137756 228200 137762 228212
rect 146806 228200 146812 228212
rect 146864 228200 146870 228252
rect 231998 228200 232004 228252
rect 232056 228240 232062 228252
rect 240738 228240 240744 228252
rect 232056 228212 240744 228240
rect 232056 228200 232062 228212
rect 240738 228200 240744 228212
rect 240796 228200 240802 228252
rect 156098 226840 156104 226892
rect 156156 226880 156162 226892
rect 157757 226883 157815 226889
rect 157757 226880 157769 226883
rect 156156 226852 157769 226880
rect 156156 226840 156162 226852
rect 157757 226849 157769 226852
rect 157803 226849 157815 226883
rect 157757 226843 157815 226849
rect 60804 225560 61108 225588
rect 56186 225412 56192 225464
rect 56244 225452 56250 225464
rect 57658 225452 57664 225464
rect 56244 225424 57664 225452
rect 56244 225412 56250 225424
rect 57658 225412 57664 225424
rect 57716 225412 57722 225464
rect 58670 225412 58676 225464
rect 58728 225452 58734 225464
rect 59498 225452 59504 225464
rect 58728 225424 59504 225452
rect 58728 225412 58734 225424
rect 59498 225412 59504 225424
rect 59556 225412 59562 225464
rect 59593 225455 59651 225461
rect 59593 225421 59605 225455
rect 59639 225452 59651 225455
rect 60804 225452 60832 225560
rect 60881 225523 60939 225529
rect 60881 225489 60893 225523
rect 60927 225520 60939 225523
rect 60973 225523 61031 225529
rect 60973 225520 60985 225523
rect 60927 225492 60985 225520
rect 60927 225489 60939 225492
rect 60881 225483 60939 225489
rect 60973 225489 60985 225492
rect 61019 225489 61031 225523
rect 60973 225483 61031 225489
rect 61080 225452 61108 225560
rect 231906 225480 231912 225532
rect 231964 225520 231970 225532
rect 234114 225520 234120 225532
rect 231964 225492 234120 225520
rect 231964 225480 231970 225492
rect 234114 225480 234120 225492
rect 234172 225480 234178 225532
rect 64282 225452 64288 225464
rect 59639 225424 60832 225452
rect 60896 225424 61016 225452
rect 61080 225424 64288 225452
rect 59639 225421 59651 225424
rect 59593 225415 59651 225421
rect 55266 225344 55272 225396
rect 55324 225384 55330 225396
rect 60896 225384 60924 225424
rect 55324 225356 60924 225384
rect 55324 225344 55330 225356
rect 51862 225276 51868 225328
rect 51920 225316 51926 225328
rect 60881 225319 60939 225325
rect 60881 225316 60893 225319
rect 51920 225288 60893 225316
rect 51920 225276 51926 225288
rect 60881 225285 60893 225288
rect 60927 225285 60939 225319
rect 60988 225316 61016 225424
rect 64282 225412 64288 225424
rect 64340 225412 64346 225464
rect 151406 225412 151412 225464
rect 151464 225452 151470 225464
rect 159686 225452 159692 225464
rect 151464 225424 159692 225452
rect 151464 225412 151470 225424
rect 159686 225412 159692 225424
rect 159744 225412 159750 225464
rect 161158 225412 161164 225464
rect 161216 225452 161222 225464
rect 163550 225452 163556 225464
rect 161216 225424 163556 225452
rect 161216 225412 161222 225424
rect 163550 225412 163556 225424
rect 163608 225412 163614 225464
rect 244418 225412 244424 225464
rect 244476 225452 244482 225464
rect 248558 225452 248564 225464
rect 244476 225424 248564 225452
rect 244476 225412 244482 225424
rect 248558 225412 248564 225424
rect 248616 225412 248622 225464
rect 250030 225412 250036 225464
rect 250088 225452 250094 225464
rect 253713 225455 253771 225461
rect 253713 225452 253725 225455
rect 250088 225424 253725 225452
rect 250088 225412 250094 225424
rect 253713 225421 253725 225424
rect 253759 225421 253771 225455
rect 253713 225415 253771 225421
rect 254722 225412 254728 225464
rect 254780 225452 254786 225464
rect 258678 225452 258684 225464
rect 254780 225424 258684 225452
rect 254780 225412 254786 225424
rect 258678 225412 258684 225424
rect 258736 225412 258742 225464
rect 61065 225387 61123 225393
rect 61065 225353 61077 225387
rect 61111 225384 61123 225387
rect 64006 225384 64012 225396
rect 61111 225356 64012 225384
rect 61111 225353 61123 225356
rect 61065 225347 61123 225353
rect 64006 225344 64012 225356
rect 64064 225344 64070 225396
rect 149842 225344 149848 225396
rect 149900 225384 149906 225396
rect 160330 225384 160336 225396
rect 149900 225356 160336 225384
rect 149900 225344 149906 225356
rect 160330 225344 160336 225356
rect 160388 225344 160394 225396
rect 160974 225344 160980 225396
rect 161032 225384 161038 225396
rect 163918 225384 163924 225396
rect 161032 225356 163924 225384
rect 161032 225344 161038 225356
rect 163918 225344 163924 225356
rect 163976 225344 163982 225396
rect 244050 225344 244056 225396
rect 244108 225384 244114 225396
rect 248006 225384 248012 225396
rect 244108 225356 248012 225384
rect 244108 225344 244114 225356
rect 248006 225344 248012 225356
rect 248064 225344 248070 225396
rect 248282 225344 248288 225396
rect 248340 225384 248346 225396
rect 252054 225384 252060 225396
rect 248340 225356 252060 225384
rect 248340 225344 248346 225356
rect 252054 225344 252060 225356
rect 252112 225344 252118 225396
rect 252698 225344 252704 225396
rect 252756 225384 252762 225396
rect 258310 225384 258316 225396
rect 252756 225356 258316 225384
rect 252756 225344 252762 225356
rect 258310 225344 258316 225356
rect 258368 225344 258374 225396
rect 65938 225316 65944 225328
rect 60988 225288 65944 225316
rect 60881 225279 60939 225285
rect 65938 225276 65944 225288
rect 65996 225276 66002 225328
rect 156190 225276 156196 225328
rect 156248 225316 156254 225328
rect 159226 225316 159232 225328
rect 156248 225288 159232 225316
rect 156248 225276 156254 225288
rect 159226 225276 159232 225288
rect 159284 225276 159290 225328
rect 159778 225276 159784 225328
rect 159836 225316 159842 225328
rect 163090 225316 163096 225328
rect 159836 225288 163096 225316
rect 159836 225276 159842 225288
rect 163090 225276 163096 225288
rect 163148 225276 163154 225328
rect 175326 225276 175332 225328
rect 175384 225316 175390 225328
rect 281862 225316 281868 225328
rect 175384 225288 281868 225316
rect 175384 225276 175390 225288
rect 281862 225276 281868 225288
rect 281920 225276 281926 225328
rect 55818 225208 55824 225260
rect 55876 225248 55882 225260
rect 59593 225251 59651 225257
rect 59593 225248 59605 225251
rect 55876 225220 59605 225248
rect 55876 225208 55882 225220
rect 59593 225217 59605 225220
rect 59639 225217 59651 225251
rect 59593 225211 59651 225217
rect 59682 225208 59688 225260
rect 59740 225248 59746 225260
rect 60970 225248 60976 225260
rect 59740 225220 60976 225248
rect 59740 225208 59746 225220
rect 60970 225208 60976 225220
rect 61028 225208 61034 225260
rect 61433 225251 61491 225257
rect 61433 225217 61445 225251
rect 61479 225248 61491 225251
rect 61479 225220 62120 225248
rect 61479 225217 61491 225220
rect 61433 225211 61491 225217
rect 54622 225140 54628 225192
rect 54680 225180 54686 225192
rect 54680 225152 56324 225180
rect 54680 225140 54686 225152
rect 52506 225072 52512 225124
rect 52564 225112 52570 225124
rect 56296 225112 56324 225152
rect 56554 225140 56560 225192
rect 56612 225180 56618 225192
rect 57934 225180 57940 225192
rect 56612 225152 57940 225180
rect 56612 225140 56618 225152
rect 57934 225140 57940 225152
rect 57992 225140 57998 225192
rect 58118 225140 58124 225192
rect 58176 225180 58182 225192
rect 61982 225180 61988 225192
rect 58176 225152 61988 225180
rect 58176 225140 58182 225152
rect 61982 225140 61988 225152
rect 62040 225140 62046 225192
rect 62092 225180 62120 225220
rect 62810 225208 62816 225260
rect 62868 225248 62874 225260
rect 70262 225248 70268 225260
rect 62868 225220 70268 225248
rect 62868 225208 62874 225220
rect 70262 225208 70268 225220
rect 70320 225208 70326 225260
rect 154810 225208 154816 225260
rect 154868 225248 154874 225260
rect 158398 225248 158404 225260
rect 154868 225220 158404 225248
rect 154868 225208 154874 225220
rect 158398 225208 158404 225220
rect 158456 225208 158462 225260
rect 245430 225208 245436 225260
rect 245488 225248 245494 225260
rect 250858 225248 250864 225260
rect 245488 225220 250864 225248
rect 245488 225208 245494 225220
rect 250858 225208 250864 225220
rect 250916 225208 250922 225260
rect 251318 225208 251324 225260
rect 251376 225248 251382 225260
rect 251376 225220 252560 225248
rect 251376 225208 251382 225220
rect 67870 225180 67876 225192
rect 62092 225152 67876 225180
rect 67870 225140 67876 225152
rect 67928 225140 67934 225192
rect 150210 225140 150216 225192
rect 150268 225180 150274 225192
rect 160422 225180 160428 225192
rect 150268 225152 160428 225180
rect 150268 225140 150274 225152
rect 160422 225140 160428 225152
rect 160480 225140 160486 225192
rect 246994 225140 247000 225192
rect 247052 225180 247058 225192
rect 251686 225180 251692 225192
rect 247052 225152 251692 225180
rect 247052 225140 247058 225152
rect 251686 225140 251692 225152
rect 251744 225140 251750 225192
rect 252532 225180 252560 225220
rect 257574 225180 257580 225192
rect 252532 225152 257580 225180
rect 257574 225140 257580 225152
rect 257632 225140 257638 225192
rect 59317 225115 59375 225121
rect 59317 225112 59329 225115
rect 52564 225084 56232 225112
rect 56296 225084 59329 225112
rect 52564 225072 52570 225084
rect 51218 225004 51224 225056
rect 51276 225044 51282 225056
rect 51276 225016 56048 225044
rect 51276 225004 51282 225016
rect 51126 224868 51132 224920
rect 51184 224908 51190 224920
rect 51184 224880 55956 224908
rect 51184 224868 51190 224880
rect 29138 224800 29144 224852
rect 29196 224840 29202 224852
rect 31622 224840 31628 224852
rect 29196 224812 31628 224840
rect 29196 224800 29202 224812
rect 31622 224800 31628 224812
rect 31680 224800 31686 224852
rect 49838 224732 49844 224784
rect 49896 224772 49902 224784
rect 49896 224744 53932 224772
rect 49896 224732 49902 224744
rect 53904 224568 53932 224744
rect 55928 224704 55956 224880
rect 56020 224772 56048 225016
rect 56204 224840 56232 225084
rect 59317 225081 59329 225084
rect 59363 225081 59375 225115
rect 59317 225075 59375 225081
rect 59406 225072 59412 225124
rect 59464 225112 59470 225124
rect 59464 225084 61660 225112
rect 59464 225072 59470 225084
rect 56281 225047 56339 225053
rect 56281 225013 56293 225047
rect 56327 225044 56339 225047
rect 58857 225047 58915 225053
rect 58857 225044 58869 225047
rect 56327 225016 58869 225044
rect 56327 225013 56339 225016
rect 56281 225007 56339 225013
rect 58857 225013 58869 225016
rect 58903 225013 58915 225047
rect 58857 225007 58915 225013
rect 58578 224936 58584 224988
rect 58636 224976 58642 224988
rect 61433 224979 61491 224985
rect 61433 224976 61445 224979
rect 58636 224948 61445 224976
rect 58636 224936 58642 224948
rect 61433 224945 61445 224948
rect 61479 224945 61491 224979
rect 61632 224976 61660 225084
rect 61890 225072 61896 225124
rect 61948 225112 61954 225124
rect 69526 225112 69532 225124
rect 61948 225084 69532 225112
rect 61948 225072 61954 225084
rect 69526 225072 69532 225084
rect 69584 225072 69590 225124
rect 148646 225072 148652 225124
rect 148704 225112 148710 225124
rect 157294 225112 157300 225124
rect 148704 225084 157300 225112
rect 148704 225072 148710 225084
rect 157294 225072 157300 225084
rect 157352 225072 157358 225124
rect 157389 225115 157447 225121
rect 157389 225081 157401 225115
rect 157435 225112 157447 225115
rect 157662 225112 157668 225124
rect 157435 225084 157668 225112
rect 157435 225081 157447 225084
rect 157389 225075 157447 225081
rect 157662 225072 157668 225084
rect 157720 225072 157726 225124
rect 157757 225115 157815 225121
rect 157757 225081 157769 225115
rect 157803 225112 157815 225115
rect 157803 225084 159548 225112
rect 157803 225081 157815 225084
rect 157757 225075 157815 225081
rect 63638 225004 63644 225056
rect 63696 225044 63702 225056
rect 69066 225044 69072 225056
rect 63696 225016 69072 225044
rect 63696 225004 63702 225016
rect 69066 225004 69072 225016
rect 69124 225004 69130 225056
rect 149474 225004 149480 225056
rect 149532 225044 149538 225056
rect 158582 225044 158588 225056
rect 149532 225016 158588 225044
rect 149532 225004 149538 225016
rect 158582 225004 158588 225016
rect 158640 225004 158646 225056
rect 159520 225044 159548 225084
rect 159594 225072 159600 225124
rect 159652 225112 159658 225124
rect 164654 225112 164660 225124
rect 159652 225084 164660 225112
rect 159652 225072 159658 225084
rect 164654 225072 164660 225084
rect 164712 225072 164718 225124
rect 247638 225072 247644 225124
rect 247696 225112 247702 225124
rect 251318 225112 251324 225124
rect 247696 225084 251324 225112
rect 247696 225072 247702 225084
rect 251318 225072 251324 225084
rect 251376 225072 251382 225124
rect 251410 225072 251416 225124
rect 251468 225112 251474 225124
rect 253986 225112 253992 225124
rect 251468 225084 253992 225112
rect 251468 225072 251474 225084
rect 253986 225072 253992 225084
rect 254044 225072 254050 225124
rect 160882 225044 160888 225056
rect 159520 225016 160888 225044
rect 160882 225004 160888 225016
rect 160940 225004 160946 225056
rect 161066 225004 161072 225056
rect 161124 225044 161130 225056
rect 164286 225044 164292 225056
rect 161124 225016 164292 225044
rect 161124 225004 161130 225016
rect 164286 225004 164292 225016
rect 164344 225004 164350 225056
rect 245614 225004 245620 225056
rect 245672 225044 245678 225056
rect 249478 225044 249484 225056
rect 245672 225016 249484 225044
rect 245672 225004 245678 225016
rect 249478 225004 249484 225016
rect 249536 225004 249542 225056
rect 251042 225004 251048 225056
rect 251100 225044 251106 225056
rect 251100 225016 253296 225044
rect 251100 225004 251106 225016
rect 68330 224976 68336 224988
rect 61632 224948 68336 224976
rect 61433 224939 61491 224945
rect 68330 224936 68336 224948
rect 68388 224936 68394 224988
rect 156282 224936 156288 224988
rect 156340 224976 156346 224988
rect 159594 224976 159600 224988
rect 156340 224948 159600 224976
rect 156340 224936 156346 224948
rect 159594 224936 159600 224948
rect 159652 224936 159658 224988
rect 159870 224936 159876 224988
rect 159928 224976 159934 224988
rect 162722 224976 162728 224988
rect 159928 224948 162728 224976
rect 159928 224936 159934 224948
rect 162722 224936 162728 224948
rect 162780 224936 162786 224988
rect 243314 224936 243320 224988
rect 243372 224976 243378 224988
rect 253158 224976 253164 224988
rect 243372 224948 253164 224976
rect 243372 224936 243378 224948
rect 253158 224936 253164 224948
rect 253216 224936 253222 224988
rect 253268 224976 253296 225016
rect 257114 224976 257120 224988
rect 253268 224948 257120 224976
rect 257114 224936 257120 224948
rect 257172 224936 257178 224988
rect 56373 224911 56431 224917
rect 56373 224877 56385 224911
rect 56419 224908 56431 224911
rect 60881 224911 60939 224917
rect 60881 224908 60893 224911
rect 56419 224880 60893 224908
rect 56419 224877 56431 224880
rect 56373 224871 56431 224877
rect 60881 224877 60893 224880
rect 60927 224877 60939 224911
rect 60881 224871 60939 224877
rect 61154 224868 61160 224920
rect 61212 224908 61218 224920
rect 61525 224911 61583 224917
rect 61525 224908 61537 224911
rect 61212 224880 61537 224908
rect 61212 224868 61218 224880
rect 61525 224877 61537 224880
rect 61571 224877 61583 224911
rect 61525 224871 61583 224877
rect 61706 224868 61712 224920
rect 61764 224908 61770 224920
rect 69894 224908 69900 224920
rect 61764 224880 69900 224908
rect 61764 224868 61770 224880
rect 69894 224868 69900 224880
rect 69952 224868 69958 224920
rect 151038 224868 151044 224920
rect 151096 224908 151102 224920
rect 159502 224908 159508 224920
rect 151096 224880 159508 224908
rect 151096 224868 151102 224880
rect 159502 224868 159508 224880
rect 159560 224868 159566 224920
rect 243682 224868 243688 224920
rect 243740 224908 243746 224920
rect 253618 224908 253624 224920
rect 243740 224880 253624 224908
rect 243740 224868 243746 224880
rect 253618 224868 253624 224880
rect 253676 224868 253682 224920
rect 253713 224911 253771 224917
rect 253713 224877 253725 224911
rect 253759 224908 253771 224911
rect 256746 224908 256752 224920
rect 253759 224880 256752 224908
rect 253759 224877 253771 224880
rect 253713 224871 253771 224877
rect 256746 224868 256752 224880
rect 256804 224868 256810 224920
rect 64374 224840 64380 224852
rect 56204 224812 64380 224840
rect 64374 224800 64380 224812
rect 64432 224800 64438 224852
rect 152602 224800 152608 224852
rect 152660 224840 152666 224852
rect 164562 224840 164568 224852
rect 152660 224812 164568 224840
rect 152660 224800 152666 224812
rect 164562 224800 164568 224812
rect 164620 224800 164626 224852
rect 247546 224800 247552 224852
rect 247604 224840 247610 224852
rect 252422 224840 252428 224852
rect 247604 224812 252428 224840
rect 247604 224800 247610 224812
rect 252422 224800 252428 224812
rect 252480 224800 252486 224852
rect 252517 224843 252575 224849
rect 252517 224809 252529 224843
rect 252563 224840 252575 224843
rect 256010 224840 256016 224852
rect 252563 224812 256016 224840
rect 252563 224809 252575 224812
rect 252517 224803 252575 224809
rect 256010 224800 256016 224812
rect 256068 224800 256074 224852
rect 63362 224772 63368 224784
rect 56020 224744 63368 224772
rect 63362 224732 63368 224744
rect 63420 224732 63426 224784
rect 149106 224732 149112 224784
rect 149164 224772 149170 224784
rect 156374 224772 156380 224784
rect 149164 224744 156380 224772
rect 149164 224732 149170 224744
rect 156374 224732 156380 224744
rect 156432 224732 156438 224784
rect 156466 224732 156472 224784
rect 156524 224772 156530 224784
rect 170174 224772 170180 224784
rect 156524 224744 170180 224772
rect 156524 224732 156530 224744
rect 170174 224732 170180 224744
rect 170232 224732 170238 224784
rect 247270 224732 247276 224784
rect 247328 224772 247334 224784
rect 250309 224775 250367 224781
rect 250309 224772 250321 224775
rect 247328 224744 250321 224772
rect 247328 224732 247334 224744
rect 250309 224741 250321 224744
rect 250355 224741 250367 224775
rect 250309 224735 250367 224741
rect 250674 224732 250680 224784
rect 250732 224772 250738 224784
rect 263830 224772 263836 224784
rect 250732 224744 263836 224772
rect 250732 224732 250738 224744
rect 263830 224732 263836 224744
rect 263888 224732 263894 224784
rect 267234 224732 267240 224784
rect 267292 224772 267298 224784
rect 289866 224772 289872 224784
rect 267292 224744 289872 224772
rect 267292 224732 267298 224744
rect 289866 224732 289872 224744
rect 289924 224732 289930 224784
rect 56281 224707 56339 224713
rect 56281 224704 56293 224707
rect 55928 224676 56293 224704
rect 56281 224673 56293 224676
rect 56327 224673 56339 224707
rect 56281 224667 56339 224673
rect 57290 224664 57296 224716
rect 57348 224704 57354 224716
rect 62166 224704 62172 224716
rect 57348 224676 62172 224704
rect 57348 224664 57354 224676
rect 62166 224664 62172 224676
rect 62224 224664 62230 224716
rect 62350 224664 62356 224716
rect 62408 224704 62414 224716
rect 64834 224704 64840 224716
rect 62408 224676 64840 224704
rect 62408 224664 62414 224676
rect 64834 224664 64840 224676
rect 64892 224664 64898 224716
rect 149198 224664 149204 224716
rect 149256 224704 149262 224716
rect 157389 224707 157447 224713
rect 157389 224704 157401 224707
rect 149256 224676 157401 224704
rect 149256 224664 149262 224676
rect 157389 224673 157401 224676
rect 157435 224673 157447 224707
rect 157389 224667 157447 224673
rect 247546 224664 247552 224716
rect 247604 224704 247610 224716
rect 249110 224704 249116 224716
rect 247604 224676 249116 224704
rect 247604 224664 247610 224676
rect 249110 224664 249116 224676
rect 249168 224664 249174 224716
rect 249202 224664 249208 224716
rect 249260 224704 249266 224716
rect 252517 224707 252575 224713
rect 252517 224704 252529 224707
rect 249260 224676 252529 224704
rect 249260 224664 249266 224676
rect 252517 224673 252529 224676
rect 252563 224673 252575 224707
rect 256378 224704 256384 224716
rect 252517 224667 252575 224673
rect 252624 224676 256384 224704
rect 53978 224596 53984 224648
rect 54036 224636 54042 224648
rect 65202 224636 65208 224648
rect 54036 224608 65208 224636
rect 54036 224596 54042 224608
rect 65202 224596 65208 224608
rect 65260 224596 65266 224648
rect 147818 224596 147824 224648
rect 147876 224636 147882 224648
rect 156834 224636 156840 224648
rect 147876 224608 156840 224636
rect 147876 224596 147882 224608
rect 156834 224596 156840 224608
rect 156892 224596 156898 224648
rect 158214 224596 158220 224648
rect 158272 224636 158278 224648
rect 160422 224636 160428 224648
rect 158272 224608 160428 224636
rect 158272 224596 158278 224608
rect 160422 224596 160428 224608
rect 160480 224596 160486 224648
rect 244878 224596 244884 224648
rect 244936 224636 244942 224648
rect 249018 224636 249024 224648
rect 244936 224608 249024 224636
rect 244936 224596 244942 224608
rect 249018 224596 249024 224608
rect 249076 224596 249082 224648
rect 249754 224596 249760 224648
rect 249812 224636 249818 224648
rect 252624 224636 252652 224676
rect 256378 224664 256384 224676
rect 256436 224664 256442 224716
rect 249812 224608 252652 224636
rect 249812 224596 249818 224608
rect 56373 224571 56431 224577
rect 56373 224568 56385 224571
rect 53904 224540 56385 224568
rect 56373 224537 56385 224540
rect 56419 224537 56431 224571
rect 56373 224531 56431 224537
rect 57750 224528 57756 224580
rect 57808 224568 57814 224580
rect 61522 224568 61528 224580
rect 57808 224540 61528 224568
rect 57808 224528 57814 224540
rect 61522 224528 61528 224540
rect 61580 224528 61586 224580
rect 61801 224571 61859 224577
rect 61801 224537 61813 224571
rect 61847 224568 61859 224571
rect 68698 224568 68704 224580
rect 61847 224540 68704 224568
rect 61847 224537 61859 224540
rect 61801 224531 61859 224537
rect 68698 224528 68704 224540
rect 68756 224528 68762 224580
rect 158306 224528 158312 224580
rect 158364 224568 158370 224580
rect 161526 224568 161532 224580
rect 158364 224540 161532 224568
rect 158364 224528 158370 224540
rect 161526 224528 161532 224540
rect 161584 224528 161590 224580
rect 245246 224528 245252 224580
rect 245304 224568 245310 224580
rect 248650 224568 248656 224580
rect 245304 224540 248656 224568
rect 245304 224528 245310 224540
rect 248650 224528 248656 224540
rect 248708 224528 248714 224580
rect 249662 224528 249668 224580
rect 249720 224568 249726 224580
rect 253618 224568 253624 224580
rect 249720 224540 253624 224568
rect 249720 224528 249726 224540
rect 253618 224528 253624 224540
rect 253676 224528 253682 224580
rect 253713 224571 253771 224577
rect 253713 224537 253725 224571
rect 253759 224568 253771 224571
rect 254446 224568 254452 224580
rect 253759 224540 254452 224568
rect 253759 224537 253771 224540
rect 253713 224531 253771 224537
rect 254446 224528 254452 224540
rect 254504 224528 254510 224580
rect 57382 224460 57388 224512
rect 57440 224500 57446 224512
rect 61614 224500 61620 224512
rect 57440 224472 61620 224500
rect 57440 224460 57446 224472
rect 61614 224460 61620 224472
rect 61672 224460 61678 224512
rect 61706 224460 61712 224512
rect 61764 224500 61770 224512
rect 67134 224500 67140 224512
rect 61764 224472 67140 224500
rect 61764 224460 61770 224472
rect 67134 224460 67140 224472
rect 67192 224460 67198 224512
rect 151866 224460 151872 224512
rect 151924 224500 151930 224512
rect 158030 224500 158036 224512
rect 151924 224472 158036 224500
rect 151924 224460 151930 224472
rect 158030 224460 158036 224472
rect 158088 224460 158094 224512
rect 249386 224460 249392 224512
rect 249444 224500 249450 224512
rect 253250 224500 253256 224512
rect 249444 224472 253256 224500
rect 249444 224460 249450 224472
rect 253250 224460 253256 224472
rect 253308 224460 253314 224512
rect 60881 224435 60939 224441
rect 60881 224401 60893 224435
rect 60927 224432 60939 224435
rect 62810 224432 62816 224444
rect 60927 224404 62816 224432
rect 60927 224401 60939 224404
rect 60881 224395 60939 224401
rect 62810 224392 62816 224404
rect 62868 224392 62874 224444
rect 62902 224392 62908 224444
rect 62960 224432 62966 224444
rect 67962 224432 67968 224444
rect 62960 224404 67968 224432
rect 62960 224392 62966 224404
rect 67962 224392 67968 224404
rect 68020 224392 68026 224444
rect 155178 224392 155184 224444
rect 155236 224432 155242 224444
rect 159962 224432 159968 224444
rect 155236 224404 159968 224432
rect 155236 224392 155242 224404
rect 159962 224392 159968 224404
rect 160020 224392 160026 224444
rect 246442 224392 246448 224444
rect 246500 224432 246506 224444
rect 256194 224432 256200 224444
rect 246500 224404 256200 224432
rect 246500 224392 246506 224404
rect 256194 224392 256200 224404
rect 256252 224392 256258 224444
rect 55082 224324 55088 224376
rect 55140 224364 55146 224376
rect 59501 224367 59559 224373
rect 55140 224336 59452 224364
rect 55140 224324 55146 224336
rect 55726 224256 55732 224308
rect 55784 224296 55790 224308
rect 59317 224299 59375 224305
rect 59317 224296 59329 224299
rect 55784 224268 59329 224296
rect 55784 224256 55790 224268
rect 59317 224265 59329 224268
rect 59363 224265 59375 224299
rect 59424 224296 59452 224336
rect 59501 224333 59513 224367
rect 59547 224364 59559 224367
rect 65570 224364 65576 224376
rect 59547 224336 65576 224364
rect 59547 224333 59559 224336
rect 59501 224327 59559 224333
rect 65570 224324 65576 224336
rect 65628 224324 65634 224376
rect 153430 224324 153436 224376
rect 153488 224364 153494 224376
rect 158858 224364 158864 224376
rect 153488 224336 158864 224364
rect 153488 224324 153494 224336
rect 158858 224324 158864 224336
rect 158916 224324 158922 224376
rect 249938 224324 249944 224376
rect 249996 224364 250002 224376
rect 255182 224364 255188 224376
rect 249996 224336 255188 224364
rect 249996 224324 250002 224336
rect 255182 224324 255188 224336
rect 255240 224324 255246 224376
rect 61798 224296 61804 224308
rect 59424 224268 61804 224296
rect 59317 224259 59375 224265
rect 61798 224256 61804 224268
rect 61856 224256 61862 224308
rect 61890 224256 61896 224308
rect 61948 224296 61954 224308
rect 67502 224296 67508 224308
rect 61948 224268 67508 224296
rect 61948 224256 61954 224268
rect 67502 224256 67508 224268
rect 67560 224256 67566 224308
rect 152142 224256 152148 224308
rect 152200 224296 152206 224308
rect 162262 224296 162268 224308
rect 152200 224268 162268 224296
rect 152200 224256 152206 224268
rect 162262 224256 162268 224268
rect 162320 224256 162326 224308
rect 249570 224256 249576 224308
rect 249628 224296 249634 224308
rect 253713 224299 253771 224305
rect 253713 224296 253725 224299
rect 249628 224268 253725 224296
rect 249628 224256 249634 224268
rect 253713 224265 253725 224268
rect 253759 224265 253771 224299
rect 253713 224259 253771 224265
rect 253805 224299 253863 224305
rect 253805 224265 253817 224299
rect 253851 224296 253863 224299
rect 254814 224296 254820 224308
rect 253851 224268 254820 224296
rect 253851 224265 253863 224268
rect 253805 224259 253863 224265
rect 254814 224256 254820 224268
rect 254872 224256 254878 224308
rect 58946 224188 58952 224240
rect 59004 224228 59010 224240
rect 61154 224228 61160 224240
rect 59004 224200 61160 224228
rect 59004 224188 59010 224200
rect 61154 224188 61160 224200
rect 61212 224188 61218 224240
rect 61448 224200 68100 224228
rect 38246 224120 38252 224172
rect 38304 224160 38310 224172
rect 61448 224160 61476 224200
rect 67962 224160 67968 224172
rect 38304 224132 61476 224160
rect 61540 224132 67968 224160
rect 38304 224120 38310 224132
rect 59498 224052 59504 224104
rect 59556 224092 59562 224104
rect 61540 224092 61568 224132
rect 67962 224120 67968 224132
rect 68020 224120 68026 224172
rect 68072 224160 68100 224200
rect 154994 224188 155000 224240
rect 155052 224228 155058 224240
rect 160790 224228 160796 224240
rect 155052 224200 160796 224228
rect 155052 224188 155058 224200
rect 160790 224188 160796 224200
rect 160848 224188 160854 224240
rect 248374 224188 248380 224240
rect 248432 224228 248438 224240
rect 248432 224200 253940 224228
rect 248432 224188 248438 224200
rect 70630 224160 70636 224172
rect 68072 224132 70636 224160
rect 70630 224120 70636 224132
rect 70688 224120 70694 224172
rect 155822 224120 155828 224172
rect 155880 224160 155886 224172
rect 161986 224160 161992 224172
rect 155880 224132 161992 224160
rect 155880 224120 155886 224132
rect 161986 224120 161992 224132
rect 162044 224120 162050 224172
rect 250309 224163 250367 224169
rect 250309 224129 250321 224163
rect 250355 224160 250367 224163
rect 253805 224163 253863 224169
rect 253805 224160 253817 224163
rect 250355 224132 253817 224160
rect 250355 224129 250367 224132
rect 250309 224123 250367 224129
rect 253805 224129 253817 224132
rect 253851 224129 253863 224163
rect 253912 224160 253940 224200
rect 255550 224160 255556 224172
rect 253912 224132 255556 224160
rect 253805 224123 253863 224129
rect 255550 224120 255556 224132
rect 255608 224120 255614 224172
rect 59556 224064 61568 224092
rect 59556 224052 59562 224064
rect 137698 224052 137704 224104
rect 137756 224092 137762 224104
rect 146714 224092 146720 224104
rect 137756 224064 146720 224092
rect 137756 224052 137762 224064
rect 146714 224052 146720 224064
rect 146772 224052 146778 224104
rect 155914 224052 155920 224104
rect 155972 224092 155978 224104
rect 162354 224092 162360 224104
rect 155972 224064 162360 224092
rect 155972 224052 155978 224064
rect 162354 224052 162360 224064
rect 162412 224052 162418 224104
rect 231998 224052 232004 224104
rect 232056 224092 232062 224104
rect 240370 224092 240376 224104
rect 232056 224064 240376 224092
rect 232056 224052 232062 224064
rect 240370 224052 240376 224064
rect 240428 224052 240434 224104
rect 247362 224052 247368 224104
rect 247420 224092 247426 224104
rect 252790 224092 252796 224104
rect 247420 224064 252796 224092
rect 247420 224052 247426 224064
rect 252790 224052 252796 224064
rect 252848 224052 252854 224104
rect 59317 224027 59375 224033
rect 59317 223993 59329 224027
rect 59363 224024 59375 224027
rect 63730 224024 63736 224036
rect 59363 223996 63736 224024
rect 59363 223993 59375 223996
rect 59317 223987 59375 223993
rect 63730 223984 63736 223996
rect 63788 223984 63794 224036
rect 58857 223687 58915 223693
rect 58857 223653 58869 223687
rect 58903 223684 58915 223687
rect 63270 223684 63276 223696
rect 58903 223656 63276 223684
rect 58903 223653 58915 223656
rect 58857 223647 58915 223653
rect 63270 223644 63276 223656
rect 63328 223644 63334 223696
rect 257022 223032 257028 223084
rect 257080 223072 257086 223084
rect 257896 223072 257902 223084
rect 257080 223044 257902 223072
rect 257080 223032 257086 223044
rect 257896 223032 257902 223044
rect 257954 223032 257960 223084
rect 148738 221332 148744 221384
rect 148796 221372 148802 221384
rect 165114 221372 165120 221384
rect 148796 221344 165120 221372
rect 148796 221332 148802 221344
rect 165114 221332 165120 221344
rect 165172 221332 165178 221384
rect 231078 221332 231084 221384
rect 231136 221372 231142 221384
rect 239358 221372 239364 221384
rect 231136 221344 239364 221372
rect 231136 221332 231142 221344
rect 239358 221332 239364 221344
rect 239416 221332 239422 221384
rect 12946 219972 12952 220024
rect 13004 220012 13010 220024
rect 18834 220012 18840 220024
rect 13004 219984 18840 220012
rect 13004 219972 13010 219984
rect 18834 219972 18840 219984
rect 18892 219972 18898 220024
rect 230986 218816 230992 218868
rect 231044 218856 231050 218868
rect 232734 218856 232740 218868
rect 231044 218828 232740 218856
rect 231044 218816 231050 218828
rect 232734 218816 232740 218828
rect 232792 218816 232798 218868
rect 231722 218680 231728 218732
rect 231780 218720 231786 218732
rect 240922 218720 240928 218732
rect 231780 218692 240928 218720
rect 231780 218680 231786 218692
rect 240922 218680 240928 218692
rect 240980 218680 240986 218732
rect 137422 218612 137428 218664
rect 137480 218652 137486 218664
rect 145610 218652 145616 218664
rect 137480 218624 145616 218652
rect 137480 218612 137486 218624
rect 145610 218612 145616 218624
rect 145668 218612 145674 218664
rect 292810 217116 292816 217168
rect 292868 217156 292874 217168
rect 300170 217156 300176 217168
rect 292868 217128 300176 217156
rect 292868 217116 292874 217128
rect 300170 217116 300176 217128
rect 300228 217116 300234 217168
rect 231998 215960 232004 216012
rect 232056 216000 232062 216012
rect 238254 216000 238260 216012
rect 232056 215972 238260 216000
rect 232056 215960 232062 215972
rect 238254 215960 238260 215972
rect 238312 215960 238318 216012
rect 137330 215824 137336 215876
rect 137388 215864 137394 215876
rect 145610 215864 145616 215876
rect 137388 215836 145616 215864
rect 137388 215824 137394 215836
rect 145610 215824 145616 215836
rect 145668 215824 145674 215876
rect 231814 215824 231820 215876
rect 231872 215864 231878 215876
rect 240462 215864 240468 215876
rect 231872 215836 240468 215864
rect 231872 215824 231878 215836
rect 240462 215824 240468 215836
rect 240520 215824 240526 215876
rect 165114 215756 165120 215808
rect 165172 215796 165178 215808
rect 175510 215796 175516 215808
rect 165172 215768 175516 215796
rect 165172 215756 165178 215768
rect 175510 215756 175516 215768
rect 175568 215756 175574 215808
rect 137146 213104 137152 213156
rect 137204 213144 137210 213156
rect 145610 213144 145616 213156
rect 137204 213116 145616 213144
rect 137204 213104 137210 213116
rect 145610 213104 145616 213116
rect 145668 213104 145674 213156
rect 231906 213104 231912 213156
rect 231964 213144 231970 213156
rect 240922 213144 240928 213156
rect 231964 213116 240928 213144
rect 231964 213104 231970 213116
rect 240922 213104 240928 213116
rect 240980 213104 240986 213156
rect 262358 212832 262364 212884
rect 262416 212872 262422 212884
rect 265210 212872 265216 212884
rect 262416 212844 265216 212872
rect 262416 212832 262422 212844
rect 265210 212832 265216 212844
rect 265268 212832 265274 212884
rect 231998 212288 232004 212340
rect 232056 212328 232062 212340
rect 236874 212328 236880 212340
rect 232056 212300 236880 212328
rect 232056 212288 232062 212300
rect 236874 212288 236880 212300
rect 236932 212288 236938 212340
rect 137238 211676 137244 211728
rect 137296 211716 137302 211728
rect 145610 211716 145616 211728
rect 137296 211688 145616 211716
rect 137296 211676 137302 211688
rect 145610 211676 145616 211688
rect 145668 211676 145674 211728
rect 231630 211676 231636 211728
rect 231688 211716 231694 211728
rect 240922 211716 240928 211728
rect 231688 211688 240928 211716
rect 231688 211676 231694 211688
rect 240922 211676 240928 211688
rect 240980 211676 240986 211728
rect 231998 209228 232004 209280
rect 232056 209268 232062 209280
rect 235494 209268 235500 209280
rect 232056 209240 235500 209268
rect 232056 209228 232062 209240
rect 235494 209228 235500 209240
rect 235552 209228 235558 209280
rect 137054 208956 137060 209008
rect 137112 208996 137118 209008
rect 145610 208996 145616 209008
rect 137112 208968 145616 208996
rect 137112 208956 137118 208968
rect 145610 208956 145616 208968
rect 145668 208956 145674 209008
rect 231538 208956 231544 209008
rect 231596 208996 231602 209008
rect 240462 208996 240468 209008
rect 231596 208968 240468 208996
rect 231596 208956 231602 208968
rect 240462 208956 240468 208968
rect 240520 208956 240526 209008
rect 258954 208888 258960 208940
rect 259012 208928 259018 208940
rect 274870 208928 274876 208940
rect 259012 208900 274876 208928
rect 259012 208888 259018 208900
rect 274870 208888 274876 208900
rect 274928 208888 274934 208940
rect 231998 206440 232004 206492
rect 232056 206480 232062 206492
rect 234206 206480 234212 206492
rect 232056 206452 234212 206480
rect 232056 206440 232062 206452
rect 234206 206440 234212 206452
rect 234264 206440 234270 206492
rect 231998 206168 232004 206220
rect 232056 206208 232062 206220
rect 240646 206208 240652 206220
rect 232056 206180 240652 206208
rect 232056 206168 232062 206180
rect 240646 206168 240652 206180
rect 240704 206168 240710 206220
rect 136962 204808 136968 204860
rect 137020 204848 137026 204860
rect 145610 204848 145616 204860
rect 137020 204820 145616 204848
rect 137020 204808 137026 204820
rect 145610 204808 145616 204820
rect 145668 204808 145674 204860
rect 231446 204808 231452 204860
rect 231504 204848 231510 204860
rect 240922 204848 240928 204860
rect 231504 204820 240928 204848
rect 231504 204808 231510 204820
rect 240922 204808 240928 204820
rect 240980 204808 240986 204860
rect 143034 202020 143040 202072
rect 143092 202060 143098 202072
rect 145518 202060 145524 202072
rect 143092 202032 145524 202060
rect 143092 202020 143098 202032
rect 145518 202020 145524 202032
rect 145576 202020 145582 202072
rect 231262 202020 231268 202072
rect 231320 202060 231326 202072
rect 240370 202060 240376 202072
rect 231320 202032 240376 202060
rect 231320 202020 231326 202032
rect 240370 202020 240376 202032
rect 240428 202020 240434 202072
rect 231722 199300 231728 199352
rect 231780 199340 231786 199352
rect 240462 199340 240468 199352
rect 231780 199312 240468 199340
rect 231780 199300 231786 199312
rect 240462 199300 240468 199312
rect 240520 199300 240526 199352
rect 140274 197872 140280 197924
rect 140332 197912 140338 197924
rect 145610 197912 145616 197924
rect 140332 197884 145616 197912
rect 140332 197872 140338 197884
rect 145610 197872 145616 197884
rect 145668 197872 145674 197924
rect 231814 197872 231820 197924
rect 231872 197912 231878 197924
rect 240922 197912 240928 197924
rect 231872 197884 240928 197912
rect 231872 197872 231878 197884
rect 240922 197872 240928 197884
rect 240980 197872 240986 197924
rect 263738 196512 263744 196564
rect 263796 196552 263802 196564
rect 274870 196552 274876 196564
rect 263796 196524 274876 196552
rect 263796 196512 263802 196524
rect 274870 196512 274876 196524
rect 274928 196512 274934 196564
rect 140366 195152 140372 195204
rect 140424 195192 140430 195204
rect 145610 195192 145616 195204
rect 140424 195164 145616 195192
rect 140424 195152 140430 195164
rect 145610 195152 145616 195164
rect 145668 195152 145674 195204
rect 234298 195152 234304 195204
rect 234356 195192 234362 195204
rect 240922 195192 240928 195204
rect 234356 195164 240928 195192
rect 234356 195152 234362 195164
rect 240922 195152 240928 195164
rect 240980 195152 240986 195204
rect 137422 195084 137428 195136
rect 137480 195124 137486 195136
rect 145794 195124 145800 195136
rect 137480 195096 145800 195124
rect 137480 195084 137486 195096
rect 145794 195084 145800 195096
rect 145852 195084 145858 195136
rect 236966 192432 236972 192484
rect 237024 192472 237030 192484
rect 240462 192472 240468 192484
rect 237024 192444 240468 192472
rect 237024 192432 237030 192444
rect 240462 192432 240468 192444
rect 240520 192432 240526 192484
rect 143126 192364 143132 192416
rect 143184 192404 143190 192416
rect 145794 192404 145800 192416
rect 143184 192376 145800 192404
rect 143184 192364 143190 192376
rect 145794 192364 145800 192376
rect 145852 192364 145858 192416
rect 167874 192364 167880 192416
rect 167932 192404 167938 192416
rect 175510 192404 175516 192416
rect 167932 192376 175516 192404
rect 167932 192364 167938 192376
rect 175510 192364 175516 192376
rect 175568 192364 175574 192416
rect 262358 192364 262364 192416
rect 262416 192404 262422 192416
rect 275514 192404 275520 192416
rect 262416 192376 275520 192404
rect 262416 192364 262422 192376
rect 275514 192364 275520 192376
rect 275572 192364 275578 192416
rect 137422 191072 137428 191124
rect 137480 191112 137486 191124
rect 143034 191112 143040 191124
rect 137480 191084 143040 191112
rect 137480 191072 137486 191084
rect 143034 191072 143040 191084
rect 143092 191072 143098 191124
rect 74034 190936 74040 190988
rect 74092 190976 74098 190988
rect 81670 190976 81676 190988
rect 74092 190948 81676 190976
rect 74092 190936 74098 190948
rect 81670 190936 81676 190948
rect 81728 190936 81734 190988
rect 137054 189644 137060 189696
rect 137112 189684 137118 189696
rect 145150 189684 145156 189696
rect 137112 189656 145156 189684
rect 137112 189644 137118 189656
rect 145150 189644 145156 189656
rect 145208 189644 145214 189696
rect 230802 189644 230808 189696
rect 230860 189684 230866 189696
rect 240646 189684 240652 189696
rect 230860 189656 240652 189684
rect 230860 189644 230866 189656
rect 240646 189644 240652 189656
rect 240704 189644 240710 189696
rect 137422 189372 137428 189424
rect 137480 189412 137486 189424
rect 144414 189412 144420 189424
rect 137480 189384 144420 189412
rect 137480 189372 137486 189384
rect 144414 189372 144420 189384
rect 144472 189372 144478 189424
rect 292810 188896 292816 188948
rect 292868 188936 292874 188948
rect 293546 188936 293552 188948
rect 292868 188908 293552 188936
rect 292868 188896 292874 188908
rect 293546 188896 293552 188908
rect 293604 188896 293610 188948
rect 47078 188216 47084 188268
rect 47136 188256 47142 188268
rect 51310 188256 51316 188268
rect 47136 188228 51316 188256
rect 47136 188216 47142 188228
rect 51310 188216 51316 188228
rect 51368 188216 51374 188268
rect 137330 188216 137336 188268
rect 137388 188256 137394 188268
rect 145610 188256 145616 188268
rect 137388 188228 145616 188256
rect 137388 188216 137394 188228
rect 145610 188216 145616 188228
rect 145668 188216 145674 188268
rect 231262 188216 231268 188268
rect 231320 188256 231326 188268
rect 240738 188256 240744 188268
rect 231320 188228 240744 188256
rect 231320 188216 231326 188228
rect 240738 188216 240744 188228
rect 240796 188216 240802 188268
rect 137422 188148 137428 188200
rect 137480 188188 137486 188200
rect 140274 188188 140280 188200
rect 137480 188160 140280 188188
rect 137480 188148 137486 188160
rect 140274 188148 140280 188160
rect 140332 188148 140338 188200
rect 38798 186788 38804 186840
rect 38856 186828 38862 186840
rect 47078 186828 47084 186840
rect 38856 186800 47084 186828
rect 38856 186788 38862 186800
rect 47078 186788 47084 186800
rect 47136 186788 47142 186840
rect 137422 186788 137428 186840
rect 137480 186828 137486 186840
rect 140366 186828 140372 186840
rect 137480 186800 140372 186828
rect 137480 186788 137486 186800
rect 140366 186788 140372 186800
rect 140424 186788 140430 186840
rect 231814 186788 231820 186840
rect 231872 186828 231878 186840
rect 234298 186828 234304 186840
rect 231872 186800 234304 186828
rect 231872 186788 231878 186800
rect 234298 186788 234304 186800
rect 234356 186788 234362 186840
rect 237610 185496 237616 185548
rect 237668 185536 237674 185548
rect 240922 185536 240928 185548
rect 237668 185508 240928 185536
rect 237668 185496 237674 185508
rect 240922 185496 240928 185508
rect 240980 185496 240986 185548
rect 231814 185428 231820 185480
rect 231872 185468 231878 185480
rect 236966 185468 236972 185480
rect 231872 185440 236972 185468
rect 231872 185428 231878 185440
rect 236966 185428 236972 185440
rect 237024 185428 237030 185480
rect 137422 184204 137428 184256
rect 137480 184244 137486 184256
rect 143126 184244 143132 184256
rect 137480 184216 143132 184244
rect 137480 184204 137486 184216
rect 143126 184204 143132 184216
rect 143184 184204 143190 184256
rect 58857 181391 58915 181397
rect 58857 181357 58869 181391
rect 58903 181388 58915 181391
rect 63822 181388 63828 181400
rect 58903 181360 63828 181388
rect 58903 181357 58915 181360
rect 58857 181351 58915 181357
rect 63822 181348 63828 181360
rect 63880 181348 63886 181400
rect 156208 181360 157616 181388
rect 18834 181280 18840 181332
rect 18892 181320 18898 181332
rect 23710 181320 23716 181332
rect 18892 181292 23716 181320
rect 18892 181280 18898 181292
rect 23710 181280 23716 181292
rect 23768 181280 23774 181332
rect 23805 181323 23863 181329
rect 23805 181289 23817 181323
rect 23851 181320 23863 181323
rect 31622 181320 31628 181332
rect 23851 181292 31628 181320
rect 23851 181289 23863 181292
rect 23805 181283 23863 181289
rect 31622 181280 31628 181292
rect 31680 181280 31686 181332
rect 55818 181280 55824 181332
rect 55876 181320 55882 181332
rect 63730 181320 63736 181332
rect 55876 181292 63736 181320
rect 55876 181280 55882 181292
rect 63730 181280 63736 181292
rect 63788 181280 63794 181332
rect 150670 181280 150676 181332
rect 150728 181320 150734 181332
rect 151682 181320 151688 181332
rect 150728 181292 151688 181320
rect 150728 181280 150734 181292
rect 151682 181280 151688 181292
rect 151740 181280 151746 181332
rect 153062 181280 153068 181332
rect 153120 181320 153126 181332
rect 156208 181320 156236 181360
rect 153120 181292 156236 181320
rect 153120 181280 153126 181292
rect 156282 181280 156288 181332
rect 156340 181320 156346 181332
rect 157478 181320 157484 181332
rect 156340 181292 157484 181320
rect 156340 181280 156346 181292
rect 157478 181280 157484 181292
rect 157536 181280 157542 181332
rect 157588 181320 157616 181360
rect 249220 181360 250076 181388
rect 158398 181320 158404 181332
rect 157588 181292 158404 181320
rect 158398 181280 158404 181292
rect 158456 181280 158462 181332
rect 244418 181280 244424 181332
rect 244476 181320 244482 181332
rect 245430 181320 245436 181332
rect 244476 181292 245436 181320
rect 244476 181280 244482 181292
rect 245430 181280 245436 181292
rect 245488 181280 245494 181332
rect 58121 181255 58179 181261
rect 58121 181221 58133 181255
rect 58167 181252 58179 181255
rect 60881 181255 60939 181261
rect 60881 181252 60893 181255
rect 58167 181224 60893 181252
rect 58167 181221 58179 181224
rect 58121 181215 58179 181221
rect 60881 181221 60893 181224
rect 60927 181221 60939 181255
rect 60881 181215 60939 181221
rect 62074 181212 62080 181264
rect 62132 181252 62138 181264
rect 69802 181252 69808 181264
rect 62132 181224 69808 181252
rect 62132 181212 62138 181224
rect 69802 181212 69808 181224
rect 69860 181212 69866 181264
rect 149198 181212 149204 181264
rect 149256 181252 149262 181264
rect 160698 181252 160704 181264
rect 149256 181224 160704 181252
rect 149256 181212 149262 181224
rect 160698 181212 160704 181224
rect 160756 181212 160762 181264
rect 243314 181212 243320 181264
rect 243372 181252 243378 181264
rect 245154 181252 245160 181264
rect 243372 181224 245160 181252
rect 243372 181212 243378 181224
rect 245154 181212 245160 181224
rect 245212 181212 245218 181264
rect 245706 181212 245712 181264
rect 245764 181252 245770 181264
rect 249220 181252 249248 181360
rect 249570 181280 249576 181332
rect 249628 181320 249634 181332
rect 249938 181320 249944 181332
rect 249628 181292 249944 181320
rect 249628 181280 249634 181292
rect 249938 181280 249944 181292
rect 249996 181280 250002 181332
rect 250048 181320 250076 181360
rect 250490 181348 250496 181400
rect 250548 181388 250554 181400
rect 251505 181391 251563 181397
rect 251505 181388 251517 181391
rect 250548 181360 251517 181388
rect 250548 181348 250554 181360
rect 251505 181357 251517 181360
rect 251551 181357 251563 181391
rect 251505 181351 251563 181357
rect 253434 181320 253440 181332
rect 250048 181292 253440 181320
rect 253434 181280 253440 181292
rect 253492 181280 253498 181332
rect 253618 181280 253624 181332
rect 253676 181320 253682 181332
rect 255182 181320 255188 181332
rect 253676 181292 255188 181320
rect 253676 181280 253682 181292
rect 255182 181280 255188 181292
rect 255240 181280 255246 181332
rect 245764 181224 249248 181252
rect 245764 181212 245770 181224
rect 249294 181212 249300 181264
rect 249352 181252 249358 181264
rect 250766 181252 250772 181264
rect 249352 181224 250772 181252
rect 249352 181212 249358 181224
rect 250766 181212 250772 181224
rect 250824 181212 250830 181264
rect 250858 181212 250864 181264
rect 250916 181252 250922 181264
rect 253710 181252 253716 181264
rect 250916 181224 253716 181252
rect 250916 181212 250922 181224
rect 253710 181212 253716 181224
rect 253768 181212 253774 181264
rect 59866 181144 59872 181196
rect 59924 181184 59930 181196
rect 69894 181184 69900 181196
rect 59924 181156 69900 181184
rect 59924 181144 59930 181156
rect 69894 181144 69900 181156
rect 69952 181144 69958 181196
rect 145150 181144 145156 181196
rect 145208 181184 145214 181196
rect 157202 181184 157208 181196
rect 145208 181156 157208 181184
rect 145208 181144 145214 181156
rect 157202 181144 157208 181156
rect 157260 181144 157266 181196
rect 243038 181144 243044 181196
rect 243096 181184 243102 181196
rect 251410 181184 251416 181196
rect 243096 181156 251416 181184
rect 243096 181144 243102 181156
rect 251410 181144 251416 181156
rect 251468 181144 251474 181196
rect 251505 181187 251563 181193
rect 251505 181153 251517 181187
rect 251551 181184 251563 181187
rect 254265 181187 254323 181193
rect 254265 181184 254277 181187
rect 251551 181156 254277 181184
rect 251551 181153 251563 181156
rect 251505 181147 251563 181153
rect 254265 181153 254277 181156
rect 254311 181153 254323 181187
rect 254265 181147 254323 181153
rect 20214 181076 20220 181128
rect 20272 181116 20278 181128
rect 23805 181119 23863 181125
rect 23805 181116 23817 181119
rect 20272 181088 23817 181116
rect 20272 181076 20278 181088
rect 23805 181085 23817 181088
rect 23851 181085 23863 181119
rect 23805 181079 23863 181085
rect 59038 181076 59044 181128
rect 59096 181116 59102 181128
rect 69342 181116 69348 181128
rect 59096 181088 69348 181116
rect 59096 181076 59102 181088
rect 69342 181076 69348 181088
rect 69400 181076 69406 181128
rect 152234 181076 152240 181128
rect 152292 181116 152298 181128
rect 156929 181119 156987 181125
rect 156929 181116 156941 181119
rect 152292 181088 156941 181116
rect 152292 181076 152298 181088
rect 156929 181085 156941 181088
rect 156975 181085 156987 181119
rect 156929 181079 156987 181085
rect 245706 181076 245712 181128
rect 245764 181116 245770 181128
rect 248837 181119 248895 181125
rect 248837 181116 248849 181119
rect 245764 181088 248849 181116
rect 245764 181076 245770 181088
rect 248837 181085 248849 181088
rect 248883 181085 248895 181119
rect 248837 181079 248895 181085
rect 248926 181076 248932 181128
rect 248984 181116 248990 181128
rect 250674 181116 250680 181128
rect 248984 181088 250680 181116
rect 248984 181076 248990 181088
rect 250674 181076 250680 181088
rect 250732 181076 250738 181128
rect 251318 181076 251324 181128
rect 251376 181116 251382 181128
rect 257206 181116 257212 181128
rect 251376 181088 257212 181116
rect 251376 181076 251382 181088
rect 257206 181076 257212 181088
rect 257264 181076 257270 181128
rect 55450 181008 55456 181060
rect 55508 181048 55514 181060
rect 60421 181051 60479 181057
rect 60421 181048 60433 181051
rect 55508 181020 60433 181048
rect 55508 181008 55514 181020
rect 60421 181017 60433 181020
rect 60467 181017 60479 181051
rect 60421 181011 60479 181017
rect 62813 181051 62871 181057
rect 62813 181017 62825 181051
rect 62859 181048 62871 181051
rect 69250 181048 69256 181060
rect 62859 181020 69256 181048
rect 62859 181017 62871 181020
rect 62813 181011 62871 181017
rect 69250 181008 69256 181020
rect 69308 181008 69314 181060
rect 147726 181008 147732 181060
rect 147784 181048 147790 181060
rect 159502 181048 159508 181060
rect 147784 181020 159508 181048
rect 147784 181008 147790 181020
rect 159502 181008 159508 181020
rect 159560 181008 159566 181060
rect 245338 181008 245344 181060
rect 245396 181048 245402 181060
rect 249665 181051 249723 181057
rect 249665 181048 249677 181051
rect 245396 181020 249677 181048
rect 245396 181008 245402 181020
rect 249665 181017 249677 181020
rect 249711 181017 249723 181051
rect 249665 181011 249723 181017
rect 249754 181008 249760 181060
rect 249812 181048 249818 181060
rect 252422 181048 252428 181060
rect 249812 181020 252428 181048
rect 249812 181008 249818 181020
rect 252422 181008 252428 181020
rect 252480 181008 252486 181060
rect 53978 180940 53984 180992
rect 54036 180980 54042 180992
rect 65478 180980 65484 180992
rect 54036 180952 65484 180980
rect 54036 180940 54042 180952
rect 65478 180940 65484 180952
rect 65536 180940 65542 180992
rect 147818 180940 147824 180992
rect 147876 180980 147882 180992
rect 160238 180980 160244 180992
rect 147876 180952 160244 180980
rect 147876 180940 147882 180952
rect 160238 180940 160244 180952
rect 160296 180940 160302 180992
rect 242946 180940 242952 180992
rect 243004 180980 243010 180992
rect 251594 180980 251600 180992
rect 243004 180952 251600 180980
rect 243004 180940 243010 180952
rect 251594 180940 251600 180952
rect 251652 180940 251658 180992
rect 58670 180872 58676 180924
rect 58728 180912 58734 180924
rect 62813 180915 62871 180921
rect 62813 180912 62825 180915
rect 58728 180884 62825 180912
rect 58728 180872 58734 180884
rect 62813 180881 62825 180884
rect 62859 180881 62871 180915
rect 62813 180875 62871 180881
rect 62905 180915 62963 180921
rect 62905 180881 62917 180915
rect 62951 180912 62963 180915
rect 67042 180912 67048 180924
rect 62951 180884 67048 180912
rect 62951 180881 62963 180884
rect 62905 180875 62963 180881
rect 67042 180872 67048 180884
rect 67100 180872 67106 180924
rect 149474 180872 149480 180924
rect 149532 180912 149538 180924
rect 153154 180912 153160 180924
rect 149532 180884 153160 180912
rect 149532 180872 149538 180884
rect 153154 180872 153160 180884
rect 153212 180872 153218 180924
rect 153246 180872 153252 180924
rect 153304 180912 153310 180924
rect 157205 180915 157263 180921
rect 157205 180912 157217 180915
rect 153304 180884 157217 180912
rect 153304 180872 153310 180884
rect 157205 180881 157217 180884
rect 157251 180881 157263 180915
rect 157205 180875 157263 180881
rect 231630 180872 231636 180924
rect 231688 180912 231694 180924
rect 237610 180912 237616 180924
rect 231688 180884 237616 180912
rect 231688 180872 231694 180884
rect 237610 180872 237616 180884
rect 237668 180872 237674 180924
rect 242854 180872 242860 180924
rect 242912 180912 242918 180924
rect 251962 180912 251968 180924
rect 242912 180884 251968 180912
rect 242912 180872 242918 180884
rect 251962 180872 251968 180884
rect 252020 180872 252026 180924
rect 252054 180872 252060 180924
rect 252112 180912 252118 180924
rect 254814 180912 254820 180924
rect 252112 180884 254820 180912
rect 252112 180872 252118 180884
rect 254814 180872 254820 180884
rect 254872 180872 254878 180924
rect 56646 180804 56652 180856
rect 56704 180844 56710 180856
rect 65110 180844 65116 180856
rect 56704 180816 65116 180844
rect 56704 180804 56710 180816
rect 65110 180804 65116 180816
rect 65168 180804 65174 180856
rect 147634 180804 147640 180856
rect 147692 180844 147698 180856
rect 159870 180844 159876 180856
rect 147692 180816 159876 180844
rect 147692 180804 147698 180816
rect 159870 180804 159876 180816
rect 159928 180804 159934 180856
rect 244878 180804 244884 180856
rect 244936 180844 244942 180856
rect 248745 180847 248803 180853
rect 248745 180844 248757 180847
rect 244936 180816 248757 180844
rect 244936 180804 244942 180816
rect 248745 180813 248757 180816
rect 248791 180813 248803 180847
rect 248745 180807 248803 180813
rect 248837 180847 248895 180853
rect 248837 180813 248849 180847
rect 248883 180844 248895 180847
rect 254170 180844 254176 180856
rect 248883 180816 254176 180844
rect 248883 180813 248895 180816
rect 248837 180807 248895 180813
rect 254170 180804 254176 180816
rect 254228 180804 254234 180856
rect 60881 180779 60939 180785
rect 60881 180745 60893 180779
rect 60927 180776 60939 180779
rect 63454 180776 63460 180788
rect 60927 180748 63460 180776
rect 60927 180745 60939 180748
rect 60881 180739 60939 180745
rect 63454 180736 63460 180748
rect 63512 180736 63518 180788
rect 146438 180736 146444 180788
rect 146496 180776 146502 180788
rect 159042 180776 159048 180788
rect 146496 180748 159048 180776
rect 146496 180736 146502 180748
rect 159042 180736 159048 180748
rect 159100 180736 159106 180788
rect 159137 180779 159195 180785
rect 159137 180745 159149 180779
rect 159183 180776 159195 180779
rect 163090 180776 163096 180788
rect 159183 180748 163096 180776
rect 159183 180745 159195 180748
rect 159137 180739 159195 180745
rect 163090 180736 163096 180748
rect 163148 180736 163154 180788
rect 247178 180736 247184 180788
rect 247236 180776 247242 180788
rect 251045 180779 251103 180785
rect 251045 180776 251057 180779
rect 247236 180748 251057 180776
rect 247236 180736 247242 180748
rect 251045 180745 251057 180748
rect 251091 180745 251103 180779
rect 251045 180739 251103 180745
rect 251134 180736 251140 180788
rect 251192 180776 251198 180788
rect 257574 180776 257580 180788
rect 251192 180748 257580 180776
rect 251192 180736 251198 180748
rect 257574 180736 257580 180748
rect 257632 180736 257638 180788
rect 49838 180668 49844 180720
rect 49896 180708 49902 180720
rect 49896 180680 56140 180708
rect 49896 180668 49902 180680
rect 51126 180600 51132 180652
rect 51184 180640 51190 180652
rect 51184 180612 51356 180640
rect 51184 180600 51190 180612
rect 51328 180164 51356 180612
rect 56112 180572 56140 180680
rect 58210 180668 58216 180720
rect 58268 180708 58274 180720
rect 63365 180711 63423 180717
rect 63365 180708 63377 180711
rect 58268 180680 63377 180708
rect 58268 180668 58274 180680
rect 63365 180677 63377 180680
rect 63411 180677 63423 180711
rect 63365 180671 63423 180677
rect 63546 180668 63552 180720
rect 63604 180708 63610 180720
rect 70630 180708 70636 180720
rect 63604 180680 70636 180708
rect 63604 180668 63610 180680
rect 70630 180668 70636 180680
rect 70688 180668 70694 180720
rect 144874 180668 144880 180720
rect 144932 180708 144938 180720
rect 158306 180708 158312 180720
rect 144932 180680 158312 180708
rect 144932 180668 144938 180680
rect 158306 180668 158312 180680
rect 158364 180668 158370 180720
rect 246902 180668 246908 180720
rect 246960 180708 246966 180720
rect 250401 180711 250459 180717
rect 250401 180708 250413 180711
rect 246960 180680 250413 180708
rect 246960 180668 246966 180680
rect 250401 180677 250413 180680
rect 250447 180677 250459 180711
rect 250401 180671 250459 180677
rect 56278 180600 56284 180652
rect 56336 180640 56342 180652
rect 65202 180640 65208 180652
rect 56336 180612 65208 180640
rect 56336 180600 56342 180612
rect 65202 180600 65208 180612
rect 65260 180600 65266 180652
rect 144966 180600 144972 180652
rect 145024 180640 145030 180652
rect 157846 180640 157852 180652
rect 145024 180612 157852 180640
rect 145024 180600 145030 180612
rect 157846 180600 157852 180612
rect 157904 180600 157910 180652
rect 158214 180600 158220 180652
rect 158272 180640 158278 180652
rect 164654 180640 164660 180652
rect 158272 180612 164660 180640
rect 158272 180600 158278 180612
rect 164654 180600 164660 180612
rect 164712 180600 164718 180652
rect 242394 180600 242400 180652
rect 242452 180640 242458 180652
rect 251042 180640 251048 180652
rect 242452 180612 251048 180640
rect 242452 180600 242458 180612
rect 251042 180600 251048 180612
rect 251100 180600 251106 180652
rect 253158 180640 253164 180652
rect 251152 180612 253164 180640
rect 63086 180572 63092 180584
rect 56112 180544 63092 180572
rect 63086 180532 63092 180544
rect 63144 180532 63150 180584
rect 63365 180575 63423 180581
rect 63365 180541 63377 180575
rect 63411 180572 63423 180575
rect 65754 180572 65760 180584
rect 63411 180544 65760 180572
rect 63411 180541 63423 180544
rect 63365 180535 63423 180541
rect 65754 180532 65760 180544
rect 65812 180532 65818 180584
rect 153430 180532 153436 180584
rect 153488 180572 153494 180584
rect 163826 180572 163832 180584
rect 153488 180544 163832 180572
rect 153488 180532 153494 180544
rect 163826 180532 163832 180544
rect 163884 180532 163890 180584
rect 245798 180532 245804 180584
rect 245856 180572 245862 180584
rect 251152 180572 251180 180612
rect 253158 180600 253164 180612
rect 253216 180600 253222 180652
rect 254265 180643 254323 180649
rect 254265 180609 254277 180643
rect 254311 180640 254323 180643
rect 261070 180640 261076 180652
rect 254311 180612 261076 180640
rect 254311 180609 254323 180612
rect 254265 180603 254323 180609
rect 261070 180600 261076 180612
rect 261128 180600 261134 180652
rect 245856 180544 251180 180572
rect 245856 180532 245862 180544
rect 251226 180532 251232 180584
rect 251284 180572 251290 180584
rect 258310 180572 258316 180584
rect 251284 180544 258316 180572
rect 251284 180532 251290 180544
rect 258310 180532 258316 180544
rect 258368 180532 258374 180584
rect 52506 180464 52512 180516
rect 52564 180504 52570 180516
rect 64282 180504 64288 180516
rect 52564 180476 64288 180504
rect 52564 180464 52570 180476
rect 64282 180464 64288 180476
rect 64340 180464 64346 180516
rect 150302 180464 150308 180516
rect 150360 180504 150366 180516
rect 152970 180504 152976 180516
rect 150360 180476 152976 180504
rect 150360 180464 150366 180476
rect 152970 180464 152976 180476
rect 153028 180464 153034 180516
rect 155454 180464 155460 180516
rect 155512 180504 155518 180516
rect 156098 180504 156104 180516
rect 155512 180476 156104 180504
rect 155512 180464 155518 180476
rect 156098 180464 156104 180476
rect 156156 180464 156162 180516
rect 156929 180507 156987 180513
rect 156929 180473 156941 180507
rect 156975 180504 156987 180507
rect 162446 180504 162452 180516
rect 156975 180476 162452 180504
rect 156975 180473 156987 180476
rect 156929 180467 156987 180473
rect 162446 180464 162452 180476
rect 162504 180464 162510 180516
rect 243682 180464 243688 180516
rect 243740 180504 243746 180516
rect 245246 180504 245252 180516
rect 243740 180476 245252 180504
rect 243740 180464 243746 180476
rect 245246 180464 245252 180476
rect 245304 180464 245310 180516
rect 246074 180464 246080 180516
rect 246132 180504 246138 180516
rect 249202 180504 249208 180516
rect 246132 180476 249208 180504
rect 246132 180464 246138 180476
rect 249202 180464 249208 180476
rect 249260 180464 249266 180516
rect 249294 180464 249300 180516
rect 249352 180504 249358 180516
rect 252790 180504 252796 180516
rect 249352 180476 252796 180504
rect 249352 180464 249358 180476
rect 252790 180464 252796 180476
rect 252848 180464 252854 180516
rect 52598 180396 52604 180448
rect 52656 180436 52662 180448
rect 64650 180436 64656 180448
rect 52656 180408 64656 180436
rect 52656 180396 52662 180408
rect 64650 180396 64656 180408
rect 64708 180396 64714 180448
rect 151774 180396 151780 180448
rect 151832 180436 151838 180448
rect 162630 180436 162636 180448
rect 151832 180408 162636 180436
rect 151832 180396 151838 180408
rect 162630 180396 162636 180408
rect 162688 180396 162694 180448
rect 247178 180396 247184 180448
rect 247236 180436 247242 180448
rect 254354 180436 254360 180448
rect 247236 180408 254360 180436
rect 247236 180396 247242 180408
rect 254354 180396 254360 180408
rect 254412 180396 254418 180448
rect 57014 180328 57020 180380
rect 57072 180368 57078 180380
rect 60602 180368 60608 180380
rect 57072 180340 60608 180368
rect 57072 180328 57078 180340
rect 60602 180328 60608 180340
rect 60660 180328 60666 180380
rect 63086 180328 63092 180380
rect 63144 180368 63150 180380
rect 68606 180368 68612 180380
rect 63144 180340 68612 180368
rect 63144 180328 63150 180340
rect 68606 180328 68612 180340
rect 68664 180328 68670 180380
rect 146346 180328 146352 180380
rect 146404 180368 146410 180380
rect 146404 180340 153844 180368
rect 146404 180328 146410 180340
rect 63917 180303 63975 180309
rect 63917 180269 63929 180303
rect 63963 180300 63975 180303
rect 70262 180300 70268 180312
rect 63963 180272 70268 180300
rect 63963 180269 63975 180272
rect 63917 180263 63975 180269
rect 70262 180260 70268 180272
rect 70320 180260 70326 180312
rect 152050 180260 152056 180312
rect 152108 180300 152114 180312
rect 153341 180303 153399 180309
rect 153341 180300 153353 180303
rect 152108 180272 153353 180300
rect 152108 180260 152114 180272
rect 153341 180269 153353 180272
rect 153387 180269 153399 180303
rect 153816 180300 153844 180340
rect 153890 180328 153896 180380
rect 153948 180368 153954 180380
rect 163734 180368 163740 180380
rect 153948 180340 163740 180368
rect 153948 180328 153954 180340
rect 163734 180328 163740 180340
rect 163792 180328 163798 180380
rect 249846 180328 249852 180380
rect 249904 180368 249910 180380
rect 256378 180368 256384 180380
rect 249904 180340 256384 180368
rect 249904 180328 249910 180340
rect 256378 180328 256384 180340
rect 256436 180328 256442 180380
rect 158674 180300 158680 180312
rect 153816 180272 158680 180300
rect 153341 180263 153399 180269
rect 158674 180260 158680 180272
rect 158732 180260 158738 180312
rect 248745 180303 248803 180309
rect 248745 180269 248757 180303
rect 248791 180300 248803 180303
rect 253710 180300 253716 180312
rect 248791 180272 253716 180300
rect 248791 180269 248803 180272
rect 248745 180263 248803 180269
rect 253710 180260 253716 180272
rect 253768 180260 253774 180312
rect 55082 180192 55088 180244
rect 55140 180232 55146 180244
rect 60142 180232 60148 180244
rect 55140 180204 60148 180232
rect 55140 180192 55146 180204
rect 60142 180192 60148 180204
rect 60200 180192 60206 180244
rect 60418 180192 60424 180244
rect 60476 180232 60482 180244
rect 66674 180232 66680 180244
rect 60476 180204 66680 180232
rect 60476 180192 60482 180204
rect 66674 180192 66680 180204
rect 66732 180192 66738 180244
rect 153157 180235 153215 180241
rect 153157 180201 153169 180235
rect 153203 180232 153215 180235
rect 157110 180232 157116 180244
rect 153203 180204 157116 180232
rect 153203 180201 153215 180204
rect 153157 180195 153215 180201
rect 157110 180192 157116 180204
rect 157168 180192 157174 180244
rect 157205 180235 157263 180241
rect 157205 180201 157217 180235
rect 157251 180232 157263 180235
rect 162354 180232 162360 180244
rect 157251 180204 162360 180232
rect 157251 180201 157263 180204
rect 157205 180195 157263 180201
rect 162354 180192 162360 180204
rect 162412 180192 162418 180244
rect 247730 180192 247736 180244
rect 247788 180232 247794 180244
rect 249570 180232 249576 180244
rect 247788 180204 249576 180232
rect 247788 180192 247794 180204
rect 249570 180192 249576 180204
rect 249628 180192 249634 180244
rect 249665 180235 249723 180241
rect 249665 180201 249677 180235
rect 249711 180232 249723 180235
rect 253526 180232 253532 180244
rect 249711 180204 253532 180232
rect 249711 180201 249723 180204
rect 249665 180195 249723 180201
rect 253526 180192 253532 180204
rect 253584 180192 253590 180244
rect 58857 180167 58915 180173
rect 58857 180164 58869 180167
rect 51328 180136 58869 180164
rect 58857 180133 58869 180136
rect 58903 180133 58915 180167
rect 58857 180127 58915 180133
rect 60050 180124 60056 180176
rect 60108 180164 60114 180176
rect 62905 180167 62963 180173
rect 62905 180164 62917 180167
rect 60108 180136 62917 180164
rect 60108 180124 60114 180136
rect 62905 180133 62917 180136
rect 62951 180133 62963 180167
rect 62905 180127 62963 180133
rect 62994 180124 63000 180176
rect 63052 180164 63058 180176
rect 68238 180164 68244 180176
rect 63052 180136 68244 180164
rect 63052 180124 63058 180136
rect 68238 180124 68244 180136
rect 68296 180124 68302 180176
rect 149106 180124 149112 180176
rect 149164 180164 149170 180176
rect 152878 180164 152884 180176
rect 149164 180136 152884 180164
rect 149164 180124 149170 180136
rect 152878 180124 152884 180136
rect 152936 180124 152942 180176
rect 156834 180164 156840 180176
rect 153080 180136 156840 180164
rect 57566 180056 57572 180108
rect 57624 180096 57630 180108
rect 65018 180096 65024 180108
rect 57624 180068 65024 180096
rect 57624 180056 57630 180068
rect 65018 180056 65024 180068
rect 65076 180056 65082 180108
rect 149842 180056 149848 180108
rect 149900 180096 149906 180108
rect 152786 180096 152792 180108
rect 149900 180068 152792 180096
rect 149900 180056 149906 180068
rect 152786 180056 152792 180068
rect 152844 180056 152850 180108
rect 57474 179988 57480 180040
rect 57532 180028 57538 180040
rect 60234 180028 60240 180040
rect 57532 180000 60240 180028
rect 57532 179988 57538 180000
rect 60234 179988 60240 180000
rect 60292 179988 60298 180040
rect 60421 180031 60479 180037
rect 60421 179997 60433 180031
rect 60467 180028 60479 180031
rect 63730 180028 63736 180040
rect 60467 180000 63736 180028
rect 60467 179997 60479 180000
rect 60421 179991 60479 179997
rect 63730 179988 63736 180000
rect 63788 179988 63794 180040
rect 64466 179988 64472 180040
rect 64524 180028 64530 180040
rect 69434 180028 69440 180040
rect 64524 180000 69440 180028
rect 64524 179988 64530 180000
rect 69434 179988 69440 180000
rect 69492 179988 69498 180040
rect 137422 179988 137428 180040
rect 137480 180028 137486 180040
rect 144782 180028 144788 180040
rect 137480 180000 144788 180028
rect 137480 179988 137486 180000
rect 144782 179988 144788 180000
rect 144840 179988 144846 180040
rect 151038 179988 151044 180040
rect 151096 180028 151102 180040
rect 153080 180028 153108 180136
rect 156834 180124 156840 180136
rect 156892 180124 156898 180176
rect 159137 180167 159195 180173
rect 159137 180164 159149 180167
rect 156944 180136 159149 180164
rect 153341 180099 153399 180105
rect 153341 180065 153353 180099
rect 153387 180096 153399 180099
rect 156944 180096 156972 180136
rect 159137 180133 159149 180136
rect 159183 180133 159195 180167
rect 159137 180127 159195 180133
rect 248834 180124 248840 180176
rect 248892 180164 248898 180176
rect 250401 180167 250459 180173
rect 248892 180136 249524 180164
rect 248892 180124 248898 180136
rect 153387 180068 156972 180096
rect 157481 180099 157539 180105
rect 153387 180065 153399 180068
rect 153341 180059 153399 180065
rect 157481 180065 157493 180099
rect 157527 180096 157539 180099
rect 163458 180096 163464 180108
rect 157527 180068 163464 180096
rect 157527 180065 157539 180068
rect 157481 180059 157539 180065
rect 163458 180056 163464 180068
rect 163516 180056 163522 180108
rect 244142 180056 244148 180108
rect 244200 180096 244206 180108
rect 245338 180096 245344 180108
rect 244200 180068 245344 180096
rect 244200 180056 244206 180068
rect 245338 180056 245344 180068
rect 245396 180056 245402 180108
rect 246534 180056 246540 180108
rect 246592 180096 246598 180108
rect 248926 180096 248932 180108
rect 246592 180068 248932 180096
rect 246592 180056 246598 180068
rect 248926 180056 248932 180068
rect 248984 180056 248990 180108
rect 151096 180000 153108 180028
rect 151096 179988 151102 180000
rect 153246 179988 153252 180040
rect 153304 180028 153310 180040
rect 154905 180031 154963 180037
rect 154905 180028 154917 180031
rect 153304 180000 154917 180028
rect 153304 179988 153310 180000
rect 154905 179997 154917 180000
rect 154951 179997 154963 180031
rect 154905 179991 154963 179997
rect 157018 179988 157024 180040
rect 157076 180028 157082 180040
rect 164286 180028 164292 180040
rect 157076 180000 164292 180028
rect 157076 179988 157082 180000
rect 164286 179988 164292 180000
rect 164344 179988 164350 180040
rect 248098 179988 248104 180040
rect 248156 180028 248162 180040
rect 249386 180028 249392 180040
rect 248156 180000 249392 180028
rect 248156 179988 248162 180000
rect 249386 179988 249392 180000
rect 249444 179988 249450 180040
rect 57842 179920 57848 179972
rect 57900 179960 57906 179972
rect 57900 179932 59912 179960
rect 57900 179920 57906 179932
rect 59884 179824 59912 179932
rect 61062 179920 61068 179972
rect 61120 179960 61126 179972
rect 61798 179960 61804 179972
rect 61120 179932 61804 179960
rect 61120 179920 61126 179932
rect 61798 179920 61804 179932
rect 61856 179920 61862 179972
rect 61890 179920 61896 179972
rect 61948 179960 61954 179972
rect 62258 179960 62264 179972
rect 61948 179932 62264 179960
rect 61948 179920 61954 179932
rect 62258 179920 62264 179932
rect 62316 179920 62322 179972
rect 62626 179920 62632 179972
rect 62684 179960 62690 179972
rect 63638 179960 63644 179972
rect 62684 179932 63644 179960
rect 62684 179920 62690 179932
rect 63638 179920 63644 179932
rect 63696 179920 63702 179972
rect 63917 179963 63975 179969
rect 63917 179960 63929 179963
rect 63748 179932 63929 179960
rect 60510 179824 60516 179836
rect 59884 179796 60516 179824
rect 60510 179784 60516 179796
rect 60568 179784 60574 179836
rect 62258 179784 62264 179836
rect 62316 179824 62322 179836
rect 63748 179824 63776 179932
rect 63917 179929 63929 179932
rect 63963 179929 63975 179963
rect 63917 179923 63975 179929
rect 64374 179920 64380 179972
rect 64432 179960 64438 179972
rect 69066 179960 69072 179972
rect 64432 179932 69072 179960
rect 64432 179920 64438 179932
rect 69066 179920 69072 179932
rect 69124 179920 69130 179972
rect 143678 179920 143684 179972
rect 143736 179960 143742 179972
rect 153157 179963 153215 179969
rect 153157 179960 153169 179963
rect 143736 179932 153169 179960
rect 143736 179920 143742 179932
rect 153157 179929 153169 179932
rect 153203 179929 153215 179963
rect 153157 179923 153215 179929
rect 153338 179920 153344 179972
rect 153396 179960 153402 179972
rect 155273 179963 155331 179969
rect 155273 179960 155285 179963
rect 153396 179932 155285 179960
rect 153396 179920 153402 179932
rect 155273 179929 155285 179932
rect 155319 179929 155331 179963
rect 157481 179963 157539 179969
rect 157481 179960 157493 179963
rect 155273 179923 155331 179929
rect 155840 179932 157493 179960
rect 137422 179852 137428 179904
rect 137480 179892 137486 179904
rect 145794 179892 145800 179904
rect 137480 179864 145800 179892
rect 137480 179852 137486 179864
rect 145794 179852 145800 179864
rect 145852 179852 145858 179904
rect 154905 179895 154963 179901
rect 154905 179861 154917 179895
rect 154951 179892 154963 179895
rect 155840 179892 155868 179932
rect 157481 179929 157493 179932
rect 157527 179929 157539 179963
rect 163550 179960 163556 179972
rect 157481 179923 157539 179929
rect 157588 179932 163556 179960
rect 154951 179864 155868 179892
rect 154951 179861 154963 179864
rect 154905 179855 154963 179861
rect 62316 179796 63776 179824
rect 155273 179827 155331 179833
rect 62316 179784 62322 179796
rect 155273 179793 155285 179827
rect 155319 179824 155331 179827
rect 157588 179824 157616 179932
rect 163550 179920 163556 179932
rect 163608 179920 163614 179972
rect 248374 179920 248380 179972
rect 248432 179960 248438 179972
rect 249018 179960 249024 179972
rect 248432 179932 249024 179960
rect 248432 179920 248438 179932
rect 249018 179920 249024 179932
rect 249076 179920 249082 179972
rect 249496 179960 249524 180136
rect 250401 180133 250413 180167
rect 250447 180164 250459 180167
rect 257022 180164 257028 180176
rect 250447 180136 257028 180164
rect 250447 180133 250459 180136
rect 250401 180127 250459 180133
rect 257022 180124 257028 180136
rect 257080 180124 257086 180176
rect 250582 180056 250588 180108
rect 250640 180096 250646 180108
rect 250950 180096 250956 180108
rect 250640 180068 250956 180096
rect 250640 180056 250646 180068
rect 250950 180056 250956 180068
rect 251008 180056 251014 180108
rect 252698 180056 252704 180108
rect 252756 180096 252762 180108
rect 258402 180096 258408 180108
rect 252756 180068 258408 180096
rect 252756 180056 252762 180068
rect 258402 180056 258408 180068
rect 258460 180056 258466 180108
rect 251045 180031 251103 180037
rect 251045 179997 251057 180031
rect 251091 180028 251103 180031
rect 256930 180028 256936 180040
rect 251091 180000 256936 180028
rect 251091 179997 251103 180000
rect 251045 179991 251103 179997
rect 256930 179988 256936 180000
rect 256988 179988 256994 180040
rect 257114 179960 257120 179972
rect 249496 179932 257120 179960
rect 257114 179920 257120 179932
rect 257172 179920 257178 179972
rect 231630 179852 231636 179904
rect 231688 179892 231694 179904
rect 239634 179892 239640 179904
rect 231688 179864 239640 179892
rect 231688 179852 231694 179864
rect 239634 179852 239640 179864
rect 239692 179852 239698 179904
rect 155319 179796 157616 179824
rect 155319 179793 155331 179796
rect 155273 179787 155331 179793
rect 88202 177948 88208 178000
rect 88260 177948 88266 178000
rect 86822 177880 86828 177932
rect 86880 177920 86886 177932
rect 86880 177892 87144 177920
rect 86880 177880 86886 177892
rect 87116 177796 87144 177892
rect 87098 177744 87104 177796
rect 87156 177744 87162 177796
rect 88220 177784 88248 177948
rect 90870 177880 90876 177932
rect 90928 177920 90934 177932
rect 90928 177892 91284 177920
rect 90928 177880 90934 177892
rect 91256 177796 91284 177892
rect 88478 177784 88484 177796
rect 88220 177756 88484 177784
rect 88478 177744 88484 177756
rect 88536 177744 88542 177796
rect 91238 177744 91244 177796
rect 91296 177744 91302 177796
rect 249570 176248 249576 176300
rect 249628 176248 249634 176300
rect 249588 176096 249616 176248
rect 249570 176044 249576 176096
rect 249628 176044 249634 176096
rect 85534 175772 85540 175824
rect 85592 175812 85598 175824
rect 179558 175812 179564 175824
rect 85592 175784 179564 175812
rect 85592 175772 85598 175784
rect 179558 175772 179564 175784
rect 179616 175772 179622 175824
rect 188942 175772 188948 175824
rect 189000 175812 189006 175824
rect 198234 175812 198240 175824
rect 189000 175784 198240 175812
rect 189000 175772 189006 175784
rect 198234 175772 198240 175784
rect 198292 175772 198298 175824
rect 200353 175815 200411 175821
rect 200353 175781 200365 175815
rect 200399 175812 200411 175815
rect 205137 175815 205195 175821
rect 205137 175812 205149 175815
rect 200399 175784 205149 175812
rect 200399 175781 200411 175784
rect 200353 175775 200411 175781
rect 205137 175781 205149 175784
rect 205183 175781 205195 175815
rect 205137 175775 205195 175781
rect 228686 175772 228692 175824
rect 228744 175812 228750 175824
rect 261162 175812 261168 175824
rect 228744 175784 261168 175812
rect 228744 175772 228750 175784
rect 261162 175772 261168 175784
rect 261220 175772 261226 175824
rect 94918 175704 94924 175756
rect 94976 175744 94982 175756
rect 104210 175744 104216 175756
rect 94976 175716 104216 175744
rect 94976 175704 94982 175716
rect 104210 175704 104216 175716
rect 104268 175704 104274 175756
rect 132730 175704 132736 175756
rect 132788 175744 132794 175756
rect 226754 175744 226760 175756
rect 132788 175716 226760 175744
rect 132788 175704 132794 175716
rect 226754 175704 226760 175716
rect 226812 175704 226818 175756
rect 103753 175679 103811 175685
rect 103753 175645 103765 175679
rect 103799 175676 103811 175679
rect 115158 175676 115164 175688
rect 103799 175648 115164 175676
rect 103799 175645 103811 175648
rect 103753 175639 103811 175645
rect 115158 175636 115164 175648
rect 115216 175636 115222 175688
rect 173394 175636 173400 175688
rect 173452 175676 173458 175688
rect 203846 175676 203852 175688
rect 173452 175648 203852 175676
rect 173452 175636 173458 175648
rect 203846 175636 203852 175648
rect 203904 175636 203910 175688
rect 205137 175679 205195 175685
rect 205137 175645 205149 175679
rect 205183 175676 205195 175679
rect 211942 175676 211948 175688
rect 205183 175648 211948 175676
rect 205183 175645 205195 175648
rect 205137 175639 205195 175645
rect 211942 175636 211948 175648
rect 212000 175636 212006 175688
rect 79738 175568 79744 175620
rect 79796 175608 79802 175620
rect 109822 175608 109828 175620
rect 79796 175580 109828 175608
rect 79796 175568 79802 175580
rect 109822 175568 109828 175580
rect 109880 175568 109886 175620
rect 111110 175568 111116 175620
rect 111168 175608 111174 175620
rect 140274 175608 140280 175620
rect 111168 175580 140280 175608
rect 111168 175568 111174 175580
rect 140274 175568 140280 175580
rect 140332 175568 140338 175620
rect 173854 175568 173860 175620
rect 173912 175608 173918 175620
rect 206514 175608 206520 175620
rect 173912 175580 206520 175608
rect 173912 175568 173918 175580
rect 206514 175568 206520 175580
rect 206572 175568 206578 175620
rect 228134 175568 228140 175620
rect 228192 175608 228198 175620
rect 228686 175608 228692 175620
rect 228192 175580 228692 175608
rect 228192 175568 228198 175580
rect 228686 175568 228692 175580
rect 228744 175568 228750 175620
rect 79554 175500 79560 175552
rect 79612 175540 79618 175552
rect 112490 175540 112496 175552
rect 79612 175512 112496 175540
rect 79612 175500 79618 175512
rect 112490 175500 112496 175512
rect 112548 175500 112554 175552
rect 173670 175500 173676 175552
rect 173728 175540 173734 175552
rect 209182 175540 209188 175552
rect 173728 175512 209188 175540
rect 173728 175500 173734 175512
rect 209182 175500 209188 175512
rect 209240 175500 209246 175552
rect 213230 175500 213236 175552
rect 213288 175540 213294 175552
rect 213288 175512 221464 175540
rect 213288 175500 213294 175512
rect 51218 175432 51224 175484
rect 51276 175472 51282 175484
rect 58121 175475 58179 175481
rect 58121 175472 58133 175475
rect 51276 175444 58133 175472
rect 51276 175432 51282 175444
rect 58121 175441 58133 175444
rect 58167 175441 58179 175475
rect 58121 175435 58179 175441
rect 65570 175432 65576 175484
rect 65628 175472 65634 175484
rect 65846 175472 65852 175484
rect 65628 175444 65852 175472
rect 65628 175432 65634 175444
rect 65846 175432 65852 175444
rect 65904 175432 65910 175484
rect 79646 175432 79652 175484
rect 79704 175472 79710 175484
rect 103753 175475 103811 175481
rect 103753 175472 103765 175475
rect 79704 175444 103765 175472
rect 79704 175432 79710 175444
rect 103753 175441 103765 175444
rect 103799 175441 103811 175475
rect 103753 175435 103811 175441
rect 152694 175432 152700 175484
rect 152752 175472 152758 175484
rect 152970 175472 152976 175484
rect 152752 175444 152976 175472
rect 152752 175432 152758 175444
rect 152970 175432 152976 175444
rect 153028 175432 153034 175484
rect 173486 175432 173492 175484
rect 173544 175472 173550 175484
rect 200353 175475 200411 175481
rect 200353 175472 200365 175475
rect 173544 175444 200365 175472
rect 173544 175432 173550 175444
rect 200353 175441 200365 175444
rect 200399 175441 200411 175475
rect 221436 175472 221464 175512
rect 232826 175472 232832 175484
rect 221436 175444 232832 175472
rect 200353 175435 200411 175441
rect 232826 175432 232832 175444
rect 232884 175432 232890 175484
rect 79830 175364 79836 175416
rect 79888 175404 79894 175416
rect 117918 175404 117924 175416
rect 79888 175376 117924 175404
rect 79888 175364 79894 175376
rect 117918 175364 117924 175376
rect 117976 175364 117982 175416
rect 173762 175364 173768 175416
rect 173820 175404 173826 175416
rect 214610 175404 214616 175416
rect 173820 175376 214616 175404
rect 173820 175364 173826 175376
rect 214610 175364 214616 175376
rect 214668 175364 214674 175416
rect 215990 175364 215996 175416
rect 216048 175404 216054 175416
rect 224454 175404 224460 175416
rect 216048 175376 224460 175404
rect 216048 175364 216054 175376
rect 224454 175364 224460 175376
rect 224512 175364 224518 175416
rect 79922 175296 79928 175348
rect 79980 175336 79986 175348
rect 123254 175336 123260 175348
rect 79980 175308 123260 175336
rect 79980 175296 79986 175308
rect 123254 175296 123260 175308
rect 123312 175296 123318 175348
rect 173578 175296 173584 175348
rect 173636 175336 173642 175348
rect 217278 175336 217284 175348
rect 173636 175308 217284 175336
rect 173636 175296 173642 175308
rect 217278 175296 217284 175308
rect 217336 175296 217342 175348
rect 80198 175228 80204 175280
rect 80256 175268 80262 175280
rect 126014 175268 126020 175280
rect 80256 175240 126020 175268
rect 80256 175228 80262 175240
rect 126014 175228 126020 175240
rect 126072 175228 126078 175280
rect 176154 175228 176160 175280
rect 176212 175268 176218 175280
rect 220038 175268 220044 175280
rect 176212 175240 220044 175268
rect 176212 175228 176218 175240
rect 220038 175228 220044 175240
rect 220096 175228 220102 175280
rect 221326 175228 221332 175280
rect 221384 175268 221390 175280
rect 264842 175268 264848 175280
rect 221384 175240 264848 175268
rect 221384 175228 221390 175240
rect 264842 175228 264848 175240
rect 264900 175228 264906 175280
rect 80014 175160 80020 175212
rect 80072 175200 80078 175212
rect 128682 175200 128688 175212
rect 80072 175172 128688 175200
rect 80072 175160 80078 175172
rect 128682 175160 128688 175172
rect 128740 175160 128746 175212
rect 174774 175160 174780 175212
rect 174832 175200 174838 175212
rect 222706 175200 222712 175212
rect 174832 175172 222712 175200
rect 174832 175160 174838 175172
rect 222706 175160 222712 175172
rect 222764 175160 222770 175212
rect 65110 175092 65116 175144
rect 65168 175132 65174 175144
rect 65846 175132 65852 175144
rect 65168 175104 65852 175132
rect 65168 175092 65174 175104
rect 65846 175092 65852 175104
rect 65904 175092 65910 175144
rect 80106 175092 80112 175144
rect 80164 175132 80170 175144
rect 120586 175132 120592 175144
rect 80164 175104 120592 175132
rect 80164 175092 80170 175104
rect 120586 175092 120592 175104
rect 120644 175092 120650 175144
rect 121966 175092 121972 175144
rect 122024 175132 122030 175144
rect 170634 175132 170640 175144
rect 122024 175104 170640 175132
rect 122024 175092 122030 175104
rect 170634 175092 170640 175104
rect 170692 175092 170698 175144
rect 190322 175092 190328 175144
rect 190380 175132 190386 175144
rect 199614 175132 199620 175144
rect 190380 175104 199620 175132
rect 190380 175092 190386 175104
rect 199614 175092 199620 175104
rect 199672 175092 199678 175144
rect 202466 175092 202472 175144
rect 202524 175132 202530 175144
rect 264750 175132 264756 175144
rect 202524 175104 264756 175132
rect 202524 175092 202530 175104
rect 264750 175092 264756 175104
rect 264808 175092 264814 175144
rect 92250 175024 92256 175076
rect 92308 175064 92314 175076
rect 97494 175064 97500 175076
rect 92308 175036 97500 175064
rect 92308 175024 92314 175036
rect 97494 175024 97500 175036
rect 97552 175024 97558 175076
rect 105682 175064 105688 175076
rect 99996 175036 105688 175064
rect 93630 174956 93636 175008
rect 93688 174996 93694 175008
rect 98874 174996 98880 175008
rect 93688 174968 98880 174996
rect 93688 174956 93694 174968
rect 98874 174956 98880 174968
rect 98932 174956 98938 175008
rect 89582 174888 89588 174940
rect 89640 174928 89646 174940
rect 95470 174928 95476 174940
rect 89640 174900 95476 174928
rect 89640 174888 89646 174900
rect 95470 174888 95476 174900
rect 95528 174888 95534 174940
rect 96298 174820 96304 174872
rect 96356 174860 96362 174872
rect 99996 174860 100024 175036
rect 105682 175024 105688 175036
rect 105740 175024 105746 175076
rect 256930 175024 256936 175076
rect 256988 175064 256994 175076
rect 257574 175064 257580 175076
rect 256988 175036 257580 175064
rect 256988 175024 256994 175036
rect 257574 175024 257580 175036
rect 257632 175024 257638 175076
rect 96356 174832 100024 174860
rect 96356 174820 96362 174832
rect 186274 174752 186280 174804
rect 186332 174792 186338 174804
rect 191334 174792 191340 174804
rect 186332 174764 191340 174792
rect 186332 174752 186338 174764
rect 191334 174752 191340 174764
rect 191392 174752 191398 174804
rect 187654 174616 187660 174668
rect 187712 174656 187718 174668
rect 192714 174656 192720 174668
rect 187712 174628 192720 174656
rect 187712 174616 187718 174628
rect 192714 174616 192720 174628
rect 192772 174616 192778 174668
rect 97678 174412 97684 174464
rect 97736 174452 97742 174464
rect 98138 174452 98144 174464
rect 97736 174424 98144 174452
rect 97736 174412 97742 174424
rect 98138 174412 98144 174424
rect 98196 174412 98202 174464
rect 98966 174412 98972 174464
rect 99024 174452 99030 174464
rect 99518 174452 99524 174464
rect 99024 174424 99524 174452
rect 99024 174412 99030 174424
rect 99518 174412 99524 174424
rect 99576 174412 99582 174464
rect 100346 174412 100352 174464
rect 100404 174452 100410 174464
rect 100898 174452 100904 174464
rect 100404 174424 100904 174452
rect 100404 174412 100410 174424
rect 100898 174412 100904 174424
rect 100956 174412 100962 174464
rect 101726 174412 101732 174464
rect 101784 174452 101790 174464
rect 102278 174452 102284 174464
rect 101784 174424 102284 174452
rect 101784 174412 101790 174424
rect 102278 174412 102284 174424
rect 102336 174412 102342 174464
rect 103014 174412 103020 174464
rect 103072 174452 103078 174464
rect 103658 174452 103664 174464
rect 103072 174424 103664 174452
rect 103072 174412 103078 174424
rect 103658 174412 103664 174424
rect 103716 174412 103722 174464
rect 104394 174412 104400 174464
rect 104452 174452 104458 174464
rect 105038 174452 105044 174464
rect 104452 174424 105044 174452
rect 104452 174412 104458 174424
rect 105038 174412 105044 174424
rect 105096 174412 105102 174464
rect 105774 174412 105780 174464
rect 105832 174452 105838 174464
rect 106418 174452 106424 174464
rect 105832 174424 106424 174452
rect 105832 174412 105838 174424
rect 106418 174412 106424 174424
rect 106476 174412 106482 174464
rect 107062 174412 107068 174464
rect 107120 174452 107126 174464
rect 107798 174452 107804 174464
rect 107120 174424 107804 174452
rect 107120 174412 107126 174424
rect 107798 174412 107804 174424
rect 107856 174412 107862 174464
rect 116538 174412 116544 174464
rect 116596 174452 116602 174464
rect 117458 174452 117464 174464
rect 116596 174424 117464 174452
rect 116596 174412 116602 174424
rect 117458 174412 117464 174424
rect 117516 174412 117522 174464
rect 119206 174412 119212 174464
rect 119264 174452 119270 174464
rect 120218 174452 120224 174464
rect 119264 174424 120224 174452
rect 119264 174412 119270 174424
rect 120218 174412 120224 174424
rect 120276 174412 120282 174464
rect 124634 174412 124640 174464
rect 124692 174452 124698 174464
rect 125738 174452 125744 174464
rect 124692 174424 125744 174452
rect 124692 174412 124698 174424
rect 125738 174412 125744 174424
rect 125796 174412 125802 174464
rect 134110 174412 134116 174464
rect 134168 174452 134174 174464
rect 134754 174452 134760 174464
rect 134168 174424 134760 174452
rect 134168 174412 134174 174424
rect 134754 174412 134760 174424
rect 134812 174452 134818 174464
rect 171370 174452 171376 174464
rect 134812 174424 171376 174452
rect 134812 174412 134818 174424
rect 171370 174412 171376 174424
rect 171428 174412 171434 174464
rect 183606 174412 183612 174464
rect 183664 174452 183670 174464
rect 189310 174452 189316 174464
rect 183664 174424 189316 174452
rect 183664 174412 183670 174424
rect 189310 174412 189316 174424
rect 189368 174412 189374 174464
rect 197038 174412 197044 174464
rect 197096 174452 197102 174464
rect 197498 174452 197504 174464
rect 197096 174424 197504 174452
rect 197096 174412 197102 174424
rect 197498 174412 197504 174424
rect 197556 174412 197562 174464
rect 198418 174412 198424 174464
rect 198476 174452 198482 174464
rect 198878 174452 198884 174464
rect 198476 174424 198884 174452
rect 198476 174412 198482 174424
rect 198878 174412 198884 174424
rect 198936 174412 198942 174464
rect 199798 174412 199804 174464
rect 199856 174452 199862 174464
rect 200258 174452 200264 174464
rect 199856 174424 200264 174452
rect 199856 174412 199862 174424
rect 200258 174412 200264 174424
rect 200316 174412 200322 174464
rect 201086 174412 201092 174464
rect 201144 174452 201150 174464
rect 201638 174452 201644 174464
rect 201144 174424 201644 174452
rect 201144 174412 201150 174424
rect 201638 174412 201644 174424
rect 201696 174412 201702 174464
rect 205134 174412 205140 174464
rect 205192 174452 205198 174464
rect 205778 174452 205784 174464
rect 205192 174424 205784 174452
rect 205192 174412 205198 174424
rect 205778 174412 205784 174424
rect 205836 174412 205842 174464
rect 210562 174412 210568 174464
rect 210620 174452 210626 174464
rect 211298 174452 211304 174464
rect 210620 174424 211304 174452
rect 210620 174412 210626 174424
rect 211298 174412 211304 174424
rect 211356 174412 211362 174464
rect 243038 173120 243044 173172
rect 243096 173120 243102 173172
rect 151406 173052 151412 173104
rect 151464 173092 151470 173104
rect 152053 173095 152111 173101
rect 151464 173064 152004 173092
rect 151464 173052 151470 173064
rect 60786 172984 60792 173036
rect 60844 173024 60850 173036
rect 64466 173024 64472 173036
rect 60844 172996 64472 173024
rect 60844 172984 60850 172996
rect 64466 172984 64472 172996
rect 64524 172984 64530 173036
rect 65938 172984 65944 173036
rect 65996 173024 66002 173036
rect 68974 173024 68980 173036
rect 65996 172996 68980 173024
rect 65996 172984 66002 172996
rect 68974 172984 68980 172996
rect 69032 172984 69038 173036
rect 69894 172984 69900 173036
rect 69952 173024 69958 173036
rect 71642 173024 71648 173036
rect 69952 172996 71648 173024
rect 69952 172984 69958 172996
rect 71642 172984 71648 172996
rect 71700 172984 71706 173036
rect 144598 172984 144604 173036
rect 144656 173024 144662 173036
rect 144966 173024 144972 173036
rect 144656 172996 144972 173024
rect 144656 172984 144662 172996
rect 144966 172984 144972 172996
rect 145024 172984 145030 173036
rect 145702 172984 145708 173036
rect 145760 173024 145766 173036
rect 146346 173024 146352 173036
rect 145760 172996 146352 173024
rect 145760 172984 145766 172996
rect 146346 172984 146352 172996
rect 146404 172984 146410 173036
rect 148462 172984 148468 173036
rect 148520 173024 148526 173036
rect 149198 173024 149204 173036
rect 148520 172996 149204 173024
rect 148520 172984 148526 172996
rect 149198 172984 149204 172996
rect 149256 172984 149262 173036
rect 151314 172984 151320 173036
rect 151372 173024 151378 173036
rect 151774 173024 151780 173036
rect 151372 172996 151780 173024
rect 151372 172984 151378 172996
rect 151774 172984 151780 172996
rect 151832 172984 151838 173036
rect 151976 173024 152004 173064
rect 152053 173061 152065 173095
rect 152099 173092 152111 173095
rect 153065 173095 153123 173101
rect 153065 173092 153077 173095
rect 152099 173064 153077 173092
rect 152099 173061 152111 173064
rect 152053 173055 152111 173061
rect 153065 173061 153077 173064
rect 153111 173061 153123 173095
rect 243056 173092 243084 173120
rect 153065 173055 153123 173061
rect 242780 173064 243084 173092
rect 161802 173024 161808 173036
rect 151976 172996 161808 173024
rect 161802 172984 161808 172996
rect 161860 172984 161866 173036
rect 162446 172984 162452 173036
rect 162504 173024 162510 173036
rect 163182 173024 163188 173036
rect 162504 172996 163188 173024
rect 162504 172984 162510 172996
rect 163182 172984 163188 172996
rect 163240 172984 163246 173036
rect 163826 172984 163832 173036
rect 163884 173024 163890 173036
rect 164654 173024 164660 173036
rect 163884 172996 164660 173024
rect 163884 172984 163890 172996
rect 164654 172984 164660 172996
rect 164712 172984 164718 173036
rect 231354 172984 231360 173036
rect 231412 173024 231418 173036
rect 236782 173024 236788 173036
rect 231412 172996 236788 173024
rect 231412 172984 231418 172996
rect 236782 172984 236788 172996
rect 236840 172984 236846 173036
rect 236874 172984 236880 173036
rect 236932 173024 236938 173036
rect 238346 173024 238352 173036
rect 236932 172996 238352 173024
rect 236932 172984 236938 172996
rect 238346 172984 238352 172996
rect 238404 172984 238410 173036
rect 242302 172984 242308 173036
rect 242360 173024 242366 173036
rect 242780 173024 242808 173064
rect 242360 172996 242808 173024
rect 242360 172984 242366 172996
rect 242854 172984 242860 173036
rect 242912 173024 242918 173036
rect 243038 173024 243044 173036
rect 242912 172996 243044 173024
rect 242912 172984 242918 172996
rect 243038 172984 243044 172996
rect 243096 172984 243102 173036
rect 246718 172984 246724 173036
rect 246776 173024 246782 173036
rect 247178 173024 247184 173036
rect 246776 172996 247184 173024
rect 246776 172984 246782 172996
rect 247178 172984 247184 172996
rect 247236 172984 247242 173036
rect 248834 172984 248840 173036
rect 248892 173024 248898 173036
rect 249846 173024 249852 173036
rect 248892 172996 249852 173024
rect 248892 172984 248898 172996
rect 249846 172984 249852 172996
rect 249904 172984 249910 173036
rect 250582 172984 250588 173036
rect 250640 173024 250646 173036
rect 251318 173024 251324 173036
rect 250640 172996 251324 173024
rect 250640 172984 250646 172996
rect 251318 172984 251324 172996
rect 251376 172984 251382 173036
rect 252146 172984 252152 173036
rect 252204 173024 252210 173036
rect 252698 173024 252704 173036
rect 252204 172996 252704 173024
rect 252204 172984 252210 172996
rect 252698 172984 252704 172996
rect 252756 172984 252762 173036
rect 253710 172984 253716 173036
rect 253768 173024 253774 173036
rect 254262 173024 254268 173036
rect 253768 172996 254268 173024
rect 253768 172984 253774 172996
rect 254262 172984 254268 172996
rect 254320 172984 254326 173036
rect 59406 172916 59412 172968
rect 59464 172956 59470 172968
rect 63086 172956 63092 172968
rect 59464 172928 63092 172956
rect 59464 172916 59470 172928
rect 63086 172916 63092 172928
rect 63144 172916 63150 172968
rect 143862 172916 143868 172968
rect 143920 172956 143926 172968
rect 145058 172956 145064 172968
rect 143920 172928 145064 172956
rect 143920 172916 143926 172928
rect 145058 172916 145064 172928
rect 145116 172916 145122 172968
rect 152053 172959 152111 172965
rect 152053 172956 152065 172959
rect 151884 172928 152065 172956
rect 58670 172848 58676 172900
rect 58728 172888 58734 172900
rect 62994 172888 63000 172900
rect 58728 172860 63000 172888
rect 58728 172848 58734 172860
rect 62994 172848 63000 172860
rect 63052 172848 63058 172900
rect 150118 172848 150124 172900
rect 150176 172888 150182 172900
rect 151884 172888 151912 172928
rect 152053 172925 152065 172928
rect 152099 172925 152111 172959
rect 152053 172919 152111 172925
rect 162354 172916 162360 172968
rect 162412 172956 162418 172968
rect 163458 172956 163464 172968
rect 162412 172928 163464 172956
rect 162412 172916 162418 172928
rect 163458 172916 163464 172928
rect 163516 172916 163522 172968
rect 163734 172916 163740 172968
rect 163792 172956 163798 172968
rect 165206 172956 165212 172968
rect 163792 172928 165212 172956
rect 163792 172916 163798 172928
rect 165206 172916 165212 172928
rect 165264 172916 165270 172968
rect 235494 172916 235500 172968
rect 235552 172956 235558 172968
rect 237794 172956 237800 172968
rect 235552 172928 237800 172956
rect 235552 172916 235558 172928
rect 237794 172916 237800 172928
rect 237852 172916 237858 172968
rect 245338 172916 245344 172968
rect 245396 172956 245402 172968
rect 253158 172956 253164 172968
rect 245396 172928 253164 172956
rect 245396 172916 245402 172928
rect 253158 172916 253164 172928
rect 253216 172916 253222 172968
rect 253526 172916 253532 172968
rect 253584 172956 253590 172968
rect 254814 172956 254820 172968
rect 253584 172928 254820 172956
rect 253584 172916 253590 172928
rect 254814 172916 254820 172928
rect 254872 172916 254878 172968
rect 150176 172860 151912 172888
rect 151961 172891 152019 172897
rect 150176 172848 150182 172860
rect 151961 172857 151973 172891
rect 152007 172888 152019 172891
rect 152329 172891 152387 172897
rect 152329 172888 152341 172891
rect 152007 172860 152341 172888
rect 152007 172857 152019 172860
rect 151961 172851 152019 172857
rect 152329 172857 152341 172860
rect 152375 172857 152387 172891
rect 152329 172851 152387 172857
rect 152418 172848 152424 172900
rect 152476 172888 152482 172900
rect 152970 172888 152976 172900
rect 152476 172860 152976 172888
rect 152476 172848 152482 172860
rect 152970 172848 152976 172860
rect 153028 172848 153034 172900
rect 153065 172891 153123 172897
rect 153065 172857 153077 172891
rect 153111 172888 153123 172891
rect 156745 172891 156803 172897
rect 156745 172888 156757 172891
rect 153111 172860 156757 172888
rect 153111 172857 153123 172860
rect 153065 172851 153123 172857
rect 156745 172857 156757 172860
rect 156791 172857 156803 172891
rect 156745 172851 156803 172857
rect 156834 172848 156840 172900
rect 156892 172888 156898 172900
rect 161250 172888 161256 172900
rect 156892 172860 161256 172888
rect 156892 172848 156898 172860
rect 161250 172848 161256 172860
rect 161308 172848 161314 172900
rect 161345 172891 161403 172897
rect 161345 172857 161357 172891
rect 161391 172888 161403 172891
rect 161894 172888 161900 172900
rect 161391 172860 161900 172888
rect 161391 172857 161403 172860
rect 161345 172851 161403 172857
rect 161894 172848 161900 172860
rect 161952 172848 161958 172900
rect 234206 172848 234212 172900
rect 234264 172888 234270 172900
rect 237242 172888 237248 172900
rect 234264 172860 237248 172888
rect 234264 172848 234270 172860
rect 237242 172848 237248 172860
rect 237300 172848 237306 172900
rect 245430 172848 245436 172900
rect 245488 172888 245494 172900
rect 245488 172860 252928 172888
rect 245488 172848 245494 172860
rect 60510 172780 60516 172832
rect 60568 172820 60574 172832
rect 68238 172820 68244 172832
rect 60568 172792 68244 172820
rect 60568 172780 60574 172792
rect 68238 172780 68244 172792
rect 68296 172780 68302 172832
rect 150578 172780 150584 172832
rect 150636 172820 150642 172832
rect 162262 172820 162268 172832
rect 150636 172792 162268 172820
rect 150636 172780 150642 172792
rect 162262 172780 162268 172792
rect 162320 172780 162326 172832
rect 245246 172780 245252 172832
rect 245304 172820 245310 172832
rect 252790 172820 252796 172832
rect 245304 172792 252796 172820
rect 245304 172780 245310 172792
rect 252790 172780 252796 172792
rect 252848 172780 252854 172832
rect 252900 172820 252928 172860
rect 253434 172848 253440 172900
rect 253492 172888 253498 172900
rect 255550 172888 255556 172900
rect 253492 172860 255556 172888
rect 253492 172848 253498 172860
rect 255550 172848 255556 172860
rect 255608 172848 255614 172900
rect 253802 172820 253808 172832
rect 252900 172792 253808 172820
rect 253802 172780 253808 172792
rect 253860 172780 253866 172832
rect 57290 172712 57296 172764
rect 57348 172752 57354 172764
rect 67410 172752 67416 172764
rect 57348 172724 67416 172752
rect 57348 172712 57354 172724
rect 67410 172712 67416 172724
rect 67468 172712 67474 172764
rect 151682 172712 151688 172764
rect 151740 172752 151746 172764
rect 153249 172755 153307 172761
rect 153249 172752 153261 172755
rect 151740 172724 153261 172752
rect 151740 172712 151746 172724
rect 153249 172721 153261 172724
rect 153295 172721 153307 172755
rect 153249 172715 153307 172721
rect 153338 172712 153344 172764
rect 153396 172752 153402 172764
rect 157018 172752 157024 172764
rect 153396 172724 157024 172752
rect 153396 172712 153402 172724
rect 157018 172712 157024 172724
rect 157076 172712 157082 172764
rect 248374 172712 248380 172764
rect 248432 172752 248438 172764
rect 255918 172752 255924 172764
rect 248432 172724 255924 172752
rect 248432 172712 248438 172724
rect 255918 172712 255924 172724
rect 255976 172712 255982 172764
rect 58026 172644 58032 172696
rect 58084 172684 58090 172696
rect 67870 172684 67876 172696
rect 58084 172656 67876 172684
rect 58084 172644 58090 172656
rect 67870 172644 67876 172656
rect 67928 172644 67934 172696
rect 138066 172644 138072 172696
rect 138124 172684 138130 172696
rect 154810 172684 154816 172696
rect 138124 172656 154816 172684
rect 138124 172644 138130 172656
rect 154810 172644 154816 172656
rect 154868 172644 154874 172696
rect 156745 172687 156803 172693
rect 156745 172653 156757 172687
rect 156791 172684 156803 172687
rect 161345 172687 161403 172693
rect 161345 172684 161357 172687
rect 156791 172656 161357 172684
rect 156791 172653 156803 172656
rect 156745 172647 156803 172653
rect 161345 172653 161357 172656
rect 161391 172653 161403 172687
rect 161345 172647 161403 172653
rect 248558 172644 248564 172696
rect 248616 172684 248622 172696
rect 256286 172684 256292 172696
rect 248616 172656 256292 172684
rect 248616 172644 248622 172656
rect 256286 172644 256292 172656
rect 256344 172644 256350 172696
rect 54622 172576 54628 172628
rect 54680 172616 54686 172628
rect 65570 172616 65576 172628
rect 54680 172588 65576 172616
rect 54680 172576 54686 172588
rect 65570 172576 65576 172588
rect 65628 172576 65634 172628
rect 138158 172576 138164 172628
rect 138216 172616 138222 172628
rect 154166 172616 154172 172628
rect 138216 172588 154172 172616
rect 138216 172576 138222 172588
rect 154166 172576 154172 172588
rect 154224 172576 154230 172628
rect 156098 172576 156104 172628
rect 156156 172616 156162 172628
rect 167414 172616 167420 172628
rect 156156 172588 167420 172616
rect 156156 172576 156162 172588
rect 167414 172576 167420 172588
rect 167472 172576 167478 172628
rect 245062 172576 245068 172628
rect 245120 172616 245126 172628
rect 245798 172616 245804 172628
rect 245120 172588 245804 172616
rect 245120 172576 245126 172588
rect 245798 172576 245804 172588
rect 245856 172576 245862 172628
rect 249570 172576 249576 172628
rect 249628 172616 249634 172628
rect 258310 172616 258316 172628
rect 249628 172588 258316 172616
rect 249628 172576 249634 172588
rect 258310 172576 258316 172588
rect 258368 172576 258374 172628
rect 50482 172508 50488 172560
rect 50540 172548 50546 172560
rect 51218 172548 51224 172560
rect 50540 172520 51224 172548
rect 50540 172508 50546 172520
rect 51218 172508 51224 172520
rect 51276 172508 51282 172560
rect 61982 172508 61988 172560
rect 62040 172548 62046 172560
rect 74402 172548 74408 172560
rect 62040 172520 74408 172548
rect 62040 172508 62046 172520
rect 74402 172508 74408 172520
rect 74460 172508 74466 172560
rect 137882 172508 137888 172560
rect 137940 172548 137946 172560
rect 155638 172548 155644 172560
rect 137940 172520 155644 172548
rect 137940 172508 137946 172520
rect 155638 172508 155644 172520
rect 155696 172508 155702 172560
rect 155822 172508 155828 172560
rect 155880 172548 155886 172560
rect 167966 172548 167972 172560
rect 155880 172520 167972 172548
rect 155880 172508 155886 172520
rect 167966 172508 167972 172520
rect 168024 172508 168030 172560
rect 250766 172508 250772 172560
rect 250824 172548 250830 172560
rect 260334 172548 260340 172560
rect 250824 172520 260340 172548
rect 250824 172508 250830 172520
rect 260334 172508 260340 172520
rect 260392 172508 260398 172560
rect 137790 172440 137796 172492
rect 137848 172480 137854 172492
rect 156190 172480 156196 172492
rect 137848 172452 156196 172480
rect 137848 172440 137854 172452
rect 156190 172440 156196 172452
rect 156248 172440 156254 172492
rect 157478 172440 157484 172492
rect 157536 172480 157542 172492
rect 168610 172480 168616 172492
rect 157536 172452 168616 172480
rect 157536 172440 157542 172452
rect 168610 172440 168616 172452
rect 168668 172440 168674 172492
rect 241566 172440 241572 172492
rect 241624 172480 241630 172492
rect 242394 172480 242400 172492
rect 241624 172452 242400 172480
rect 241624 172440 241630 172452
rect 242394 172440 242400 172452
rect 242452 172440 242458 172492
rect 249386 172440 249392 172492
rect 249444 172480 249450 172492
rect 258678 172480 258684 172492
rect 249444 172452 258684 172480
rect 249444 172440 249450 172452
rect 258678 172440 258684 172452
rect 258736 172440 258742 172492
rect 61798 172372 61804 172424
rect 61856 172412 61862 172424
rect 73666 172412 73672 172424
rect 61856 172384 73672 172412
rect 61856 172372 61862 172384
rect 73666 172372 73672 172384
rect 73724 172372 73730 172424
rect 137974 172372 137980 172424
rect 138032 172412 138038 172424
rect 155086 172412 155092 172424
rect 138032 172384 155092 172412
rect 138032 172372 138038 172384
rect 155086 172372 155092 172384
rect 155144 172372 155150 172424
rect 155730 172372 155736 172424
rect 155788 172412 155794 172424
rect 167230 172412 167236 172424
rect 155788 172384 167236 172412
rect 155788 172372 155794 172384
rect 167230 172372 167236 172384
rect 167288 172372 167294 172424
rect 250674 172372 250680 172424
rect 250732 172412 250738 172424
rect 259782 172412 259788 172424
rect 250732 172384 259788 172412
rect 250732 172372 250738 172384
rect 259782 172372 259788 172384
rect 259840 172372 259846 172424
rect 38154 172304 38160 172356
rect 38212 172344 38218 172356
rect 49194 172344 49200 172356
rect 38212 172316 49200 172344
rect 38212 172304 38218 172316
rect 49194 172304 49200 172316
rect 49252 172304 49258 172356
rect 63638 172304 63644 172356
rect 63696 172344 63702 172356
rect 76426 172344 76432 172356
rect 63696 172316 76432 172344
rect 63696 172304 63702 172316
rect 76426 172304 76432 172316
rect 76484 172304 76490 172356
rect 137606 172304 137612 172356
rect 137664 172344 137670 172356
rect 156834 172344 156840 172356
rect 137664 172316 156840 172344
rect 137664 172304 137670 172316
rect 156834 172304 156840 172316
rect 156892 172304 156898 172356
rect 157386 172304 157392 172356
rect 157444 172344 157450 172356
rect 169070 172344 169076 172356
rect 157444 172316 169076 172344
rect 157444 172304 157450 172316
rect 169070 172304 169076 172316
rect 169128 172304 169134 172356
rect 249202 172304 249208 172356
rect 249260 172344 249266 172356
rect 255918 172344 255924 172356
rect 249260 172316 255924 172344
rect 249260 172304 249266 172316
rect 255918 172304 255924 172316
rect 255976 172304 255982 172356
rect 256013 172347 256071 172353
rect 256013 172313 256025 172347
rect 256059 172344 256071 172347
rect 259230 172344 259236 172356
rect 256059 172316 259236 172344
rect 256059 172313 256071 172316
rect 256013 172307 256071 172313
rect 259230 172304 259236 172316
rect 259288 172304 259294 172356
rect 60326 172236 60332 172288
rect 60384 172276 60390 172288
rect 60384 172248 63776 172276
rect 60384 172236 60390 172248
rect 60234 172168 60240 172220
rect 60292 172208 60298 172220
rect 63638 172208 63644 172220
rect 60292 172180 63644 172208
rect 60292 172168 60298 172180
rect 63638 172168 63644 172180
rect 63696 172168 63702 172220
rect 63748 172208 63776 172248
rect 65110 172236 65116 172288
rect 65168 172276 65174 172288
rect 66214 172276 66220 172288
rect 65168 172248 66220 172276
rect 65168 172236 65174 172248
rect 66214 172236 66220 172248
rect 66272 172236 66278 172288
rect 151866 172236 151872 172288
rect 151924 172276 151930 172288
rect 162538 172276 162544 172288
rect 151924 172248 162544 172276
rect 151924 172236 151930 172248
rect 162538 172236 162544 172248
rect 162596 172236 162602 172288
rect 67594 172208 67600 172220
rect 63748 172180 67600 172208
rect 67594 172168 67600 172180
rect 67652 172168 67658 172220
rect 149014 172168 149020 172220
rect 149072 172208 149078 172220
rect 151961 172211 152019 172217
rect 151961 172208 151973 172211
rect 149072 172180 151973 172208
rect 149072 172168 149078 172180
rect 151961 172177 151973 172180
rect 152007 172177 152019 172211
rect 151961 172171 152019 172177
rect 154074 172168 154080 172220
rect 154132 172208 154138 172220
rect 158214 172208 158220 172220
rect 154132 172180 158220 172208
rect 154132 172168 154138 172180
rect 158214 172168 158220 172180
rect 158272 172168 158278 172220
rect 248926 172168 248932 172220
rect 248984 172208 248990 172220
rect 256470 172208 256476 172220
rect 248984 172180 256476 172208
rect 248984 172168 248990 172180
rect 256470 172168 256476 172180
rect 256528 172168 256534 172220
rect 65110 172140 65116 172152
rect 60252 172112 65116 172140
rect 55266 172032 55272 172084
rect 55324 172072 55330 172084
rect 60252 172072 60280 172112
rect 65110 172100 65116 172112
rect 65168 172100 65174 172152
rect 153249 172143 153307 172149
rect 153249 172109 153261 172143
rect 153295 172140 153307 172143
rect 160698 172140 160704 172152
rect 153295 172112 160704 172140
rect 153295 172109 153307 172112
rect 153249 172103 153307 172109
rect 160698 172100 160704 172112
rect 160756 172100 160762 172152
rect 245154 172100 245160 172152
rect 245212 172140 245218 172152
rect 252238 172140 252244 172152
rect 245212 172112 252244 172140
rect 245212 172100 245218 172112
rect 252238 172100 252244 172112
rect 252296 172100 252302 172152
rect 55324 172044 60280 172072
rect 55324 172032 55330 172044
rect 60602 172032 60608 172084
rect 60660 172072 60666 172084
rect 66858 172072 66864 172084
rect 60660 172044 66864 172072
rect 60660 172032 60666 172044
rect 66858 172032 66864 172044
rect 66916 172032 66922 172084
rect 152878 172032 152884 172084
rect 152936 172072 152942 172084
rect 159042 172072 159048 172084
rect 152936 172044 159048 172072
rect 152936 172032 152942 172044
rect 159042 172032 159048 172044
rect 159100 172032 159106 172084
rect 247822 172032 247828 172084
rect 247880 172072 247886 172084
rect 253618 172072 253624 172084
rect 247880 172044 253624 172072
rect 247880 172032 247886 172044
rect 253618 172032 253624 172044
rect 253676 172032 253682 172084
rect 56002 171964 56008 172016
rect 56060 172004 56066 172016
rect 60418 172004 60424 172016
rect 56060 171976 60424 172004
rect 56060 171964 56066 171976
rect 60418 171964 60424 171976
rect 60476 171964 60482 172016
rect 152329 172007 152387 172013
rect 152329 171973 152341 172007
rect 152375 172004 152387 172007
rect 161066 172004 161072 172016
rect 152375 171976 161072 172004
rect 152375 171973 152387 171976
rect 152329 171967 152387 171973
rect 161066 171964 161072 171976
rect 161124 171964 161130 172016
rect 232734 171964 232740 172016
rect 232792 172004 232798 172016
rect 239266 172004 239272 172016
rect 232792 171976 239272 172004
rect 232792 171964 232798 171976
rect 239266 171964 239272 171976
rect 239324 171964 239330 172016
rect 247086 171964 247092 172016
rect 247144 172004 247150 172016
rect 252054 172004 252060 172016
rect 247144 171976 252060 172004
rect 247144 171964 247150 171976
rect 252054 171964 252060 171976
rect 252112 171964 252118 172016
rect 146530 171896 146536 171948
rect 146588 171936 146594 171948
rect 147726 171936 147732 171948
rect 146588 171908 147732 171936
rect 146588 171896 146594 171908
rect 147726 171896 147732 171908
rect 147784 171896 147790 171948
rect 152786 171896 152792 171948
rect 152844 171936 152850 171948
rect 158490 171936 158496 171948
rect 152844 171908 158496 171936
rect 152844 171896 152850 171908
rect 158490 171896 158496 171908
rect 158548 171896 158554 171948
rect 234114 171896 234120 171948
rect 234172 171936 234178 171948
rect 240554 171936 240560 171948
rect 234172 171908 240560 171936
rect 234172 171896 234178 171908
rect 240554 171896 240560 171908
rect 240612 171896 240618 171948
rect 245614 171896 245620 171948
rect 245672 171936 245678 171948
rect 250858 171936 250864 171948
rect 245672 171908 250864 171936
rect 245672 171896 245678 171908
rect 250858 171896 250864 171908
rect 250916 171896 250922 171948
rect 152694 171828 152700 171880
rect 152752 171868 152758 171880
rect 160330 171868 160336 171880
rect 152752 171840 160336 171868
rect 152752 171828 152758 171840
rect 160330 171828 160336 171840
rect 160388 171828 160394 171880
rect 243958 171828 243964 171880
rect 244016 171868 244022 171880
rect 249662 171868 249668 171880
rect 244016 171840 249668 171868
rect 244016 171828 244022 171840
rect 249662 171828 249668 171840
rect 249720 171828 249726 171880
rect 56646 171760 56652 171812
rect 56704 171800 56710 171812
rect 60050 171800 60056 171812
rect 56704 171772 60056 171800
rect 56704 171760 56710 171772
rect 60050 171760 60056 171772
rect 60108 171760 60114 171812
rect 152602 171760 152608 171812
rect 152660 171800 152666 171812
rect 159594 171800 159600 171812
rect 152660 171772 159600 171800
rect 152660 171760 152666 171772
rect 159594 171760 159600 171772
rect 159652 171760 159658 171812
rect 244418 171760 244424 171812
rect 244476 171800 244482 171812
rect 249294 171800 249300 171812
rect 244476 171772 249300 171800
rect 244476 171760 244482 171772
rect 249294 171760 249300 171772
rect 249352 171760 249358 171812
rect 53242 171692 53248 171744
rect 53300 171732 53306 171744
rect 57566 171732 57572 171744
rect 53300 171704 57572 171732
rect 53300 171692 53306 171704
rect 57566 171692 57572 171704
rect 57624 171692 57630 171744
rect 64374 171732 64380 171744
rect 60068 171704 64380 171732
rect 60068 171676 60096 171704
rect 64374 171692 64380 171704
rect 64432 171692 64438 171744
rect 149566 171692 149572 171744
rect 149624 171732 149630 171744
rect 161434 171732 161440 171744
rect 149624 171704 161440 171732
rect 149624 171692 149630 171704
rect 161434 171692 161440 171704
rect 161492 171692 161498 171744
rect 238254 171692 238260 171744
rect 238312 171732 238318 171744
rect 238990 171732 238996 171744
rect 238312 171704 238996 171732
rect 238312 171692 238318 171704
rect 238990 171692 238996 171704
rect 239048 171692 239054 171744
rect 249018 171692 249024 171744
rect 249076 171732 249082 171744
rect 256013 171735 256071 171741
rect 256013 171732 256025 171735
rect 249076 171704 256025 171732
rect 249076 171692 249082 171704
rect 256013 171701 256025 171704
rect 256059 171701 256071 171735
rect 256013 171695 256071 171701
rect 60050 171624 60056 171676
rect 60108 171624 60114 171676
rect 120218 170196 120224 170248
rect 120276 170236 120282 170248
rect 170726 170236 170732 170248
rect 120276 170208 170732 170236
rect 120276 170196 120282 170208
rect 170726 170196 170732 170208
rect 170784 170196 170790 170248
rect 211298 170196 211304 170248
rect 211356 170236 211362 170248
rect 233470 170236 233476 170248
rect 211356 170208 233476 170236
rect 211356 170196 211362 170208
rect 233470 170196 233476 170208
rect 233528 170196 233534 170248
rect 125738 170128 125744 170180
rect 125796 170168 125802 170180
rect 139630 170168 139636 170180
rect 125796 170140 139636 170168
rect 125796 170128 125802 170140
rect 139630 170128 139636 170140
rect 139688 170128 139694 170180
rect 239358 169992 239364 170044
rect 239416 170032 239422 170044
rect 240002 170032 240008 170044
rect 239416 170004 240008 170032
rect 239416 169992 239422 170004
rect 240002 169992 240008 170004
rect 240060 169992 240066 170044
rect 117458 168836 117464 168888
rect 117516 168876 117522 168888
rect 139630 168876 139636 168888
rect 117516 168848 139636 168876
rect 117516 168836 117522 168848
rect 139630 168836 139636 168848
rect 139688 168836 139694 168888
rect 205778 168836 205784 168888
rect 205836 168876 205842 168888
rect 233470 168876 233476 168888
rect 205836 168848 233476 168876
rect 205836 168836 205842 168848
rect 233470 168836 233476 168848
rect 233528 168836 233534 168888
rect 236690 168836 236696 168888
rect 236748 168876 236754 168888
rect 292626 168876 292632 168888
rect 236748 168848 292632 168876
rect 236748 168836 236754 168848
rect 292626 168836 292632 168848
rect 292684 168836 292690 168888
rect 228686 168156 228692 168208
rect 228744 168196 228750 168208
rect 228870 168196 228876 168208
rect 228744 168168 228876 168196
rect 228744 168156 228750 168168
rect 228870 168156 228876 168168
rect 228928 168156 228934 168208
rect 174038 167816 174044 167868
rect 174096 167856 174102 167868
rect 177534 167856 177540 167868
rect 174096 167828 177540 167856
rect 174096 167816 174102 167828
rect 177534 167816 177540 167828
rect 177592 167816 177598 167868
rect 173302 167680 173308 167732
rect 173360 167720 173366 167732
rect 180294 167720 180300 167732
rect 173360 167692 180300 167720
rect 173360 167680 173366 167692
rect 180294 167680 180300 167692
rect 180352 167680 180358 167732
rect 265854 167544 265860 167596
rect 265912 167584 265918 167596
rect 300170 167584 300176 167596
rect 265912 167556 300176 167584
rect 265912 167544 265918 167556
rect 300170 167544 300176 167556
rect 300228 167544 300234 167596
rect 98138 167272 98144 167324
rect 98196 167312 98202 167324
rect 109454 167312 109460 167324
rect 98196 167284 109460 167312
rect 98196 167272 98202 167284
rect 109454 167272 109460 167284
rect 109512 167272 109518 167324
rect 191978 167272 191984 167324
rect 192036 167312 192042 167324
rect 203754 167312 203760 167324
rect 192036 167284 203760 167312
rect 192036 167272 192042 167284
rect 203754 167272 203760 167284
rect 203812 167272 203818 167324
rect 100898 167204 100904 167256
rect 100956 167244 100962 167256
rect 114146 167244 114152 167256
rect 100956 167216 114152 167244
rect 100956 167204 100962 167216
rect 114146 167204 114152 167216
rect 114204 167204 114210 167256
rect 194738 167204 194744 167256
rect 194796 167244 194802 167256
rect 208446 167244 208452 167256
rect 194796 167216 208452 167244
rect 194796 167204 194802 167216
rect 208446 167204 208452 167216
rect 208504 167204 208510 167256
rect 99518 167136 99524 167188
rect 99576 167176 99582 167188
rect 112030 167176 112036 167188
rect 99576 167148 112036 167176
rect 99576 167136 99582 167148
rect 112030 167136 112036 167148
rect 112088 167136 112094 167188
rect 193358 167136 193364 167188
rect 193416 167176 193422 167188
rect 206146 167176 206152 167188
rect 193416 167148 206152 167176
rect 193416 167136 193422 167148
rect 206146 167136 206152 167148
rect 206204 167136 206210 167188
rect 102278 167068 102284 167120
rect 102336 167108 102342 167120
rect 116538 167108 116544 167120
rect 102336 167080 116544 167108
rect 102336 167068 102342 167080
rect 116538 167068 116544 167080
rect 116596 167068 116602 167120
rect 196118 167068 196124 167120
rect 196176 167108 196182 167120
rect 210838 167108 210844 167120
rect 196176 167080 210844 167108
rect 196176 167068 196182 167080
rect 210838 167068 210844 167080
rect 210896 167068 210902 167120
rect 105038 167000 105044 167052
rect 105096 167040 105102 167052
rect 121230 167040 121236 167052
rect 105096 167012 121236 167040
rect 105096 167000 105102 167012
rect 121230 167000 121236 167012
rect 121288 167000 121294 167052
rect 197498 167000 197504 167052
rect 197556 167040 197562 167052
rect 213230 167040 213236 167052
rect 197556 167012 213236 167040
rect 197556 167000 197562 167012
rect 213230 167000 213236 167012
rect 213288 167000 213294 167052
rect 103658 166932 103664 166984
rect 103716 166972 103722 166984
rect 118930 166972 118936 166984
rect 103716 166944 118936 166972
rect 103716 166932 103722 166944
rect 118930 166932 118936 166944
rect 118988 166932 118994 166984
rect 184986 166932 184992 166984
rect 185044 166972 185050 166984
rect 191978 166972 191984 166984
rect 185044 166944 191984 166972
rect 185044 166932 185050 166944
rect 191978 166932 191984 166944
rect 192036 166932 192042 166984
rect 198878 166932 198884 166984
rect 198936 166972 198942 166984
rect 215530 166972 215536 166984
rect 198936 166944 215536 166972
rect 198936 166932 198942 166944
rect 215530 166932 215536 166944
rect 215588 166932 215594 166984
rect 106418 166864 106424 166916
rect 106476 166904 106482 166916
rect 123622 166904 123628 166916
rect 106476 166876 123628 166904
rect 106476 166864 106482 166876
rect 123622 166864 123628 166876
rect 123680 166864 123686 166916
rect 182226 166864 182232 166916
rect 182284 166904 182290 166916
rect 187286 166904 187292 166916
rect 182284 166876 187292 166904
rect 182284 166864 182290 166876
rect 187286 166864 187292 166876
rect 187344 166864 187350 166916
rect 200258 166864 200264 166916
rect 200316 166904 200322 166916
rect 217922 166904 217928 166916
rect 200316 166876 217928 166904
rect 200316 166864 200322 166876
rect 217922 166864 217928 166876
rect 217980 166864 217986 166916
rect 87098 166796 87104 166848
rect 87156 166836 87162 166848
rect 90686 166836 90692 166848
rect 87156 166808 90692 166836
rect 87156 166796 87162 166808
rect 90686 166796 90692 166808
rect 90744 166796 90750 166848
rect 91238 166796 91244 166848
rect 91296 166836 91302 166848
rect 97678 166836 97684 166848
rect 91296 166808 97684 166836
rect 91296 166796 91302 166808
rect 97678 166796 97684 166808
rect 97736 166796 97742 166848
rect 98874 166796 98880 166848
rect 98932 166836 98938 166848
rect 102370 166836 102376 166848
rect 98932 166808 102376 166836
rect 98932 166796 98938 166808
rect 102370 166796 102376 166808
rect 102428 166796 102434 166848
rect 104394 166796 104400 166848
rect 104452 166836 104458 166848
rect 105130 166836 105136 166848
rect 104452 166808 105136 166836
rect 104452 166796 104458 166808
rect 105130 166796 105136 166808
rect 105188 166796 105194 166848
rect 107798 166796 107804 166848
rect 107856 166836 107862 166848
rect 125922 166836 125928 166848
rect 107856 166808 125928 166836
rect 107856 166796 107862 166808
rect 125922 166796 125928 166808
rect 125980 166796 125986 166848
rect 180846 166796 180852 166848
rect 180904 166836 180910 166848
rect 184986 166836 184992 166848
rect 180904 166808 184992 166836
rect 180904 166796 180910 166808
rect 184986 166796 184992 166808
rect 185044 166796 185050 166848
rect 198234 166796 198240 166848
rect 198292 166836 198298 166848
rect 199062 166836 199068 166848
rect 198292 166808 199068 166836
rect 198292 166796 198298 166808
rect 199062 166796 199068 166808
rect 199120 166796 199126 166848
rect 201638 166796 201644 166848
rect 201696 166836 201702 166848
rect 220222 166836 220228 166848
rect 201696 166808 220228 166836
rect 201696 166796 201702 166808
rect 220222 166796 220228 166808
rect 220280 166796 220286 166848
rect 192714 166660 192720 166712
rect 192772 166700 192778 166712
rect 196670 166700 196676 166712
rect 192772 166672 196676 166700
rect 192772 166660 192778 166672
rect 196670 166660 196676 166672
rect 196728 166660 196734 166712
rect 199614 166660 199620 166712
rect 199672 166700 199678 166712
rect 201454 166700 201460 166712
rect 199672 166672 201460 166700
rect 199672 166660 199678 166672
rect 201454 166660 201460 166672
rect 201512 166660 201518 166712
rect 97494 166592 97500 166644
rect 97552 166632 97558 166644
rect 100070 166632 100076 166644
rect 97552 166604 100076 166632
rect 97552 166592 97558 166604
rect 100070 166592 100076 166604
rect 100128 166592 100134 166644
rect 173118 166592 173124 166644
rect 173176 166632 173182 166644
rect 178914 166632 178920 166644
rect 173176 166604 178920 166632
rect 173176 166592 173182 166604
rect 178914 166592 178920 166604
rect 178972 166592 178978 166644
rect 191334 166524 191340 166576
rect 191392 166564 191398 166576
rect 194370 166564 194376 166576
rect 191392 166536 194376 166564
rect 191392 166524 191398 166536
rect 194370 166524 194376 166536
rect 194428 166524 194434 166576
rect 231814 166524 231820 166576
rect 231872 166564 231878 166576
rect 233470 166564 233476 166576
rect 231872 166536 233476 166564
rect 231872 166524 231878 166536
rect 233470 166524 233476 166536
rect 233528 166524 233534 166576
rect 88478 166456 88484 166508
rect 88536 166496 88542 166508
rect 92986 166496 92992 166508
rect 88536 166468 92992 166496
rect 88536 166456 88542 166468
rect 92986 166456 92992 166468
rect 93044 166456 93050 166508
rect 105774 166456 105780 166508
rect 105832 166496 105838 166508
rect 107154 166496 107160 166508
rect 105832 166468 107160 166496
rect 105832 166456 105838 166468
rect 107154 166456 107160 166468
rect 107212 166456 107218 166508
rect 135030 166252 135036 166304
rect 135088 166292 135094 166304
rect 139722 166292 139728 166304
rect 135088 166264 139728 166292
rect 135088 166252 135094 166264
rect 139722 166252 139728 166264
rect 139780 166252 139786 166304
rect 76702 166184 76708 166236
rect 76760 166224 76766 166236
rect 128682 166224 128688 166236
rect 76760 166196 128688 166224
rect 76760 166184 76766 166196
rect 128682 166184 128688 166196
rect 128740 166184 128746 166236
rect 132086 166184 132092 166236
rect 132144 166224 132150 166236
rect 139630 166224 139636 166236
rect 132144 166196 139636 166224
rect 132144 166184 132150 166196
rect 139630 166184 139636 166196
rect 139688 166184 139694 166236
rect 170726 166184 170732 166236
rect 170784 166224 170790 166236
rect 222614 166224 222620 166236
rect 170784 166196 222620 166224
rect 170784 166184 170790 166196
rect 222614 166184 222620 166196
rect 222672 166184 222678 166236
rect 230894 166184 230900 166236
rect 230952 166224 230958 166236
rect 233470 166224 233476 166236
rect 230952 166196 233476 166224
rect 230952 166184 230958 166196
rect 233470 166184 233476 166196
rect 233528 166184 233534 166236
rect 80198 164756 80204 164808
rect 80256 164796 80262 164808
rect 80256 164768 85396 164796
rect 80256 164756 80262 164768
rect 85368 164728 85396 164768
rect 174038 164756 174044 164808
rect 174096 164796 174102 164808
rect 181582 164796 181588 164808
rect 174096 164768 181588 164796
rect 174096 164756 174102 164768
rect 181582 164756 181588 164768
rect 181640 164756 181646 164808
rect 87190 164728 87196 164740
rect 85368 164700 87196 164728
rect 87190 164688 87196 164700
rect 87248 164688 87254 164740
rect 225926 164688 225932 164740
rect 225984 164728 225990 164740
rect 233654 164728 233660 164740
rect 225984 164700 233660 164728
rect 225984 164688 225990 164700
rect 233654 164688 233660 164700
rect 233712 164688 233718 164740
rect 80198 163872 80204 163924
rect 80256 163912 80262 163924
rect 85442 163912 85448 163924
rect 80256 163884 85448 163912
rect 80256 163872 80262 163884
rect 85442 163872 85448 163884
rect 85500 163872 85506 163924
rect 131902 163532 131908 163584
rect 131960 163572 131966 163584
rect 140550 163572 140556 163584
rect 131960 163544 140556 163572
rect 131960 163532 131966 163544
rect 140550 163532 140556 163544
rect 140608 163532 140614 163584
rect 177902 163532 177908 163584
rect 177960 163572 177966 163584
rect 181766 163572 181772 163584
rect 177960 163544 181772 163572
rect 177960 163532 177966 163544
rect 181766 163532 181772 163544
rect 181824 163532 181830 163584
rect 80198 163464 80204 163516
rect 80256 163504 80262 163516
rect 80256 163476 84384 163504
rect 80256 163464 80262 163476
rect 84356 163368 84384 163476
rect 132270 163464 132276 163516
rect 132328 163504 132334 163516
rect 140642 163504 140648 163516
rect 132328 163476 140648 163504
rect 132328 163464 132334 163476
rect 140642 163464 140648 163476
rect 140700 163464 140706 163516
rect 132362 163396 132368 163448
rect 132420 163436 132426 163448
rect 140366 163436 140372 163448
rect 132420 163408 140372 163436
rect 132420 163396 132426 163408
rect 140366 163396 140372 163408
rect 140424 163396 140430 163448
rect 174038 163396 174044 163448
rect 174096 163436 174102 163448
rect 181766 163436 181772 163448
rect 174096 163408 181772 163436
rect 174096 163396 174102 163408
rect 181766 163396 181772 163408
rect 181824 163396 181830 163448
rect 87190 163368 87196 163380
rect 84356 163340 87196 163368
rect 87190 163328 87196 163340
rect 87248 163328 87254 163380
rect 226386 163328 226392 163380
rect 226444 163368 226450 163380
rect 231814 163368 231820 163380
rect 226444 163340 231820 163368
rect 226444 163328 226450 163340
rect 231814 163328 231820 163340
rect 231872 163328 231878 163380
rect 85442 163260 85448 163312
rect 85500 163300 85506 163312
rect 87282 163300 87288 163312
rect 85500 163272 87288 163300
rect 85500 163260 85506 163272
rect 87282 163260 87288 163272
rect 87340 163260 87346 163312
rect 226478 163260 226484 163312
rect 226536 163300 226542 163312
rect 230894 163300 230900 163312
rect 226536 163272 230900 163300
rect 226536 163260 226542 163272
rect 230894 163260 230900 163272
rect 230952 163260 230958 163312
rect 225558 163192 225564 163244
rect 225616 163232 225622 163244
rect 233562 163232 233568 163244
rect 225616 163204 233568 163232
rect 225616 163192 225622 163204
rect 233562 163192 233568 163204
rect 233620 163192 233626 163244
rect 225926 162988 225932 163040
rect 225984 163028 225990 163040
rect 233470 163028 233476 163040
rect 225984 163000 233476 163028
rect 225984 162988 225990 163000
rect 233470 162988 233476 163000
rect 233528 162988 233534 163040
rect 172934 162784 172940 162836
rect 172992 162824 172998 162836
rect 179098 162824 179104 162836
rect 172992 162796 179104 162824
rect 172992 162784 172998 162796
rect 179098 162784 179104 162796
rect 179156 162784 179162 162836
rect 80106 162716 80112 162768
rect 80164 162756 80170 162768
rect 87190 162756 87196 162768
rect 80164 162728 87196 162756
rect 80164 162716 80170 162728
rect 87190 162716 87196 162728
rect 87248 162716 87254 162768
rect 80198 162648 80204 162700
rect 80256 162688 80262 162700
rect 87282 162688 87288 162700
rect 80256 162660 87288 162688
rect 80256 162648 80262 162660
rect 87282 162648 87288 162660
rect 87340 162648 87346 162700
rect 132638 162308 132644 162360
rect 132696 162348 132702 162360
rect 139722 162348 139728 162360
rect 132696 162320 139728 162348
rect 132696 162308 132702 162320
rect 139722 162308 139728 162320
rect 139780 162308 139786 162360
rect 172934 162240 172940 162292
rect 172992 162280 172998 162292
rect 179006 162280 179012 162292
rect 172992 162252 179012 162280
rect 172992 162240 172998 162252
rect 179006 162240 179012 162252
rect 179064 162240 179070 162292
rect 132638 162172 132644 162224
rect 132696 162212 132702 162224
rect 139906 162212 139912 162224
rect 132696 162184 139912 162212
rect 132696 162172 132702 162184
rect 139906 162172 139912 162184
rect 139964 162172 139970 162224
rect 132454 162104 132460 162156
rect 132512 162144 132518 162156
rect 135306 162144 135312 162156
rect 132512 162116 135312 162144
rect 132512 162104 132518 162116
rect 135306 162104 135312 162116
rect 135364 162104 135370 162156
rect 136226 162104 136232 162156
rect 136284 162144 136290 162156
rect 140458 162144 140464 162156
rect 136284 162116 140464 162144
rect 136284 162104 136290 162116
rect 140458 162104 140464 162116
rect 140516 162104 140522 162156
rect 132546 162036 132552 162088
rect 132604 162076 132610 162088
rect 134110 162076 134116 162088
rect 132604 162048 134116 162076
rect 132604 162036 132610 162048
rect 134110 162036 134116 162048
rect 134168 162036 134174 162088
rect 136318 162036 136324 162088
rect 136376 162076 136382 162088
rect 140550 162076 140556 162088
rect 136376 162048 140556 162076
rect 136376 162036 136382 162048
rect 140550 162036 140556 162048
rect 140608 162036 140614 162088
rect 179650 162036 179656 162088
rect 179708 162076 179714 162088
rect 182318 162076 182324 162088
rect 179708 162048 182324 162076
rect 179708 162036 179714 162048
rect 182318 162036 182324 162048
rect 182376 162036 182382 162088
rect 229330 162036 229336 162088
rect 229388 162076 229394 162088
rect 233470 162076 233476 162088
rect 229388 162048 233476 162076
rect 229388 162036 229394 162048
rect 233470 162036 233476 162048
rect 233528 162036 233534 162088
rect 226478 161628 226484 161680
rect 226536 161668 226542 161680
rect 233746 161668 233752 161680
rect 226536 161640 233752 161668
rect 226536 161628 226542 161640
rect 233746 161628 233752 161640
rect 233804 161628 233810 161680
rect 226478 161492 226484 161544
rect 226536 161532 226542 161544
rect 233838 161532 233844 161544
rect 226536 161504 233844 161532
rect 226536 161492 226542 161504
rect 233838 161492 233844 161504
rect 233896 161492 233902 161544
rect 80198 161424 80204 161476
rect 80256 161464 80262 161476
rect 87190 161464 87196 161476
rect 80256 161436 87196 161464
rect 80256 161424 80262 161436
rect 87190 161424 87196 161436
rect 87248 161424 87254 161476
rect 80106 161356 80112 161408
rect 80164 161396 80170 161408
rect 87374 161396 87380 161408
rect 80164 161368 87380 161396
rect 80164 161356 80170 161368
rect 87374 161356 87380 161368
rect 87432 161356 87438 161408
rect 80014 161288 80020 161340
rect 80072 161328 80078 161340
rect 87282 161328 87288 161340
rect 80072 161300 87288 161328
rect 80072 161288 80078 161300
rect 87282 161288 87288 161300
rect 87340 161288 87346 161340
rect 225926 161152 225932 161204
rect 225984 161192 225990 161204
rect 233562 161192 233568 161204
rect 225984 161164 233568 161192
rect 225984 161152 225990 161164
rect 233562 161152 233568 161164
rect 233620 161152 233626 161204
rect 181030 160948 181036 161000
rect 181088 160988 181094 161000
rect 181858 160988 181864 161000
rect 181088 160960 181864 160988
rect 181088 160948 181094 160960
rect 181858 160948 181864 160960
rect 181916 160948 181922 161000
rect 132638 160880 132644 160932
rect 132696 160920 132702 160932
rect 139998 160920 140004 160932
rect 132696 160892 140004 160920
rect 132696 160880 132702 160892
rect 139998 160880 140004 160892
rect 140056 160880 140062 160932
rect 173946 160880 173952 160932
rect 174004 160920 174010 160932
rect 181950 160920 181956 160932
rect 174004 160892 181956 160920
rect 174004 160880 174010 160892
rect 181950 160880 181956 160892
rect 182008 160880 182014 160932
rect 136410 160812 136416 160864
rect 136468 160852 136474 160864
rect 139814 160852 139820 160864
rect 136468 160824 139820 160852
rect 136468 160812 136474 160824
rect 139814 160812 139820 160824
rect 139872 160812 139878 160864
rect 174038 160812 174044 160864
rect 174096 160852 174102 160864
rect 181030 160852 181036 160864
rect 174096 160824 181036 160852
rect 174096 160812 174102 160824
rect 181030 160812 181036 160824
rect 181088 160812 181094 160864
rect 173118 160744 173124 160796
rect 173176 160784 173182 160796
rect 173946 160784 173952 160796
rect 173176 160756 173952 160784
rect 173176 160744 173182 160756
rect 173946 160744 173952 160756
rect 174004 160744 174010 160796
rect 174866 160744 174872 160796
rect 174924 160784 174930 160796
rect 182318 160784 182324 160796
rect 174924 160756 182324 160784
rect 174924 160744 174930 160756
rect 182318 160744 182324 160756
rect 182376 160744 182382 160796
rect 132546 160676 132552 160728
rect 132604 160716 132610 160728
rect 140090 160716 140096 160728
rect 132604 160688 140096 160716
rect 132604 160676 132610 160688
rect 140090 160676 140096 160688
rect 140148 160676 140154 160728
rect 180110 160676 180116 160728
rect 180168 160716 180174 160728
rect 182134 160716 182140 160728
rect 180168 160688 182140 160716
rect 180168 160676 180174 160688
rect 182134 160676 182140 160688
rect 182192 160676 182198 160728
rect 136502 160608 136508 160660
rect 136560 160648 136566 160660
rect 140458 160648 140464 160660
rect 136560 160620 140464 160648
rect 136560 160608 136566 160620
rect 140458 160608 140464 160620
rect 140516 160608 140522 160660
rect 175418 160608 175424 160660
rect 175476 160648 175482 160660
rect 181398 160648 181404 160660
rect 175476 160620 181404 160648
rect 175476 160608 175482 160620
rect 181398 160608 181404 160620
rect 181456 160608 181462 160660
rect 226478 160540 226484 160592
rect 226536 160580 226542 160592
rect 229330 160580 229336 160592
rect 226536 160552 229336 160580
rect 226536 160540 226542 160552
rect 229330 160540 229336 160552
rect 229388 160540 229394 160592
rect 225926 160472 225932 160524
rect 225984 160512 225990 160524
rect 233470 160512 233476 160524
rect 225984 160484 233476 160512
rect 225984 160472 225990 160484
rect 233470 160472 233476 160484
rect 233528 160472 233534 160524
rect 173026 160376 173032 160388
rect 172987 160348 173032 160376
rect 173026 160336 173032 160348
rect 173084 160336 173090 160388
rect 225558 160268 225564 160320
rect 225616 160308 225622 160320
rect 233654 160308 233660 160320
rect 225616 160280 233660 160308
rect 225616 160268 225622 160280
rect 233654 160268 233660 160280
rect 233712 160268 233718 160320
rect 80106 159928 80112 159980
rect 80164 159968 80170 159980
rect 87190 159968 87196 159980
rect 80164 159940 87196 159968
rect 80164 159928 80170 159940
rect 87190 159928 87196 159940
rect 87248 159928 87254 159980
rect 173302 159928 173308 159980
rect 173360 159968 173366 159980
rect 180478 159968 180484 159980
rect 173360 159940 180484 159968
rect 173360 159928 173366 159940
rect 180478 159928 180484 159940
rect 180536 159928 180542 159980
rect 80198 159860 80204 159912
rect 80256 159900 80262 159912
rect 87282 159900 87288 159912
rect 80256 159872 87288 159900
rect 80256 159860 80262 159872
rect 87282 159860 87288 159872
rect 87340 159860 87346 159912
rect 226478 159724 226484 159776
rect 226536 159764 226542 159776
rect 233562 159764 233568 159776
rect 226536 159736 233568 159764
rect 226536 159724 226542 159736
rect 233562 159724 233568 159736
rect 233620 159724 233626 159776
rect 172750 159588 172756 159640
rect 172808 159628 172814 159640
rect 180662 159628 180668 159640
rect 172808 159600 180668 159628
rect 172808 159588 172814 159600
rect 180662 159588 180668 159600
rect 180720 159588 180726 159640
rect 173210 159520 173216 159572
rect 173268 159560 173274 159572
rect 174038 159560 174044 159572
rect 173268 159532 174044 159560
rect 173268 159520 173274 159532
rect 174038 159520 174044 159532
rect 174096 159520 174102 159572
rect 132638 159452 132644 159504
rect 132696 159492 132702 159504
rect 140918 159492 140924 159504
rect 132696 159464 140924 159492
rect 132696 159452 132702 159464
rect 140918 159452 140924 159464
rect 140976 159452 140982 159504
rect 176062 159452 176068 159504
rect 176120 159492 176126 159504
rect 181398 159492 181404 159504
rect 176120 159464 181404 159492
rect 176120 159452 176126 159464
rect 181398 159452 181404 159464
rect 181456 159452 181462 159504
rect 132454 159384 132460 159436
rect 132512 159424 132518 159436
rect 139262 159424 139268 159436
rect 132512 159396 139268 159424
rect 132512 159384 132518 159396
rect 139262 159384 139268 159396
rect 139320 159384 139326 159436
rect 174038 159384 174044 159436
rect 174096 159424 174102 159436
rect 180386 159424 180392 159436
rect 174096 159396 180392 159424
rect 174096 159384 174102 159396
rect 180386 159384 180392 159396
rect 180444 159384 180450 159436
rect 132546 159316 132552 159368
rect 132604 159356 132610 159368
rect 140734 159356 140740 159368
rect 132604 159328 140740 159356
rect 132604 159316 132610 159328
rect 140734 159316 140740 159328
rect 140792 159316 140798 159368
rect 176890 159316 176896 159368
rect 176948 159356 176954 159368
rect 181306 159356 181312 159368
rect 176948 159328 181312 159356
rect 176948 159316 176954 159328
rect 181306 159316 181312 159328
rect 181364 159316 181370 159368
rect 132638 159248 132644 159300
rect 132696 159288 132702 159300
rect 134938 159288 134944 159300
rect 132696 159260 134944 159288
rect 132696 159248 132702 159260
rect 134938 159248 134944 159260
rect 134996 159248 135002 159300
rect 176982 159248 176988 159300
rect 177040 159288 177046 159300
rect 181030 159288 181036 159300
rect 177040 159260 181036 159288
rect 177040 159248 177046 159260
rect 181030 159248 181036 159260
rect 181088 159248 181094 159300
rect 80198 159180 80204 159232
rect 80256 159220 80262 159232
rect 87190 159220 87196 159232
rect 80256 159192 87196 159220
rect 80256 159180 80262 159192
rect 87190 159180 87196 159192
rect 87248 159180 87254 159232
rect 226478 158908 226484 158960
rect 226536 158948 226542 158960
rect 233470 158948 233476 158960
rect 226536 158920 233476 158948
rect 226536 158908 226542 158920
rect 233470 158908 233476 158920
rect 233528 158908 233534 158960
rect 225558 158636 225564 158688
rect 225616 158676 225622 158688
rect 233562 158676 233568 158688
rect 225616 158648 233568 158676
rect 225616 158636 225622 158648
rect 233562 158636 233568 158648
rect 233620 158636 233626 158688
rect 80198 158500 80204 158552
rect 80256 158540 80262 158552
rect 87282 158540 87288 158552
rect 80256 158512 87288 158540
rect 80256 158500 80262 158512
rect 87282 158500 87288 158512
rect 87340 158500 87346 158552
rect 226386 158228 226392 158280
rect 226444 158268 226450 158280
rect 233470 158268 233476 158280
rect 226444 158240 233476 158268
rect 226444 158228 226450 158240
rect 233470 158228 233476 158240
rect 233528 158228 233534 158280
rect 173302 158160 173308 158212
rect 173360 158200 173366 158212
rect 176338 158200 176344 158212
rect 173360 158172 176344 158200
rect 173360 158160 173366 158172
rect 176338 158160 176344 158172
rect 176396 158160 176402 158212
rect 132546 158092 132552 158144
rect 132604 158132 132610 158144
rect 140642 158132 140648 158144
rect 132604 158104 140648 158132
rect 132604 158092 132610 158104
rect 140642 158092 140648 158104
rect 140700 158092 140706 158144
rect 132638 158024 132644 158076
rect 132696 158064 132702 158076
rect 140550 158064 140556 158076
rect 132696 158036 140556 158064
rect 132696 158024 132702 158036
rect 140550 158024 140556 158036
rect 140608 158024 140614 158076
rect 135214 157956 135220 158008
rect 135272 157996 135278 158008
rect 140366 157996 140372 158008
rect 135272 157968 140372 157996
rect 135272 157956 135278 157968
rect 140366 157956 140372 157968
rect 140424 157956 140430 158008
rect 132362 157928 132368 157940
rect 132288 157900 132368 157928
rect 80106 157820 80112 157872
rect 80164 157860 80170 157872
rect 87190 157860 87196 157872
rect 80164 157832 87196 157860
rect 80164 157820 80170 157832
rect 87190 157820 87196 157832
rect 87248 157820 87254 157872
rect 80198 157752 80204 157804
rect 80256 157792 80262 157804
rect 87282 157792 87288 157804
rect 80256 157764 87288 157792
rect 80256 157752 80262 157764
rect 87282 157752 87288 157764
rect 87340 157752 87346 157804
rect 132288 157736 132316 157900
rect 132362 157888 132368 157900
rect 132420 157888 132426 157940
rect 132454 157888 132460 157940
rect 132512 157928 132518 157940
rect 136134 157928 136140 157940
rect 132512 157900 136140 157928
rect 132512 157888 132518 157900
rect 136134 157888 136140 157900
rect 136192 157888 136198 157940
rect 173118 157888 173124 157940
rect 173176 157928 173182 157940
rect 176246 157928 176252 157940
rect 173176 157900 176252 157928
rect 173176 157888 173182 157900
rect 176246 157888 176252 157900
rect 176304 157888 176310 157940
rect 178270 157888 178276 157940
rect 178328 157928 178334 157940
rect 181490 157928 181496 157940
rect 178328 157900 181496 157928
rect 178328 157888 178334 157900
rect 181490 157888 181496 157900
rect 181548 157888 181554 157940
rect 79462 157684 79468 157736
rect 79520 157724 79526 157736
rect 87374 157724 87380 157736
rect 79520 157696 87380 157724
rect 79520 157684 79526 157696
rect 87374 157684 87380 157696
rect 87432 157684 87438 157736
rect 132270 157684 132276 157736
rect 132328 157684 132334 157736
rect 226294 157684 226300 157736
rect 226352 157724 226358 157736
rect 233470 157724 233476 157736
rect 226352 157696 233476 157724
rect 226352 157684 226358 157696
rect 233470 157684 233476 157696
rect 233528 157684 233534 157736
rect 173118 157616 173124 157668
rect 173176 157656 173182 157668
rect 180938 157656 180944 157668
rect 173176 157628 180944 157656
rect 173176 157616 173182 157628
rect 180938 157616 180944 157628
rect 180996 157616 181002 157668
rect 173210 157548 173216 157600
rect 173268 157588 173274 157600
rect 177902 157588 177908 157600
rect 173268 157560 177908 157588
rect 173268 157548 173274 157560
rect 177902 157548 177908 157560
rect 177960 157548 177966 157600
rect 226478 157412 226484 157464
rect 226536 157452 226542 157464
rect 233470 157452 233476 157464
rect 226536 157424 233476 157452
rect 226536 157412 226542 157424
rect 233470 157412 233476 157424
rect 233528 157412 233534 157464
rect 131534 157140 131540 157192
rect 131592 157180 131598 157192
rect 140826 157180 140832 157192
rect 131592 157152 140832 157180
rect 131592 157140 131598 157152
rect 140826 157140 140832 157152
rect 140884 157140 140890 157192
rect 173029 157183 173087 157189
rect 173029 157149 173041 157183
rect 173075 157180 173087 157183
rect 173210 157180 173216 157192
rect 173075 157152 173216 157180
rect 173075 157149 173087 157152
rect 173029 157143 173087 157149
rect 173210 157140 173216 157152
rect 173268 157140 173274 157192
rect 132546 157072 132552 157124
rect 132604 157112 132610 157124
rect 137514 157112 137520 157124
rect 132604 157084 137520 157112
rect 132604 157072 132610 157084
rect 137514 157072 137520 157084
rect 137572 157072 137578 157124
rect 172934 157072 172940 157124
rect 172992 157112 172998 157124
rect 177626 157112 177632 157124
rect 172992 157084 177632 157112
rect 172992 157072 172998 157084
rect 177626 157072 177632 157084
rect 177684 157072 177690 157124
rect 138802 156936 138808 156988
rect 138860 156976 138866 156988
rect 140182 156976 140188 156988
rect 138860 156948 140188 156976
rect 138860 156936 138866 156948
rect 140182 156936 140188 156948
rect 140240 156936 140246 156988
rect 226478 156936 226484 156988
rect 226536 156976 226542 156988
rect 233470 156976 233476 156988
rect 226536 156948 233476 156976
rect 226536 156936 226542 156948
rect 233470 156936 233476 156948
rect 233528 156936 233534 156988
rect 132638 156732 132644 156784
rect 132696 156772 132702 156784
rect 140458 156772 140464 156784
rect 132696 156744 140464 156772
rect 132696 156732 132702 156744
rect 140458 156732 140464 156744
rect 140516 156732 140522 156784
rect 139722 156664 139728 156716
rect 139780 156704 139786 156716
rect 140090 156704 140096 156716
rect 139780 156676 140096 156704
rect 139780 156664 139786 156676
rect 140090 156664 140096 156676
rect 140148 156664 140154 156716
rect 132546 156596 132552 156648
rect 132604 156636 132610 156648
rect 138894 156636 138900 156648
rect 132604 156608 138900 156636
rect 132604 156596 132610 156608
rect 138894 156596 138900 156608
rect 138952 156596 138958 156648
rect 132638 156528 132644 156580
rect 132696 156568 132702 156580
rect 140366 156568 140372 156580
rect 132696 156540 140372 156568
rect 132696 156528 132702 156540
rect 140366 156528 140372 156540
rect 140424 156528 140430 156580
rect 225374 156528 225380 156580
rect 225432 156568 225438 156580
rect 233470 156568 233476 156580
rect 225432 156540 233476 156568
rect 225432 156528 225438 156540
rect 233470 156528 233476 156540
rect 233528 156528 233534 156580
rect 131902 156460 131908 156512
rect 131960 156500 131966 156512
rect 132546 156500 132552 156512
rect 131960 156472 132552 156500
rect 131960 156460 131966 156472
rect 132546 156460 132552 156472
rect 132604 156460 132610 156512
rect 180202 156460 180208 156512
rect 180260 156500 180266 156512
rect 182042 156500 182048 156512
rect 180260 156472 182048 156500
rect 180260 156460 180266 156472
rect 182042 156460 182048 156472
rect 182100 156460 182106 156512
rect 80106 156392 80112 156444
rect 80164 156432 80170 156444
rect 87190 156432 87196 156444
rect 80164 156404 87196 156432
rect 80164 156392 80170 156404
rect 87190 156392 87196 156404
rect 87248 156392 87254 156444
rect 177534 156392 177540 156444
rect 177592 156432 177598 156444
rect 181030 156432 181036 156444
rect 177592 156404 181036 156432
rect 177592 156392 177598 156404
rect 181030 156392 181036 156404
rect 181088 156392 181094 156444
rect 80198 156324 80204 156376
rect 80256 156364 80262 156376
rect 87282 156364 87288 156376
rect 80256 156336 87288 156364
rect 80256 156324 80262 156336
rect 87282 156324 87288 156336
rect 87340 156324 87346 156376
rect 174038 156324 174044 156376
rect 174096 156364 174102 156376
rect 181122 156364 181128 156376
rect 174096 156336 181128 156364
rect 174096 156324 174102 156336
rect 181122 156324 181128 156336
rect 181180 156324 181186 156376
rect 173946 156188 173952 156240
rect 174004 156228 174010 156240
rect 181214 156228 181220 156240
rect 174004 156200 181220 156228
rect 174004 156188 174010 156200
rect 181214 156188 181220 156200
rect 181272 156188 181278 156240
rect 226478 155984 226484 156036
rect 226536 156024 226542 156036
rect 233470 156024 233476 156036
rect 226536 155996 233476 156024
rect 226536 155984 226542 155996
rect 233470 155984 233476 155996
rect 233528 155984 233534 156036
rect 226478 155576 226484 155628
rect 226536 155616 226542 155628
rect 233562 155616 233568 155628
rect 226536 155588 233568 155616
rect 226536 155576 226542 155588
rect 233562 155576 233568 155588
rect 233620 155576 233626 155628
rect 225558 155304 225564 155356
rect 225616 155344 225622 155356
rect 233470 155344 233476 155356
rect 225616 155316 233476 155344
rect 225616 155304 225622 155316
rect 233470 155304 233476 155316
rect 233528 155304 233534 155356
rect 131810 155100 131816 155152
rect 131868 155140 131874 155152
rect 134846 155140 134852 155152
rect 131868 155112 134852 155140
rect 131868 155100 131874 155112
rect 134846 155100 134852 155112
rect 134904 155100 134910 155152
rect 135122 155100 135128 155152
rect 135180 155140 135186 155152
rect 139722 155140 139728 155152
rect 135180 155112 139728 155140
rect 135180 155100 135186 155112
rect 139722 155100 139728 155112
rect 139780 155100 139786 155152
rect 80106 155032 80112 155084
rect 80164 155072 80170 155084
rect 87374 155072 87380 155084
rect 80164 155044 87380 155072
rect 80164 155032 80170 155044
rect 87374 155032 87380 155044
rect 87432 155032 87438 155084
rect 131350 155032 131356 155084
rect 131408 155072 131414 155084
rect 135030 155072 135036 155084
rect 131408 155044 135036 155072
rect 131408 155032 131414 155044
rect 135030 155032 135036 155044
rect 135088 155032 135094 155084
rect 135306 155032 135312 155084
rect 135364 155072 135370 155084
rect 139630 155072 139636 155084
rect 135364 155044 139636 155072
rect 135364 155032 135370 155044
rect 139630 155032 139636 155044
rect 139688 155032 139694 155084
rect 172934 155032 172940 155084
rect 172992 155072 172998 155084
rect 175418 155072 175424 155084
rect 172992 155044 175424 155072
rect 172992 155032 172998 155044
rect 175418 155032 175424 155044
rect 175476 155032 175482 155084
rect 178914 155032 178920 155084
rect 178972 155072 178978 155084
rect 181214 155072 181220 155084
rect 178972 155044 181220 155072
rect 178972 155032 178978 155044
rect 181214 155032 181220 155044
rect 181272 155032 181278 155084
rect 80014 154964 80020 155016
rect 80072 155004 80078 155016
rect 87190 155004 87196 155016
rect 80072 154976 87196 155004
rect 80072 154964 80078 154976
rect 87190 154964 87196 154976
rect 87248 154964 87254 155016
rect 131442 154964 131448 155016
rect 131500 155004 131506 155016
rect 134021 155007 134079 155013
rect 134021 155004 134033 155007
rect 131500 154976 134033 155004
rect 131500 154964 131506 154976
rect 134021 154973 134033 154976
rect 134067 154973 134079 155007
rect 134021 154967 134079 154973
rect 134110 154964 134116 155016
rect 134168 155004 134174 155016
rect 139722 155004 139728 155016
rect 134168 154976 139728 155004
rect 134168 154964 134174 154976
rect 139722 154964 139728 154976
rect 139780 154964 139786 155016
rect 173946 154964 173952 155016
rect 174004 155004 174010 155016
rect 179650 155004 179656 155016
rect 174004 154976 179656 155004
rect 174004 154964 174010 154976
rect 179650 154964 179656 154976
rect 179708 154964 179714 155016
rect 181030 155004 181036 155016
rect 179760 154976 181036 155004
rect 173026 154896 173032 154948
rect 173084 154936 173090 154948
rect 179760 154936 179788 154976
rect 181030 154964 181036 154976
rect 181088 154964 181094 155016
rect 173084 154908 179788 154936
rect 173084 154896 173090 154908
rect 131350 154828 131356 154880
rect 131408 154868 131414 154880
rect 138986 154868 138992 154880
rect 131408 154840 138992 154868
rect 131408 154828 131414 154840
rect 138986 154828 138992 154840
rect 139044 154828 139050 154880
rect 174038 154828 174044 154880
rect 174096 154868 174102 154880
rect 181122 154868 181128 154880
rect 174096 154840 181128 154868
rect 174096 154828 174102 154840
rect 181122 154828 181128 154840
rect 181180 154828 181186 154880
rect 134021 154803 134079 154809
rect 134021 154769 134033 154803
rect 134067 154800 134079 154803
rect 139078 154800 139084 154812
rect 134067 154772 139084 154800
rect 134067 154769 134079 154772
rect 134021 154763 134079 154769
rect 139078 154760 139084 154772
rect 139136 154760 139142 154812
rect 80198 154556 80204 154608
rect 80256 154596 80262 154608
rect 87098 154596 87104 154608
rect 80256 154568 87104 154596
rect 80256 154556 80262 154568
rect 87098 154556 87104 154568
rect 87156 154556 87162 154608
rect 225742 154488 225748 154540
rect 225800 154528 225806 154540
rect 233562 154528 233568 154540
rect 225800 154500 233568 154528
rect 225800 154488 225806 154500
rect 233562 154488 233568 154500
rect 233620 154488 233626 154540
rect 173118 154420 173124 154472
rect 173176 154460 173182 154472
rect 174866 154460 174872 154472
rect 173176 154432 174872 154460
rect 173176 154420 173182 154432
rect 174866 154420 174872 154432
rect 174924 154420 174930 154472
rect 225834 154080 225840 154132
rect 225892 154120 225898 154132
rect 233654 154120 233660 154132
rect 225892 154092 233660 154120
rect 225892 154080 225898 154092
rect 233654 154080 233660 154092
rect 233712 154080 233718 154132
rect 79922 153876 79928 153928
rect 79980 153916 79986 153928
rect 87190 153916 87196 153928
rect 79980 153888 87196 153916
rect 79980 153876 79986 153888
rect 87190 153876 87196 153888
rect 87248 153876 87254 153928
rect 226110 153808 226116 153860
rect 226168 153848 226174 153860
rect 233470 153848 233476 153860
rect 226168 153820 233476 153848
rect 226168 153808 226174 153820
rect 233470 153808 233476 153820
rect 233528 153808 233534 153860
rect 226478 153740 226484 153792
rect 226536 153780 226542 153792
rect 233746 153780 233752 153792
rect 226536 153752 233752 153780
rect 226536 153740 226542 153752
rect 233746 153740 233752 153752
rect 233804 153740 233810 153792
rect 173210 153604 173216 153656
rect 173268 153644 173274 153656
rect 181214 153644 181220 153656
rect 173268 153616 181220 153644
rect 173268 153604 173274 153616
rect 181214 153604 181220 153616
rect 181272 153604 181278 153656
rect 173302 153536 173308 153588
rect 173360 153576 173366 153588
rect 181030 153576 181036 153588
rect 173360 153548 181036 153576
rect 173360 153536 173366 153548
rect 181030 153536 181036 153548
rect 181088 153536 181094 153588
rect 172842 153468 172848 153520
rect 172900 153508 172906 153520
rect 172900 153480 176752 153508
rect 172900 153468 172906 153480
rect 173302 153400 173308 153452
rect 173360 153440 173366 153452
rect 176062 153440 176068 153452
rect 173360 153412 176068 153440
rect 173360 153400 173366 153412
rect 176062 153400 176068 153412
rect 176120 153400 176126 153452
rect 176724 153440 176752 153480
rect 181122 153440 181128 153452
rect 176724 153412 181128 153440
rect 181122 153400 181128 153412
rect 181180 153400 181186 153452
rect 226110 153400 226116 153452
rect 226168 153440 226174 153452
rect 233562 153440 233568 153452
rect 226168 153412 233568 153440
rect 226168 153400 226174 153412
rect 233562 153400 233568 153412
rect 233620 153400 233626 153452
rect 174038 153332 174044 153384
rect 174096 153372 174102 153384
rect 180110 153372 180116 153384
rect 174096 153344 180116 153372
rect 174096 153332 174102 153344
rect 180110 153332 180116 153344
rect 180168 153332 180174 153384
rect 80198 153196 80204 153248
rect 80256 153236 80262 153248
rect 87006 153236 87012 153248
rect 80256 153208 87012 153236
rect 80256 153196 80262 153208
rect 87006 153196 87012 153208
rect 87064 153196 87070 153248
rect 80198 152924 80204 152976
rect 80256 152964 80262 152976
rect 86914 152964 86920 152976
rect 80256 152936 86920 152964
rect 80256 152924 80262 152936
rect 86914 152924 86920 152936
rect 86972 152924 86978 152976
rect 225374 152584 225380 152636
rect 225432 152624 225438 152636
rect 233838 152624 233844 152636
rect 225432 152596 233844 152624
rect 225432 152584 225438 152596
rect 233838 152584 233844 152596
rect 233896 152584 233902 152636
rect 85810 152448 85816 152500
rect 85868 152488 85874 152500
rect 87926 152488 87932 152500
rect 85868 152460 87932 152488
rect 85868 152448 85874 152460
rect 87926 152448 87932 152460
rect 87984 152448 87990 152500
rect 85902 152380 85908 152432
rect 85960 152420 85966 152432
rect 87558 152420 87564 152432
rect 85960 152392 87564 152420
rect 85960 152380 85966 152392
rect 87558 152380 87564 152392
rect 87616 152380 87622 152432
rect 225742 152380 225748 152432
rect 225800 152420 225806 152432
rect 233470 152420 233476 152432
rect 225800 152392 233476 152420
rect 225800 152380 225806 152392
rect 233470 152380 233476 152392
rect 233528 152380 233534 152432
rect 80106 152312 80112 152364
rect 80164 152352 80170 152364
rect 87098 152352 87104 152364
rect 80164 152324 87104 152352
rect 80164 152312 80170 152324
rect 87098 152312 87104 152324
rect 87156 152312 87162 152364
rect 131534 152312 131540 152364
rect 131592 152352 131598 152364
rect 136502 152352 136508 152364
rect 131592 152324 136508 152352
rect 131592 152312 131598 152324
rect 136502 152312 136508 152324
rect 136560 152312 136566 152364
rect 179098 152312 179104 152364
rect 179156 152352 179162 152364
rect 181030 152352 181036 152364
rect 179156 152324 181036 152352
rect 179156 152312 179162 152324
rect 181030 152312 181036 152324
rect 181088 152312 181094 152364
rect 131350 152244 131356 152296
rect 131408 152284 131414 152296
rect 136226 152284 136232 152296
rect 131408 152256 136232 152284
rect 131408 152244 131414 152256
rect 136226 152244 136232 152256
rect 136284 152244 136290 152296
rect 174038 152244 174044 152296
rect 174096 152284 174102 152296
rect 176890 152284 176896 152296
rect 174096 152256 176896 152284
rect 174096 152244 174102 152256
rect 176890 152244 176896 152256
rect 176948 152244 176954 152296
rect 179006 152244 179012 152296
rect 179064 152284 179070 152296
rect 181122 152284 181128 152296
rect 179064 152256 181128 152284
rect 179064 152244 179070 152256
rect 181122 152244 181128 152256
rect 181180 152244 181186 152296
rect 131442 152176 131448 152228
rect 131500 152216 131506 152228
rect 136410 152216 136416 152228
rect 131500 152188 136416 152216
rect 131500 152176 131506 152188
rect 136410 152176 136416 152188
rect 136468 152176 136474 152228
rect 131350 152108 131356 152160
rect 131408 152148 131414 152160
rect 136318 152148 136324 152160
rect 131408 152120 136324 152148
rect 131408 152108 131414 152120
rect 136318 152108 136324 152120
rect 136376 152108 136382 152160
rect 173302 151836 173308 151888
rect 173360 151876 173366 151888
rect 176982 151876 176988 151888
rect 173360 151848 176988 151876
rect 173360 151836 173366 151848
rect 176982 151836 176988 151848
rect 177040 151836 177046 151888
rect 225926 151700 225932 151752
rect 225984 151740 225990 151752
rect 227950 151740 227956 151752
rect 225984 151712 227956 151740
rect 225984 151700 225990 151712
rect 227950 151700 227956 151712
rect 228008 151700 228014 151752
rect 80198 151496 80204 151548
rect 80256 151536 80262 151548
rect 86822 151536 86828 151548
rect 80256 151508 86828 151536
rect 80256 151496 80262 151508
rect 86822 151496 86828 151508
rect 86880 151496 86886 151548
rect 173946 151428 173952 151480
rect 174004 151468 174010 151480
rect 178270 151468 178276 151480
rect 174004 151440 178276 151468
rect 174004 151428 174010 151440
rect 178270 151428 178276 151440
rect 178328 151428 178334 151480
rect 225374 151360 225380 151412
rect 225432 151400 225438 151412
rect 229238 151400 229244 151412
rect 225432 151372 229244 151400
rect 225432 151360 225438 151372
rect 229238 151360 229244 151372
rect 229296 151360 229302 151412
rect 79370 151088 79376 151140
rect 79428 151128 79434 151140
rect 87282 151128 87288 151140
rect 79428 151100 87288 151128
rect 79428 151088 79434 151100
rect 87282 151088 87288 151100
rect 87340 151088 87346 151140
rect 226478 151088 226484 151140
rect 226536 151128 226542 151140
rect 228042 151128 228048 151140
rect 226536 151100 228048 151128
rect 226536 151088 226542 151100
rect 228042 151088 228048 151100
rect 228100 151088 228106 151140
rect 79738 151020 79744 151072
rect 79796 151060 79802 151072
rect 87374 151060 87380 151072
rect 79796 151032 87380 151060
rect 79796 151020 79802 151032
rect 87374 151020 87380 151032
rect 87432 151020 87438 151072
rect 79278 150952 79284 151004
rect 79336 150992 79342 151004
rect 87190 150992 87196 151004
rect 79336 150964 87196 150992
rect 79336 150952 79342 150964
rect 87190 150952 87196 150964
rect 87248 150952 87254 151004
rect 226110 150952 226116 151004
rect 226168 150992 226174 151004
rect 229146 150992 229152 151004
rect 226168 150964 229152 150992
rect 226168 150952 226174 150964
rect 229146 150952 229152 150964
rect 229204 150952 229210 151004
rect 133374 150884 133380 150936
rect 133432 150924 133438 150936
rect 139630 150924 139636 150936
rect 133432 150896 139636 150924
rect 133432 150884 133438 150896
rect 139630 150884 139636 150896
rect 139688 150884 139694 150936
rect 131350 150816 131356 150868
rect 131408 150856 131414 150868
rect 139354 150856 139360 150868
rect 131408 150828 139360 150856
rect 131408 150816 131414 150828
rect 139354 150816 139360 150828
rect 139412 150816 139418 150868
rect 172934 150816 172940 150868
rect 172992 150856 172998 150868
rect 182318 150856 182324 150868
rect 172992 150828 182324 150856
rect 172992 150816 172998 150828
rect 182318 150816 182324 150828
rect 182376 150816 182382 150868
rect 174038 150748 174044 150800
rect 174096 150788 174102 150800
rect 182134 150788 182140 150800
rect 174096 150760 182140 150788
rect 174096 150748 174102 150760
rect 182134 150748 182140 150760
rect 182192 150748 182198 150800
rect 131442 150680 131448 150732
rect 131500 150720 131506 150732
rect 139446 150720 139452 150732
rect 131500 150692 139452 150720
rect 131500 150680 131506 150692
rect 139446 150680 139452 150692
rect 139504 150680 139510 150732
rect 131350 150476 131356 150528
rect 131408 150516 131414 150528
rect 135214 150516 135220 150528
rect 131408 150488 135220 150516
rect 131408 150476 131414 150488
rect 135214 150476 135220 150488
rect 135272 150476 135278 150528
rect 80106 150340 80112 150392
rect 80164 150380 80170 150392
rect 85902 150380 85908 150392
rect 80164 150352 85908 150380
rect 80164 150340 80170 150352
rect 85902 150340 85908 150352
rect 85960 150340 85966 150392
rect 80198 150136 80204 150188
rect 80256 150176 80262 150188
rect 85810 150176 85816 150188
rect 80256 150148 85816 150176
rect 80256 150136 80262 150148
rect 85810 150136 85816 150148
rect 85868 150136 85874 150188
rect 225558 150068 225564 150120
rect 225616 150108 225622 150120
rect 230618 150108 230624 150120
rect 225616 150080 230624 150108
rect 225616 150068 225622 150080
rect 230618 150068 230624 150080
rect 230676 150068 230682 150120
rect 80014 149728 80020 149780
rect 80072 149768 80078 149780
rect 87374 149768 87380 149780
rect 80072 149740 87380 149768
rect 80072 149728 80078 149740
rect 87374 149728 87380 149740
rect 87432 149728 87438 149780
rect 79922 149660 79928 149712
rect 79980 149700 79986 149712
rect 87282 149700 87288 149712
rect 79980 149672 87288 149700
rect 79980 149660 79986 149672
rect 87282 149660 87288 149672
rect 87340 149660 87346 149712
rect 79830 149592 79836 149644
rect 79888 149632 79894 149644
rect 87190 149632 87196 149644
rect 79888 149604 87196 149632
rect 79888 149592 79894 149604
rect 87190 149592 87196 149604
rect 87248 149592 87254 149644
rect 225742 149592 225748 149644
rect 225800 149632 225806 149644
rect 230342 149632 230348 149644
rect 225800 149604 230348 149632
rect 225800 149592 225806 149604
rect 230342 149592 230348 149604
rect 230400 149592 230406 149644
rect 80198 149524 80204 149576
rect 80256 149564 80262 149576
rect 87742 149564 87748 149576
rect 80256 149536 87748 149564
rect 80256 149524 80262 149536
rect 87742 149524 87748 149536
rect 87800 149524 87806 149576
rect 131626 149524 131632 149576
rect 131684 149564 131690 149576
rect 139538 149564 139544 149576
rect 131684 149536 139544 149564
rect 131684 149524 131690 149536
rect 139538 149524 139544 149536
rect 139596 149524 139602 149576
rect 176246 149524 176252 149576
rect 176304 149564 176310 149576
rect 182318 149564 182324 149576
rect 176304 149536 182324 149564
rect 176304 149524 176310 149536
rect 182318 149524 182324 149536
rect 182376 149524 182382 149576
rect 227950 149524 227956 149576
rect 228008 149564 228014 149576
rect 233470 149564 233476 149576
rect 228008 149536 233476 149564
rect 228008 149524 228014 149536
rect 233470 149524 233476 149536
rect 233528 149524 233534 149576
rect 80106 149456 80112 149508
rect 80164 149496 80170 149508
rect 88110 149496 88116 149508
rect 80164 149468 88116 149496
rect 80164 149456 80170 149468
rect 88110 149456 88116 149468
rect 88168 149456 88174 149508
rect 131534 149456 131540 149508
rect 131592 149496 131598 149508
rect 139814 149496 139820 149508
rect 131592 149468 139820 149496
rect 131592 149456 131598 149468
rect 139814 149456 139820 149468
rect 139872 149456 139878 149508
rect 173302 149456 173308 149508
rect 173360 149496 173366 149508
rect 173854 149496 173860 149508
rect 173360 149468 173860 149496
rect 173360 149456 173366 149468
rect 173854 149456 173860 149468
rect 173912 149456 173918 149508
rect 176338 149456 176344 149508
rect 176396 149496 176402 149508
rect 181766 149496 181772 149508
rect 176396 149468 181772 149496
rect 176396 149456 176402 149468
rect 181766 149456 181772 149468
rect 181824 149456 181830 149508
rect 229146 149456 229152 149508
rect 229204 149496 229210 149508
rect 233562 149496 233568 149508
rect 229204 149468 233568 149496
rect 229204 149456 229210 149468
rect 233562 149456 233568 149468
rect 233620 149456 233626 149508
rect 131442 149388 131448 149440
rect 131500 149428 131506 149440
rect 139170 149428 139176 149440
rect 131500 149400 139176 149428
rect 131500 149388 131506 149400
rect 139170 149388 139176 149400
rect 139228 149388 139234 149440
rect 174038 149388 174044 149440
rect 174096 149428 174102 149440
rect 180754 149428 180760 149440
rect 174096 149400 180760 149428
rect 174096 149388 174102 149400
rect 180754 149388 180760 149400
rect 180812 149388 180818 149440
rect 131350 149320 131356 149372
rect 131408 149360 131414 149372
rect 138802 149360 138808 149372
rect 131408 149332 138808 149360
rect 131408 149320 131414 149332
rect 138802 149320 138808 149332
rect 138860 149320 138866 149372
rect 173854 149320 173860 149372
rect 173912 149360 173918 149372
rect 180202 149360 180208 149372
rect 173912 149332 180208 149360
rect 173912 149320 173918 149332
rect 180202 149320 180208 149332
rect 180260 149320 180266 149372
rect 225374 149048 225380 149100
rect 225432 149088 225438 149100
rect 233746 149088 233752 149100
rect 225432 149060 233752 149088
rect 225432 149048 225438 149060
rect 233746 149048 233752 149060
rect 233804 149048 233810 149100
rect 132270 148844 132276 148896
rect 132328 148884 132334 148896
rect 139630 148884 139636 148896
rect 132328 148856 139636 148884
rect 132328 148844 132334 148856
rect 139630 148844 139636 148856
rect 139688 148844 139694 148896
rect 174038 148844 174044 148896
rect 174096 148884 174102 148896
rect 180938 148884 180944 148896
rect 174096 148856 180944 148884
rect 174096 148844 174102 148856
rect 180938 148844 180944 148856
rect 180996 148844 181002 148896
rect 226478 148640 226484 148692
rect 226536 148680 226542 148692
rect 233930 148680 233936 148692
rect 226536 148652 233936 148680
rect 226536 148640 226542 148652
rect 233930 148640 233936 148652
rect 233988 148640 233994 148692
rect 225558 148300 225564 148352
rect 225616 148340 225622 148352
rect 233654 148340 233660 148352
rect 225616 148312 233660 148340
rect 225616 148300 225622 148312
rect 233654 148300 233660 148312
rect 233712 148300 233718 148352
rect 226478 148232 226484 148284
rect 226536 148272 226542 148284
rect 233838 148272 233844 148284
rect 226536 148244 233844 148272
rect 226536 148232 226542 148244
rect 233838 148232 233844 148244
rect 233896 148232 233902 148284
rect 134938 148164 134944 148216
rect 134996 148204 135002 148216
rect 139722 148204 139728 148216
rect 134996 148176 139728 148204
rect 134996 148164 135002 148176
rect 139722 148164 139728 148176
rect 139780 148164 139786 148216
rect 229238 148164 229244 148216
rect 229296 148204 229302 148216
rect 233470 148204 233476 148216
rect 229296 148176 233476 148204
rect 229296 148164 229302 148176
rect 233470 148164 233476 148176
rect 233528 148164 233534 148216
rect 131350 148096 131356 148148
rect 131408 148136 131414 148148
rect 135122 148136 135128 148148
rect 131408 148108 135128 148136
rect 131408 148096 131414 148108
rect 135122 148096 135128 148108
rect 135180 148096 135186 148148
rect 228042 148096 228048 148148
rect 228100 148136 228106 148148
rect 233562 148136 233568 148148
rect 228100 148108 233568 148136
rect 228100 148096 228106 148108
rect 233562 148096 233568 148108
rect 233620 148096 233626 148148
rect 177626 148028 177632 148080
rect 177684 148068 177690 148080
rect 182318 148068 182324 148080
rect 177684 148040 182324 148068
rect 177684 148028 177690 148040
rect 182318 148028 182324 148040
rect 182376 148028 182382 148080
rect 172750 147824 172756 147876
rect 172808 147864 172814 147876
rect 180846 147864 180852 147876
rect 172808 147836 180852 147864
rect 172808 147824 172814 147836
rect 180846 147824 180852 147836
rect 180904 147824 180910 147876
rect 174038 147756 174044 147808
rect 174096 147796 174102 147808
rect 180570 147796 180576 147808
rect 174096 147768 180576 147796
rect 174096 147756 174102 147768
rect 180570 147756 180576 147768
rect 180628 147756 180634 147808
rect 225558 147348 225564 147400
rect 225616 147388 225622 147400
rect 231998 147388 232004 147400
rect 225616 147360 232004 147388
rect 225616 147348 225622 147360
rect 231998 147348 232004 147360
rect 232056 147348 232062 147400
rect 136134 146736 136140 146788
rect 136192 146776 136198 146788
rect 139722 146776 139728 146788
rect 136192 146748 139728 146776
rect 136192 146736 136198 146748
rect 139722 146736 139728 146748
rect 139780 146736 139786 146788
rect 174038 146668 174044 146720
rect 174096 146708 174102 146720
rect 181950 146708 181956 146720
rect 174096 146680 181956 146708
rect 174096 146668 174102 146680
rect 181950 146668 181956 146680
rect 182008 146668 182014 146720
rect 230618 146668 230624 146720
rect 230676 146708 230682 146720
rect 233470 146708 233476 146720
rect 230676 146680 233476 146708
rect 230676 146668 230682 146680
rect 233470 146668 233476 146680
rect 233528 146668 233534 146720
rect 172750 146328 172756 146380
rect 172808 146368 172814 146380
rect 174774 146368 174780 146380
rect 172808 146340 174780 146368
rect 172808 146328 172814 146340
rect 174774 146328 174780 146340
rect 174832 146328 174838 146380
rect 230342 146328 230348 146380
rect 230400 146368 230406 146380
rect 233470 146368 233476 146380
rect 230400 146340 233476 146368
rect 230400 146328 230406 146340
rect 233470 146328 233476 146340
rect 233528 146328 233534 146380
rect 228318 145960 228324 145972
rect 228279 145932 228324 145960
rect 228318 145920 228324 145932
rect 228376 145920 228382 145972
rect 80198 145376 80204 145428
rect 80256 145416 80262 145428
rect 87466 145416 87472 145428
rect 80256 145388 87472 145416
rect 80256 145376 80262 145388
rect 87466 145376 87472 145388
rect 87524 145376 87530 145428
rect 137514 145376 137520 145428
rect 137572 145416 137578 145428
rect 139906 145416 139912 145428
rect 137572 145388 139912 145416
rect 137572 145376 137578 145388
rect 139906 145376 139912 145388
rect 139964 145376 139970 145428
rect 173670 145376 173676 145428
rect 173728 145416 173734 145428
rect 176154 145416 176160 145428
rect 173728 145388 176160 145416
rect 173728 145376 173734 145388
rect 176154 145376 176160 145388
rect 176212 145376 176218 145428
rect 176249 145419 176307 145425
rect 176249 145385 176261 145419
rect 176295 145416 176307 145419
rect 203846 145416 203852 145428
rect 176295 145388 203852 145416
rect 176295 145385 176307 145388
rect 176249 145379 176307 145385
rect 203846 145376 203852 145388
rect 203904 145416 203910 145428
rect 228321 145419 228379 145425
rect 228321 145416 228333 145419
rect 203904 145388 228333 145416
rect 203904 145376 203910 145388
rect 228321 145385 228333 145388
rect 228367 145385 228379 145419
rect 228321 145379 228379 145385
rect 226570 145308 226576 145360
rect 226628 145348 226634 145360
rect 233470 145348 233476 145360
rect 226628 145320 233476 145348
rect 226628 145308 226634 145320
rect 233470 145308 233476 145320
rect 233528 145308 233534 145360
rect 228318 145280 228324 145292
rect 228279 145252 228324 145280
rect 228318 145240 228324 145252
rect 228376 145240 228382 145292
rect 170818 144696 170824 144748
rect 170876 144736 170882 144748
rect 171370 144736 171376 144748
rect 170876 144708 171376 144736
rect 170876 144696 170882 144708
rect 171370 144696 171376 144708
rect 171428 144736 171434 144748
rect 176249 144739 176307 144745
rect 176249 144736 176261 144739
rect 171428 144708 176261 144736
rect 171428 144696 171434 144708
rect 176249 144705 176261 144708
rect 176295 144705 176307 144739
rect 176249 144699 176307 144705
rect 80014 144016 80020 144068
rect 80072 144056 80078 144068
rect 87190 144056 87196 144068
rect 80072 144028 87196 144056
rect 80072 144016 80078 144028
rect 87190 144016 87196 144028
rect 87248 144016 87254 144068
rect 109546 144016 109552 144068
rect 109604 144056 109610 144068
rect 134754 144056 134760 144068
rect 109604 144028 134760 144056
rect 109604 144016 109610 144028
rect 134754 144016 134760 144028
rect 134812 144016 134818 144068
rect 134846 144016 134852 144068
rect 134904 144056 134910 144068
rect 139722 144056 139728 144068
rect 134904 144028 139728 144056
rect 134904 144016 134910 144028
rect 139722 144016 139728 144028
rect 139780 144016 139786 144068
rect 296214 144016 296220 144068
rect 296272 144056 296278 144068
rect 300170 144056 300176 144068
rect 296272 144028 300176 144056
rect 296272 144016 296278 144028
rect 300170 144016 300176 144028
rect 300228 144016 300234 144068
rect 80198 143948 80204 144000
rect 80256 143988 80262 144000
rect 87558 143988 87564 144000
rect 80256 143960 87564 143988
rect 80256 143948 80262 143960
rect 87558 143948 87564 143960
rect 87616 143948 87622 144000
rect 80106 143880 80112 143932
rect 80164 143920 80170 143932
rect 87282 143920 87288 143932
rect 80164 143892 87288 143920
rect 80164 143880 80170 143892
rect 87282 143880 87288 143892
rect 87340 143880 87346 143932
rect 80198 142656 80204 142708
rect 80256 142696 80262 142708
rect 87374 142696 87380 142708
rect 80256 142668 87380 142696
rect 80256 142656 80262 142668
rect 87374 142656 87380 142668
rect 87432 142656 87438 142708
rect 231998 142656 232004 142708
rect 232056 142696 232062 142708
rect 233470 142696 233476 142708
rect 232056 142668 233476 142696
rect 232056 142656 232062 142668
rect 233470 142656 233476 142668
rect 233528 142656 233534 142708
rect 169990 141704 169996 141756
rect 170048 141744 170054 141756
rect 170634 141744 170640 141756
rect 170048 141716 170640 141744
rect 170048 141704 170054 141716
rect 170634 141704 170640 141716
rect 170692 141704 170698 141756
rect 168426 141636 168432 141688
rect 168484 141676 168490 141688
rect 170726 141676 170732 141688
rect 168484 141648 170732 141676
rect 168484 141636 168490 141648
rect 170726 141636 170732 141648
rect 170784 141636 170790 141688
rect 250033 139979 250091 139985
rect 59976 139948 61200 139976
rect 56738 139868 56744 139920
rect 56796 139908 56802 139920
rect 59976 139908 60004 139948
rect 56796 139880 60004 139908
rect 56796 139868 56802 139880
rect 60050 139868 60056 139920
rect 60108 139908 60114 139920
rect 61172 139908 61200 139948
rect 250033 139945 250045 139979
rect 250079 139976 250091 139979
rect 250079 139948 250904 139976
rect 250079 139945 250091 139948
rect 250033 139939 250091 139945
rect 65110 139908 65116 139920
rect 60108 139880 61108 139908
rect 61172 139880 65116 139908
rect 60108 139868 60114 139880
rect 56462 139800 56468 139852
rect 56520 139840 56526 139852
rect 60970 139840 60976 139852
rect 56520 139812 60976 139840
rect 56520 139800 56526 139812
rect 60970 139800 60976 139812
rect 61028 139800 61034 139852
rect 61080 139840 61108 139880
rect 65110 139868 65116 139880
rect 65168 139868 65174 139920
rect 131994 139868 132000 139920
rect 132052 139908 132058 139920
rect 168978 139908 168984 139920
rect 132052 139880 168984 139908
rect 132052 139868 132058 139880
rect 168978 139868 168984 139880
rect 169036 139868 169042 139920
rect 224454 139868 224460 139920
rect 224512 139908 224518 139920
rect 250677 139911 250735 139917
rect 250677 139908 250689 139911
rect 224512 139880 250689 139908
rect 224512 139868 224518 139880
rect 250677 139877 250689 139880
rect 250723 139877 250735 139911
rect 250677 139871 250735 139877
rect 67134 139840 67140 139852
rect 61080 139812 67140 139840
rect 67134 139800 67140 139812
rect 67192 139800 67198 139852
rect 140274 139800 140280 139852
rect 140332 139840 140338 139852
rect 169438 139840 169444 139852
rect 140332 139812 169444 139840
rect 140332 139800 140338 139812
rect 169438 139800 169444 139812
rect 169496 139800 169502 139852
rect 250766 139840 250772 139852
rect 244712 139812 250772 139840
rect 59958 139732 59964 139784
rect 60016 139772 60022 139784
rect 71826 139772 71832 139784
rect 60016 139744 71832 139772
rect 60016 139732 60022 139744
rect 71826 139732 71832 139744
rect 71884 139732 71890 139784
rect 149382 139732 149388 139784
rect 149440 139772 149446 139784
rect 157846 139772 157852 139784
rect 149440 139744 157852 139772
rect 149440 139732 149446 139744
rect 157846 139732 157852 139744
rect 157904 139732 157910 139784
rect 57106 139664 57112 139716
rect 57164 139704 57170 139716
rect 61249 139707 61307 139713
rect 61249 139704 61261 139707
rect 57164 139676 61261 139704
rect 57164 139664 57170 139676
rect 61249 139673 61261 139676
rect 61295 139673 61307 139707
rect 61249 139667 61307 139673
rect 61706 139664 61712 139716
rect 61764 139704 61770 139716
rect 63822 139704 63828 139716
rect 61764 139676 63828 139704
rect 61764 139664 61770 139676
rect 63822 139664 63828 139676
rect 63880 139664 63886 139716
rect 150486 139664 150492 139716
rect 150544 139704 150550 139716
rect 150544 139676 155040 139704
rect 150544 139664 150550 139676
rect 59866 139596 59872 139648
rect 59924 139636 59930 139648
rect 71090 139636 71096 139648
rect 59924 139608 71096 139636
rect 59924 139596 59930 139608
rect 71090 139596 71096 139608
rect 71148 139596 71154 139648
rect 155012 139636 155040 139676
rect 155270 139664 155276 139716
rect 155328 139704 155334 139716
rect 165758 139704 165764 139716
rect 155328 139676 165764 139704
rect 155328 139664 155334 139676
rect 165758 139664 165764 139676
rect 165816 139664 165822 139716
rect 242762 139664 242768 139716
rect 242820 139704 242826 139716
rect 244605 139707 244663 139713
rect 244605 139704 244617 139707
rect 242820 139676 244617 139704
rect 242820 139664 242826 139676
rect 244605 139673 244617 139676
rect 244651 139673 244663 139707
rect 244605 139667 244663 139673
rect 159226 139636 159232 139648
rect 155012 139608 159232 139636
rect 159226 139596 159232 139608
rect 159284 139596 159290 139648
rect 54438 139528 54444 139580
rect 54496 139568 54502 139580
rect 57566 139568 57572 139580
rect 54496 139540 57572 139568
rect 54496 139528 54502 139540
rect 57566 139528 57572 139540
rect 57624 139528 57630 139580
rect 59682 139528 59688 139580
rect 59740 139568 59746 139580
rect 60510 139568 60516 139580
rect 59740 139540 60516 139568
rect 59740 139528 59746 139540
rect 60510 139528 60516 139540
rect 60568 139528 60574 139580
rect 61154 139528 61160 139580
rect 61212 139568 61218 139580
rect 61982 139568 61988 139580
rect 61212 139540 61988 139568
rect 61212 139528 61218 139540
rect 61982 139528 61988 139540
rect 62040 139528 62046 139580
rect 62442 139528 62448 139580
rect 62500 139568 62506 139580
rect 65754 139568 65760 139580
rect 62500 139540 65760 139568
rect 62500 139528 62506 139540
rect 65754 139528 65760 139540
rect 65812 139528 65818 139580
rect 67226 139528 67232 139580
rect 67284 139568 67290 139580
rect 70446 139568 70452 139580
rect 67284 139540 70452 139568
rect 67284 139528 67290 139540
rect 70446 139528 70452 139540
rect 70504 139528 70510 139580
rect 70541 139571 70599 139577
rect 70541 139537 70553 139571
rect 70587 139568 70599 139571
rect 73758 139568 73764 139580
rect 70587 139540 73764 139568
rect 70587 139537 70599 139540
rect 70541 139531 70599 139537
rect 73758 139528 73764 139540
rect 73816 139528 73822 139580
rect 154994 139528 155000 139580
rect 155052 139568 155058 139580
rect 166310 139568 166316 139580
rect 155052 139540 166316 139568
rect 155052 139528 155058 139540
rect 166310 139528 166316 139540
rect 166368 139528 166374 139580
rect 243038 139528 243044 139580
rect 243096 139568 243102 139580
rect 244712 139568 244740 139812
rect 250766 139800 250772 139812
rect 250824 139800 250830 139852
rect 250876 139840 250904 139948
rect 250953 139911 251011 139917
rect 250953 139877 250965 139911
rect 250999 139908 251011 139911
rect 263830 139908 263836 139920
rect 250999 139880 263836 139908
rect 250999 139877 251011 139880
rect 250953 139871 251011 139877
rect 263830 139868 263836 139880
rect 263888 139868 263894 139920
rect 254170 139840 254176 139852
rect 250876 139812 254176 139840
rect 254170 139800 254176 139812
rect 254228 139800 254234 139852
rect 247638 139732 247644 139784
rect 247696 139772 247702 139784
rect 250858 139772 250864 139784
rect 247696 139744 250864 139772
rect 247696 139732 247702 139744
rect 250858 139732 250864 139744
rect 250916 139732 250922 139784
rect 250953 139775 251011 139781
rect 250953 139741 250965 139775
rect 250999 139772 251011 139775
rect 254446 139772 254452 139784
rect 250999 139744 254452 139772
rect 250999 139741 251011 139744
rect 250953 139735 251011 139741
rect 254446 139732 254452 139744
rect 254504 139732 254510 139784
rect 249662 139664 249668 139716
rect 249720 139704 249726 139716
rect 249720 139676 255688 139704
rect 249720 139664 249726 139676
rect 244878 139596 244884 139648
rect 244936 139636 244942 139648
rect 249386 139636 249392 139648
rect 244936 139608 249392 139636
rect 244936 139596 244942 139608
rect 249386 139596 249392 139608
rect 249444 139596 249450 139648
rect 250030 139596 250036 139648
rect 250088 139636 250094 139648
rect 251962 139636 251968 139648
rect 250088 139608 251968 139636
rect 250088 139596 250094 139608
rect 251962 139596 251968 139608
rect 252020 139596 252026 139648
rect 252057 139639 252115 139645
rect 252057 139605 252069 139639
rect 252103 139636 252115 139639
rect 255550 139636 255556 139648
rect 252103 139608 255556 139636
rect 252103 139605 252115 139608
rect 252057 139599 252115 139605
rect 255550 139596 255556 139608
rect 255608 139596 255614 139648
rect 255660 139636 255688 139676
rect 260426 139636 260432 139648
rect 255660 139608 260432 139636
rect 260426 139596 260432 139608
rect 260484 139596 260490 139648
rect 243096 139540 244740 139568
rect 243096 139528 243102 139540
rect 245798 139528 245804 139580
rect 245856 139568 245862 139580
rect 249110 139568 249116 139580
rect 245856 139540 249116 139568
rect 245856 139528 245862 139540
rect 249110 139528 249116 139540
rect 249168 139528 249174 139580
rect 249202 139528 249208 139580
rect 249260 139568 249266 139580
rect 250674 139568 250680 139580
rect 249260 139540 250680 139568
rect 249260 139528 249266 139540
rect 250674 139528 250680 139540
rect 250732 139528 250738 139580
rect 251870 139528 251876 139580
rect 251928 139568 251934 139580
rect 252698 139568 252704 139580
rect 251928 139540 252704 139568
rect 251928 139528 251934 139540
rect 252698 139528 252704 139540
rect 252756 139528 252762 139580
rect 58486 139460 58492 139512
rect 58544 139500 58550 139512
rect 60602 139500 60608 139512
rect 58544 139472 60608 139500
rect 58544 139460 58550 139472
rect 60602 139460 60608 139472
rect 60660 139460 60666 139512
rect 60694 139460 60700 139512
rect 60752 139500 60758 139512
rect 72470 139500 72476 139512
rect 60752 139472 72476 139500
rect 60752 139460 60758 139472
rect 72470 139460 72476 139472
rect 72528 139460 72534 139512
rect 149106 139460 149112 139512
rect 149164 139500 149170 139512
rect 157570 139500 157576 139512
rect 149164 139472 157576 139500
rect 149164 139460 149170 139472
rect 157570 139460 157576 139472
rect 157628 139460 157634 139512
rect 157665 139503 157723 139509
rect 157665 139469 157677 139503
rect 157711 139500 157723 139503
rect 160514 139500 160520 139512
rect 157711 139472 160520 139500
rect 157711 139469 157723 139472
rect 157665 139463 157723 139469
rect 160514 139460 160520 139472
rect 160572 139460 160578 139512
rect 242210 139460 242216 139512
rect 242268 139500 242274 139512
rect 247914 139500 247920 139512
rect 242268 139472 247920 139500
rect 242268 139460 242274 139472
rect 247914 139460 247920 139472
rect 247972 139460 247978 139512
rect 251042 139500 251048 139512
rect 248024 139472 251048 139500
rect 59130 139392 59136 139444
rect 59188 139432 59194 139444
rect 60418 139432 60424 139444
rect 59188 139404 60424 139432
rect 59188 139392 59194 139404
rect 60418 139392 60424 139404
rect 60476 139392 60482 139444
rect 63178 139432 63184 139444
rect 60528 139404 63184 139432
rect 59038 139324 59044 139376
rect 59096 139364 59102 139376
rect 60528 139364 60556 139404
rect 63178 139392 63184 139404
rect 63236 139392 63242 139444
rect 63638 139392 63644 139444
rect 63696 139432 63702 139444
rect 75782 139432 75788 139444
rect 63696 139404 75788 139432
rect 63696 139392 63702 139404
rect 75782 139392 75788 139404
rect 75840 139392 75846 139444
rect 153246 139392 153252 139444
rect 153304 139432 153310 139444
rect 156101 139435 156159 139441
rect 153304 139404 156052 139432
rect 153304 139392 153310 139404
rect 59096 139336 60556 139364
rect 59096 139324 59102 139336
rect 60786 139324 60792 139376
rect 60844 139364 60850 139376
rect 73114 139364 73120 139376
rect 60844 139336 73120 139364
rect 60844 139324 60850 139336
rect 73114 139324 73120 139336
rect 73172 139324 73178 139376
rect 137974 139324 137980 139376
rect 138032 139364 138038 139376
rect 145150 139364 145156 139376
rect 138032 139336 145156 139364
rect 138032 139324 138038 139336
rect 145150 139324 145156 139336
rect 145208 139324 145214 139376
rect 155178 139324 155184 139376
rect 155236 139364 155242 139376
rect 155914 139364 155920 139376
rect 155236 139336 155920 139364
rect 155236 139324 155242 139336
rect 155914 139324 155920 139336
rect 155972 139324 155978 139376
rect 156024 139364 156052 139404
rect 156101 139401 156113 139435
rect 156147 139432 156159 139435
rect 166862 139432 166868 139444
rect 156147 139404 166868 139432
rect 156147 139401 156159 139404
rect 156101 139395 156159 139401
rect 166862 139392 166868 139404
rect 166920 139392 166926 139444
rect 244605 139435 244663 139441
rect 244605 139401 244617 139435
rect 244651 139432 244663 139435
rect 248024 139432 248052 139472
rect 251042 139460 251048 139472
rect 251100 139460 251106 139512
rect 251318 139460 251324 139512
rect 251376 139500 251382 139512
rect 261438 139500 261444 139512
rect 251376 139472 261444 139500
rect 251376 139460 251382 139472
rect 261438 139460 261444 139472
rect 261496 139460 261502 139512
rect 250033 139435 250091 139441
rect 250033 139432 250045 139435
rect 244651 139404 248052 139432
rect 248116 139404 250045 139432
rect 244651 139401 244663 139404
rect 244605 139395 244663 139401
rect 163642 139364 163648 139376
rect 156024 139336 163648 139364
rect 163642 139324 163648 139336
rect 163700 139324 163706 139376
rect 245338 139324 245344 139376
rect 245396 139364 245402 139376
rect 248116 139364 248144 139404
rect 250033 139401 250045 139404
rect 250079 139401 250091 139435
rect 250033 139395 250091 139401
rect 250122 139392 250128 139444
rect 250180 139432 250186 139444
rect 253434 139432 253440 139444
rect 250180 139404 253440 139432
rect 250180 139392 250186 139404
rect 253434 139392 253440 139404
rect 253492 139392 253498 139444
rect 253529 139435 253587 139441
rect 253529 139401 253541 139435
rect 253575 139432 253587 139435
rect 259874 139432 259880 139444
rect 253575 139404 259880 139432
rect 253575 139401 253587 139404
rect 253529 139395 253587 139401
rect 259874 139392 259880 139404
rect 259932 139392 259938 139444
rect 245396 139336 248144 139364
rect 245396 139324 245402 139336
rect 249754 139324 249760 139376
rect 249812 139364 249818 139376
rect 252146 139364 252152 139376
rect 249812 139336 252152 139364
rect 249812 139324 249818 139336
rect 252146 139324 252152 139336
rect 252204 139324 252210 139376
rect 252241 139367 252299 139373
rect 252241 139333 252253 139367
rect 252287 139364 252299 139367
rect 258770 139364 258776 139376
rect 252287 139336 258776 139364
rect 252287 139333 252299 139336
rect 252241 139327 252299 139333
rect 258770 139324 258776 139336
rect 258828 139324 258834 139376
rect 55174 139256 55180 139308
rect 55232 139296 55238 139308
rect 57474 139296 57480 139308
rect 55232 139268 57480 139296
rect 55232 139256 55238 139268
rect 57474 139256 57480 139268
rect 57532 139256 57538 139308
rect 59774 139256 59780 139308
rect 59832 139296 59838 139308
rect 60878 139296 60884 139308
rect 59832 139268 60884 139296
rect 59832 139256 59838 139268
rect 60878 139256 60884 139268
rect 60936 139256 60942 139308
rect 61338 139256 61344 139308
rect 61396 139296 61402 139308
rect 74494 139296 74500 139308
rect 61396 139268 74500 139296
rect 61396 139256 61402 139268
rect 74494 139256 74500 139268
rect 74552 139256 74558 139308
rect 138986 139256 138992 139308
rect 139044 139296 139050 139308
rect 146254 139296 146260 139308
rect 139044 139268 146260 139296
rect 139044 139256 139050 139268
rect 146254 139256 146260 139268
rect 146312 139256 146318 139308
rect 158858 139296 158864 139308
rect 152804 139268 158864 139296
rect 38246 139188 38252 139240
rect 38304 139228 38310 139240
rect 49194 139228 49200 139240
rect 38304 139200 49200 139228
rect 38304 139188 38310 139200
rect 49194 139188 49200 139200
rect 49252 139188 49258 139240
rect 53150 139188 53156 139240
rect 53208 139228 53214 139240
rect 61798 139228 61804 139240
rect 53208 139200 61804 139228
rect 53208 139188 53214 139200
rect 61798 139188 61804 139200
rect 61856 139188 61862 139240
rect 66490 139228 66496 139240
rect 61908 139200 66496 139228
rect 60142 139120 60148 139172
rect 60200 139160 60206 139172
rect 60973 139163 61031 139169
rect 60973 139160 60985 139163
rect 60200 139132 60985 139160
rect 60200 139120 60206 139132
rect 60973 139129 60985 139132
rect 61019 139129 61031 139163
rect 60973 139123 61031 139129
rect 61157 139163 61215 139169
rect 61157 139129 61169 139163
rect 61203 139160 61215 139163
rect 61908 139160 61936 139200
rect 66490 139188 66496 139200
rect 66548 139188 66554 139240
rect 67134 139188 67140 139240
rect 67192 139228 67198 139240
rect 69802 139228 69808 139240
rect 67192 139200 69808 139228
rect 67192 139188 67198 139200
rect 69802 139188 69808 139200
rect 69860 139188 69866 139240
rect 69897 139231 69955 139237
rect 69897 139197 69909 139231
rect 69943 139228 69955 139231
rect 75138 139228 75144 139240
rect 69943 139200 75144 139228
rect 69943 139197 69955 139200
rect 69897 139191 69955 139197
rect 75138 139188 75144 139200
rect 75196 139188 75202 139240
rect 137882 139188 137888 139240
rect 137940 139228 137946 139240
rect 145702 139228 145708 139240
rect 137940 139200 145708 139228
rect 137940 139188 137946 139200
rect 145702 139188 145708 139200
rect 145760 139188 145766 139240
rect 61203 139132 61936 139160
rect 61203 139129 61215 139132
rect 61157 139123 61215 139129
rect 60234 139052 60240 139104
rect 60292 139092 60298 139104
rect 61065 139095 61123 139101
rect 61065 139092 61077 139095
rect 60292 139064 61077 139092
rect 60292 139052 60298 139064
rect 61065 139061 61077 139064
rect 61111 139061 61123 139095
rect 61065 139055 61123 139061
rect 61246 139052 61252 139104
rect 61304 139092 61310 139104
rect 65478 139092 65484 139104
rect 61304 139064 65484 139092
rect 61304 139052 61310 139064
rect 65478 139052 65484 139064
rect 65536 139052 65542 139104
rect 149934 139052 149940 139104
rect 149992 139092 149998 139104
rect 152804 139092 152832 139268
rect 158858 139256 158864 139268
rect 158916 139256 158922 139308
rect 158953 139299 159011 139305
rect 158953 139265 158965 139299
rect 158999 139296 159011 139299
rect 163090 139296 163096 139308
rect 158999 139268 163096 139296
rect 158999 139265 159011 139268
rect 158953 139259 159011 139265
rect 163090 139256 163096 139268
rect 163148 139256 163154 139308
rect 231814 139256 231820 139308
rect 231872 139296 231878 139308
rect 238990 139296 238996 139308
rect 231872 139268 238996 139296
rect 231872 139256 231878 139268
rect 238990 139256 238996 139268
rect 239048 139256 239054 139308
rect 245430 139256 245436 139308
rect 245488 139296 245494 139308
rect 249294 139296 249300 139308
rect 245488 139268 249300 139296
rect 245488 139256 245494 139268
rect 249294 139256 249300 139268
rect 249352 139256 249358 139308
rect 250401 139299 250459 139305
rect 250401 139296 250413 139299
rect 249404 139268 250413 139296
rect 154166 139188 154172 139240
rect 154224 139228 154230 139240
rect 155546 139228 155552 139240
rect 154224 139200 155552 139228
rect 154224 139188 154230 139200
rect 155546 139188 155552 139200
rect 155604 139188 155610 139240
rect 155822 139188 155828 139240
rect 155880 139228 155886 139240
rect 167322 139228 167328 139240
rect 155880 139200 167328 139228
rect 155880 139188 155886 139200
rect 167322 139188 167328 139200
rect 167380 139188 167386 139240
rect 231722 139188 231728 139240
rect 231780 139228 231786 139240
rect 239450 139228 239456 139240
rect 231780 139200 239456 139228
rect 231780 139188 231786 139200
rect 239450 139188 239456 139200
rect 239508 139188 239514 139240
rect 245706 139188 245712 139240
rect 245764 139228 245770 139240
rect 249404 139228 249432 139268
rect 250401 139265 250413 139268
rect 250447 139265 250459 139299
rect 250401 139259 250459 139265
rect 250490 139256 250496 139308
rect 250548 139296 250554 139308
rect 259322 139296 259328 139308
rect 250548 139268 259328 139296
rect 250548 139256 250554 139268
rect 259322 139256 259328 139268
rect 259380 139256 259386 139308
rect 245764 139200 249432 139228
rect 245764 139188 245770 139200
rect 249570 139188 249576 139240
rect 249628 139228 249634 139240
rect 256930 139228 256936 139240
rect 249628 139200 256936 139228
rect 249628 139188 249634 139200
rect 256930 139188 256936 139200
rect 256988 139188 256994 139240
rect 261162 139228 261168 139240
rect 257040 139200 261168 139228
rect 155362 139120 155368 139172
rect 155420 139160 155426 139172
rect 159410 139160 159416 139172
rect 155420 139132 159416 139160
rect 155420 139120 155426 139132
rect 159410 139120 159416 139132
rect 159468 139120 159474 139172
rect 248926 139120 248932 139172
rect 248984 139160 248990 139172
rect 253529 139163 253587 139169
rect 253529 139160 253541 139163
rect 248984 139132 253541 139160
rect 248984 139120 248990 139132
rect 253529 139129 253541 139132
rect 253575 139129 253587 139163
rect 253529 139123 253587 139129
rect 253621 139163 253679 139169
rect 253621 139129 253633 139163
rect 253667 139160 253679 139163
rect 254998 139160 255004 139172
rect 253667 139132 255004 139160
rect 253667 139129 253679 139132
rect 253621 139123 253679 139129
rect 254998 139120 255004 139132
rect 255056 139120 255062 139172
rect 149992 139064 152832 139092
rect 149992 139052 149998 139064
rect 154718 139052 154724 139104
rect 154776 139092 154782 139104
rect 155454 139092 155460 139104
rect 154776 139064 155460 139092
rect 154776 139052 154782 139064
rect 155454 139052 155460 139064
rect 155512 139052 155518 139104
rect 155730 139052 155736 139104
rect 155788 139092 155794 139104
rect 159962 139092 159968 139104
rect 155788 139064 159968 139092
rect 155788 139052 155794 139064
rect 159962 139052 159968 139064
rect 160020 139052 160026 139104
rect 249846 139052 249852 139104
rect 249904 139092 249910 139104
rect 257040 139092 257068 139200
rect 261162 139188 261168 139200
rect 261220 139188 261226 139240
rect 249904 139064 257068 139092
rect 249904 139052 249910 139064
rect 55818 138984 55824 139036
rect 55876 139024 55882 139036
rect 58854 139024 58860 139036
rect 55876 138996 58860 139024
rect 55876 138984 55882 138996
rect 58854 138984 58860 138996
rect 58912 138984 58918 139036
rect 59498 138984 59504 139036
rect 59556 139024 59562 139036
rect 61341 139027 61399 139033
rect 61341 139024 61353 139027
rect 59556 138996 61353 139024
rect 59556 138984 59562 138996
rect 61341 138993 61353 138996
rect 61387 138993 61399 139027
rect 61341 138987 61399 138993
rect 61430 138984 61436 139036
rect 61488 139024 61494 139036
rect 70541 139027 70599 139033
rect 70541 139024 70553 139027
rect 61488 138996 70553 139024
rect 61488 138984 61494 138996
rect 70541 138993 70553 138996
rect 70587 138993 70599 139027
rect 70541 138987 70599 138993
rect 152694 138984 152700 139036
rect 152752 139024 152758 139036
rect 152752 138996 154856 139024
rect 152752 138984 152758 138996
rect 60326 138916 60332 138968
rect 60384 138956 60390 138968
rect 61157 138959 61215 138965
rect 61157 138956 61169 138959
rect 60384 138928 61169 138956
rect 60384 138916 60390 138928
rect 61157 138925 61169 138928
rect 61203 138925 61215 138959
rect 61157 138919 61215 138925
rect 61522 138916 61528 138968
rect 61580 138956 61586 138968
rect 64466 138956 64472 138968
rect 61580 138928 64472 138956
rect 61580 138916 61586 138928
rect 64466 138916 64472 138928
rect 64524 138916 64530 138968
rect 153614 138916 153620 138968
rect 153672 138956 153678 138968
rect 154718 138956 154724 138968
rect 153672 138928 154724 138956
rect 153672 138916 153678 138928
rect 154718 138916 154724 138928
rect 154776 138916 154782 138968
rect 154828 138956 154856 138996
rect 156006 138984 156012 139036
rect 156064 139024 156070 139036
rect 156101 139027 156159 139033
rect 156101 139024 156113 139027
rect 156064 138996 156113 139024
rect 156064 138984 156070 138996
rect 156101 138993 156113 138996
rect 156147 138993 156159 139027
rect 156101 138987 156159 138993
rect 156742 138984 156748 139036
rect 156800 139024 156806 139036
rect 165206 139024 165212 139036
rect 156800 138996 165212 139024
rect 156800 138984 156806 138996
rect 165206 138984 165212 138996
rect 165264 138984 165270 139036
rect 246534 138984 246540 139036
rect 246592 139024 246598 139036
rect 249478 139024 249484 139036
rect 246592 138996 249484 139024
rect 246592 138984 246598 138996
rect 249478 138984 249484 138996
rect 249536 138984 249542 139036
rect 250214 138984 250220 139036
rect 250272 139024 250278 139036
rect 252882 139024 252888 139036
rect 250272 138996 252888 139024
rect 250272 138984 250278 138996
rect 252882 138984 252888 138996
rect 252940 138984 252946 139036
rect 156837 138959 156895 138965
rect 156837 138956 156849 138959
rect 154828 138928 156849 138956
rect 156837 138925 156849 138928
rect 156883 138925 156895 138959
rect 156837 138919 156895 138925
rect 156926 138916 156932 138968
rect 156984 138956 156990 138968
rect 164746 138956 164752 138968
rect 156984 138928 164752 138956
rect 156984 138916 156990 138928
rect 164746 138916 164752 138928
rect 164804 138916 164810 138968
rect 243866 138916 243872 138968
rect 243924 138956 243930 138968
rect 249018 138956 249024 138968
rect 243924 138928 249024 138956
rect 243924 138916 243930 138928
rect 249018 138916 249024 138928
rect 249076 138916 249082 138968
rect 253621 138959 253679 138965
rect 253621 138956 253633 138959
rect 249128 138928 253633 138956
rect 57842 138848 57848 138900
rect 57900 138888 57906 138900
rect 61890 138888 61896 138900
rect 57900 138860 61896 138888
rect 57900 138848 57906 138860
rect 61890 138848 61896 138860
rect 61948 138848 61954 138900
rect 61985 138891 62043 138897
rect 61985 138857 61997 138891
rect 62031 138888 62043 138891
rect 69158 138888 69164 138900
rect 62031 138860 69164 138888
rect 62031 138857 62043 138860
rect 61985 138851 62043 138857
rect 69158 138848 69164 138860
rect 69216 138848 69222 138900
rect 151038 138848 151044 138900
rect 151096 138888 151102 138900
rect 157570 138888 157576 138900
rect 151096 138860 157576 138888
rect 151096 138848 151102 138860
rect 157570 138848 157576 138860
rect 157628 138848 157634 138900
rect 158398 138848 158404 138900
rect 158456 138888 158462 138900
rect 161066 138888 161072 138900
rect 158456 138860 161072 138888
rect 158456 138848 158462 138860
rect 161066 138848 161072 138860
rect 161124 138848 161130 138900
rect 231354 138848 231360 138900
rect 231412 138888 231418 138900
rect 237242 138888 237248 138900
rect 231412 138860 237248 138888
rect 231412 138848 231418 138860
rect 237242 138848 237248 138860
rect 237300 138848 237306 138900
rect 245614 138848 245620 138900
rect 245672 138888 245678 138900
rect 249128 138888 249156 138928
rect 253621 138925 253633 138928
rect 253667 138925 253679 138959
rect 253621 138919 253679 138925
rect 245672 138860 249156 138888
rect 245672 138848 245678 138860
rect 249202 138848 249208 138900
rect 249260 138888 249266 138900
rect 256102 138888 256108 138900
rect 249260 138860 256108 138888
rect 249260 138848 249266 138860
rect 256102 138848 256108 138860
rect 256160 138848 256166 138900
rect 61065 138823 61123 138829
rect 61065 138789 61077 138823
rect 61111 138820 61123 138823
rect 67778 138820 67784 138832
rect 61111 138792 67784 138820
rect 61111 138789 61123 138792
rect 61065 138783 61123 138789
rect 67778 138780 67784 138792
rect 67836 138780 67842 138832
rect 137790 138780 137796 138832
rect 137848 138820 137854 138832
rect 144690 138820 144696 138832
rect 137848 138792 144696 138820
rect 137848 138780 137854 138792
rect 144690 138780 144696 138792
rect 144748 138780 144754 138832
rect 151498 138780 151504 138832
rect 151556 138820 151562 138832
rect 158214 138820 158220 138832
rect 151556 138792 158220 138820
rect 151556 138780 151562 138792
rect 158214 138780 158220 138792
rect 158272 138780 158278 138832
rect 158306 138780 158312 138832
rect 158364 138820 158370 138832
rect 161526 138820 161532 138832
rect 158364 138792 161532 138820
rect 158364 138780 158370 138792
rect 161526 138780 161532 138792
rect 161584 138780 161590 138832
rect 164194 138820 164200 138832
rect 162924 138792 164200 138820
rect 60973 138755 61031 138761
rect 60973 138721 60985 138755
rect 61019 138752 61031 138755
rect 68422 138752 68428 138764
rect 61019 138724 68428 138752
rect 61019 138721 61031 138724
rect 60973 138715 61031 138721
rect 68422 138712 68428 138724
rect 68480 138712 68486 138764
rect 137698 138712 137704 138764
rect 137756 138752 137762 138764
rect 144138 138752 144144 138764
rect 137756 138724 144144 138752
rect 137756 138712 137762 138724
rect 144138 138712 144144 138724
rect 144196 138712 144202 138764
rect 147818 138712 147824 138764
rect 147876 138752 147882 138764
rect 154258 138752 154264 138764
rect 147876 138724 154264 138752
rect 147876 138712 147882 138724
rect 154258 138712 154264 138724
rect 154316 138712 154322 138764
rect 155638 138712 155644 138764
rect 155696 138752 155702 138764
rect 158950 138752 158956 138764
rect 155696 138724 158956 138752
rect 155696 138712 155702 138724
rect 158950 138712 158956 138724
rect 159008 138712 159014 138764
rect 161066 138712 161072 138764
rect 161124 138752 161130 138764
rect 162924 138752 162952 138792
rect 164194 138780 164200 138792
rect 164252 138780 164258 138832
rect 231630 138780 231636 138832
rect 231688 138820 231694 138832
rect 238346 138820 238352 138832
rect 231688 138792 238352 138820
rect 231688 138780 231694 138792
rect 238346 138780 238352 138792
rect 238404 138780 238410 138832
rect 248374 138780 248380 138832
rect 248432 138820 248438 138832
rect 252241 138823 252299 138829
rect 252241 138820 252253 138823
rect 248432 138792 252253 138820
rect 248432 138780 248438 138792
rect 252241 138789 252253 138792
rect 252287 138789 252299 138823
rect 252241 138783 252299 138789
rect 254814 138780 254820 138832
rect 254872 138820 254878 138832
rect 258310 138820 258316 138832
rect 254872 138792 258316 138820
rect 254872 138780 254878 138792
rect 258310 138780 258316 138792
rect 258368 138780 258374 138832
rect 161124 138724 162952 138752
rect 161124 138712 161130 138724
rect 163734 138712 163740 138764
rect 163792 138752 163798 138764
rect 167874 138752 167880 138764
rect 163792 138724 167880 138752
rect 163792 138712 163798 138724
rect 167874 138712 167880 138724
rect 167932 138712 167938 138764
rect 231538 138712 231544 138764
rect 231596 138752 231602 138764
rect 237794 138752 237800 138764
rect 231596 138724 237800 138752
rect 231596 138712 231602 138724
rect 237794 138712 237800 138724
rect 237852 138712 237858 138764
rect 250398 138712 250404 138764
rect 250456 138752 250462 138764
rect 250456 138724 257896 138752
rect 250456 138712 250462 138724
rect 61249 138687 61307 138693
rect 61249 138653 61261 138687
rect 61295 138684 61307 138687
rect 66674 138684 66680 138696
rect 61295 138656 66680 138684
rect 61295 138653 61307 138656
rect 61249 138647 61307 138653
rect 66674 138644 66680 138656
rect 66732 138644 66738 138696
rect 137606 138644 137612 138696
rect 137664 138684 137670 138696
rect 143586 138684 143592 138696
rect 137664 138656 143592 138684
rect 137664 138644 137670 138656
rect 143586 138644 143592 138656
rect 143644 138644 143650 138696
rect 147266 138644 147272 138696
rect 147324 138684 147330 138696
rect 154074 138684 154080 138696
rect 147324 138656 154080 138684
rect 147324 138644 147330 138656
rect 154074 138644 154080 138656
rect 154132 138644 154138 138696
rect 154184 138656 155684 138684
rect 60970 138576 60976 138628
rect 61028 138616 61034 138628
rect 62994 138616 63000 138628
rect 61028 138588 63000 138616
rect 61028 138576 61034 138588
rect 62994 138576 63000 138588
rect 63052 138576 63058 138628
rect 69897 138619 69955 138625
rect 69897 138616 69909 138619
rect 63104 138588 69909 138616
rect 62258 138508 62264 138560
rect 62316 138548 62322 138560
rect 63104 138548 63132 138588
rect 69897 138585 69909 138588
rect 69943 138585 69955 138619
rect 69897 138579 69955 138585
rect 137514 138576 137520 138628
rect 137572 138616 137578 138628
rect 142758 138616 142764 138628
rect 137572 138588 142764 138616
rect 137572 138576 137578 138588
rect 142758 138576 142764 138588
rect 142816 138576 142822 138628
rect 148370 138576 148376 138628
rect 148428 138616 148434 138628
rect 149014 138616 149020 138628
rect 148428 138588 149020 138616
rect 148428 138576 148434 138588
rect 149014 138576 149020 138588
rect 149072 138576 149078 138628
rect 152050 138576 152056 138628
rect 152108 138616 152114 138628
rect 153154 138616 153160 138628
rect 152108 138588 153160 138616
rect 152108 138576 152114 138588
rect 153154 138576 153160 138588
rect 153212 138576 153218 138628
rect 154184 138616 154212 138656
rect 153264 138588 154212 138616
rect 155656 138616 155684 138656
rect 156282 138644 156288 138696
rect 156340 138684 156346 138696
rect 157478 138684 157484 138696
rect 156340 138656 157484 138684
rect 156340 138644 156346 138656
rect 157478 138644 157484 138656
rect 157536 138644 157542 138696
rect 157570 138644 157576 138696
rect 157628 138684 157634 138696
rect 158490 138684 158496 138696
rect 157628 138656 158496 138684
rect 157628 138644 157634 138656
rect 158490 138644 158496 138656
rect 158548 138644 158554 138696
rect 160974 138644 160980 138696
rect 161032 138684 161038 138696
rect 162630 138684 162636 138696
rect 161032 138656 162636 138684
rect 161032 138644 161038 138656
rect 162630 138644 162636 138656
rect 162688 138644 162694 138696
rect 231446 138644 231452 138696
rect 231504 138684 231510 138696
rect 236782 138684 236788 138696
rect 231504 138656 236788 138684
rect 231504 138644 231510 138656
rect 236782 138644 236788 138656
rect 236840 138644 236846 138696
rect 244418 138644 244424 138696
rect 244476 138684 244482 138696
rect 246534 138684 246540 138696
rect 244476 138656 246540 138684
rect 244476 138644 244482 138656
rect 246534 138644 246540 138656
rect 246592 138644 246598 138696
rect 247086 138644 247092 138696
rect 247144 138684 247150 138696
rect 253434 138684 253440 138696
rect 247144 138656 253440 138684
rect 247144 138644 247150 138656
rect 253434 138644 253440 138656
rect 253492 138644 253498 138696
rect 254906 138644 254912 138696
rect 254964 138684 254970 138696
rect 257758 138684 257764 138696
rect 254964 138656 257764 138684
rect 254964 138644 254970 138656
rect 257758 138644 257764 138656
rect 257816 138644 257822 138696
rect 155656 138588 156788 138616
rect 62316 138520 63132 138548
rect 62316 138508 62322 138520
rect 152878 138508 152884 138560
rect 152936 138548 152942 138560
rect 153264 138548 153292 138588
rect 152936 138520 153292 138548
rect 156760 138548 156788 138588
rect 156834 138576 156840 138628
rect 156892 138616 156898 138628
rect 157294 138616 157300 138628
rect 156892 138588 157300 138616
rect 156892 138576 156898 138588
rect 157294 138576 157300 138588
rect 157352 138576 157358 138628
rect 158953 138619 159011 138625
rect 158953 138616 158965 138619
rect 157404 138588 158965 138616
rect 157404 138548 157432 138588
rect 158953 138585 158965 138588
rect 158999 138585 159011 138619
rect 158953 138579 159011 138585
rect 161158 138576 161164 138628
rect 161216 138616 161222 138628
rect 162078 138616 162084 138628
rect 161216 138588 162084 138616
rect 161216 138576 161222 138588
rect 162078 138576 162084 138588
rect 162136 138576 162142 138628
rect 167874 138576 167880 138628
rect 167932 138616 167938 138628
rect 170818 138616 170824 138628
rect 167932 138588 170824 138616
rect 167932 138576 167938 138588
rect 170818 138576 170824 138588
rect 170876 138576 170882 138628
rect 232918 138576 232924 138628
rect 232976 138616 232982 138628
rect 240002 138616 240008 138628
rect 232976 138588 240008 138616
rect 232976 138576 232982 138588
rect 240002 138576 240008 138588
rect 240060 138576 240066 138628
rect 245798 138576 245804 138628
rect 245856 138616 245862 138628
rect 252057 138619 252115 138625
rect 252057 138616 252069 138619
rect 245856 138588 252069 138616
rect 245856 138576 245862 138588
rect 252057 138585 252069 138588
rect 252103 138585 252115 138619
rect 252057 138579 252115 138585
rect 254998 138576 255004 138628
rect 255056 138616 255062 138628
rect 257206 138616 257212 138628
rect 255056 138588 257212 138616
rect 255056 138576 255062 138588
rect 257206 138576 257212 138588
rect 257264 138576 257270 138628
rect 257868 138616 257896 138724
rect 261990 138616 261996 138628
rect 257868 138588 261996 138616
rect 261990 138576 261996 138588
rect 262048 138576 262054 138628
rect 263186 138576 263192 138628
rect 263244 138616 263250 138628
rect 263738 138616 263744 138628
rect 263244 138588 263744 138616
rect 263244 138576 263250 138588
rect 263738 138576 263744 138588
rect 263796 138576 263802 138628
rect 156760 138520 157432 138548
rect 152936 138508 152942 138520
rect 126474 135788 126480 135840
rect 126532 135828 126538 135840
rect 159594 135828 159600 135840
rect 126532 135800 159600 135828
rect 126532 135788 126538 135800
rect 159594 135788 159600 135800
rect 159652 135788 159658 135840
rect 220498 135788 220504 135840
rect 220556 135828 220562 135840
rect 255458 135828 255464 135840
rect 220556 135800 255464 135828
rect 220556 135788 220562 135800
rect 255458 135788 255464 135800
rect 255516 135788 255522 135840
rect 136870 132932 136876 132984
rect 136928 132972 136934 132984
rect 146806 132972 146812 132984
rect 136928 132944 146812 132972
rect 136928 132932 136934 132944
rect 146806 132932 146812 132944
rect 146864 132932 146870 132984
rect 231906 132932 231912 132984
rect 231964 132972 231970 132984
rect 240554 132972 240560 132984
rect 231964 132944 240560 132972
rect 231964 132932 231970 132944
rect 240554 132932 240560 132944
rect 240612 132932 240618 132984
rect 249389 131751 249447 131757
rect 249389 131717 249401 131751
rect 249435 131748 249447 131751
rect 250030 131748 250036 131760
rect 249435 131720 250036 131748
rect 249435 131717 249447 131720
rect 249389 131711 249447 131717
rect 250030 131708 250036 131720
rect 250088 131708 250094 131760
rect 148922 131640 148928 131692
rect 148980 131680 148986 131692
rect 149198 131680 149204 131692
rect 148980 131652 149204 131680
rect 148980 131640 148986 131652
rect 149198 131640 149204 131652
rect 149256 131640 149262 131692
rect 157849 131683 157907 131689
rect 157849 131680 157861 131683
rect 155472 131652 157861 131680
rect 155472 131624 155500 131652
rect 157849 131649 157861 131652
rect 157895 131649 157907 131683
rect 252149 131683 252207 131689
rect 252149 131680 252161 131683
rect 157849 131643 157907 131649
rect 248484 131652 252161 131680
rect 56186 131572 56192 131624
rect 56244 131612 56250 131624
rect 56738 131612 56744 131624
rect 56244 131584 56744 131612
rect 56244 131572 56250 131584
rect 56738 131572 56744 131584
rect 56796 131572 56802 131624
rect 57382 131572 57388 131624
rect 57440 131612 57446 131624
rect 60050 131612 60056 131624
rect 57440 131584 60056 131612
rect 57440 131572 57446 131584
rect 60050 131572 60056 131584
rect 60108 131572 60114 131624
rect 60418 131572 60424 131624
rect 60476 131612 60482 131624
rect 68330 131612 68336 131624
rect 60476 131584 68336 131612
rect 60476 131572 60482 131584
rect 68330 131572 68336 131584
rect 68388 131572 68394 131624
rect 150210 131572 150216 131624
rect 150268 131612 150274 131624
rect 155362 131612 155368 131624
rect 150268 131584 155368 131612
rect 150268 131572 150274 131584
rect 155362 131572 155368 131584
rect 155420 131572 155426 131624
rect 155454 131572 155460 131624
rect 155512 131572 155518 131624
rect 157294 131572 157300 131624
rect 157352 131612 157358 131624
rect 163918 131612 163924 131624
rect 157352 131584 163924 131612
rect 157352 131572 157358 131584
rect 163918 131572 163924 131584
rect 163976 131572 163982 131624
rect 244878 131572 244884 131624
rect 244936 131612 244942 131624
rect 245338 131612 245344 131624
rect 244936 131584 245344 131612
rect 244936 131572 244942 131584
rect 245338 131572 245344 131584
rect 245396 131572 245402 131624
rect 248006 131572 248012 131624
rect 248064 131612 248070 131624
rect 248484 131612 248512 131652
rect 252149 131649 252161 131652
rect 252195 131649 252207 131683
rect 252149 131643 252207 131649
rect 248064 131584 248512 131612
rect 248064 131572 248070 131584
rect 248558 131572 248564 131624
rect 248616 131612 248622 131624
rect 250490 131612 250496 131624
rect 248616 131584 250496 131612
rect 248616 131572 248622 131584
rect 250490 131572 250496 131584
rect 250548 131572 250554 131624
rect 254262 131612 254268 131624
rect 250600 131584 254268 131612
rect 55082 131504 55088 131556
rect 55140 131544 55146 131556
rect 59038 131544 59044 131556
rect 55140 131516 59044 131544
rect 55140 131504 55146 131516
rect 59038 131504 59044 131516
rect 59096 131504 59102 131556
rect 65570 131544 65576 131556
rect 59148 131516 65576 131544
rect 57566 131436 57572 131488
rect 57624 131476 57630 131488
rect 59148 131476 59176 131516
rect 65570 131504 65576 131516
rect 65628 131504 65634 131556
rect 149842 131504 149848 131556
rect 149900 131544 149906 131556
rect 155638 131544 155644 131556
rect 149900 131516 155644 131544
rect 149900 131504 149906 131516
rect 155638 131504 155644 131516
rect 155696 131504 155702 131556
rect 155733 131547 155791 131553
rect 155733 131513 155745 131547
rect 155779 131544 155791 131547
rect 157205 131547 157263 131553
rect 157205 131544 157217 131547
rect 155779 131516 157217 131544
rect 155779 131513 155791 131516
rect 155733 131507 155791 131513
rect 157205 131513 157217 131516
rect 157251 131513 157263 131547
rect 157205 131507 157263 131513
rect 157386 131504 157392 131556
rect 157444 131544 157450 131556
rect 164286 131544 164292 131556
rect 157444 131516 164292 131544
rect 157444 131504 157450 131516
rect 164286 131504 164292 131516
rect 164344 131504 164350 131556
rect 243314 131504 243320 131556
rect 243372 131544 243378 131556
rect 249389 131547 249447 131553
rect 249389 131544 249401 131547
rect 243372 131516 249401 131544
rect 243372 131504 243378 131516
rect 249389 131513 249401 131516
rect 249435 131513 249447 131547
rect 249389 131507 249447 131513
rect 249478 131504 249484 131556
rect 249536 131544 249542 131556
rect 250600 131544 250628 131584
rect 254262 131572 254268 131584
rect 254320 131572 254326 131624
rect 255458 131572 255464 131624
rect 255516 131612 255522 131624
rect 258402 131612 258408 131624
rect 255516 131584 258408 131612
rect 255516 131572 255522 131584
rect 258402 131572 258408 131584
rect 258460 131572 258466 131624
rect 249536 131516 250628 131544
rect 250769 131547 250827 131553
rect 249536 131504 249542 131516
rect 250769 131513 250781 131547
rect 250815 131544 250827 131547
rect 254998 131544 255004 131556
rect 250815 131516 255004 131544
rect 250815 131513 250827 131516
rect 250769 131507 250827 131513
rect 254998 131504 255004 131516
rect 255056 131504 255062 131556
rect 57624 131448 59176 131476
rect 57624 131436 57630 131448
rect 59682 131436 59688 131488
rect 59740 131476 59746 131488
rect 60418 131476 60424 131488
rect 59740 131448 60424 131476
rect 59740 131436 59746 131448
rect 60418 131436 60424 131448
rect 60476 131436 60482 131488
rect 65202 131476 65208 131488
rect 60620 131448 65208 131476
rect 57474 131368 57480 131420
rect 57532 131408 57538 131420
rect 60510 131408 60516 131420
rect 57532 131380 60516 131408
rect 57532 131368 57538 131380
rect 60510 131368 60516 131380
rect 60568 131368 60574 131420
rect 53978 131300 53984 131352
rect 54036 131340 54042 131352
rect 60620 131340 60648 131448
rect 65202 131436 65208 131448
rect 65260 131436 65266 131488
rect 153154 131436 153160 131488
rect 153212 131476 153218 131488
rect 160422 131476 160428 131488
rect 153212 131448 160428 131476
rect 153212 131436 153218 131448
rect 160422 131436 160428 131448
rect 160480 131436 160486 131488
rect 246353 131479 246411 131485
rect 246353 131445 246365 131479
rect 246399 131476 246411 131479
rect 250030 131476 250036 131488
rect 246399 131448 250036 131476
rect 246399 131445 246411 131448
rect 246353 131439 246411 131445
rect 250030 131436 250036 131448
rect 250088 131436 250094 131488
rect 255642 131476 255648 131488
rect 250140 131448 255648 131476
rect 60789 131411 60847 131417
rect 60789 131377 60801 131411
rect 60835 131408 60847 131411
rect 61522 131408 61528 131420
rect 60835 131380 61528 131408
rect 60835 131377 60847 131380
rect 60789 131371 60847 131377
rect 61522 131368 61528 131380
rect 61580 131368 61586 131420
rect 61614 131368 61620 131420
rect 61672 131408 61678 131420
rect 64929 131411 64987 131417
rect 64929 131408 64941 131411
rect 61672 131380 64941 131408
rect 61672 131368 61678 131380
rect 64929 131377 64941 131380
rect 64975 131377 64987 131411
rect 67226 131408 67232 131420
rect 64929 131371 64987 131377
rect 65036 131380 67232 131408
rect 54036 131312 60648 131340
rect 60697 131343 60755 131349
rect 54036 131300 54042 131312
rect 60697 131309 60709 131343
rect 60743 131340 60755 131343
rect 64374 131340 64380 131352
rect 60743 131312 64380 131340
rect 60743 131309 60755 131312
rect 60697 131303 60755 131309
rect 64374 131300 64380 131312
rect 64432 131300 64438 131352
rect 60878 131232 60884 131284
rect 60936 131272 60942 131284
rect 63362 131272 63368 131284
rect 60936 131244 63368 131272
rect 60936 131232 60942 131244
rect 63362 131232 63368 131244
rect 63420 131232 63426 131284
rect 65036 131272 65064 131380
rect 67226 131368 67232 131380
rect 67284 131368 67290 131420
rect 151038 131368 151044 131420
rect 151096 131408 151102 131420
rect 152694 131408 152700 131420
rect 151096 131380 152700 131408
rect 151096 131368 151102 131380
rect 152694 131368 152700 131380
rect 152752 131368 152758 131420
rect 152970 131368 152976 131420
rect 153028 131408 153034 131420
rect 157389 131411 157447 131417
rect 157389 131408 157401 131411
rect 153028 131380 157401 131408
rect 153028 131368 153034 131380
rect 157389 131377 157401 131380
rect 157435 131377 157447 131411
rect 157389 131371 157447 131377
rect 157478 131368 157484 131420
rect 157536 131408 157542 131420
rect 163550 131408 163556 131420
rect 157536 131380 163556 131408
rect 157536 131368 157542 131380
rect 163550 131368 163556 131380
rect 163608 131368 163614 131420
rect 248466 131368 248472 131420
rect 248524 131408 248530 131420
rect 250140 131408 250168 131448
rect 255642 131436 255648 131448
rect 255700 131436 255706 131488
rect 248524 131380 250168 131408
rect 250217 131411 250275 131417
rect 248524 131368 248530 131380
rect 250217 131377 250229 131411
rect 250263 131408 250275 131411
rect 252054 131408 252060 131420
rect 250263 131380 252060 131408
rect 250263 131377 250275 131380
rect 250217 131371 250275 131377
rect 252054 131368 252060 131380
rect 252112 131368 252118 131420
rect 252698 131368 252704 131420
rect 252756 131408 252762 131420
rect 258310 131408 258316 131420
rect 252756 131380 258316 131408
rect 252756 131368 252762 131380
rect 258310 131368 258316 131380
rect 258368 131368 258374 131420
rect 154718 131300 154724 131352
rect 154776 131340 154782 131352
rect 161526 131340 161532 131352
rect 154776 131312 161532 131340
rect 154776 131300 154782 131312
rect 161526 131300 161532 131312
rect 161584 131300 161590 131352
rect 248006 131300 248012 131352
rect 248064 131340 248070 131352
rect 254814 131340 254820 131352
rect 248064 131312 254820 131340
rect 248064 131300 248070 131312
rect 254814 131300 254820 131312
rect 254872 131300 254878 131352
rect 157662 131272 157668 131284
rect 63472 131244 65064 131272
rect 152528 131244 157668 131272
rect 52414 131164 52420 131216
rect 52472 131204 52478 131216
rect 59225 131207 59283 131213
rect 59225 131204 59237 131207
rect 52472 131176 59237 131204
rect 52472 131164 52478 131176
rect 59225 131173 59237 131176
rect 59271 131173 59283 131207
rect 59225 131167 59283 131173
rect 59314 131164 59320 131216
rect 59372 131204 59378 131216
rect 63472 131204 63500 131244
rect 59372 131176 63500 131204
rect 59372 131164 59378 131176
rect 149474 131164 149480 131216
rect 149532 131204 149538 131216
rect 152528 131204 152556 131244
rect 157662 131232 157668 131244
rect 157720 131232 157726 131284
rect 157757 131275 157815 131281
rect 157757 131241 157769 131275
rect 157803 131272 157815 131275
rect 160974 131272 160980 131284
rect 157803 131244 160980 131272
rect 157803 131241 157815 131244
rect 157757 131235 157815 131241
rect 160974 131232 160980 131244
rect 161032 131232 161038 131284
rect 175418 131232 175424 131284
rect 175476 131272 175482 131284
rect 281862 131272 281868 131284
rect 175476 131244 281868 131272
rect 175476 131232 175482 131244
rect 281862 131232 281868 131244
rect 281920 131232 281926 131284
rect 149532 131176 152556 131204
rect 149532 131164 149538 131176
rect 152602 131164 152608 131216
rect 152660 131204 152666 131216
rect 155733 131207 155791 131213
rect 155733 131204 155745 131207
rect 152660 131176 155745 131204
rect 152660 131164 152666 131176
rect 155733 131173 155745 131176
rect 155779 131173 155791 131207
rect 155733 131167 155791 131173
rect 156466 131164 156472 131216
rect 156524 131204 156530 131216
rect 163734 131204 163740 131216
rect 156524 131176 163740 131204
rect 156524 131164 156530 131176
rect 163734 131164 163740 131176
rect 163792 131164 163798 131216
rect 249386 131164 249392 131216
rect 249444 131204 249450 131216
rect 252974 131204 252980 131216
rect 249444 131176 252980 131204
rect 249444 131164 249450 131176
rect 252974 131164 252980 131176
rect 253032 131164 253038 131216
rect 51034 131096 51040 131148
rect 51092 131136 51098 131148
rect 51092 131108 51448 131136
rect 51092 131096 51098 131108
rect 51420 131068 51448 131108
rect 57014 131096 57020 131148
rect 57072 131136 57078 131148
rect 60326 131136 60332 131148
rect 57072 131108 60332 131136
rect 57072 131096 57078 131108
rect 60326 131096 60332 131108
rect 60384 131096 60390 131148
rect 60418 131096 60424 131148
rect 60476 131136 60482 131148
rect 69066 131136 69072 131148
rect 60476 131108 69072 131136
rect 60476 131096 60482 131108
rect 69066 131096 69072 131108
rect 69124 131096 69130 131148
rect 149198 131096 149204 131148
rect 149256 131136 149262 131148
rect 158030 131136 158036 131148
rect 149256 131108 158036 131136
rect 149256 131096 149262 131108
rect 158030 131096 158036 131108
rect 158088 131096 158094 131148
rect 159594 131096 159600 131148
rect 159652 131136 159658 131148
rect 164654 131136 164660 131148
rect 159652 131108 164660 131136
rect 159652 131096 159658 131108
rect 164654 131096 164660 131108
rect 164712 131096 164718 131148
rect 246534 131096 246540 131148
rect 246592 131136 246598 131148
rect 249849 131139 249907 131145
rect 249849 131136 249861 131139
rect 246592 131108 249861 131136
rect 246592 131096 246598 131108
rect 249849 131105 249861 131108
rect 249895 131105 249907 131139
rect 249849 131099 249907 131105
rect 249938 131096 249944 131148
rect 249996 131136 250002 131148
rect 256930 131136 256936 131148
rect 249996 131108 256936 131136
rect 249996 131096 250002 131108
rect 256930 131096 256936 131108
rect 256988 131096 256994 131148
rect 63270 131068 63276 131080
rect 51420 131040 63276 131068
rect 63270 131028 63276 131040
rect 63328 131028 63334 131080
rect 153706 131028 153712 131080
rect 153764 131068 153770 131080
rect 157849 131071 157907 131077
rect 153764 131040 157800 131068
rect 153764 131028 153770 131040
rect 51218 130960 51224 131012
rect 51276 131000 51282 131012
rect 58762 131000 58768 131012
rect 51276 130972 58768 131000
rect 51276 130960 51282 130972
rect 58762 130960 58768 130972
rect 58820 130960 58826 131012
rect 58854 130960 58860 131012
rect 58912 131000 58918 131012
rect 60329 131003 60387 131009
rect 60329 131000 60341 131003
rect 58912 130972 60341 131000
rect 58912 130960 58918 130972
rect 60329 130969 60341 130972
rect 60375 130969 60387 131003
rect 60329 130963 60387 130969
rect 60602 130960 60608 131012
rect 60660 131000 60666 131012
rect 67962 131000 67968 131012
rect 60660 130972 67968 131000
rect 60660 130960 60666 130972
rect 67962 130960 67968 130972
rect 68020 130960 68026 131012
rect 149014 130960 149020 131012
rect 149072 131000 149078 131012
rect 157662 131000 157668 131012
rect 149072 130972 157668 131000
rect 149072 130960 149078 130972
rect 157662 130960 157668 130972
rect 157720 130960 157726 131012
rect 157772 131000 157800 131040
rect 157849 131037 157861 131071
rect 157895 131068 157907 131071
rect 162354 131068 162360 131080
rect 157895 131040 162360 131068
rect 157895 131037 157907 131040
rect 157849 131031 157907 131037
rect 162354 131028 162360 131040
rect 162412 131028 162418 131080
rect 249018 131028 249024 131080
rect 249076 131068 249082 131080
rect 252238 131068 252244 131080
rect 249076 131040 252244 131068
rect 249076 131028 249082 131040
rect 252238 131028 252244 131040
rect 252296 131028 252302 131080
rect 161066 131000 161072 131012
rect 157772 130972 161072 131000
rect 161066 130960 161072 130972
rect 161124 130960 161130 131012
rect 245065 131003 245123 131009
rect 245065 130969 245077 131003
rect 245111 131000 245123 131003
rect 250217 131003 250275 131009
rect 250217 131000 250229 131003
rect 245111 130972 250229 131000
rect 245111 130969 245123 130972
rect 245065 130963 245123 130969
rect 250217 130969 250229 130972
rect 250263 130969 250275 131003
rect 250217 130963 250275 130969
rect 250306 130960 250312 131012
rect 250364 131000 250370 131012
rect 257206 131000 257212 131012
rect 250364 130972 257212 131000
rect 250364 130960 250370 130972
rect 257206 130960 257212 130972
rect 257264 130960 257270 131012
rect 49838 130892 49844 130944
rect 49896 130932 49902 130944
rect 62810 130932 62816 130944
rect 49896 130904 62816 130932
rect 49896 130892 49902 130904
rect 62810 130892 62816 130904
rect 62868 130892 62874 130944
rect 64006 130932 64012 130944
rect 62920 130904 64012 130932
rect 52598 130824 52604 130876
rect 52656 130864 52662 130876
rect 60697 130867 60755 130873
rect 60697 130864 60709 130867
rect 52656 130836 60709 130864
rect 52656 130824 52662 130836
rect 60697 130833 60709 130836
rect 60743 130833 60755 130867
rect 60697 130827 60755 130833
rect 60881 130867 60939 130873
rect 60881 130833 60893 130867
rect 60927 130864 60939 130867
rect 62920 130864 62948 130904
rect 64006 130892 64012 130904
rect 64064 130892 64070 130944
rect 65754 130892 65760 130944
rect 65812 130932 65818 130944
rect 70262 130932 70268 130944
rect 65812 130904 70268 130932
rect 65812 130892 65818 130904
rect 70262 130892 70268 130904
rect 70320 130892 70326 130944
rect 158306 130932 158312 130944
rect 155196 130904 158312 130932
rect 60927 130836 62948 130864
rect 60927 130833 60939 130836
rect 60881 130827 60939 130833
rect 62994 130824 63000 130876
rect 63052 130864 63058 130876
rect 66766 130864 66772 130876
rect 63052 130836 66772 130864
rect 63052 130824 63058 130836
rect 66766 130824 66772 130836
rect 66824 130824 66830 130876
rect 151406 130824 151412 130876
rect 151464 130864 151470 130876
rect 155089 130867 155147 130873
rect 155089 130864 155101 130867
rect 151464 130836 155101 130864
rect 151464 130824 151470 130836
rect 155089 130833 155101 130836
rect 155135 130833 155147 130867
rect 155089 130827 155147 130833
rect 56554 130756 56560 130808
rect 56612 130796 56618 130808
rect 61246 130796 61252 130808
rect 56612 130768 61252 130796
rect 56612 130756 56618 130768
rect 61246 130756 61252 130768
rect 61304 130756 61310 130808
rect 61982 130756 61988 130808
rect 62040 130796 62046 130808
rect 69526 130796 69532 130808
rect 62040 130768 69532 130796
rect 62040 130756 62046 130768
rect 69526 130756 69532 130768
rect 69584 130756 69590 130808
rect 151774 130756 151780 130808
rect 151832 130796 151838 130808
rect 155196 130796 155224 130904
rect 158306 130892 158312 130904
rect 158364 130892 158370 130944
rect 241658 130892 241664 130944
rect 241716 130932 241722 130944
rect 250582 130932 250588 130944
rect 241716 130904 250588 130932
rect 241716 130892 241722 130904
rect 250582 130892 250588 130904
rect 250640 130892 250646 130944
rect 250677 130935 250735 130941
rect 250677 130901 250689 130935
rect 250723 130932 250735 130935
rect 252882 130932 252888 130944
rect 250723 130904 252888 130932
rect 250723 130901 250735 130904
rect 250677 130895 250735 130901
rect 252882 130892 252888 130904
rect 252940 130892 252946 130944
rect 155273 130867 155331 130873
rect 155273 130833 155285 130867
rect 155319 130864 155331 130867
rect 158398 130864 158404 130876
rect 155319 130836 158404 130864
rect 155319 130833 155331 130836
rect 155273 130827 155331 130833
rect 158398 130824 158404 130836
rect 158456 130824 158462 130876
rect 247178 130824 247184 130876
rect 247236 130864 247242 130876
rect 250769 130867 250827 130873
rect 250769 130864 250781 130867
rect 247236 130836 250781 130864
rect 247236 130824 247242 130836
rect 250769 130833 250781 130836
rect 250815 130833 250827 130867
rect 250769 130827 250827 130833
rect 251137 130867 251195 130873
rect 251137 130833 251149 130867
rect 251183 130864 251195 130867
rect 253710 130864 253716 130876
rect 251183 130836 253716 130864
rect 251183 130833 251195 130836
rect 251137 130827 251195 130833
rect 253710 130824 253716 130836
rect 253768 130824 253774 130876
rect 151832 130768 155224 130796
rect 151832 130756 151838 130768
rect 155546 130756 155552 130808
rect 155604 130796 155610 130808
rect 157021 130799 157079 130805
rect 157021 130796 157033 130799
rect 155604 130768 157033 130796
rect 155604 130756 155610 130768
rect 157021 130765 157033 130768
rect 157067 130765 157079 130799
rect 157021 130759 157079 130765
rect 157389 130799 157447 130805
rect 157389 130765 157401 130799
rect 157435 130796 157447 130799
rect 160790 130796 160796 130808
rect 157435 130768 160796 130796
rect 157435 130765 157447 130768
rect 157389 130759 157447 130765
rect 160790 130756 160796 130768
rect 160848 130756 160854 130808
rect 243682 130756 243688 130808
rect 243740 130796 243746 130808
rect 245065 130799 245123 130805
rect 245065 130796 245077 130799
rect 243740 130768 245077 130796
rect 243740 130756 243746 130768
rect 245065 130765 245077 130768
rect 245111 130765 245123 130799
rect 250214 130796 250220 130808
rect 245065 130759 245123 130765
rect 245172 130768 250220 130796
rect 58118 130688 58124 130740
rect 58176 130728 58182 130740
rect 60142 130728 60148 130740
rect 58176 130700 60148 130728
rect 58176 130688 58182 130700
rect 60142 130688 60148 130700
rect 60200 130688 60206 130740
rect 61706 130728 61712 130740
rect 60252 130700 61712 130728
rect 58578 130620 58584 130672
rect 58636 130660 58642 130672
rect 59498 130660 59504 130672
rect 58636 130632 59504 130660
rect 58636 130620 58642 130632
rect 59498 130620 59504 130632
rect 59556 130620 59562 130672
rect 60252 130660 60280 130700
rect 61706 130688 61712 130700
rect 61764 130688 61770 130740
rect 61890 130688 61896 130740
rect 61948 130728 61954 130740
rect 67502 130728 67508 130740
rect 61948 130700 67508 130728
rect 61948 130688 61954 130700
rect 67502 130688 67508 130700
rect 67560 130688 67566 130740
rect 153062 130688 153068 130740
rect 153120 130728 153126 130740
rect 153120 130700 155868 130728
rect 153120 130688 153126 130700
rect 59608 130632 60280 130660
rect 55450 130552 55456 130604
rect 55508 130592 55514 130604
rect 59608 130592 59636 130632
rect 62166 130620 62172 130672
rect 62224 130660 62230 130672
rect 69894 130660 69900 130672
rect 62224 130632 69900 130660
rect 62224 130620 62230 130632
rect 69894 130620 69900 130632
rect 69952 130620 69958 130672
rect 155730 130660 155736 130672
rect 153908 130632 155736 130660
rect 55508 130564 59636 130592
rect 59685 130595 59743 130601
rect 55508 130552 55514 130564
rect 59685 130561 59697 130595
rect 59731 130592 59743 130595
rect 60881 130595 60939 130601
rect 60881 130592 60893 130595
rect 59731 130564 60893 130592
rect 59731 130561 59743 130564
rect 59685 130555 59743 130561
rect 60881 130561 60893 130564
rect 60927 130561 60939 130595
rect 60881 130555 60939 130561
rect 60970 130552 60976 130604
rect 61028 130592 61034 130604
rect 68698 130592 68704 130604
rect 61028 130564 68704 130592
rect 61028 130552 61034 130564
rect 68698 130552 68704 130564
rect 68756 130552 68762 130604
rect 150578 130552 150584 130604
rect 150636 130592 150642 130604
rect 153908 130592 153936 130632
rect 155730 130620 155736 130632
rect 155788 130620 155794 130672
rect 155840 130660 155868 130700
rect 155914 130688 155920 130740
rect 155972 130728 155978 130740
rect 155972 130700 161296 130728
rect 155972 130688 155978 130700
rect 156009 130663 156067 130669
rect 156009 130660 156021 130663
rect 155840 130632 156021 130660
rect 156009 130629 156021 130632
rect 156055 130629 156067 130663
rect 156009 130623 156067 130629
rect 156098 130620 156104 130672
rect 156156 130660 156162 130672
rect 158309 130663 158367 130669
rect 156156 130632 158260 130660
rect 156156 130620 156162 130632
rect 150636 130564 153936 130592
rect 150636 130552 150642 130564
rect 154258 130552 154264 130604
rect 154316 130592 154322 130604
rect 157294 130592 157300 130604
rect 154316 130564 157300 130592
rect 154316 130552 154322 130564
rect 157294 130552 157300 130564
rect 157352 130552 157358 130604
rect 158232 130592 158260 130632
rect 158309 130629 158321 130663
rect 158355 130660 158367 130663
rect 161158 130660 161164 130672
rect 158355 130632 161164 130660
rect 158355 130629 158367 130632
rect 158309 130623 158367 130629
rect 161158 130620 161164 130632
rect 161216 130620 161222 130672
rect 161268 130660 161296 130700
rect 244050 130688 244056 130740
rect 244108 130728 244114 130740
rect 245172 130728 245200 130768
rect 250214 130756 250220 130768
rect 250272 130756 250278 130808
rect 250674 130756 250680 130808
rect 250732 130796 250738 130808
rect 250732 130768 252100 130796
rect 250732 130756 250738 130768
rect 244108 130700 245200 130728
rect 244108 130688 244114 130700
rect 245246 130688 245252 130740
rect 245304 130728 245310 130740
rect 245706 130728 245712 130740
rect 245304 130700 245712 130728
rect 245304 130688 245310 130700
rect 245706 130688 245712 130700
rect 245764 130688 245770 130740
rect 246810 130688 246816 130740
rect 246868 130728 246874 130740
rect 249570 130728 249576 130740
rect 246868 130700 249576 130728
rect 246868 130688 246874 130700
rect 249570 130688 249576 130700
rect 249628 130688 249634 130740
rect 249849 130731 249907 130737
rect 249849 130697 249861 130731
rect 249895 130728 249907 130731
rect 249895 130700 250260 130728
rect 249895 130697 249907 130700
rect 249849 130691 249907 130697
rect 162722 130660 162728 130672
rect 161268 130632 162728 130660
rect 162722 130620 162728 130632
rect 162780 130620 162786 130672
rect 250232 130660 250260 130700
rect 250306 130688 250312 130740
rect 250364 130728 250370 130740
rect 251318 130728 251324 130740
rect 250364 130700 251324 130728
rect 250364 130688 250370 130700
rect 251318 130688 251324 130700
rect 251376 130688 251382 130740
rect 250585 130663 250643 130669
rect 250585 130660 250597 130663
rect 250232 130632 250597 130660
rect 250585 130629 250597 130632
rect 250631 130629 250643 130663
rect 251137 130663 251195 130669
rect 251137 130660 251149 130663
rect 250585 130623 250643 130629
rect 250692 130632 251149 130660
rect 163090 130592 163096 130604
rect 158232 130564 163096 130592
rect 163090 130552 163096 130564
rect 163148 130552 163154 130604
rect 244326 130552 244332 130604
rect 244384 130592 244390 130604
rect 246353 130595 246411 130601
rect 246353 130592 246365 130595
rect 244384 130564 246365 130592
rect 244384 130552 244390 130564
rect 246353 130561 246365 130564
rect 246399 130561 246411 130595
rect 246353 130555 246411 130561
rect 246442 130552 246448 130604
rect 246500 130592 246506 130604
rect 249202 130592 249208 130604
rect 246500 130564 249208 130592
rect 246500 130552 246506 130564
rect 249202 130552 249208 130564
rect 249260 130552 249266 130604
rect 58946 130484 58952 130536
rect 59004 130524 59010 130536
rect 67134 130524 67140 130536
rect 59004 130496 67140 130524
rect 59004 130484 59010 130496
rect 67134 130484 67140 130496
rect 67192 130484 67198 130536
rect 154166 130484 154172 130536
rect 154224 130524 154230 130536
rect 156926 130524 156932 130536
rect 154224 130496 156932 130524
rect 154224 130484 154230 130496
rect 156926 130484 156932 130496
rect 156984 130484 156990 130536
rect 157021 130527 157079 130533
rect 157021 130493 157033 130527
rect 157067 130524 157079 130527
rect 161986 130524 161992 130536
rect 157067 130496 161992 130524
rect 157067 130493 157079 130496
rect 157021 130487 157079 130493
rect 161986 130484 161992 130496
rect 162044 130484 162050 130536
rect 249110 130484 249116 130536
rect 249168 130524 249174 130536
rect 250692 130524 250720 130632
rect 251137 130629 251149 130632
rect 251183 130629 251195 130663
rect 251137 130623 251195 130629
rect 251226 130620 251232 130672
rect 251284 130660 251290 130672
rect 252072 130660 252100 130768
rect 252149 130731 252207 130737
rect 252149 130697 252161 130731
rect 252195 130728 252207 130731
rect 255550 130728 255556 130740
rect 252195 130700 255556 130728
rect 252195 130697 252207 130700
rect 252149 130691 252207 130697
rect 255550 130688 255556 130700
rect 255608 130688 255614 130740
rect 256102 130660 256108 130672
rect 251284 130632 251916 130660
rect 252072 130632 256108 130660
rect 251284 130620 251290 130632
rect 250766 130552 250772 130604
rect 250824 130592 250830 130604
rect 251778 130592 251784 130604
rect 250824 130564 251784 130592
rect 250824 130552 250830 130564
rect 251778 130552 251784 130564
rect 251836 130552 251842 130604
rect 251888 130592 251916 130632
rect 256102 130620 256108 130632
rect 256160 130620 256166 130672
rect 257666 130592 257672 130604
rect 251888 130564 257672 130592
rect 257666 130552 257672 130564
rect 257724 130552 257730 130604
rect 249168 130496 250720 130524
rect 249168 130484 249174 130496
rect 250858 130484 250864 130536
rect 250916 130524 250922 130536
rect 254906 130524 254912 130536
rect 250916 130496 254912 130524
rect 250916 130484 250922 130496
rect 254906 130484 254912 130496
rect 254964 130484 254970 130536
rect 57750 130416 57756 130468
rect 57808 130456 57814 130468
rect 60234 130456 60240 130468
rect 57808 130428 60240 130456
rect 57808 130416 57814 130428
rect 60234 130416 60240 130428
rect 60292 130416 60298 130468
rect 60329 130459 60387 130465
rect 60329 130425 60341 130459
rect 60375 130456 60387 130459
rect 60375 130428 61844 130456
rect 60375 130425 60387 130428
rect 60329 130419 60387 130425
rect 55818 130348 55824 130400
rect 55876 130388 55882 130400
rect 60789 130391 60847 130397
rect 60789 130388 60801 130391
rect 55876 130360 60801 130388
rect 55876 130348 55882 130360
rect 60789 130357 60801 130360
rect 60835 130357 60847 130391
rect 60789 130351 60847 130357
rect 61338 130348 61344 130400
rect 61396 130388 61402 130400
rect 61706 130388 61712 130400
rect 61396 130360 61712 130388
rect 61396 130348 61402 130360
rect 61706 130348 61712 130360
rect 61764 130348 61770 130400
rect 61816 130388 61844 130428
rect 61890 130416 61896 130468
rect 61948 130456 61954 130468
rect 64834 130456 64840 130468
rect 61948 130428 64840 130456
rect 61948 130416 61954 130428
rect 64834 130416 64840 130428
rect 64892 130416 64898 130468
rect 66398 130456 66404 130468
rect 64944 130428 66404 130456
rect 62353 130391 62411 130397
rect 62353 130388 62365 130391
rect 61816 130360 62365 130388
rect 62353 130357 62365 130360
rect 62399 130357 62411 130391
rect 62353 130351 62411 130357
rect 62442 130348 62448 130400
rect 62500 130388 62506 130400
rect 63638 130388 63644 130400
rect 62500 130360 63644 130388
rect 62500 130348 62506 130360
rect 63638 130348 63644 130360
rect 63696 130348 63702 130400
rect 64944 130388 64972 130428
rect 66398 130416 66404 130428
rect 66456 130416 66462 130468
rect 154074 130416 154080 130468
rect 154132 130456 154138 130468
rect 156558 130456 156564 130468
rect 154132 130428 156564 130456
rect 154132 130416 154138 130428
rect 156558 130416 156564 130428
rect 156616 130416 156622 130468
rect 161158 130456 161164 130468
rect 158140 130428 161164 130456
rect 63840 130360 64972 130388
rect 65021 130391 65079 130397
rect 13774 130280 13780 130332
rect 13832 130320 13838 130332
rect 31898 130320 31904 130332
rect 13832 130292 31904 130320
rect 13832 130280 13838 130292
rect 31898 130280 31904 130292
rect 31956 130280 31962 130332
rect 38338 130280 38344 130332
rect 38396 130320 38402 130332
rect 63733 130323 63791 130329
rect 63733 130320 63745 130323
rect 38396 130292 63745 130320
rect 38396 130280 38402 130292
rect 63733 130289 63745 130292
rect 63779 130289 63791 130323
rect 63733 130283 63791 130289
rect 62353 130255 62411 130261
rect 62353 130221 62365 130255
rect 62399 130252 62411 130255
rect 63840 130252 63868 130360
rect 65021 130357 65033 130391
rect 65067 130388 65079 130391
rect 65938 130388 65944 130400
rect 65067 130360 65944 130388
rect 65067 130357 65079 130360
rect 65021 130351 65079 130357
rect 65938 130348 65944 130360
rect 65996 130348 66002 130400
rect 70630 130388 70636 130400
rect 66048 130360 70636 130388
rect 63917 130323 63975 130329
rect 63917 130289 63929 130323
rect 63963 130320 63975 130323
rect 63963 130292 65708 130320
rect 63963 130289 63975 130292
rect 63917 130283 63975 130289
rect 62399 130224 63868 130252
rect 65680 130252 65708 130292
rect 66048 130252 66076 130360
rect 70630 130348 70636 130360
rect 70688 130348 70694 130400
rect 154534 130348 154540 130400
rect 154592 130388 154598 130400
rect 156834 130388 156840 130400
rect 154592 130360 156840 130388
rect 154592 130348 154598 130360
rect 156834 130348 156840 130360
rect 156892 130348 156898 130400
rect 152142 130280 152148 130332
rect 152200 130320 152206 130332
rect 152200 130292 154856 130320
rect 152200 130280 152206 130292
rect 65680 130224 66076 130252
rect 62399 130221 62411 130224
rect 62353 130215 62411 130221
rect 136870 130212 136876 130264
rect 136928 130252 136934 130264
rect 138986 130252 138992 130264
rect 136928 130224 138992 130252
rect 136928 130212 136934 130224
rect 138986 130212 138992 130224
rect 139044 130212 139050 130264
rect 154828 130252 154856 130292
rect 154902 130280 154908 130332
rect 154960 130320 154966 130332
rect 155270 130320 155276 130332
rect 154960 130292 155276 130320
rect 154960 130280 154966 130292
rect 155270 130280 155276 130292
rect 155328 130280 155334 130332
rect 155730 130280 155736 130332
rect 155788 130320 155794 130332
rect 156006 130320 156012 130332
rect 155788 130292 156012 130320
rect 155788 130280 155794 130292
rect 156006 130280 156012 130292
rect 156064 130280 156070 130332
rect 156101 130323 156159 130329
rect 156101 130289 156113 130323
rect 156147 130320 156159 130323
rect 158140 130320 158168 130428
rect 161158 130416 161164 130428
rect 161216 130416 161222 130468
rect 247546 130416 247552 130468
rect 247604 130456 247610 130468
rect 254814 130456 254820 130468
rect 247604 130428 254820 130456
rect 247604 130416 247610 130428
rect 254814 130416 254820 130428
rect 254872 130416 254878 130468
rect 158214 130348 158220 130400
rect 158272 130388 158278 130400
rect 159962 130388 159968 130400
rect 158272 130360 159968 130388
rect 158272 130348 158278 130360
rect 159962 130348 159968 130360
rect 160020 130348 160026 130400
rect 247914 130348 247920 130400
rect 247972 130388 247978 130400
rect 250950 130388 250956 130400
rect 247972 130360 250956 130388
rect 247972 130348 247978 130360
rect 250950 130348 250956 130360
rect 251008 130348 251014 130400
rect 251042 130348 251048 130400
rect 251100 130388 251106 130400
rect 251410 130388 251416 130400
rect 251100 130360 251416 130388
rect 251100 130348 251106 130360
rect 251410 130348 251416 130360
rect 251468 130348 251474 130400
rect 252146 130348 252152 130400
rect 252204 130388 252210 130400
rect 256470 130388 256476 130400
rect 252204 130360 256476 130388
rect 252204 130348 252210 130360
rect 256470 130348 256476 130360
rect 256528 130348 256534 130400
rect 158309 130323 158367 130329
rect 158309 130320 158321 130323
rect 156147 130292 158168 130320
rect 158232 130292 158321 130320
rect 156147 130289 156159 130292
rect 156101 130283 156159 130289
rect 158232 130252 158260 130292
rect 158309 130289 158321 130292
rect 158355 130289 158367 130323
rect 158309 130283 158367 130289
rect 158490 130280 158496 130332
rect 158548 130320 158554 130332
rect 159594 130320 159600 130332
rect 158548 130292 159600 130320
rect 158548 130280 158554 130292
rect 159594 130280 159600 130292
rect 159652 130280 159658 130332
rect 249294 130280 249300 130332
rect 249352 130320 249358 130332
rect 253342 130320 253348 130332
rect 249352 130292 253348 130320
rect 249352 130280 249358 130292
rect 253342 130280 253348 130292
rect 253400 130280 253406 130332
rect 253434 130280 253440 130332
rect 253492 130320 253498 130332
rect 254538 130320 254544 130332
rect 253492 130292 254544 130320
rect 253492 130280 253498 130292
rect 254538 130280 254544 130292
rect 254596 130280 254602 130332
rect 154828 130224 158260 130252
rect 231998 130212 232004 130264
rect 232056 130252 232062 130264
rect 232918 130252 232924 130264
rect 232056 130224 232924 130252
rect 232056 130212 232062 130224
rect 232918 130212 232924 130224
rect 232976 130212 232982 130264
rect 228502 127600 228508 127612
rect 228428 127572 228508 127600
rect 136870 127492 136876 127544
rect 136928 127532 136934 127544
rect 145334 127532 145340 127544
rect 136928 127504 145340 127532
rect 136928 127492 136934 127504
rect 145334 127492 145340 127504
rect 145392 127492 145398 127544
rect 228428 127476 228456 127572
rect 228502 127560 228508 127572
rect 228560 127560 228566 127612
rect 230710 127492 230716 127544
rect 230768 127532 230774 127544
rect 239634 127532 239640 127544
rect 230768 127504 239640 127532
rect 230768 127492 230774 127504
rect 239634 127492 239640 127504
rect 239692 127492 239698 127544
rect 228410 127424 228416 127476
rect 228468 127424 228474 127476
rect 148738 126608 148744 126660
rect 148796 126648 148802 126660
rect 165114 126648 165120 126660
rect 148796 126620 165120 126648
rect 148796 126608 148802 126620
rect 165114 126608 165120 126620
rect 165172 126608 165178 126660
rect 231630 124976 231636 125028
rect 231688 125016 231694 125028
rect 238254 125016 238260 125028
rect 231688 124988 238260 125016
rect 231688 124976 231694 124988
rect 238254 124976 238260 124988
rect 238312 124976 238318 125028
rect 138158 124840 138164 124892
rect 138216 124880 138222 124892
rect 144414 124880 144420 124892
rect 138216 124852 144420 124880
rect 138216 124840 138222 124852
rect 144414 124840 144420 124852
rect 144472 124840 144478 124892
rect 137882 124772 137888 124824
rect 137940 124812 137946 124824
rect 145610 124812 145616 124824
rect 137940 124784 145616 124812
rect 137940 124772 137946 124784
rect 145610 124772 145616 124784
rect 145668 124772 145674 124824
rect 231906 124772 231912 124824
rect 231964 124812 231970 124824
rect 240922 124812 240928 124824
rect 231964 124784 240928 124812
rect 231964 124772 231970 124784
rect 240922 124772 240928 124784
rect 240980 124772 240986 124824
rect 228410 124744 228416 124756
rect 228371 124716 228416 124744
rect 228410 124704 228416 124716
rect 228468 124704 228474 124756
rect 47814 122188 47820 122240
rect 47872 122228 47878 122240
rect 51310 122228 51316 122240
rect 47872 122200 51316 122228
rect 47872 122188 47878 122200
rect 51310 122188 51316 122200
rect 51368 122188 51374 122240
rect 138158 122052 138164 122104
rect 138216 122092 138222 122104
rect 143034 122092 143040 122104
rect 138216 122064 143040 122092
rect 138216 122052 138222 122064
rect 143034 122052 143040 122064
rect 143092 122052 143098 122104
rect 231630 122052 231636 122104
rect 231688 122092 231694 122104
rect 236874 122092 236880 122104
rect 231688 122064 236880 122092
rect 231688 122052 231694 122064
rect 236874 122052 236880 122064
rect 236932 122052 236938 122104
rect 137974 121984 137980 122036
rect 138032 122024 138038 122036
rect 145610 122024 145616 122036
rect 138032 121996 145616 122024
rect 138032 121984 138038 121996
rect 145610 121984 145616 121996
rect 145668 121984 145674 122036
rect 231998 121984 232004 122036
rect 232056 122024 232062 122036
rect 240922 122024 240928 122036
rect 232056 121996 240928 122024
rect 232056 121984 232062 121996
rect 240922 121984 240928 121996
rect 240980 121984 240986 122036
rect 165114 121916 165120 121968
rect 165172 121956 165178 121968
rect 175510 121956 175516 121968
rect 165172 121928 175516 121956
rect 165172 121916 165178 121928
rect 175510 121916 175516 121928
rect 175568 121916 175574 121968
rect 228413 120531 228471 120537
rect 228413 120497 228425 120531
rect 228459 120528 228471 120531
rect 228502 120528 228508 120540
rect 228459 120500 228508 120528
rect 228459 120497 228471 120500
rect 228413 120491 228471 120497
rect 228502 120488 228508 120500
rect 228560 120488 228566 120540
rect 138066 119264 138072 119316
rect 138124 119304 138130 119316
rect 145610 119304 145616 119316
rect 138124 119276 145616 119304
rect 138124 119264 138130 119276
rect 145610 119264 145616 119276
rect 145668 119264 145674 119316
rect 231906 119264 231912 119316
rect 231964 119304 231970 119316
rect 240922 119304 240928 119316
rect 231964 119276 240928 119304
rect 231964 119264 231970 119276
rect 240922 119264 240928 119276
rect 240980 119264 240986 119316
rect 231630 118448 231636 118500
rect 231688 118488 231694 118500
rect 235494 118488 235500 118500
rect 231688 118460 235500 118488
rect 231688 118448 231694 118460
rect 235494 118448 235500 118460
rect 235552 118448 235558 118500
rect 138158 117904 138164 117956
rect 138216 117944 138222 117956
rect 141654 117944 141660 117956
rect 138216 117916 141660 117944
rect 138216 117904 138222 117916
rect 141654 117904 141660 117916
rect 141712 117904 141718 117956
rect 137790 117836 137796 117888
rect 137848 117876 137854 117888
rect 145610 117876 145616 117888
rect 137848 117848 145616 117876
rect 137848 117836 137854 117848
rect 145610 117836 145616 117848
rect 145668 117836 145674 117888
rect 231630 117836 231636 117888
rect 231688 117876 231694 117888
rect 240922 117876 240928 117888
rect 231688 117848 240928 117876
rect 231688 117836 231694 117848
rect 240922 117836 240928 117848
rect 240980 117836 240986 117888
rect 292810 117836 292816 117888
rect 292868 117876 292874 117888
rect 300170 117876 300176 117888
rect 292868 117848 300176 117876
rect 292868 117836 292874 117848
rect 300170 117836 300176 117848
rect 300228 117836 300234 117888
rect 137330 115184 137336 115236
rect 137388 115224 137394 115236
rect 140274 115224 140280 115236
rect 137388 115196 140280 115224
rect 137388 115184 137394 115196
rect 140274 115184 140280 115196
rect 140332 115184 140338 115236
rect 231262 115184 231268 115236
rect 231320 115224 231326 115236
rect 234114 115224 234120 115236
rect 231320 115196 234120 115224
rect 231320 115184 231326 115196
rect 234114 115184 234120 115196
rect 234172 115184 234178 115236
rect 137698 115116 137704 115168
rect 137756 115156 137762 115168
rect 145610 115156 145616 115168
rect 137756 115128 145616 115156
rect 137756 115116 137762 115128
rect 145610 115116 145616 115128
rect 145668 115116 145674 115168
rect 231538 115116 231544 115168
rect 231596 115156 231602 115168
rect 240922 115156 240928 115168
rect 231596 115128 240928 115156
rect 231596 115116 231602 115128
rect 240922 115116 240928 115128
rect 240980 115116 240986 115168
rect 263738 115048 263744 115100
rect 263796 115088 263802 115100
rect 274870 115088 274876 115100
rect 263796 115060 274876 115088
rect 263796 115048 263802 115060
rect 274870 115048 274876 115060
rect 274928 115048 274934 115100
rect 138158 112532 138164 112584
rect 138216 112572 138222 112584
rect 138986 112572 138992 112584
rect 138216 112544 138992 112572
rect 138216 112532 138222 112544
rect 138986 112532 138992 112544
rect 139044 112532 139050 112584
rect 292810 112504 292816 112516
rect 292771 112476 292816 112504
rect 292810 112464 292816 112476
rect 292868 112464 292874 112516
rect 137422 112328 137428 112380
rect 137480 112368 137486 112380
rect 145610 112368 145616 112380
rect 137480 112340 145616 112368
rect 137480 112328 137486 112340
rect 145610 112328 145616 112340
rect 145668 112328 145674 112380
rect 231262 112328 231268 112380
rect 231320 112368 231326 112380
rect 240738 112368 240744 112380
rect 231320 112340 240744 112368
rect 231320 112328 231326 112340
rect 240738 112328 240744 112340
rect 240796 112328 240802 112380
rect 292810 111920 292816 111972
rect 292868 111960 292874 111972
rect 293546 111960 293552 111972
rect 292868 111932 293552 111960
rect 292868 111920 292874 111932
rect 293546 111920 293552 111932
rect 293604 111920 293610 111972
rect 138158 110968 138164 111020
rect 138216 111008 138222 111020
rect 145610 111008 145616 111020
rect 138216 110980 145616 111008
rect 138216 110968 138222 110980
rect 145610 110968 145616 110980
rect 145668 110968 145674 111020
rect 231998 110968 232004 111020
rect 232056 111008 232062 111020
rect 240922 111008 240928 111020
rect 232056 110980 240928 111008
rect 232056 110968 232062 110980
rect 240922 110968 240928 110980
rect 240980 110968 240986 111020
rect 292810 110260 292816 110272
rect 292771 110232 292816 110260
rect 292810 110220 292816 110232
rect 292868 110220 292874 110272
rect 231538 109540 231544 109592
rect 231596 109580 231602 109592
rect 232826 109580 232832 109592
rect 231596 109552 232832 109580
rect 231596 109540 231602 109552
rect 232826 109540 232832 109552
rect 232884 109540 232890 109592
rect 47078 109472 47084 109524
rect 47136 109512 47142 109524
rect 51310 109512 51316 109524
rect 47136 109484 51316 109512
rect 47136 109472 47142 109484
rect 51310 109472 51316 109484
rect 51368 109472 51374 109524
rect 137330 108180 137336 108232
rect 137388 108220 137394 108232
rect 145610 108220 145616 108232
rect 137388 108192 145616 108220
rect 137388 108180 137394 108192
rect 145610 108180 145616 108192
rect 145668 108180 145674 108232
rect 228502 108180 228508 108232
rect 228560 108180 228566 108232
rect 231446 108180 231452 108232
rect 231504 108220 231510 108232
rect 240830 108220 240836 108232
rect 231504 108192 240836 108220
rect 231504 108180 231510 108192
rect 240830 108180 240836 108192
rect 240888 108180 240894 108232
rect 228520 108096 228548 108180
rect 228502 108044 228508 108096
rect 228560 108044 228566 108096
rect 140366 105460 140372 105512
rect 140424 105500 140430 105512
rect 145610 105500 145616 105512
rect 140424 105472 145616 105500
rect 140424 105460 140430 105472
rect 145610 105460 145616 105472
rect 145668 105460 145674 105512
rect 231722 105460 231728 105512
rect 231780 105500 231786 105512
rect 240922 105500 240928 105512
rect 231780 105472 240928 105500
rect 231780 105460 231786 105472
rect 240922 105460 240928 105472
rect 240980 105460 240986 105512
rect 143126 103080 143132 103132
rect 143184 103120 143190 103132
rect 145426 103120 145432 103132
rect 143184 103092 145432 103120
rect 143184 103080 143190 103092
rect 145426 103080 145432 103092
rect 145484 103080 145490 103132
rect 236966 102672 236972 102724
rect 237024 102712 237030 102724
rect 240738 102712 240744 102724
rect 237024 102684 240744 102712
rect 237024 102672 237030 102684
rect 240738 102672 240744 102684
rect 240796 102672 240802 102724
rect 265118 102672 265124 102724
rect 265176 102712 265182 102724
rect 274870 102712 274876 102724
rect 265176 102684 274876 102712
rect 265176 102672 265182 102684
rect 274870 102672 274876 102684
rect 274928 102672 274934 102724
rect 140458 101312 140464 101364
rect 140516 101352 140522 101364
rect 145610 101352 145616 101364
rect 140516 101324 145616 101352
rect 140516 101312 140522 101324
rect 145610 101312 145616 101324
rect 145668 101312 145674 101364
rect 234206 101312 234212 101364
rect 234264 101352 234270 101364
rect 240370 101352 240376 101364
rect 234264 101324 240376 101352
rect 234264 101312 234270 101324
rect 240370 101312 240376 101324
rect 240428 101312 240434 101364
rect 140550 98524 140556 98576
rect 140608 98564 140614 98576
rect 145610 98564 145616 98576
rect 140608 98536 145616 98564
rect 140608 98524 140614 98536
rect 145610 98524 145616 98536
rect 145668 98524 145674 98576
rect 167874 98524 167880 98576
rect 167932 98564 167938 98576
rect 175510 98564 175516 98576
rect 167932 98536 175516 98564
rect 167932 98524 167938 98536
rect 175510 98524 175516 98536
rect 175568 98524 175574 98576
rect 234298 98524 234304 98576
rect 234356 98564 234362 98576
rect 240830 98564 240836 98576
rect 234356 98536 240836 98564
rect 234356 98524 234362 98536
rect 240830 98524 240836 98536
rect 240888 98524 240894 98576
rect 262358 98524 262364 98576
rect 262416 98564 262422 98576
rect 272754 98564 272760 98576
rect 262416 98536 272760 98564
rect 262416 98524 262422 98536
rect 272754 98524 272760 98536
rect 272812 98524 272818 98576
rect 74034 97096 74040 97148
rect 74092 97136 74098 97148
rect 81670 97136 81676 97148
rect 74092 97108 81676 97136
rect 74092 97096 74098 97108
rect 81670 97096 81676 97108
rect 81728 97096 81734 97148
rect 238346 95804 238352 95856
rect 238404 95844 238410 95856
rect 240922 95844 240928 95856
rect 238404 95816 240928 95844
rect 238404 95804 238410 95816
rect 240922 95804 240928 95816
rect 240980 95804 240986 95856
rect 138158 95736 138164 95788
rect 138216 95776 138222 95788
rect 140366 95776 140372 95788
rect 138216 95748 140372 95776
rect 138216 95736 138222 95748
rect 140366 95736 140372 95748
rect 140424 95736 140430 95788
rect 228502 95776 228508 95788
rect 228463 95748 228508 95776
rect 228502 95736 228508 95748
rect 228560 95736 228566 95788
rect 45790 94376 45796 94428
rect 45848 94416 45854 94428
rect 51310 94416 51316 94428
rect 45848 94388 51316 94416
rect 45848 94376 45854 94388
rect 51310 94376 51316 94388
rect 51368 94376 51374 94428
rect 143770 94376 143776 94428
rect 143828 94416 143834 94428
rect 146346 94416 146352 94428
rect 143828 94388 146352 94416
rect 143828 94376 143834 94388
rect 146346 94376 146352 94388
rect 146404 94376 146410 94428
rect 237610 94376 237616 94428
rect 237668 94416 237674 94428
rect 240922 94416 240928 94428
rect 237668 94388 240928 94416
rect 237668 94376 237674 94388
rect 240922 94376 240928 94388
rect 240980 94376 240986 94428
rect 292810 94376 292816 94428
rect 292868 94416 292874 94428
rect 299710 94416 299716 94428
rect 292868 94388 299716 94416
rect 292868 94376 292874 94388
rect 299710 94376 299716 94388
rect 299768 94376 299774 94428
rect 272754 94308 272760 94360
rect 272812 94348 272818 94360
rect 274870 94348 274876 94360
rect 272812 94320 274876 94348
rect 272812 94308 272818 94320
rect 274870 94308 274876 94320
rect 274928 94308 274934 94360
rect 231814 94172 231820 94224
rect 231872 94212 231878 94224
rect 236966 94212 236972 94224
rect 231872 94184 236972 94212
rect 231872 94172 231878 94184
rect 236966 94172 236972 94184
rect 237024 94172 237030 94224
rect 138158 93832 138164 93884
rect 138216 93872 138222 93884
rect 143126 93872 143132 93884
rect 138216 93844 143132 93872
rect 138216 93832 138222 93844
rect 143126 93832 143132 93844
rect 143184 93832 143190 93884
rect 38798 92948 38804 93000
rect 38856 92988 38862 93000
rect 45790 92988 45796 93000
rect 38856 92960 45796 92988
rect 38856 92948 38862 92960
rect 45790 92948 45796 92960
rect 45848 92948 45854 93000
rect 231446 92948 231452 93000
rect 231504 92988 231510 93000
rect 234206 92988 234212 93000
rect 231504 92960 234212 92988
rect 231504 92948 231510 92960
rect 234206 92948 234212 92960
rect 234264 92948 234270 93000
rect 137790 92676 137796 92728
rect 137848 92716 137854 92728
rect 140458 92716 140464 92728
rect 137848 92688 140464 92716
rect 137848 92676 137854 92688
rect 140458 92676 140464 92688
rect 140516 92676 140522 92728
rect 143678 91656 143684 91708
rect 143736 91696 143742 91708
rect 145242 91696 145248 91708
rect 143736 91668 145248 91696
rect 143736 91656 143742 91668
rect 145242 91656 145248 91668
rect 145300 91656 145306 91708
rect 236322 91656 236328 91708
rect 236380 91696 236386 91708
rect 240922 91696 240928 91708
rect 236380 91668 240928 91696
rect 236380 91656 236386 91668
rect 240922 91656 240928 91668
rect 240980 91656 240986 91708
rect 137606 91588 137612 91640
rect 137664 91628 137670 91640
rect 140550 91628 140556 91640
rect 137664 91600 140556 91628
rect 137664 91588 137670 91600
rect 140550 91588 140556 91600
rect 140608 91588 140614 91640
rect 231446 91588 231452 91640
rect 231504 91628 231510 91640
rect 234298 91628 234304 91640
rect 231504 91600 234304 91628
rect 231504 91588 231510 91600
rect 234298 91588 234304 91600
rect 234356 91588 234362 91640
rect 228502 90880 228508 90892
rect 228463 90852 228508 90880
rect 228502 90840 228508 90852
rect 228560 90840 228566 90892
rect 231630 90024 231636 90076
rect 231688 90064 231694 90076
rect 238346 90064 238352 90076
rect 231688 90036 238352 90064
rect 231688 90024 231694 90036
rect 238346 90024 238352 90036
rect 238404 90024 238410 90076
rect 138158 89140 138164 89192
rect 138216 89180 138222 89192
rect 144598 89180 144604 89192
rect 138216 89152 144604 89180
rect 138216 89140 138222 89152
rect 144598 89140 144604 89152
rect 144656 89140 144662 89192
rect 155270 88936 155276 88988
rect 155328 88976 155334 88988
rect 155546 88976 155552 88988
rect 155328 88948 155552 88976
rect 155328 88936 155334 88948
rect 155546 88936 155552 88948
rect 155604 88936 155610 88988
rect 143494 88868 143500 88920
rect 143552 88908 143558 88920
rect 145242 88908 145248 88920
rect 143552 88880 145248 88908
rect 143552 88868 143558 88880
rect 145242 88868 145248 88880
rect 145300 88868 145306 88920
rect 236230 88868 236236 88920
rect 236288 88908 236294 88920
rect 240922 88908 240928 88920
rect 236288 88880 240928 88908
rect 236288 88868 236294 88880
rect 240922 88868 240928 88880
rect 240980 88868 240986 88920
rect 137606 88800 137612 88852
rect 137664 88840 137670 88852
rect 143770 88840 143776 88852
rect 137664 88812 143776 88840
rect 137664 88800 137670 88812
rect 143770 88800 143776 88812
rect 143828 88800 143834 88852
rect 231630 88460 231636 88512
rect 231688 88500 231694 88512
rect 237610 88500 237616 88512
rect 231688 88472 237616 88500
rect 231688 88460 231694 88472
rect 237610 88460 237616 88472
rect 237668 88460 237674 88512
rect 292534 88120 292540 88172
rect 292592 88160 292598 88172
rect 292718 88160 292724 88172
rect 292592 88132 292724 88160
rect 292592 88120 292598 88132
rect 292718 88120 292724 88132
rect 292776 88120 292782 88172
rect 60145 87551 60203 87557
rect 60145 87517 60157 87551
rect 60191 87548 60203 87551
rect 155549 87551 155607 87557
rect 60191 87520 61108 87548
rect 60191 87517 60203 87520
rect 60145 87511 60203 87517
rect 23894 87440 23900 87492
rect 23952 87480 23958 87492
rect 23952 87452 30564 87480
rect 23952 87440 23958 87452
rect 30536 87344 30564 87452
rect 31898 87440 31904 87492
rect 31956 87480 31962 87492
rect 34566 87480 34572 87492
rect 31956 87452 34572 87480
rect 31956 87440 31962 87452
rect 34566 87440 34572 87452
rect 34624 87440 34630 87492
rect 55082 87440 55088 87492
rect 55140 87480 55146 87492
rect 56094 87480 56100 87492
rect 55140 87452 56100 87480
rect 55140 87440 55146 87452
rect 56094 87440 56100 87452
rect 56152 87440 56158 87492
rect 58670 87440 58676 87492
rect 58728 87480 58734 87492
rect 60973 87483 61031 87489
rect 60973 87480 60985 87483
rect 58728 87452 60985 87480
rect 58728 87440 58734 87452
rect 60973 87449 60985 87452
rect 61019 87449 61031 87483
rect 61080 87480 61108 87520
rect 155549 87517 155561 87551
rect 155595 87548 155607 87551
rect 250769 87551 250827 87557
rect 155595 87520 157524 87548
rect 155595 87517 155607 87520
rect 155549 87511 155607 87517
rect 65478 87480 65484 87492
rect 61080 87452 65484 87480
rect 60973 87443 61031 87449
rect 65478 87440 65484 87452
rect 65536 87440 65542 87492
rect 154166 87440 154172 87492
rect 154224 87480 154230 87492
rect 157386 87480 157392 87492
rect 154224 87452 157392 87480
rect 154224 87440 154230 87452
rect 157386 87440 157392 87452
rect 157444 87440 157450 87492
rect 157496 87480 157524 87520
rect 250769 87517 250781 87551
rect 250815 87548 250827 87551
rect 250815 87520 251180 87548
rect 250815 87517 250827 87520
rect 250769 87511 250827 87517
rect 160698 87480 160704 87492
rect 157496 87452 160704 87480
rect 160698 87440 160704 87452
rect 160756 87440 160762 87492
rect 160974 87440 160980 87492
rect 161032 87480 161038 87492
rect 162262 87480 162268 87492
rect 161032 87452 162268 87480
rect 161032 87440 161038 87452
rect 162262 87440 162268 87452
rect 162320 87440 162326 87492
rect 251152 87480 251180 87520
rect 254354 87480 254360 87492
rect 251152 87452 254360 87480
rect 254354 87440 254360 87452
rect 254412 87440 254418 87492
rect 59866 87372 59872 87424
rect 59924 87412 59930 87424
rect 70722 87412 70728 87424
rect 59924 87384 70728 87412
rect 59924 87372 59930 87384
rect 70722 87372 70728 87384
rect 70780 87372 70786 87424
rect 152694 87372 152700 87424
rect 152752 87412 152758 87424
rect 158398 87412 158404 87424
rect 152752 87384 158404 87412
rect 152752 87372 152758 87384
rect 158398 87372 158404 87384
rect 158456 87372 158462 87424
rect 159594 87372 159600 87424
rect 159652 87412 159658 87424
rect 161066 87412 161072 87424
rect 159652 87384 161072 87412
rect 159652 87372 159658 87384
rect 161066 87372 161072 87384
rect 161124 87372 161130 87424
rect 249938 87372 249944 87424
rect 249996 87412 250002 87424
rect 256930 87412 256936 87424
rect 249996 87384 256936 87412
rect 249996 87372 250002 87384
rect 256930 87372 256936 87384
rect 256988 87372 256994 87424
rect 34658 87344 34664 87356
rect 30536 87316 34664 87344
rect 34658 87304 34664 87316
rect 34716 87304 34722 87356
rect 58210 87304 58216 87356
rect 58268 87344 58274 87356
rect 67134 87344 67140 87356
rect 58268 87316 67140 87344
rect 58268 87304 58274 87316
rect 67134 87304 67140 87316
rect 67192 87304 67198 87356
rect 153062 87304 153068 87356
rect 153120 87344 153126 87356
rect 158214 87344 158220 87356
rect 153120 87316 158220 87344
rect 153120 87304 153126 87316
rect 158214 87304 158220 87316
rect 158272 87304 158278 87356
rect 246074 87304 246080 87356
rect 246132 87344 246138 87356
rect 255734 87344 255740 87356
rect 246132 87316 255740 87344
rect 246132 87304 246138 87316
rect 255734 87304 255740 87316
rect 255792 87304 255798 87356
rect 53978 87236 53984 87288
rect 54036 87276 54042 87288
rect 60145 87279 60203 87285
rect 60145 87276 60157 87279
rect 54036 87248 60157 87276
rect 54036 87236 54042 87248
rect 60145 87245 60157 87248
rect 60191 87245 60203 87279
rect 60145 87239 60203 87245
rect 60234 87236 60240 87288
rect 60292 87276 60298 87288
rect 70814 87276 70820 87288
rect 60292 87248 70820 87276
rect 60292 87236 60298 87248
rect 70814 87236 70820 87248
rect 70872 87236 70878 87288
rect 152694 87236 152700 87288
rect 152752 87276 152758 87288
rect 157478 87276 157484 87288
rect 152752 87248 157484 87276
rect 152752 87236 152758 87248
rect 157478 87236 157484 87248
rect 157536 87236 157542 87288
rect 161066 87236 161072 87288
rect 161124 87276 161130 87288
rect 161894 87276 161900 87288
rect 161124 87248 161900 87276
rect 161124 87236 161130 87248
rect 161894 87236 161900 87248
rect 161952 87236 161958 87288
rect 246534 87236 246540 87288
rect 246592 87276 246598 87288
rect 256930 87276 256936 87288
rect 246592 87248 256936 87276
rect 246592 87236 246598 87248
rect 256930 87236 256936 87248
rect 256988 87236 256994 87288
rect 60973 87211 61031 87217
rect 60973 87177 60985 87211
rect 61019 87208 61031 87211
rect 67226 87208 67232 87220
rect 61019 87180 67232 87208
rect 61019 87177 61031 87180
rect 60973 87171 61031 87177
rect 67226 87168 67232 87180
rect 67284 87168 67290 87220
rect 150302 87168 150308 87220
rect 150360 87208 150366 87220
rect 159318 87208 159324 87220
rect 150360 87180 159324 87208
rect 150360 87168 150366 87180
rect 159318 87168 159324 87180
rect 159376 87168 159382 87220
rect 246902 87168 246908 87220
rect 246960 87208 246966 87220
rect 257022 87208 257028 87220
rect 246960 87180 257028 87208
rect 246960 87168 246966 87180
rect 257022 87168 257028 87180
rect 257080 87168 257086 87220
rect 58949 87143 59007 87149
rect 58949 87109 58961 87143
rect 58995 87140 59007 87143
rect 63822 87140 63828 87152
rect 58995 87112 63828 87140
rect 58995 87109 59007 87112
rect 58949 87103 59007 87109
rect 63822 87100 63828 87112
rect 63880 87100 63886 87152
rect 154074 87100 154080 87152
rect 154132 87140 154138 87152
rect 157389 87143 157447 87149
rect 157389 87140 157401 87143
rect 154132 87112 157401 87140
rect 154132 87100 154138 87112
rect 157389 87109 157401 87112
rect 157435 87109 157447 87143
rect 157389 87103 157447 87109
rect 157478 87100 157484 87152
rect 157536 87140 157542 87152
rect 158306 87140 158312 87152
rect 157536 87112 158312 87140
rect 157536 87100 157542 87112
rect 158306 87100 158312 87112
rect 158364 87100 158370 87152
rect 248098 87100 248104 87152
rect 248156 87140 248162 87152
rect 256286 87140 256292 87152
rect 248156 87112 256292 87140
rect 248156 87100 248162 87112
rect 256286 87100 256292 87112
rect 256344 87100 256350 87152
rect 52598 87032 52604 87084
rect 52656 87072 52662 87084
rect 64650 87072 64656 87084
rect 52656 87044 64656 87072
rect 52656 87032 52662 87044
rect 64650 87032 64656 87044
rect 64708 87032 64714 87084
rect 149842 87032 149848 87084
rect 149900 87072 149906 87084
rect 158950 87072 158956 87084
rect 149900 87044 158956 87072
rect 149900 87032 149906 87044
rect 158950 87032 158956 87044
rect 159008 87032 159014 87084
rect 247730 87032 247736 87084
rect 247788 87072 247794 87084
rect 256470 87072 256476 87084
rect 247788 87044 256476 87072
rect 247788 87032 247794 87044
rect 256470 87032 256476 87044
rect 256528 87032 256534 87084
rect 51218 86964 51224 87016
rect 51276 87004 51282 87016
rect 63454 87004 63460 87016
rect 51276 86976 63460 87004
rect 51276 86964 51282 86976
rect 63454 86964 63460 86976
rect 63512 86964 63518 87016
rect 151314 86964 151320 87016
rect 151372 87004 151378 87016
rect 157110 87004 157116 87016
rect 151372 86976 157116 87004
rect 151372 86964 151378 86976
rect 157110 86964 157116 86976
rect 157168 86964 157174 87016
rect 157205 87007 157263 87013
rect 157205 86973 157217 87007
rect 157251 87004 157263 87007
rect 159042 87004 159048 87016
rect 157251 86976 159048 87004
rect 157251 86973 157263 86976
rect 157205 86967 157263 86973
rect 159042 86964 159048 86976
rect 159100 86964 159106 87016
rect 247178 86964 247184 87016
rect 247236 87004 247242 87016
rect 250769 87007 250827 87013
rect 250769 87004 250781 87007
rect 247236 86976 250781 87004
rect 247236 86964 247242 86976
rect 250769 86973 250781 86976
rect 250815 86973 250827 87007
rect 250769 86967 250827 86973
rect 251042 86964 251048 87016
rect 251100 87004 251106 87016
rect 257206 87004 257212 87016
rect 251100 86976 257212 87004
rect 251100 86964 251106 86976
rect 257206 86964 257212 86976
rect 257264 86964 257270 87016
rect 52506 86896 52512 86948
rect 52564 86936 52570 86948
rect 64282 86936 64288 86948
rect 52564 86908 64288 86936
rect 52564 86896 52570 86908
rect 64282 86896 64288 86908
rect 64340 86896 64346 86948
rect 152234 86896 152240 86948
rect 152292 86936 152298 86948
rect 157389 86939 157447 86945
rect 157389 86936 157401 86939
rect 152292 86908 157401 86936
rect 152292 86896 152298 86908
rect 157389 86905 157401 86908
rect 157435 86905 157447 86939
rect 157389 86899 157447 86905
rect 157481 86939 157539 86945
rect 157481 86905 157493 86939
rect 157527 86936 157539 86939
rect 157846 86936 157852 86948
rect 157527 86908 157852 86936
rect 157527 86905 157539 86908
rect 157481 86899 157539 86905
rect 157846 86896 157852 86908
rect 157904 86896 157910 86948
rect 246994 86896 247000 86948
rect 247052 86936 247058 86948
rect 251229 86939 251287 86945
rect 251229 86936 251241 86939
rect 247052 86908 251241 86936
rect 247052 86896 247058 86908
rect 251229 86905 251241 86908
rect 251275 86905 251287 86939
rect 251229 86899 251287 86905
rect 251318 86896 251324 86948
rect 251376 86936 251382 86948
rect 257574 86936 257580 86948
rect 251376 86908 257580 86936
rect 251376 86896 251382 86908
rect 257574 86896 257580 86908
rect 257632 86896 257638 86948
rect 49838 86828 49844 86880
rect 49896 86868 49902 86880
rect 63086 86868 63092 86880
rect 49896 86840 63092 86868
rect 49896 86828 49902 86840
rect 63086 86828 63092 86840
rect 63144 86828 63150 86880
rect 63638 86828 63644 86880
rect 63696 86868 63702 86880
rect 70630 86868 70636 86880
rect 63696 86840 70636 86868
rect 63696 86828 63702 86840
rect 70630 86828 70636 86840
rect 70688 86828 70694 86880
rect 149106 86828 149112 86880
rect 149164 86868 149170 86880
rect 157754 86868 157760 86880
rect 149164 86840 157760 86868
rect 149164 86828 149170 86840
rect 157754 86828 157760 86840
rect 157812 86828 157818 86880
rect 158858 86828 158864 86880
rect 158916 86868 158922 86880
rect 164654 86868 164660 86880
rect 158916 86840 164660 86868
rect 158916 86828 158922 86840
rect 164654 86828 164660 86840
rect 164712 86828 164718 86880
rect 245706 86828 245712 86880
rect 245764 86868 245770 86880
rect 256194 86868 256200 86880
rect 245764 86840 256200 86868
rect 245764 86828 245770 86840
rect 256194 86828 256200 86840
rect 256252 86828 256258 86880
rect 51126 86760 51132 86812
rect 51184 86800 51190 86812
rect 58949 86803 59007 86809
rect 58949 86800 58961 86803
rect 51184 86772 58961 86800
rect 51184 86760 51190 86772
rect 58949 86769 58961 86772
rect 58995 86769 59007 86803
rect 58949 86763 59007 86769
rect 59038 86760 59044 86812
rect 59096 86800 59102 86812
rect 66766 86800 66772 86812
rect 59096 86772 66772 86800
rect 59096 86760 59102 86772
rect 66766 86760 66772 86772
rect 66824 86760 66830 86812
rect 156006 86760 156012 86812
rect 156064 86800 156070 86812
rect 158674 86800 158680 86812
rect 156064 86772 158680 86800
rect 156064 86760 156070 86772
rect 158674 86760 158680 86772
rect 158732 86760 158738 86812
rect 245338 86760 245344 86812
rect 245396 86800 245402 86812
rect 256102 86800 256108 86812
rect 245396 86772 256108 86800
rect 245396 86760 245402 86772
rect 256102 86760 256108 86772
rect 256160 86760 256166 86812
rect 57474 86692 57480 86744
rect 57532 86732 57538 86744
rect 61798 86732 61804 86744
rect 57532 86704 61804 86732
rect 57532 86692 57538 86704
rect 61798 86692 61804 86704
rect 61856 86692 61862 86744
rect 153338 86692 153344 86744
rect 153396 86732 153402 86744
rect 155549 86735 155607 86741
rect 155549 86732 155561 86735
rect 153396 86704 155561 86732
rect 153396 86692 153402 86704
rect 155549 86701 155561 86704
rect 155595 86701 155607 86735
rect 155549 86695 155607 86701
rect 155638 86692 155644 86744
rect 155696 86732 155702 86744
rect 159502 86732 159508 86744
rect 155696 86704 159508 86732
rect 155696 86692 155702 86704
rect 159502 86692 159508 86704
rect 159560 86692 159566 86744
rect 245154 86692 245160 86744
rect 245212 86732 245218 86744
rect 251134 86732 251140 86744
rect 245212 86704 251140 86732
rect 245212 86692 245218 86704
rect 251134 86692 251140 86704
rect 251192 86692 251198 86744
rect 251505 86735 251563 86741
rect 251505 86701 251517 86735
rect 251551 86732 251563 86735
rect 254262 86732 254268 86744
rect 251551 86704 254268 86732
rect 251551 86701 251563 86704
rect 251505 86695 251563 86701
rect 254262 86692 254268 86704
rect 254320 86692 254326 86744
rect 61338 86624 61344 86676
rect 61396 86664 61402 86676
rect 69802 86664 69808 86676
rect 61396 86636 69808 86664
rect 61396 86624 61402 86636
rect 69802 86624 69808 86636
rect 69860 86624 69866 86676
rect 150578 86624 150584 86676
rect 150636 86664 150642 86676
rect 150636 86636 155776 86664
rect 150636 86624 150642 86636
rect 60878 86556 60884 86608
rect 60936 86596 60942 86608
rect 69434 86596 69440 86608
rect 60936 86568 69440 86596
rect 60936 86556 60942 86568
rect 69434 86556 69440 86568
rect 69492 86556 69498 86608
rect 150670 86556 150676 86608
rect 150728 86596 150734 86608
rect 155362 86596 155368 86608
rect 150728 86568 155368 86596
rect 150728 86556 150734 86568
rect 155362 86556 155368 86568
rect 155420 86556 155426 86608
rect 57014 86488 57020 86540
rect 57072 86528 57078 86540
rect 61706 86528 61712 86540
rect 57072 86500 61712 86528
rect 57072 86488 57078 86500
rect 61706 86488 61712 86500
rect 61764 86488 61770 86540
rect 61982 86488 61988 86540
rect 62040 86528 62046 86540
rect 69894 86528 69900 86540
rect 62040 86500 69900 86528
rect 62040 86488 62046 86500
rect 69894 86488 69900 86500
rect 69952 86488 69958 86540
rect 155178 86488 155184 86540
rect 155236 86528 155242 86540
rect 155748 86528 155776 86636
rect 156098 86624 156104 86676
rect 156156 86664 156162 86676
rect 162630 86664 162636 86676
rect 156156 86636 162636 86664
rect 156156 86624 156162 86636
rect 162630 86624 162636 86636
rect 162688 86624 162694 86676
rect 247914 86624 247920 86676
rect 247972 86664 247978 86676
rect 251594 86664 251600 86676
rect 247972 86636 251600 86664
rect 247972 86624 247978 86636
rect 251594 86624 251600 86636
rect 251652 86624 251658 86676
rect 252698 86624 252704 86676
rect 252756 86664 252762 86676
rect 258310 86664 258316 86676
rect 252756 86636 258316 86664
rect 252756 86624 252762 86636
rect 258310 86624 258316 86636
rect 258368 86624 258374 86676
rect 155914 86556 155920 86608
rect 155972 86596 155978 86608
rect 163090 86596 163096 86608
rect 155972 86568 163096 86596
rect 155972 86556 155978 86568
rect 163090 86556 163096 86568
rect 163148 86556 163154 86608
rect 247822 86556 247828 86608
rect 247880 86596 247886 86608
rect 251502 86596 251508 86608
rect 247880 86568 251508 86596
rect 247880 86556 247886 86568
rect 251502 86556 251508 86568
rect 251560 86556 251566 86608
rect 156561 86531 156619 86537
rect 156561 86528 156573 86531
rect 155236 86500 155684 86528
rect 155748 86500 156573 86528
rect 155236 86488 155242 86500
rect 59406 86420 59412 86472
rect 59464 86460 59470 86472
rect 67318 86460 67324 86472
rect 59464 86432 67324 86460
rect 59464 86420 59470 86432
rect 67318 86420 67324 86432
rect 67376 86420 67382 86472
rect 151038 86420 151044 86472
rect 151096 86460 151102 86472
rect 155546 86460 155552 86472
rect 151096 86432 155552 86460
rect 151096 86420 151102 86432
rect 155546 86420 155552 86432
rect 155604 86420 155610 86472
rect 155656 86460 155684 86500
rect 156561 86497 156573 86500
rect 156607 86497 156619 86531
rect 156561 86491 156619 86497
rect 156650 86488 156656 86540
rect 156708 86528 156714 86540
rect 159778 86528 159784 86540
rect 156708 86500 159784 86528
rect 156708 86488 156714 86500
rect 159778 86488 159784 86500
rect 159836 86488 159842 86540
rect 244878 86488 244884 86540
rect 244936 86528 244942 86540
rect 249478 86528 249484 86540
rect 244936 86500 249484 86528
rect 244936 86488 244942 86500
rect 249478 86488 249484 86500
rect 249536 86488 249542 86540
rect 250950 86488 250956 86540
rect 251008 86528 251014 86540
rect 251226 86528 251232 86540
rect 251008 86500 251232 86528
rect 251008 86488 251014 86500
rect 251226 86488 251232 86500
rect 251284 86488 251290 86540
rect 156837 86463 156895 86469
rect 155656 86432 156788 86460
rect 57842 86352 57848 86404
rect 57900 86392 57906 86404
rect 61614 86392 61620 86404
rect 57900 86364 61620 86392
rect 57900 86352 57906 86364
rect 61614 86352 61620 86364
rect 61672 86352 61678 86404
rect 61890 86352 61896 86404
rect 61948 86392 61954 86404
rect 65846 86392 65852 86404
rect 61948 86364 65852 86392
rect 61948 86352 61954 86364
rect 65846 86352 65852 86364
rect 65904 86352 65910 86404
rect 153430 86352 153436 86404
rect 153488 86392 153494 86404
rect 156650 86392 156656 86404
rect 153488 86364 156656 86392
rect 153488 86352 153494 86364
rect 156650 86352 156656 86364
rect 156708 86352 156714 86404
rect 55818 86284 55824 86336
rect 55876 86324 55882 86336
rect 60510 86324 60516 86336
rect 55876 86296 60516 86324
rect 55876 86284 55882 86296
rect 60510 86284 60516 86296
rect 60568 86284 60574 86336
rect 61062 86284 61068 86336
rect 61120 86324 61126 86336
rect 61982 86324 61988 86336
rect 61120 86296 61988 86324
rect 61120 86284 61126 86296
rect 61982 86284 61988 86296
rect 62040 86284 62046 86336
rect 62258 86284 62264 86336
rect 62316 86324 62322 86336
rect 70262 86324 70268 86336
rect 62316 86296 70268 86324
rect 62316 86284 62322 86296
rect 70262 86284 70268 86296
rect 70320 86284 70326 86336
rect 151498 86284 151504 86336
rect 151556 86324 151562 86336
rect 155454 86324 155460 86336
rect 151556 86296 155460 86324
rect 151556 86284 151562 86296
rect 155454 86284 155460 86296
rect 155512 86284 155518 86336
rect 156760 86324 156788 86432
rect 156837 86429 156849 86463
rect 156883 86460 156895 86463
rect 157205 86463 157263 86469
rect 157205 86460 157217 86463
rect 156883 86432 157217 86460
rect 156883 86429 156895 86432
rect 156837 86423 156895 86429
rect 157205 86429 157217 86432
rect 157251 86429 157263 86463
rect 157205 86423 157263 86429
rect 157386 86420 157392 86472
rect 157444 86460 157450 86472
rect 163826 86460 163832 86472
rect 157444 86432 163832 86460
rect 157444 86420 157450 86432
rect 163826 86420 163832 86432
rect 163884 86420 163890 86472
rect 248926 86420 248932 86472
rect 248984 86460 248990 86472
rect 251410 86460 251416 86472
rect 248984 86432 251416 86460
rect 248984 86420 248990 86432
rect 251410 86420 251416 86432
rect 251468 86420 251474 86472
rect 157478 86352 157484 86404
rect 157536 86392 157542 86404
rect 164286 86392 164292 86404
rect 157536 86364 164292 86392
rect 157536 86352 157542 86364
rect 164286 86352 164292 86364
rect 164344 86352 164350 86404
rect 249386 86352 249392 86404
rect 249444 86392 249450 86404
rect 252422 86392 252428 86404
rect 249444 86364 252428 86392
rect 249444 86352 249450 86364
rect 252422 86352 252428 86364
rect 252480 86352 252486 86404
rect 163458 86324 163464 86336
rect 156760 86296 163464 86324
rect 163458 86284 163464 86296
rect 163516 86284 163522 86336
rect 243314 86284 243320 86336
rect 243372 86324 243378 86336
rect 248374 86324 248380 86336
rect 243372 86296 248380 86324
rect 243372 86284 243378 86296
rect 248374 86284 248380 86296
rect 248432 86284 248438 86336
rect 249110 86284 249116 86336
rect 249168 86324 249174 86336
rect 249846 86324 249852 86336
rect 249168 86296 249852 86324
rect 249168 86284 249174 86296
rect 249846 86284 249852 86296
rect 249904 86284 249910 86336
rect 250674 86284 250680 86336
rect 250732 86324 250738 86336
rect 253618 86324 253624 86336
rect 250732 86296 253624 86324
rect 250732 86284 250738 86296
rect 253618 86284 253624 86296
rect 253676 86284 253682 86336
rect 55450 86216 55456 86268
rect 55508 86256 55514 86268
rect 60326 86256 60332 86268
rect 55508 86228 60332 86256
rect 55508 86216 55514 86228
rect 60326 86216 60332 86228
rect 60384 86216 60390 86268
rect 64374 86216 64380 86268
rect 64432 86256 64438 86268
rect 67410 86256 67416 86268
rect 64432 86228 67416 86256
rect 64432 86216 64438 86228
rect 67410 86216 67416 86228
rect 67468 86216 67474 86268
rect 154258 86216 154264 86268
rect 154316 86256 154322 86268
rect 157018 86256 157024 86268
rect 154316 86228 157024 86256
rect 154316 86216 154322 86228
rect 157018 86216 157024 86228
rect 157076 86216 157082 86268
rect 157110 86216 157116 86268
rect 157168 86256 157174 86268
rect 159870 86256 159876 86268
rect 157168 86228 159876 86256
rect 157168 86216 157174 86228
rect 159870 86216 159876 86228
rect 159928 86216 159934 86268
rect 244418 86216 244424 86268
rect 244476 86256 244482 86268
rect 248282 86256 248288 86268
rect 244476 86228 248288 86256
rect 244476 86216 244482 86228
rect 248282 86216 248288 86228
rect 248340 86216 248346 86268
rect 249570 86216 249576 86268
rect 249628 86256 249634 86268
rect 251962 86256 251968 86268
rect 249628 86228 251968 86256
rect 249628 86216 249634 86228
rect 251962 86216 251968 86228
rect 252020 86216 252026 86268
rect 252606 86216 252612 86268
rect 252664 86256 252670 86268
rect 258402 86256 258408 86268
rect 252664 86228 258408 86256
rect 252664 86216 252670 86228
rect 258402 86216 258408 86228
rect 258460 86216 258466 86268
rect 56278 86148 56284 86200
rect 56336 86188 56342 86200
rect 60418 86188 60424 86200
rect 56336 86160 60424 86188
rect 56336 86148 56342 86160
rect 60418 86148 60424 86160
rect 60476 86148 60482 86200
rect 61982 86148 61988 86200
rect 62040 86188 62046 86200
rect 65018 86188 65024 86200
rect 62040 86160 65024 86188
rect 62040 86148 62046 86160
rect 65018 86148 65024 86160
rect 65076 86148 65082 86200
rect 65754 86148 65760 86200
rect 65812 86188 65818 86200
rect 67042 86188 67048 86200
rect 65812 86160 67048 86188
rect 65812 86148 65818 86160
rect 67042 86148 67048 86160
rect 67100 86148 67106 86200
rect 154626 86148 154632 86200
rect 154684 86188 154690 86200
rect 156926 86188 156932 86200
rect 154684 86160 156932 86188
rect 154684 86148 154690 86160
rect 156926 86148 156932 86160
rect 156984 86148 156990 86200
rect 157202 86148 157208 86200
rect 157260 86188 157266 86200
rect 160238 86188 160244 86200
rect 157260 86160 160244 86188
rect 157260 86148 157266 86160
rect 160238 86148 160244 86160
rect 160296 86148 160302 86200
rect 243682 86148 243688 86200
rect 243740 86188 243746 86200
rect 248006 86188 248012 86200
rect 243740 86160 248012 86188
rect 243740 86148 243746 86160
rect 248006 86148 248012 86160
rect 248064 86148 248070 86200
rect 249294 86148 249300 86200
rect 249352 86188 249358 86200
rect 249846 86188 249852 86200
rect 249352 86160 249852 86188
rect 249352 86148 249358 86160
rect 249846 86148 249852 86160
rect 249904 86148 249910 86200
rect 252790 86188 252796 86200
rect 249956 86160 252796 86188
rect 56646 86080 56652 86132
rect 56704 86120 56710 86132
rect 60234 86120 60240 86132
rect 56704 86092 60240 86120
rect 56704 86080 56710 86092
rect 60234 86080 60240 86092
rect 60292 86080 60298 86132
rect 62626 86080 62632 86132
rect 62684 86120 62690 86132
rect 63546 86120 63552 86132
rect 62684 86092 63552 86120
rect 62684 86080 62690 86092
rect 63546 86080 63552 86092
rect 63604 86080 63610 86132
rect 65846 86080 65852 86132
rect 65904 86120 65910 86132
rect 66674 86120 66680 86132
rect 65904 86092 66680 86120
rect 65904 86080 65910 86092
rect 66674 86080 66680 86092
rect 66732 86080 66738 86132
rect 66766 86080 66772 86132
rect 66824 86120 66830 86132
rect 67410 86120 67416 86132
rect 66824 86092 67416 86120
rect 66824 86080 66830 86092
rect 67410 86080 67416 86092
rect 67468 86080 67474 86132
rect 67502 86080 67508 86132
rect 67560 86120 67566 86132
rect 69066 86120 69072 86132
rect 67560 86092 69072 86120
rect 67560 86080 67566 86092
rect 69066 86080 69072 86092
rect 69124 86080 69130 86132
rect 149474 86080 149480 86132
rect 149532 86120 149538 86132
rect 150486 86120 150492 86132
rect 149532 86092 150492 86120
rect 149532 86080 149538 86092
rect 150486 86080 150492 86092
rect 150544 86080 150550 86132
rect 153890 86080 153896 86132
rect 153948 86120 153954 86132
rect 154718 86120 154724 86132
rect 153948 86092 154724 86120
rect 153948 86080 153954 86092
rect 154718 86080 154724 86092
rect 154776 86080 154782 86132
rect 155086 86080 155092 86132
rect 155144 86120 155150 86132
rect 155822 86120 155828 86132
rect 155144 86092 155828 86120
rect 155144 86080 155150 86092
rect 155822 86080 155828 86092
rect 155880 86080 155886 86132
rect 156282 86080 156288 86132
rect 156340 86120 156346 86132
rect 157294 86120 157300 86132
rect 156340 86092 157300 86120
rect 156340 86080 156346 86092
rect 157294 86080 157300 86092
rect 157352 86080 157358 86132
rect 157389 86123 157447 86129
rect 157389 86089 157401 86123
rect 157435 86120 157447 86123
rect 158306 86120 158312 86132
rect 157435 86092 158312 86120
rect 157435 86089 157447 86092
rect 157389 86083 157447 86089
rect 158306 86080 158312 86092
rect 158364 86080 158370 86132
rect 159686 86080 159692 86132
rect 159744 86120 159750 86132
rect 161434 86120 161440 86132
rect 159744 86092 161440 86120
rect 159744 86080 159750 86092
rect 161434 86080 161440 86092
rect 161492 86080 161498 86132
rect 244142 86080 244148 86132
rect 244200 86120 244206 86132
rect 248190 86120 248196 86132
rect 244200 86092 248196 86120
rect 244200 86080 244206 86092
rect 248190 86080 248196 86092
rect 248248 86080 248254 86132
rect 249956 86120 249984 86160
rect 252790 86148 252796 86160
rect 252848 86148 252854 86200
rect 253434 86148 253440 86200
rect 253492 86188 253498 86200
rect 255182 86188 255188 86200
rect 253492 86160 255188 86188
rect 253492 86148 253498 86160
rect 255182 86148 255188 86160
rect 255240 86148 255246 86200
rect 249312 86092 249984 86120
rect 249312 86064 249340 86092
rect 250766 86080 250772 86132
rect 250824 86120 250830 86132
rect 253158 86120 253164 86132
rect 250824 86092 253164 86120
rect 250824 86080 250830 86092
rect 253158 86080 253164 86092
rect 253216 86080 253222 86132
rect 253526 86080 253532 86132
rect 253584 86120 253590 86132
rect 254814 86120 254820 86132
rect 253584 86092 254820 86120
rect 253584 86080 253590 86092
rect 254814 86080 254820 86092
rect 254872 86080 254878 86132
rect 255550 86080 255556 86132
rect 255608 86120 255614 86132
rect 256378 86120 256384 86132
rect 255608 86092 256384 86120
rect 255608 86080 255614 86092
rect 256378 86080 256384 86092
rect 256436 86080 256442 86132
rect 231630 86012 231636 86064
rect 231688 86052 231694 86064
rect 236322 86052 236328 86064
rect 231688 86024 236328 86052
rect 231688 86012 231694 86024
rect 236322 86012 236328 86024
rect 236380 86012 236386 86064
rect 249294 86012 249300 86064
rect 249352 86012 249358 86064
rect 256010 85876 256016 85928
rect 256068 85916 256074 85928
rect 256194 85916 256200 85928
rect 256068 85888 256200 85916
rect 256068 85876 256074 85888
rect 256194 85876 256200 85888
rect 256252 85876 256258 85928
rect 256286 85604 256292 85656
rect 256344 85644 256350 85656
rect 256562 85644 256568 85656
rect 256344 85616 256568 85644
rect 256344 85604 256350 85616
rect 256562 85604 256568 85616
rect 256620 85604 256626 85656
rect 136870 85196 136876 85248
rect 136928 85236 136934 85248
rect 143678 85236 143684 85248
rect 136928 85208 143684 85236
rect 136928 85196 136934 85208
rect 143678 85196 143684 85208
rect 143736 85196 143742 85248
rect 136870 84652 136876 84704
rect 136928 84692 136934 84704
rect 143494 84692 143500 84704
rect 136928 84664 143500 84692
rect 136928 84652 136934 84664
rect 143494 84652 143500 84664
rect 143552 84652 143558 84704
rect 231630 84652 231636 84704
rect 231688 84692 231694 84704
rect 236230 84692 236236 84704
rect 231688 84664 236236 84692
rect 231688 84652 231694 84664
rect 236230 84652 236236 84664
rect 236288 84652 236294 84704
rect 155546 84244 155552 84296
rect 155604 84284 155610 84296
rect 160422 84284 160428 84296
rect 155604 84256 160428 84284
rect 155604 84244 155610 84256
rect 160422 84244 160428 84256
rect 160480 84244 160486 84296
rect 300354 84284 300360 84296
rect 182152 84256 300360 84284
rect 92250 83972 92256 84024
rect 92308 84012 92314 84024
rect 96669 84015 96727 84021
rect 96669 84012 96681 84015
rect 92308 83984 96681 84012
rect 92308 83972 92314 83984
rect 96669 83981 96681 83984
rect 96715 83981 96727 84015
rect 96669 83975 96727 83981
rect 89582 83904 89588 83956
rect 89640 83944 89646 83956
rect 89769 83947 89827 83953
rect 89769 83944 89781 83947
rect 89640 83916 89781 83944
rect 89640 83904 89646 83916
rect 89769 83913 89781 83916
rect 89815 83913 89827 83947
rect 89769 83907 89827 83913
rect 90870 83904 90876 83956
rect 90928 83944 90934 83956
rect 90928 83916 96160 83944
rect 90928 83904 90934 83916
rect 67870 83836 67876 83888
rect 67928 83876 67934 83888
rect 68238 83876 68244 83888
rect 67928 83848 68244 83876
rect 67928 83836 67934 83848
rect 68238 83836 68244 83848
rect 68296 83836 68302 83888
rect 86822 83876 86828 83888
rect 86783 83848 86828 83876
rect 86822 83836 86828 83848
rect 86880 83836 86886 83888
rect 88202 83836 88208 83888
rect 88260 83876 88266 83888
rect 93630 83876 93636 83888
rect 88260 83848 92020 83876
rect 93591 83848 93636 83876
rect 88260 83836 88266 83848
rect 91992 83820 92020 83848
rect 93630 83836 93636 83848
rect 93688 83836 93694 83888
rect 94918 83876 94924 83888
rect 94879 83848 94924 83876
rect 94918 83836 94924 83848
rect 94976 83836 94982 83888
rect 96132 83820 96160 83916
rect 116538 83904 116544 83956
rect 116596 83904 116602 83956
rect 120586 83944 120592 83956
rect 120547 83916 120592 83944
rect 120586 83904 120592 83916
rect 120644 83904 120650 83956
rect 124634 83904 124640 83956
rect 124692 83944 124698 83956
rect 124729 83947 124787 83953
rect 124729 83944 124741 83947
rect 124692 83916 124741 83944
rect 124692 83904 124698 83916
rect 124729 83913 124741 83916
rect 124775 83913 124787 83947
rect 124729 83907 124787 83913
rect 127302 83904 127308 83956
rect 127360 83944 127366 83956
rect 134846 83944 134852 83956
rect 127360 83916 134852 83944
rect 127360 83904 127366 83916
rect 134846 83904 134852 83916
rect 134904 83904 134910 83956
rect 96298 83836 96304 83888
rect 96356 83836 96362 83888
rect 97678 83836 97684 83888
rect 97736 83876 97742 83888
rect 97736 83848 97816 83876
rect 97736 83836 97742 83848
rect 91974 83768 91980 83820
rect 92032 83768 92038 83820
rect 96114 83768 96120 83820
rect 96172 83768 96178 83820
rect 96316 83740 96344 83836
rect 97788 83752 97816 83848
rect 98966 83836 98972 83888
rect 99024 83876 99030 83888
rect 99024 83848 99564 83876
rect 99024 83836 99030 83848
rect 99536 83820 99564 83848
rect 100346 83836 100352 83888
rect 100404 83876 100410 83888
rect 100404 83848 100944 83876
rect 100404 83836 100410 83848
rect 100916 83820 100944 83848
rect 101726 83836 101732 83888
rect 101784 83876 101790 83888
rect 101784 83848 102324 83876
rect 101784 83836 101790 83848
rect 102296 83820 102324 83848
rect 103014 83836 103020 83888
rect 103072 83876 103078 83888
rect 103072 83848 103704 83876
rect 103072 83836 103078 83848
rect 103676 83820 103704 83848
rect 104394 83836 104400 83888
rect 104452 83876 104458 83888
rect 104452 83848 105084 83876
rect 104452 83836 104458 83848
rect 105056 83820 105084 83848
rect 105774 83836 105780 83888
rect 105832 83876 105838 83888
rect 105832 83848 106464 83876
rect 105832 83836 105838 83848
rect 106436 83820 106464 83848
rect 107062 83836 107068 83888
rect 107120 83876 107126 83888
rect 107120 83848 107844 83876
rect 107120 83836 107126 83848
rect 107816 83820 107844 83848
rect 108442 83836 108448 83888
rect 108500 83836 108506 83888
rect 109822 83876 109828 83888
rect 109783 83848 109828 83876
rect 109822 83836 109828 83848
rect 109880 83836 109886 83888
rect 111110 83836 111116 83888
rect 111168 83876 111174 83888
rect 111205 83879 111263 83885
rect 111205 83876 111217 83879
rect 111168 83848 111217 83876
rect 111168 83836 111174 83848
rect 111205 83845 111217 83848
rect 111251 83845 111263 83879
rect 112490 83876 112496 83888
rect 112451 83848 112496 83876
rect 111205 83839 111263 83845
rect 112490 83836 112496 83848
rect 112548 83836 112554 83888
rect 113870 83836 113876 83888
rect 113928 83876 113934 83888
rect 115158 83876 115164 83888
rect 113928 83848 114008 83876
rect 115119 83848 115164 83876
rect 113928 83836 113934 83848
rect 99518 83768 99524 83820
rect 99576 83768 99582 83820
rect 100898 83768 100904 83820
rect 100956 83768 100962 83820
rect 102278 83768 102284 83820
rect 102336 83768 102342 83820
rect 103658 83768 103664 83820
rect 103716 83768 103722 83820
rect 105038 83768 105044 83820
rect 105096 83768 105102 83820
rect 106418 83768 106424 83820
rect 106476 83768 106482 83820
rect 107798 83768 107804 83820
rect 107856 83768 107862 83820
rect 108460 83808 108488 83836
rect 112950 83808 112956 83820
rect 108460 83780 112956 83808
rect 112950 83768 112956 83780
rect 113008 83768 113014 83820
rect 113980 83752 114008 83848
rect 115158 83836 115164 83848
rect 115216 83836 115222 83888
rect 96390 83740 96396 83752
rect 96316 83712 96396 83740
rect 96390 83700 96396 83712
rect 96448 83700 96454 83752
rect 97770 83700 97776 83752
rect 97828 83700 97834 83752
rect 113962 83700 113968 83752
rect 114020 83700 114026 83752
rect 116556 83740 116584 83904
rect 117918 83876 117924 83888
rect 117879 83848 117924 83876
rect 117918 83836 117924 83848
rect 117976 83836 117982 83888
rect 119206 83836 119212 83888
rect 119264 83876 119270 83888
rect 119264 83848 119344 83876
rect 119264 83836 119270 83848
rect 119316 83752 119344 83848
rect 121966 83836 121972 83888
rect 122024 83836 122030 83888
rect 123254 83876 123260 83888
rect 123215 83848 123260 83876
rect 123254 83836 123260 83848
rect 123312 83836 123318 83888
rect 126014 83876 126020 83888
rect 125975 83848 126020 83876
rect 126014 83836 126020 83848
rect 126072 83836 126078 83888
rect 128682 83876 128688 83888
rect 128643 83848 128688 83876
rect 128682 83836 128688 83848
rect 128740 83836 128746 83888
rect 132730 83836 132736 83888
rect 132788 83876 132794 83888
rect 132788 83848 133420 83876
rect 132788 83836 132794 83848
rect 121984 83808 122012 83836
rect 133392 83820 133420 83848
rect 182152 83820 182180 84256
rect 300354 84244 300360 84256
rect 300412 84244 300418 84296
rect 250490 83836 250496 83888
rect 250548 83876 250554 83888
rect 251134 83876 251140 83888
rect 250548 83848 251140 83876
rect 250548 83836 250554 83848
rect 251134 83836 251140 83848
rect 251192 83836 251198 83888
rect 125554 83808 125560 83820
rect 121984 83780 125560 83808
rect 125554 83768 125560 83780
rect 125612 83768 125618 83820
rect 133374 83768 133380 83820
rect 133432 83768 133438 83820
rect 182134 83768 182140 83820
rect 182192 83768 182198 83820
rect 116630 83740 116636 83752
rect 116556 83712 116636 83740
rect 116630 83700 116636 83712
rect 116688 83700 116694 83752
rect 119298 83700 119304 83752
rect 119356 83700 119362 83752
rect 85074 81932 85080 81984
rect 85132 81972 85138 81984
rect 179558 81972 179564 81984
rect 85132 81944 179564 81972
rect 85132 81932 85138 81944
rect 179558 81932 179564 81944
rect 179616 81932 179622 81984
rect 186274 81932 186280 81984
rect 186332 81972 186338 81984
rect 194094 81972 194100 81984
rect 186332 81944 194100 81972
rect 186332 81932 186338 81944
rect 194094 81932 194100 81944
rect 194152 81932 194158 81984
rect 196949 81975 197007 81981
rect 196949 81941 196961 81975
rect 196995 81972 197007 81975
rect 203846 81972 203852 81984
rect 196995 81944 203852 81972
rect 196995 81941 197007 81944
rect 196949 81935 197007 81941
rect 203846 81932 203852 81944
rect 203904 81932 203910 81984
rect 96669 81907 96727 81913
rect 96669 81873 96681 81907
rect 96715 81904 96727 81907
rect 99610 81904 99616 81916
rect 96715 81876 99616 81904
rect 96715 81873 96727 81876
rect 96669 81867 96727 81873
rect 99610 81864 99616 81876
rect 99668 81864 99674 81916
rect 99705 81907 99763 81913
rect 99705 81873 99717 81907
rect 99751 81904 99763 81907
rect 109825 81907 109883 81913
rect 109825 81904 109837 81907
rect 99751 81876 109837 81904
rect 99751 81873 99763 81876
rect 99705 81867 99763 81873
rect 109825 81873 109837 81876
rect 109871 81873 109883 81907
rect 109825 81867 109883 81873
rect 133374 81864 133380 81916
rect 133432 81904 133438 81916
rect 226754 81904 226760 81916
rect 133432 81876 226760 81904
rect 133432 81864 133438 81876
rect 226754 81864 226760 81876
rect 226812 81864 226818 81916
rect 86825 81839 86883 81845
rect 86825 81805 86837 81839
rect 86871 81836 86883 81839
rect 89214 81836 89220 81848
rect 86871 81808 89220 81836
rect 86871 81805 86883 81808
rect 86825 81799 86883 81805
rect 89214 81796 89220 81808
rect 89272 81796 89278 81848
rect 93633 81839 93691 81845
rect 93633 81805 93645 81839
rect 93679 81836 93691 81839
rect 100165 81839 100223 81845
rect 100165 81836 100177 81839
rect 93679 81808 100177 81836
rect 93679 81805 93691 81808
rect 93633 81799 93691 81805
rect 100165 81805 100177 81808
rect 100211 81805 100223 81839
rect 112493 81839 112551 81845
rect 112493 81836 112505 81839
rect 100165 81799 100223 81805
rect 100272 81808 112505 81836
rect 79554 81728 79560 81780
rect 79612 81768 79618 81780
rect 99613 81771 99671 81777
rect 99613 81768 99625 81771
rect 79612 81740 99625 81768
rect 79612 81728 79618 81740
rect 99613 81737 99625 81740
rect 99659 81737 99671 81771
rect 99613 81731 99671 81737
rect 79738 81660 79744 81712
rect 79796 81700 79802 81712
rect 100272 81700 100300 81808
rect 112493 81805 112505 81808
rect 112539 81805 112551 81839
rect 112493 81799 112551 81805
rect 174038 81728 174044 81780
rect 174096 81768 174102 81780
rect 196949 81771 197007 81777
rect 196949 81768 196961 81771
rect 174096 81740 196961 81768
rect 174096 81728 174102 81740
rect 196949 81737 196961 81740
rect 196995 81737 197007 81771
rect 196949 81731 197007 81737
rect 197038 81728 197044 81780
rect 197096 81768 197102 81780
rect 197498 81768 197504 81780
rect 197096 81740 197504 81768
rect 197096 81728 197102 81740
rect 197498 81728 197504 81740
rect 197556 81728 197562 81780
rect 198418 81728 198424 81780
rect 198476 81768 198482 81780
rect 198878 81768 198884 81780
rect 198476 81740 198884 81768
rect 198476 81728 198482 81740
rect 198878 81728 198884 81740
rect 198936 81728 198942 81780
rect 199798 81728 199804 81780
rect 199856 81768 199862 81780
rect 200258 81768 200264 81780
rect 199856 81740 200264 81768
rect 199856 81728 199862 81740
rect 200258 81728 200264 81740
rect 200316 81728 200322 81780
rect 201086 81728 201092 81780
rect 201144 81768 201150 81780
rect 201638 81768 201644 81780
rect 201144 81740 201644 81768
rect 201144 81728 201150 81740
rect 201638 81728 201644 81740
rect 201696 81728 201702 81780
rect 79796 81672 100300 81700
rect 79796 81660 79802 81672
rect 173762 81660 173768 81712
rect 173820 81700 173826 81712
rect 209182 81700 209188 81712
rect 173820 81672 209188 81700
rect 173820 81660 173826 81672
rect 209182 81660 209188 81672
rect 209240 81660 209246 81712
rect 79830 81592 79836 81644
rect 79888 81632 79894 81644
rect 115161 81635 115219 81641
rect 115161 81632 115173 81635
rect 79888 81604 115173 81632
rect 79888 81592 79894 81604
rect 115161 81601 115173 81604
rect 115207 81601 115219 81635
rect 115161 81595 115219 81601
rect 173486 81592 173492 81644
rect 173544 81632 173550 81644
rect 211942 81632 211948 81644
rect 173544 81604 211948 81632
rect 173544 81592 173550 81604
rect 211942 81592 211948 81604
rect 212000 81592 212006 81644
rect 79646 81524 79652 81576
rect 79704 81564 79710 81576
rect 117921 81567 117979 81573
rect 117921 81564 117933 81567
rect 79704 81536 117933 81564
rect 79704 81524 79710 81536
rect 117921 81533 117933 81536
rect 117967 81533 117979 81567
rect 117921 81527 117979 81533
rect 173854 81524 173860 81576
rect 173912 81564 173918 81576
rect 214610 81564 214616 81576
rect 173912 81536 214616 81564
rect 173912 81524 173918 81536
rect 214610 81524 214616 81536
rect 214668 81524 214674 81576
rect 79922 81456 79928 81508
rect 79980 81496 79986 81508
rect 120589 81499 120647 81505
rect 120589 81496 120601 81499
rect 79980 81468 120601 81496
rect 79980 81456 79986 81468
rect 120589 81465 120601 81468
rect 120635 81465 120647 81499
rect 120589 81459 120647 81465
rect 173670 81456 173676 81508
rect 173728 81496 173734 81508
rect 217278 81496 217284 81508
rect 173728 81468 217284 81496
rect 173728 81456 173734 81468
rect 217278 81456 217284 81468
rect 217336 81456 217342 81508
rect 80014 81388 80020 81440
rect 80072 81428 80078 81440
rect 123257 81431 123315 81437
rect 123257 81428 123269 81431
rect 80072 81400 123269 81428
rect 80072 81388 80078 81400
rect 123257 81397 123269 81400
rect 123303 81397 123315 81431
rect 123257 81391 123315 81397
rect 173946 81388 173952 81440
rect 174004 81428 174010 81440
rect 220038 81428 220044 81440
rect 174004 81400 220044 81428
rect 174004 81388 174010 81400
rect 220038 81388 220044 81400
rect 220096 81388 220102 81440
rect 221326 81388 221332 81440
rect 221384 81428 221390 81440
rect 264842 81428 264848 81440
rect 221384 81400 264848 81428
rect 221384 81388 221390 81400
rect 264842 81388 264848 81400
rect 264900 81388 264906 81440
rect 80106 81320 80112 81372
rect 80164 81360 80170 81372
rect 126017 81363 126075 81369
rect 126017 81360 126029 81363
rect 80164 81332 126029 81360
rect 80164 81320 80170 81332
rect 126017 81329 126029 81332
rect 126063 81329 126075 81363
rect 126017 81323 126075 81329
rect 173302 81320 173308 81372
rect 173360 81360 173366 81372
rect 222706 81360 222712 81372
rect 173360 81332 222712 81360
rect 173360 81320 173366 81332
rect 222706 81320 222712 81332
rect 222764 81320 222770 81372
rect 80198 81252 80204 81304
rect 80256 81292 80262 81304
rect 128685 81295 128743 81301
rect 128685 81292 128697 81295
rect 80256 81264 128697 81292
rect 80256 81252 80262 81264
rect 128685 81261 128697 81264
rect 128731 81261 128743 81295
rect 128685 81255 128743 81261
rect 173578 81252 173584 81304
rect 173636 81292 173642 81304
rect 206514 81292 206520 81304
rect 173636 81264 206520 81292
rect 173636 81252 173642 81264
rect 206514 81252 206520 81264
rect 206572 81252 206578 81304
rect 207894 81252 207900 81304
rect 207952 81292 207958 81304
rect 264750 81292 264756 81304
rect 207952 81264 264756 81292
rect 207952 81252 207958 81264
rect 264750 81252 264756 81264
rect 264808 81252 264814 81304
rect 99610 81184 99616 81236
rect 99668 81224 99674 81236
rect 100254 81224 100260 81236
rect 99668 81196 100260 81224
rect 99668 81184 99674 81196
rect 100254 81184 100260 81196
rect 100312 81184 100318 81236
rect 187654 81184 187660 81236
rect 187712 81224 187718 81236
rect 195566 81224 195572 81236
rect 187712 81196 195572 81224
rect 187712 81184 187718 81196
rect 195566 81184 195572 81196
rect 195624 81184 195630 81236
rect 100165 81159 100223 81165
rect 100165 81125 100177 81159
rect 100211 81156 100223 81159
rect 101726 81156 101732 81168
rect 100211 81128 101732 81156
rect 100211 81125 100223 81128
rect 100165 81119 100223 81125
rect 101726 81116 101732 81128
rect 101784 81116 101790 81168
rect 188942 81116 188948 81168
rect 189000 81156 189006 81168
rect 195474 81156 195480 81168
rect 189000 81128 195480 81156
rect 189000 81116 189006 81128
rect 195474 81116 195480 81128
rect 195532 81116 195538 81168
rect 94921 80751 94979 80757
rect 94921 80717 94933 80751
rect 94967 80748 94979 80751
rect 101634 80748 101640 80760
rect 94967 80720 101640 80748
rect 94967 80717 94979 80720
rect 94921 80711 94979 80717
rect 101634 80708 101640 80720
rect 101692 80708 101698 80760
rect 182226 80640 182232 80692
rect 182284 80680 182290 80692
rect 185814 80680 185820 80692
rect 182284 80652 185820 80680
rect 182284 80640 182290 80652
rect 185814 80640 185820 80652
rect 185872 80640 185878 80692
rect 180846 80572 180852 80624
rect 180904 80612 180910 80624
rect 183054 80612 183060 80624
rect 180904 80584 183060 80612
rect 180904 80572 180910 80584
rect 183054 80572 183060 80584
rect 183112 80572 183118 80624
rect 184894 80572 184900 80624
rect 184952 80612 184958 80624
rect 191334 80612 191340 80624
rect 184952 80584 191340 80612
rect 184952 80572 184958 80584
rect 191334 80572 191340 80584
rect 191392 80572 191398 80624
rect 134754 80504 134760 80556
rect 134812 80544 134818 80556
rect 167230 80544 167236 80556
rect 134812 80516 167236 80544
rect 134812 80504 134818 80516
rect 167230 80504 167236 80516
rect 167288 80504 167294 80556
rect 111202 80136 111208 80148
rect 111163 80108 111208 80136
rect 111202 80096 111208 80108
rect 111260 80096 111266 80148
rect 124726 80136 124732 80148
rect 124687 80108 124732 80136
rect 124726 80096 124732 80108
rect 124784 80096 124790 80148
rect 167230 79756 167236 79808
rect 167288 79796 167294 79808
rect 170174 79796 170180 79808
rect 167288 79768 170180 79796
rect 167288 79756 167294 79768
rect 170174 79756 170180 79768
rect 170232 79756 170238 79808
rect 155730 79416 155736 79468
rect 155788 79456 155794 79468
rect 156009 79459 156067 79465
rect 156009 79456 156021 79459
rect 155788 79428 156021 79456
rect 155788 79416 155794 79428
rect 156009 79425 156021 79428
rect 156055 79425 156067 79459
rect 156009 79419 156067 79425
rect 145334 79348 145340 79400
rect 145392 79388 145398 79400
rect 145978 79388 145984 79400
rect 145392 79360 145984 79388
rect 145392 79348 145398 79360
rect 145978 79348 145984 79360
rect 146036 79348 146042 79400
rect 257022 79348 257028 79400
rect 257080 79388 257086 79400
rect 257482 79388 257488 79400
rect 257080 79360 257488 79388
rect 257080 79348 257086 79360
rect 257482 79348 257488 79360
rect 257540 79348 257546 79400
rect 155362 79280 155368 79332
rect 155420 79320 155426 79332
rect 155420 79292 155684 79320
rect 155420 79280 155426 79292
rect 155656 79264 155684 79292
rect 155638 79212 155644 79264
rect 155696 79212 155702 79264
rect 50482 79144 50488 79196
rect 50540 79184 50546 79196
rect 51218 79184 51224 79196
rect 50540 79156 51224 79184
rect 50540 79144 50546 79156
rect 51218 79144 51224 79156
rect 51276 79144 51282 79196
rect 51770 79144 51776 79196
rect 51828 79184 51834 79196
rect 52506 79184 52512 79196
rect 51828 79156 52512 79184
rect 51828 79144 51834 79156
rect 52506 79144 52512 79156
rect 52564 79144 52570 79196
rect 56462 79144 56468 79196
rect 56520 79184 56526 79196
rect 56520 79156 62028 79184
rect 56520 79144 56526 79156
rect 54438 79008 54444 79060
rect 54496 79048 54502 79060
rect 61890 79048 61896 79060
rect 54496 79020 61896 79048
rect 54496 79008 54502 79020
rect 61890 79008 61896 79020
rect 61948 79008 61954 79060
rect 62000 79048 62028 79156
rect 62442 79144 62448 79196
rect 62500 79184 62506 79196
rect 63638 79184 63644 79196
rect 62500 79156 63644 79184
rect 62500 79144 62506 79156
rect 63638 79144 63644 79156
rect 63696 79144 63702 79196
rect 138986 79144 138992 79196
rect 139044 79184 139050 79196
rect 143218 79184 143224 79196
rect 139044 79156 143224 79184
rect 139044 79144 139050 79156
rect 143218 79144 143224 79156
rect 143276 79144 143282 79196
rect 158398 79144 158404 79196
rect 158456 79184 158462 79196
rect 162630 79184 162636 79196
rect 158456 79156 162636 79184
rect 158456 79144 158462 79156
rect 162630 79144 162636 79156
rect 162688 79144 162694 79196
rect 231354 79144 231360 79196
rect 231412 79184 231418 79196
rect 237610 79184 237616 79196
rect 231412 79156 237616 79184
rect 231412 79144 231418 79156
rect 237610 79144 237616 79156
rect 237668 79144 237674 79196
rect 238254 79144 238260 79196
rect 238312 79184 238318 79196
rect 239726 79184 239732 79196
rect 238312 79156 239732 79184
rect 238312 79144 238318 79156
rect 239726 79144 239732 79156
rect 239784 79144 239790 79196
rect 241566 79144 241572 79196
rect 241624 79184 241630 79196
rect 245154 79184 245160 79196
rect 241624 79156 245160 79184
rect 241624 79144 241630 79156
rect 245154 79144 245160 79156
rect 245212 79144 245218 79196
rect 246442 79144 246448 79196
rect 246500 79184 246506 79196
rect 246994 79184 247000 79196
rect 246500 79156 247000 79184
rect 246500 79144 246506 79156
rect 246994 79144 247000 79156
rect 247052 79144 247058 79196
rect 249754 79144 249760 79196
rect 249812 79184 249818 79196
rect 255550 79184 255556 79196
rect 249812 79156 255556 79184
rect 249812 79144 249818 79156
rect 255550 79144 255556 79156
rect 255608 79144 255614 79196
rect 256378 79144 256384 79196
rect 256436 79184 256442 79196
rect 258678 79184 258684 79196
rect 256436 79156 258684 79184
rect 256436 79144 256442 79156
rect 258678 79144 258684 79156
rect 258736 79144 258742 79196
rect 264290 79144 264296 79196
rect 264348 79184 264354 79196
rect 265118 79184 265124 79196
rect 264348 79156 265124 79184
rect 264348 79144 264354 79156
rect 265118 79144 265124 79156
rect 265176 79144 265182 79196
rect 137514 79076 137520 79128
rect 137572 79116 137578 79128
rect 142758 79116 142764 79128
rect 137572 79088 142764 79116
rect 137572 79076 137578 79088
rect 142758 79076 142764 79088
rect 142816 79076 142822 79128
rect 144322 79116 144328 79128
rect 142960 79088 144328 79116
rect 65754 79048 65760 79060
rect 62000 79020 65760 79048
rect 65754 79008 65760 79020
rect 65812 79008 65818 79060
rect 141654 79008 141660 79060
rect 141712 79048 141718 79060
rect 142960 79048 142988 79088
rect 144322 79076 144328 79088
rect 144380 79076 144386 79128
rect 158306 79076 158312 79128
rect 158364 79116 158370 79128
rect 162078 79116 162084 79128
rect 158364 79088 162084 79116
rect 158364 79076 158370 79088
rect 162078 79076 162084 79088
rect 162136 79076 162142 79128
rect 242486 79076 242492 79128
rect 242544 79116 242550 79128
rect 247822 79116 247828 79128
rect 242544 79088 247828 79116
rect 242544 79076 242550 79088
rect 247822 79076 247828 79088
rect 247880 79076 247886 79128
rect 249202 79076 249208 79128
rect 249260 79116 249266 79128
rect 255826 79116 255832 79128
rect 249260 79088 255832 79116
rect 249260 79076 249266 79088
rect 255826 79076 255832 79088
rect 255884 79076 255890 79128
rect 256286 79076 256292 79128
rect 256344 79116 256350 79128
rect 256344 79088 256516 79116
rect 256344 79076 256350 79088
rect 141712 79020 142988 79048
rect 141712 79008 141718 79020
rect 143034 79008 143040 79060
rect 143092 79048 143098 79060
rect 145242 79048 145248 79060
rect 143092 79020 145248 79048
rect 143092 79008 143098 79020
rect 145242 79008 145248 79020
rect 145300 79008 145306 79060
rect 153982 79008 153988 79060
rect 154040 79048 154046 79060
rect 158401 79051 158459 79057
rect 158401 79048 158413 79051
rect 154040 79020 158413 79048
rect 154040 79008 154046 79020
rect 158401 79017 158413 79020
rect 158447 79017 158459 79051
rect 158401 79011 158459 79017
rect 159778 79008 159784 79060
rect 159836 79048 159842 79060
rect 167966 79048 167972 79060
rect 159836 79020 167972 79048
rect 159836 79008 159842 79020
rect 167966 79008 167972 79020
rect 168024 79008 168030 79060
rect 236874 79008 236880 79060
rect 236932 79048 236938 79060
rect 239174 79048 239180 79060
rect 236932 79020 239180 79048
rect 236932 79008 236938 79020
rect 239174 79008 239180 79020
rect 239232 79008 239238 79060
rect 244418 79008 244424 79060
rect 244476 79048 244482 79060
rect 249294 79048 249300 79060
rect 244476 79020 249300 79048
rect 244476 79008 244482 79020
rect 249294 79008 249300 79020
rect 249352 79008 249358 79060
rect 255734 79008 255740 79060
rect 255792 79048 255798 79060
rect 256378 79048 256384 79060
rect 255792 79020 256384 79048
rect 255792 79008 255798 79020
rect 256378 79008 256384 79020
rect 256436 79008 256442 79060
rect 256488 79048 256516 79088
rect 256562 79076 256568 79128
rect 256620 79116 256626 79128
rect 259230 79116 259236 79128
rect 256620 79088 259236 79116
rect 256620 79076 256626 79088
rect 259230 79076 259236 79088
rect 259288 79076 259294 79128
rect 260334 79048 260340 79060
rect 256488 79020 260340 79048
rect 260334 79008 260340 79020
rect 260392 79008 260398 79060
rect 60510 78940 60516 78992
rect 60568 78980 60574 78992
rect 64466 78980 64472 78992
rect 60568 78952 64472 78980
rect 60568 78940 60574 78952
rect 64466 78940 64472 78952
rect 64524 78940 64530 78992
rect 140274 78940 140280 78992
rect 140332 78980 140338 78992
rect 143770 78980 143776 78992
rect 140332 78952 143776 78980
rect 140332 78940 140338 78952
rect 143770 78940 143776 78952
rect 143828 78940 143834 78992
rect 151406 78940 151412 78992
rect 151464 78980 151470 78992
rect 157110 78980 157116 78992
rect 151464 78952 157116 78980
rect 151464 78940 151470 78952
rect 157110 78940 157116 78952
rect 157168 78940 157174 78992
rect 158214 78940 158220 78992
rect 158272 78980 158278 78992
rect 163182 78980 163188 78992
rect 158272 78952 163188 78980
rect 158272 78940 158278 78952
rect 163182 78940 163188 78952
rect 163240 78940 163246 78992
rect 246902 78940 246908 78992
rect 246960 78980 246966 78992
rect 247178 78980 247184 78992
rect 246960 78952 247184 78980
rect 246960 78940 246966 78952
rect 247178 78940 247184 78952
rect 247236 78940 247242 78992
rect 248098 78940 248104 78992
rect 248156 78980 248162 78992
rect 253434 78980 253440 78992
rect 248156 78952 253440 78980
rect 248156 78940 248162 78952
rect 253434 78940 253440 78952
rect 253492 78940 253498 78992
rect 256194 78940 256200 78992
rect 256252 78980 256258 78992
rect 256562 78980 256568 78992
rect 256252 78952 256568 78980
rect 256252 78940 256258 78952
rect 256562 78940 256568 78952
rect 256620 78940 256626 78992
rect 59130 78872 59136 78924
rect 59188 78912 59194 78924
rect 59188 78884 66628 78912
rect 59188 78872 59194 78884
rect 61706 78804 61712 78856
rect 61764 78844 61770 78856
rect 66490 78844 66496 78856
rect 61764 78816 66496 78844
rect 61764 78804 61770 78816
rect 66490 78804 66496 78816
rect 66548 78804 66554 78856
rect 66600 78844 66628 78884
rect 67134 78872 67140 78924
rect 67192 78912 67198 78924
rect 68422 78912 68428 78924
rect 67192 78884 68428 78912
rect 67192 78872 67198 78884
rect 68422 78872 68428 78884
rect 68480 78872 68486 78924
rect 157018 78872 157024 78924
rect 157076 78912 157082 78924
rect 164746 78912 164752 78924
rect 157076 78884 164752 78912
rect 157076 78872 157082 78884
rect 164746 78872 164752 78884
rect 164804 78872 164810 78924
rect 232734 78872 232740 78924
rect 232792 78912 232798 78924
rect 240738 78912 240744 78924
rect 232792 78884 240744 78912
rect 232792 78872 232798 78884
rect 240738 78872 240744 78884
rect 240796 78872 240802 78924
rect 244142 78872 244148 78924
rect 244200 78912 244206 78924
rect 249386 78912 249392 78924
rect 244200 78884 249392 78912
rect 244200 78872 244206 78884
rect 249386 78872 249392 78884
rect 249444 78872 249450 78924
rect 68054 78844 68060 78856
rect 66600 78816 68060 78844
rect 68054 78804 68060 78816
rect 68112 78804 68118 78856
rect 69894 78804 69900 78856
rect 69952 78844 69958 78856
rect 73114 78844 73120 78856
rect 69952 78816 73120 78844
rect 69952 78804 69958 78816
rect 73114 78804 73120 78816
rect 73172 78804 73178 78856
rect 156926 78804 156932 78856
rect 156984 78844 156990 78856
rect 165298 78844 165304 78856
rect 156984 78816 165304 78844
rect 156984 78804 156990 78816
rect 165298 78804 165304 78816
rect 165356 78804 165362 78856
rect 61798 78736 61804 78788
rect 61856 78776 61862 78788
rect 67134 78776 67140 78788
rect 61856 78748 67140 78776
rect 61856 78736 61862 78748
rect 67134 78736 67140 78748
rect 67192 78736 67198 78788
rect 147634 78736 147640 78788
rect 147692 78776 147698 78788
rect 151314 78776 151320 78788
rect 147692 78748 151320 78776
rect 147692 78736 147698 78748
rect 151314 78736 151320 78748
rect 151372 78736 151378 78788
rect 154718 78736 154724 78788
rect 154776 78776 154782 78788
rect 164562 78776 164568 78788
rect 154776 78748 164568 78776
rect 154776 78736 154782 78748
rect 164562 78736 164568 78748
rect 164620 78736 164626 78788
rect 243038 78736 243044 78788
rect 243096 78776 243102 78788
rect 247914 78776 247920 78788
rect 243096 78748 247920 78776
rect 243096 78736 243102 78748
rect 247914 78736 247920 78748
rect 247972 78736 247978 78788
rect 249389 78779 249447 78785
rect 249389 78745 249401 78779
rect 249435 78776 249447 78779
rect 255642 78776 255648 78788
rect 249435 78748 255648 78776
rect 249435 78745 249447 78748
rect 249389 78739 249447 78745
rect 255642 78736 255648 78748
rect 255700 78736 255706 78788
rect 61614 78668 61620 78720
rect 61672 78708 61678 78720
rect 67778 78708 67784 78720
rect 61672 78680 67784 78708
rect 61672 78668 61678 78680
rect 67778 78668 67784 78680
rect 67836 78668 67842 78720
rect 156009 78711 156067 78717
rect 156009 78677 156021 78711
rect 156055 78708 156067 78711
rect 166402 78708 166408 78720
rect 156055 78680 166408 78708
rect 156055 78677 156067 78680
rect 156009 78671 156067 78677
rect 166402 78668 166408 78680
rect 166460 78668 166466 78720
rect 246994 78668 247000 78720
rect 247052 78708 247058 78720
rect 253526 78708 253532 78720
rect 247052 78680 253532 78708
rect 247052 78668 247058 78680
rect 253526 78668 253532 78680
rect 253584 78668 253590 78720
rect 58673 78643 58731 78649
rect 58673 78609 58685 78643
rect 58719 78640 58731 78643
rect 61982 78640 61988 78652
rect 58719 78612 61988 78640
rect 58719 78609 58731 78612
rect 58673 78603 58731 78609
rect 61982 78600 61988 78612
rect 62040 78600 62046 78652
rect 62077 78643 62135 78649
rect 62077 78609 62089 78643
rect 62123 78640 62135 78643
rect 68238 78640 68244 78652
rect 62123 78612 68244 78640
rect 62123 78609 62135 78612
rect 62077 78603 62135 78609
rect 68238 78600 68244 78612
rect 68296 78600 68302 78652
rect 151958 78600 151964 78652
rect 152016 78640 152022 78652
rect 161710 78640 161716 78652
rect 152016 78612 161716 78640
rect 152016 78600 152022 78612
rect 161710 78600 161716 78612
rect 161768 78600 161774 78652
rect 243590 78600 243596 78652
rect 243648 78640 243654 78652
rect 249570 78640 249576 78652
rect 243648 78612 249576 78640
rect 243648 78600 243654 78612
rect 249570 78600 249576 78612
rect 249628 78600 249634 78652
rect 251226 78600 251232 78652
rect 251284 78640 251290 78652
rect 263094 78640 263100 78652
rect 251284 78612 263100 78640
rect 251284 78600 251290 78612
rect 263094 78600 263100 78612
rect 263152 78600 263158 78652
rect 55174 78532 55180 78584
rect 55232 78572 55238 78584
rect 55232 78544 60280 78572
rect 55232 78532 55238 78544
rect 38246 78464 38252 78516
rect 38304 78504 38310 78516
rect 49194 78504 49200 78516
rect 38304 78476 49200 78504
rect 38304 78464 38310 78476
rect 49194 78464 49200 78476
rect 49252 78464 49258 78516
rect 53150 78464 53156 78516
rect 53208 78504 53214 78516
rect 58673 78507 58731 78513
rect 58673 78504 58685 78507
rect 53208 78476 58685 78504
rect 53208 78464 53214 78476
rect 58673 78473 58685 78476
rect 58719 78473 58731 78507
rect 60252 78504 60280 78544
rect 60326 78532 60332 78584
rect 60384 78572 60390 78584
rect 63822 78572 63828 78584
rect 60384 78544 63828 78572
rect 60384 78532 60390 78544
rect 63822 78532 63828 78544
rect 63880 78532 63886 78584
rect 151774 78532 151780 78584
rect 151832 78572 151838 78584
rect 157202 78572 157208 78584
rect 151832 78544 157208 78572
rect 151832 78532 151838 78544
rect 157202 78532 157208 78544
rect 157260 78532 157266 78584
rect 157294 78532 157300 78584
rect 157352 78572 157358 78584
rect 167414 78572 167420 78584
rect 157352 78544 167420 78572
rect 157352 78532 157358 78544
rect 167414 78532 167420 78544
rect 167472 78532 167478 78584
rect 248466 78532 248472 78584
rect 248524 78572 248530 78584
rect 249389 78575 249447 78581
rect 249389 78572 249401 78575
rect 248524 78544 249401 78572
rect 248524 78532 248530 78544
rect 249389 78541 249401 78544
rect 249435 78541 249447 78575
rect 249389 78535 249447 78541
rect 249478 78532 249484 78584
rect 249536 78572 249542 78584
rect 254722 78572 254728 78584
rect 249536 78544 254728 78572
rect 249536 78532 249542 78544
rect 254722 78532 254728 78544
rect 254780 78532 254786 78584
rect 62261 78507 62319 78513
rect 62261 78504 62273 78507
rect 60252 78476 62273 78504
rect 58673 78467 58731 78473
rect 62261 78473 62273 78476
rect 62307 78473 62319 78507
rect 62261 78467 62319 78473
rect 63546 78464 63552 78516
rect 63604 78504 63610 78516
rect 75782 78504 75788 78516
rect 63604 78476 75788 78504
rect 63604 78464 63610 78476
rect 75782 78464 75788 78476
rect 75840 78464 75846 78516
rect 138894 78464 138900 78516
rect 138952 78504 138958 78516
rect 146530 78504 146536 78516
rect 138952 78476 146536 78504
rect 138952 78464 138958 78476
rect 146530 78464 146536 78476
rect 146588 78464 146594 78516
rect 150486 78464 150492 78516
rect 150544 78504 150550 78516
rect 150544 78476 156328 78504
rect 150544 78464 150550 78476
rect 60418 78396 60424 78448
rect 60476 78436 60482 78448
rect 65110 78436 65116 78448
rect 60476 78408 65116 78436
rect 60476 78396 60482 78408
rect 65110 78396 65116 78408
rect 65168 78396 65174 78448
rect 67962 78436 67968 78448
rect 66508 78408 67968 78436
rect 60329 78371 60387 78377
rect 60329 78337 60341 78371
rect 60375 78368 60387 78371
rect 66508 78368 66536 78408
rect 67962 78396 67968 78408
rect 68020 78396 68026 78448
rect 156300 78436 156328 78476
rect 156650 78464 156656 78516
rect 156708 78504 156714 78516
rect 163734 78504 163740 78516
rect 156708 78476 163740 78504
rect 156708 78464 156714 78476
rect 163734 78464 163740 78476
rect 163792 78464 163798 78516
rect 234114 78464 234120 78516
rect 234172 78504 234178 78516
rect 237978 78504 237984 78516
rect 234172 78476 237984 78504
rect 234172 78464 234178 78476
rect 237978 78464 237984 78476
rect 238036 78464 238042 78516
rect 251134 78464 251140 78516
rect 251192 78504 251198 78516
rect 262542 78504 262548 78516
rect 251192 78476 262548 78504
rect 251192 78464 251198 78476
rect 262542 78464 262548 78476
rect 262600 78464 262606 78516
rect 264474 78464 264480 78516
rect 264532 78504 264538 78516
rect 295570 78504 295576 78516
rect 264532 78476 295576 78504
rect 264532 78464 264538 78476
rect 295570 78464 295576 78476
rect 295628 78464 295634 78516
rect 158306 78436 158312 78448
rect 156300 78408 158312 78436
rect 158306 78396 158312 78408
rect 158364 78396 158370 78448
rect 158401 78439 158459 78445
rect 158401 78405 158413 78439
rect 158447 78436 158459 78439
rect 161066 78436 161072 78448
rect 158447 78408 161072 78436
rect 158447 78405 158459 78408
rect 158401 78399 158459 78405
rect 161066 78396 161072 78408
rect 161124 78396 161130 78448
rect 248282 78396 248288 78448
rect 248340 78436 248346 78448
rect 254170 78436 254176 78448
rect 248340 78408 254176 78436
rect 248340 78396 248346 78408
rect 254170 78396 254176 78408
rect 254228 78396 254234 78448
rect 60375 78340 66536 78368
rect 60375 78337 60387 78340
rect 60329 78331 60387 78337
rect 67410 78328 67416 78380
rect 67468 78368 67474 78380
rect 69802 78368 69808 78380
rect 67468 78340 69808 78368
rect 67468 78328 67474 78340
rect 69802 78328 69808 78340
rect 69860 78328 69866 78380
rect 144414 78328 144420 78380
rect 144472 78368 144478 78380
rect 145426 78368 145432 78380
rect 144472 78340 145432 78368
rect 144472 78328 144478 78340
rect 145426 78328 145432 78340
rect 145484 78328 145490 78380
rect 150486 78328 150492 78380
rect 150544 78368 150550 78380
rect 155730 78368 155736 78380
rect 150544 78340 155736 78368
rect 150544 78328 150550 78340
rect 155730 78328 155736 78340
rect 155788 78328 155794 78380
rect 155822 78328 155828 78380
rect 155880 78368 155886 78380
rect 165850 78368 165856 78380
rect 155880 78340 165856 78368
rect 155880 78328 155886 78340
rect 165850 78328 165856 78340
rect 165908 78328 165914 78380
rect 235494 78328 235500 78380
rect 235552 78368 235558 78380
rect 238530 78368 238536 78380
rect 235552 78340 238536 78368
rect 235552 78328 235558 78340
rect 238530 78328 238536 78340
rect 238588 78328 238594 78380
rect 248006 78328 248012 78380
rect 248064 78368 248070 78380
rect 253066 78368 253072 78380
rect 248064 78340 253072 78368
rect 248064 78328 248070 78340
rect 253066 78328 253072 78340
rect 253124 78328 253130 78380
rect 149750 78260 149756 78312
rect 149808 78300 149814 78312
rect 155362 78300 155368 78312
rect 149808 78272 155368 78300
rect 149808 78260 149814 78272
rect 155362 78260 155368 78272
rect 155420 78260 155426 78312
rect 155638 78260 155644 78312
rect 155696 78300 155702 78312
rect 160330 78300 160336 78312
rect 155696 78272 160336 78300
rect 155696 78260 155702 78272
rect 160330 78260 160336 78272
rect 160388 78260 160394 78312
rect 248190 78260 248196 78312
rect 248248 78300 248254 78312
rect 253618 78300 253624 78312
rect 248248 78272 253624 78300
rect 248248 78260 248254 78272
rect 253618 78260 253624 78272
rect 253676 78260 253682 78312
rect 58486 78192 58492 78244
rect 58544 78232 58550 78244
rect 60329 78235 60387 78241
rect 60329 78232 60341 78235
rect 58544 78204 60341 78232
rect 58544 78192 58550 78204
rect 60329 78201 60341 78204
rect 60375 78201 60387 78235
rect 60329 78195 60387 78201
rect 60418 78192 60424 78244
rect 60476 78232 60482 78244
rect 62169 78235 62227 78241
rect 62169 78232 62181 78235
rect 60476 78204 62181 78232
rect 60476 78192 60482 78204
rect 62169 78201 62181 78204
rect 62215 78201 62227 78235
rect 62169 78195 62227 78201
rect 62261 78235 62319 78241
rect 62261 78201 62273 78235
rect 62307 78232 62319 78235
rect 65202 78232 65208 78244
rect 62307 78204 65208 78232
rect 62307 78201 62319 78204
rect 62261 78195 62319 78201
rect 65202 78192 65208 78204
rect 65260 78192 65266 78244
rect 67226 78192 67232 78244
rect 67284 78232 67290 78244
rect 69158 78232 69164 78244
rect 67284 78204 69164 78232
rect 67284 78192 67290 78204
rect 69158 78192 69164 78204
rect 69216 78192 69222 78244
rect 148738 78192 148744 78244
rect 148796 78232 148802 78244
rect 154074 78232 154080 78244
rect 148796 78204 154080 78232
rect 148796 78192 148802 78204
rect 154074 78192 154080 78204
rect 154132 78192 154138 78244
rect 157662 78192 157668 78244
rect 157720 78232 157726 78244
rect 158858 78232 158864 78244
rect 157720 78204 158864 78232
rect 157720 78192 157726 78204
rect 158858 78192 158864 78204
rect 158916 78192 158922 78244
rect 245338 78192 245344 78244
rect 245396 78232 245402 78244
rect 250766 78232 250772 78244
rect 245396 78204 250772 78232
rect 245396 78192 245402 78204
rect 250766 78192 250772 78204
rect 250824 78192 250830 78244
rect 55818 78124 55824 78176
rect 55876 78164 55882 78176
rect 65846 78164 65852 78176
rect 55876 78136 65852 78164
rect 55876 78124 55882 78136
rect 65846 78124 65852 78136
rect 65904 78124 65910 78176
rect 149198 78124 149204 78176
rect 149256 78164 149262 78176
rect 154166 78164 154172 78176
rect 149256 78136 154172 78164
rect 149256 78124 149262 78136
rect 154166 78124 154172 78136
rect 154224 78124 154230 78176
rect 155086 78124 155092 78176
rect 155144 78164 155150 78176
rect 156098 78164 156104 78176
rect 155144 78136 156104 78164
rect 155144 78124 155150 78136
rect 156098 78124 156104 78136
rect 156156 78124 156162 78176
rect 245798 78124 245804 78176
rect 245856 78164 245862 78176
rect 250674 78164 250680 78176
rect 245856 78136 250680 78164
rect 245856 78124 245862 78136
rect 250674 78124 250680 78136
rect 250732 78124 250738 78176
rect 252790 78164 252796 78176
rect 250784 78136 252796 78164
rect 57842 78056 57848 78108
rect 57900 78096 57906 78108
rect 62077 78099 62135 78105
rect 62077 78096 62089 78099
rect 57900 78068 62089 78096
rect 57900 78056 57906 78068
rect 62077 78065 62089 78068
rect 62123 78065 62135 78099
rect 62077 78059 62135 78065
rect 62169 78099 62227 78105
rect 62169 78065 62181 78099
rect 62215 78096 62227 78099
rect 65754 78096 65760 78108
rect 62215 78068 65760 78096
rect 62215 78065 62227 78068
rect 62169 78059 62227 78065
rect 65754 78056 65760 78068
rect 65812 78056 65818 78108
rect 67318 78056 67324 78108
rect 67376 78096 67382 78108
rect 70446 78096 70452 78108
rect 67376 78068 70452 78096
rect 67376 78056 67382 78068
rect 70446 78056 70452 78068
rect 70504 78056 70510 78108
rect 153154 78056 153160 78108
rect 153212 78096 153218 78108
rect 157389 78099 157447 78105
rect 157389 78096 157401 78099
rect 153212 78068 157401 78096
rect 153212 78056 153218 78068
rect 157389 78065 157401 78068
rect 157435 78065 157447 78099
rect 157389 78059 157447 78065
rect 232826 78056 232832 78108
rect 232884 78096 232890 78108
rect 236874 78096 236880 78108
rect 232884 78068 236880 78096
rect 232884 78056 232890 78068
rect 236874 78056 236880 78068
rect 236932 78056 236938 78108
rect 239634 78056 239640 78108
rect 239692 78096 239698 78108
rect 240370 78096 240376 78108
rect 239692 78068 240376 78096
rect 239692 78056 239698 78068
rect 240370 78056 240376 78068
rect 240428 78056 240434 78108
rect 248374 78056 248380 78108
rect 248432 78096 248438 78108
rect 250784 78096 250812 78136
rect 252790 78124 252796 78136
rect 252848 78124 252854 78176
rect 248432 78068 250812 78096
rect 248432 78056 248438 78068
rect 252054 78056 252060 78108
rect 252112 78096 252118 78108
rect 252698 78096 252704 78108
rect 252112 78068 252704 78096
rect 252112 78056 252118 78068
rect 252698 78056 252704 78068
rect 252756 78056 252762 78108
rect 59774 77988 59780 78040
rect 59832 78028 59838 78040
rect 67502 78028 67508 78040
rect 59832 78000 67508 78028
rect 59832 77988 59838 78000
rect 67502 77988 67508 78000
rect 67560 77988 67566 78040
rect 153062 77988 153068 78040
rect 153120 78028 153126 78040
rect 157297 78031 157355 78037
rect 157297 78028 157309 78031
rect 153120 78000 157309 78028
rect 153120 77988 153126 78000
rect 157297 77997 157309 78000
rect 157343 77997 157355 78031
rect 157297 77991 157355 77997
rect 157481 78031 157539 78037
rect 157481 77997 157493 78031
rect 157527 78028 157539 78031
rect 159686 78028 159692 78040
rect 157527 78000 159692 78028
rect 157527 77997 157539 78000
rect 157481 77991 157539 77997
rect 159686 77988 159692 78000
rect 159744 77988 159750 78040
rect 56094 77920 56100 77972
rect 56152 77960 56158 77972
rect 63178 77960 63184 77972
rect 56152 77932 63184 77960
rect 56152 77920 56158 77932
rect 63178 77920 63184 77932
rect 63236 77920 63242 77972
rect 148186 77920 148192 77972
rect 148244 77960 148250 77972
rect 152694 77960 152700 77972
rect 148244 77932 152700 77960
rect 148244 77920 148250 77932
rect 152694 77920 152700 77932
rect 152752 77920 152758 77972
rect 154626 77920 154632 77972
rect 154684 77960 154690 77972
rect 160882 77960 160888 77972
rect 154684 77932 160888 77960
rect 154684 77920 154690 77932
rect 160882 77920 160888 77932
rect 160940 77920 160946 77972
rect 57106 77852 57112 77904
rect 57164 77892 57170 77904
rect 64374 77892 64380 77904
rect 57164 77864 64380 77892
rect 57164 77852 57170 77864
rect 64374 77852 64380 77864
rect 64432 77852 64438 77904
rect 150394 77852 150400 77904
rect 150452 77892 150458 77904
rect 150578 77892 150584 77904
rect 150452 77864 150584 77892
rect 150452 77852 150458 77864
rect 150578 77852 150584 77864
rect 150636 77852 150642 77904
rect 152510 77852 152516 77904
rect 152568 77892 152574 77904
rect 153338 77892 153344 77904
rect 152568 77864 153344 77892
rect 152568 77852 152574 77864
rect 153338 77852 153344 77864
rect 153396 77852 153402 77904
rect 155178 77852 155184 77904
rect 155236 77892 155242 77904
rect 156006 77892 156012 77904
rect 155236 77864 156012 77892
rect 155236 77852 155242 77864
rect 156006 77852 156012 77864
rect 156064 77852 156070 77904
rect 156834 77852 156840 77904
rect 156892 77892 156898 77904
rect 157386 77892 157392 77904
rect 156892 77864 157392 77892
rect 156892 77852 156898 77864
rect 157386 77852 157392 77864
rect 157444 77852 157450 77904
rect 157481 77895 157539 77901
rect 157481 77861 157493 77895
rect 157527 77892 157539 77895
rect 159594 77892 159600 77904
rect 157527 77864 159600 77892
rect 157527 77861 157539 77864
rect 157481 77855 157539 77861
rect 159594 77852 159600 77864
rect 159652 77852 159658 77904
rect 155454 77784 155460 77836
rect 155512 77824 155518 77836
rect 160974 77824 160980 77836
rect 155512 77796 160980 77824
rect 155512 77784 155518 77796
rect 160974 77784 160980 77796
rect 161032 77784 161038 77836
rect 89766 77688 89772 77700
rect 89727 77660 89772 77688
rect 89766 77648 89772 77660
rect 89824 77648 89830 77700
rect 124726 76356 124732 76408
rect 124784 76396 124790 76408
rect 169990 76396 169996 76408
rect 124784 76368 169996 76396
rect 124784 76356 124790 76368
rect 169990 76356 169996 76368
rect 170048 76356 170054 76408
rect 218658 76356 218664 76408
rect 218716 76396 218722 76408
rect 233470 76396 233476 76408
rect 218716 76368 233476 76396
rect 218716 76356 218722 76368
rect 233470 76356 233476 76368
rect 233528 76356 233534 76408
rect 119298 76288 119304 76340
rect 119356 76328 119362 76340
rect 139630 76328 139636 76340
rect 119356 76300 139636 76328
rect 119356 76288 119362 76300
rect 139630 76288 139636 76300
rect 139688 76288 139694 76340
rect 111202 74996 111208 75048
rect 111260 75036 111266 75048
rect 170726 75036 170732 75048
rect 111260 75008 170732 75036
rect 111260 74996 111266 75008
rect 170726 74996 170732 75008
rect 170784 74996 170790 75048
rect 205134 74996 205140 75048
rect 205192 75036 205198 75048
rect 233654 75036 233660 75048
rect 205192 75008 233660 75036
rect 205192 74996 205198 75008
rect 233654 74996 233660 75008
rect 233712 74996 233718 75048
rect 113962 74928 113968 74980
rect 114020 74968 114026 74980
rect 170818 74968 170824 74980
rect 114020 74940 170824 74968
rect 114020 74928 114026 74940
rect 170818 74928 170824 74940
rect 170876 74928 170882 74980
rect 213230 74928 213236 74980
rect 213288 74968 213294 74980
rect 233562 74968 233568 74980
rect 213288 74940 233568 74968
rect 213288 74928 213294 74940
rect 233562 74928 233568 74940
rect 233620 74928 233626 74980
rect 116630 74860 116636 74912
rect 116688 74900 116694 74912
rect 170634 74900 170640 74912
rect 116688 74872 170640 74900
rect 116688 74860 116694 74872
rect 170634 74860 170640 74872
rect 170692 74860 170698 74912
rect 215990 74860 215996 74912
rect 216048 74900 216054 74912
rect 233470 74900 233476 74912
rect 216048 74872 233476 74900
rect 216048 74860 216054 74872
rect 233470 74860 233476 74872
rect 233528 74860 233534 74912
rect 138066 73704 138072 73756
rect 138124 73744 138130 73756
rect 139630 73744 139636 73756
rect 138124 73716 139636 73744
rect 138124 73704 138130 73716
rect 139630 73704 139636 73716
rect 139688 73704 139694 73756
rect 100254 73636 100260 73688
rect 100312 73676 100318 73688
rect 100990 73676 100996 73688
rect 100312 73648 100996 73676
rect 100312 73636 100318 73648
rect 100990 73636 100996 73648
rect 101048 73636 101054 73688
rect 183698 73636 183704 73688
rect 183756 73676 183762 73688
rect 190138 73676 190144 73688
rect 183756 73648 190144 73676
rect 183756 73636 183762 73648
rect 190138 73636 190144 73648
rect 190196 73636 190202 73688
rect 190598 73636 190604 73688
rect 190656 73636 190662 73688
rect 96390 73500 96396 73552
rect 96448 73540 96454 73552
rect 108258 73540 108264 73552
rect 96448 73512 108264 73540
rect 96448 73500 96454 73512
rect 108258 73500 108264 73512
rect 108316 73500 108322 73552
rect 190616 73540 190644 73636
rect 202650 73540 202656 73552
rect 190616 73512 202656 73540
rect 202650 73500 202656 73512
rect 202708 73500 202714 73552
rect 97770 73432 97776 73484
rect 97828 73472 97834 73484
rect 110742 73472 110748 73484
rect 97828 73444 110748 73472
rect 97828 73432 97834 73444
rect 110742 73432 110748 73444
rect 110800 73432 110806 73484
rect 191978 73432 191984 73484
rect 192036 73472 192042 73484
rect 205134 73472 205140 73484
rect 192036 73444 205140 73472
rect 192036 73432 192042 73444
rect 205134 73432 205140 73444
rect 205192 73432 205198 73484
rect 100898 73364 100904 73416
rect 100956 73404 100962 73416
rect 115710 73404 115716 73416
rect 100956 73376 115716 73404
rect 100956 73364 100962 73376
rect 115710 73364 115716 73376
rect 115768 73364 115774 73416
rect 193358 73364 193364 73416
rect 193416 73404 193422 73416
rect 207618 73404 207624 73416
rect 193416 73376 207624 73404
rect 193416 73364 193422 73376
rect 207618 73364 207624 73376
rect 207676 73364 207682 73416
rect 99518 73296 99524 73348
rect 99576 73336 99582 73348
rect 113410 73336 113416 73348
rect 99576 73308 113416 73336
rect 99576 73296 99582 73308
rect 113410 73296 113416 73308
rect 113468 73296 113474 73348
rect 194738 73296 194744 73348
rect 194796 73336 194802 73348
rect 210102 73336 210108 73348
rect 194796 73308 210108 73336
rect 194796 73296 194802 73308
rect 210102 73296 210108 73308
rect 210160 73296 210166 73348
rect 102278 73228 102284 73280
rect 102336 73268 102342 73280
rect 118286 73268 118292 73280
rect 102336 73240 118292 73268
rect 102336 73228 102342 73240
rect 118286 73228 118292 73240
rect 118344 73228 118350 73280
rect 196118 73228 196124 73280
rect 196176 73268 196182 73280
rect 212678 73268 212684 73280
rect 196176 73240 212684 73268
rect 196176 73228 196182 73240
rect 212678 73228 212684 73240
rect 212736 73228 212742 73280
rect 103658 73160 103664 73212
rect 103716 73200 103722 73212
rect 120770 73200 120776 73212
rect 103716 73172 120776 73200
rect 103716 73160 103722 73172
rect 120770 73160 120776 73172
rect 120828 73160 120834 73212
rect 197498 73160 197504 73212
rect 197556 73200 197562 73212
rect 215162 73200 215168 73212
rect 197556 73172 215168 73200
rect 197556 73160 197562 73172
rect 215162 73160 215168 73172
rect 215220 73160 215226 73212
rect 105038 73092 105044 73144
rect 105096 73132 105102 73144
rect 123254 73132 123260 73144
rect 105096 73104 123260 73132
rect 105096 73092 105102 73104
rect 123254 73092 123260 73104
rect 123312 73092 123318 73144
rect 198878 73092 198884 73144
rect 198936 73132 198942 73144
rect 217646 73132 217652 73144
rect 198936 73104 217652 73132
rect 198936 73092 198942 73104
rect 217646 73092 217652 73104
rect 217704 73092 217710 73144
rect 106418 73024 106424 73076
rect 106476 73064 106482 73076
rect 125830 73064 125836 73076
rect 106476 73036 125836 73064
rect 106476 73024 106482 73036
rect 125830 73024 125836 73036
rect 125888 73024 125894 73076
rect 200258 73024 200264 73076
rect 200316 73064 200322 73076
rect 220130 73064 220136 73076
rect 200316 73036 220136 73064
rect 200316 73024 200322 73036
rect 220130 73024 220136 73036
rect 220188 73024 220194 73076
rect 107798 72956 107804 73008
rect 107856 72996 107862 73008
rect 128590 72996 128596 73008
rect 107856 72968 128596 72996
rect 107856 72956 107862 72968
rect 128590 72956 128596 72968
rect 128648 72956 128654 73008
rect 201638 72956 201644 73008
rect 201696 72996 201702 73008
rect 222614 72996 222620 73008
rect 201696 72968 222620 72996
rect 201696 72956 201702 72968
rect 222614 72956 222620 72968
rect 222672 72956 222678 73008
rect 89766 72888 89772 72940
rect 89824 72928 89830 72940
rect 95746 72928 95752 72940
rect 89824 72900 95752 72928
rect 89824 72888 89830 72900
rect 95746 72888 95752 72900
rect 95804 72888 95810 72940
rect 96114 72888 96120 72940
rect 96172 72928 96178 72940
rect 98230 72928 98236 72940
rect 96172 72900 98236 72928
rect 96172 72888 96178 72900
rect 98230 72888 98236 72900
rect 98288 72888 98294 72940
rect 101634 72684 101640 72736
rect 101692 72724 101698 72736
rect 105774 72724 105780 72736
rect 101692 72696 105780 72724
rect 101692 72684 101698 72696
rect 105774 72684 105780 72696
rect 105832 72684 105838 72736
rect 91974 72616 91980 72668
rect 92032 72656 92038 72668
rect 93262 72656 93268 72668
rect 92032 72628 93268 72656
rect 92032 72616 92038 72628
rect 93262 72616 93268 72628
rect 93320 72616 93326 72668
rect 101726 72616 101732 72668
rect 101784 72656 101790 72668
rect 103198 72656 103204 72668
rect 101784 72628 103204 72656
rect 101784 72616 101790 72628
rect 103198 72616 103204 72628
rect 103256 72616 103262 72668
rect 136502 72412 136508 72464
rect 136560 72452 136566 72464
rect 139722 72452 139728 72464
rect 136560 72424 139728 72452
rect 136560 72412 136566 72424
rect 139722 72412 139728 72424
rect 139780 72412 139786 72464
rect 195474 72412 195480 72464
rect 195532 72452 195538 72464
rect 200166 72452 200172 72464
rect 195532 72424 200172 72452
rect 195532 72412 195538 72424
rect 200166 72412 200172 72424
rect 200224 72412 200230 72464
rect 89214 72344 89220 72396
rect 89272 72384 89278 72396
rect 90778 72384 90784 72396
rect 89272 72356 90784 72384
rect 89272 72344 89278 72356
rect 90778 72344 90784 72356
rect 90836 72344 90842 72396
rect 136778 72344 136784 72396
rect 136836 72384 136842 72396
rect 139630 72384 139636 72396
rect 136836 72356 139636 72384
rect 136836 72344 136842 72356
rect 139630 72344 139636 72356
rect 139688 72344 139694 72396
rect 183054 72344 183060 72396
rect 183112 72384 183118 72396
rect 184710 72384 184716 72396
rect 183112 72356 184716 72384
rect 183112 72344 183118 72356
rect 184710 72344 184716 72356
rect 184768 72344 184774 72396
rect 185814 72344 185820 72396
rect 185872 72384 185878 72396
rect 187654 72384 187660 72396
rect 185872 72356 187660 72384
rect 185872 72344 185878 72356
rect 187654 72344 187660 72356
rect 187712 72344 187718 72396
rect 191334 72344 191340 72396
rect 191392 72384 191398 72396
rect 192622 72384 192628 72396
rect 191392 72356 192628 72384
rect 191392 72344 191398 72356
rect 192622 72344 192628 72356
rect 192680 72344 192686 72396
rect 194094 72344 194100 72396
rect 194152 72384 194158 72396
rect 195106 72384 195112 72396
rect 194152 72356 195112 72384
rect 194152 72344 194158 72356
rect 195106 72344 195112 72356
rect 195164 72344 195170 72396
rect 195566 72344 195572 72396
rect 195624 72384 195630 72396
rect 197498 72384 197504 72396
rect 195624 72356 197504 72384
rect 195624 72344 195630 72356
rect 197498 72344 197504 72356
rect 197556 72344 197562 72396
rect 230618 72344 230624 72396
rect 230676 72384 230682 72396
rect 233470 72384 233476 72396
rect 230676 72356 233476 72384
rect 230676 72344 230682 72356
rect 233470 72344 233476 72356
rect 233528 72344 233534 72396
rect 80198 70916 80204 70968
rect 80256 70956 80262 70968
rect 84430 70956 84436 70968
rect 80256 70928 84436 70956
rect 80256 70916 80262 70928
rect 84430 70916 84436 70928
rect 84488 70916 84494 70968
rect 135950 70916 135956 70968
rect 136008 70956 136014 70968
rect 139630 70956 139636 70968
rect 136008 70928 139636 70956
rect 136008 70916 136014 70928
rect 139630 70916 139636 70928
rect 139688 70916 139694 70968
rect 131350 70848 131356 70900
rect 131408 70888 131414 70900
rect 138066 70888 138072 70900
rect 131408 70860 138072 70888
rect 131408 70848 131414 70860
rect 138066 70848 138072 70860
rect 138124 70848 138130 70900
rect 226018 70848 226024 70900
rect 226076 70888 226082 70900
rect 230618 70888 230624 70900
rect 226076 70860 230624 70888
rect 226076 70848 226082 70860
rect 230618 70848 230624 70860
rect 230676 70848 230682 70900
rect 276158 70848 276164 70900
rect 276216 70888 276222 70900
rect 300170 70888 300176 70900
rect 276216 70860 300176 70888
rect 276216 70848 276222 70860
rect 300170 70848 300176 70860
rect 300228 70848 300234 70900
rect 84430 70236 84436 70288
rect 84488 70276 84494 70288
rect 87190 70276 87196 70288
rect 84488 70248 87196 70276
rect 84488 70236 84494 70248
rect 87190 70236 87196 70248
rect 87248 70236 87254 70288
rect 136410 69692 136416 69744
rect 136468 69732 136474 69744
rect 139814 69732 139820 69744
rect 136468 69704 139820 69732
rect 136468 69692 136474 69704
rect 139814 69692 139820 69704
rect 139872 69692 139878 69744
rect 229882 69692 229888 69744
rect 229940 69732 229946 69744
rect 233654 69732 233660 69744
rect 229940 69704 233660 69732
rect 229940 69692 229946 69704
rect 233654 69692 233660 69704
rect 233712 69692 233718 69744
rect 79462 69624 79468 69676
rect 79520 69664 79526 69676
rect 79520 69636 85764 69664
rect 79520 69624 79526 69636
rect 80198 69556 80204 69608
rect 80256 69596 80262 69608
rect 80256 69568 85672 69596
rect 80256 69556 80262 69568
rect 85644 69460 85672 69568
rect 85736 69528 85764 69636
rect 136594 69624 136600 69676
rect 136652 69664 136658 69676
rect 139722 69664 139728 69676
rect 136652 69636 139728 69664
rect 136652 69624 136658 69636
rect 139722 69624 139728 69636
rect 139780 69624 139786 69676
rect 136686 69556 136692 69608
rect 136744 69596 136750 69608
rect 139630 69596 139636 69608
rect 136744 69568 139636 69596
rect 136744 69556 136750 69568
rect 139630 69556 139636 69568
rect 139688 69556 139694 69608
rect 87190 69528 87196 69540
rect 85736 69500 87196 69528
rect 87190 69488 87196 69500
rect 87248 69488 87254 69540
rect 131534 69488 131540 69540
rect 131592 69528 131598 69540
rect 135950 69528 135956 69540
rect 131592 69500 135956 69528
rect 131592 69488 131598 69500
rect 135950 69488 135956 69500
rect 136008 69488 136014 69540
rect 173302 69488 173308 69540
rect 173360 69528 173366 69540
rect 181766 69528 181772 69540
rect 173360 69500 181772 69528
rect 173360 69488 173366 69500
rect 181766 69488 181772 69500
rect 181824 69488 181830 69540
rect 226018 69488 226024 69540
rect 226076 69528 226082 69540
rect 233562 69528 233568 69540
rect 226076 69500 233568 69528
rect 226076 69488 226082 69500
rect 233562 69488 233568 69500
rect 233620 69488 233626 69540
rect 87282 69460 87288 69472
rect 85644 69432 87288 69460
rect 87282 69420 87288 69432
rect 87340 69420 87346 69472
rect 131350 69420 131356 69472
rect 131408 69460 131414 69472
rect 136502 69460 136508 69472
rect 131408 69432 136508 69460
rect 131408 69420 131414 69432
rect 136502 69420 136508 69432
rect 136560 69420 136566 69472
rect 225742 69420 225748 69472
rect 225800 69460 225806 69472
rect 233470 69460 233476 69472
rect 225800 69432 233476 69460
rect 225800 69420 225806 69432
rect 233470 69420 233476 69432
rect 233528 69420 233534 69472
rect 131442 69352 131448 69404
rect 131500 69392 131506 69404
rect 136778 69392 136784 69404
rect 131500 69364 136784 69392
rect 131500 69352 131506 69364
rect 136778 69352 136784 69364
rect 136836 69352 136842 69404
rect 80198 68808 80204 68860
rect 80256 68848 80262 68860
rect 87190 68848 87196 68860
rect 80256 68820 87196 68848
rect 80256 68808 80262 68820
rect 87190 68808 87196 68820
rect 87248 68808 87254 68860
rect 172842 68808 172848 68860
rect 172900 68848 172906 68860
rect 182318 68848 182324 68860
rect 172900 68820 182324 68848
rect 172900 68808 172906 68820
rect 182318 68808 182324 68820
rect 182376 68808 182382 68860
rect 226294 68740 226300 68792
rect 226352 68780 226358 68792
rect 229882 68780 229888 68792
rect 226352 68752 229888 68780
rect 226352 68740 226358 68752
rect 229882 68740 229888 68752
rect 229940 68740 229946 68792
rect 80106 68264 80112 68316
rect 80164 68304 80170 68316
rect 80164 68276 85580 68304
rect 80164 68264 80170 68276
rect 80198 68196 80204 68248
rect 80256 68236 80262 68248
rect 80256 68208 85488 68236
rect 80256 68196 80262 68208
rect 85460 68100 85488 68208
rect 85552 68168 85580 68276
rect 136502 68264 136508 68316
rect 136560 68304 136566 68316
rect 139722 68304 139728 68316
rect 136560 68276 139728 68304
rect 136560 68264 136566 68276
rect 139722 68264 139728 68276
rect 139780 68264 139786 68316
rect 136778 68196 136784 68248
rect 136836 68236 136842 68248
rect 139630 68236 139636 68248
rect 136836 68208 139636 68236
rect 136836 68196 136842 68208
rect 139630 68196 139636 68208
rect 139688 68196 139694 68248
rect 87190 68168 87196 68180
rect 85552 68140 87196 68168
rect 87190 68128 87196 68140
rect 87248 68128 87254 68180
rect 131994 68128 132000 68180
rect 132052 68168 132058 68180
rect 139906 68168 139912 68180
rect 132052 68140 139912 68168
rect 132052 68128 132058 68140
rect 139906 68128 139912 68140
rect 139964 68128 139970 68180
rect 174038 68128 174044 68180
rect 174096 68168 174102 68180
rect 181766 68168 181772 68180
rect 174096 68140 181772 68168
rect 174096 68128 174102 68140
rect 181766 68128 181772 68140
rect 181824 68128 181830 68180
rect 225466 68128 225472 68180
rect 225524 68168 225530 68180
rect 233562 68168 233568 68180
rect 225524 68140 233568 68168
rect 225524 68128 225530 68140
rect 233562 68128 233568 68140
rect 233620 68128 233626 68180
rect 87282 68100 87288 68112
rect 85460 68072 87288 68100
rect 87282 68060 87288 68072
rect 87340 68060 87346 68112
rect 132546 68060 132552 68112
rect 132604 68100 132610 68112
rect 136410 68100 136416 68112
rect 132604 68072 136416 68100
rect 132604 68060 132610 68072
rect 136410 68060 136416 68072
rect 136468 68060 136474 68112
rect 173946 68060 173952 68112
rect 174004 68100 174010 68112
rect 181582 68100 181588 68112
rect 174004 68072 181588 68100
rect 174004 68060 174010 68072
rect 181582 68060 181588 68072
rect 181640 68060 181646 68112
rect 225558 68060 225564 68112
rect 225616 68100 225622 68112
rect 233654 68100 233660 68112
rect 225616 68072 233660 68100
rect 225616 68060 225622 68072
rect 233654 68060 233660 68072
rect 233712 68060 233718 68112
rect 131810 67992 131816 68044
rect 131868 68032 131874 68044
rect 136594 68032 136600 68044
rect 131868 68004 136600 68032
rect 131868 67992 131874 68004
rect 136594 67992 136600 68004
rect 136652 67992 136658 68044
rect 225834 67992 225840 68044
rect 225892 68032 225898 68044
rect 233470 68032 233476 68044
rect 225892 68004 233476 68032
rect 225892 67992 225898 68004
rect 233470 67992 233476 68004
rect 233528 67992 233534 68044
rect 131350 67924 131356 67976
rect 131408 67964 131414 67976
rect 136686 67964 136692 67976
rect 131408 67936 136692 67964
rect 131408 67924 131414 67936
rect 136686 67924 136692 67936
rect 136744 67924 136750 67976
rect 226294 67924 226300 67976
rect 226352 67964 226358 67976
rect 233746 67964 233752 67976
rect 226352 67936 233752 67964
rect 226352 67924 226358 67936
rect 233746 67924 233752 67936
rect 233804 67924 233810 67976
rect 80198 67516 80204 67568
rect 80256 67556 80262 67568
rect 87190 67556 87196 67568
rect 80256 67528 87196 67556
rect 80256 67516 80262 67528
rect 87190 67516 87196 67528
rect 87248 67516 87254 67568
rect 80106 67448 80112 67500
rect 80164 67488 80170 67500
rect 87282 67488 87288 67500
rect 80164 67460 87288 67488
rect 80164 67448 80170 67460
rect 87282 67448 87288 67460
rect 87340 67448 87346 67500
rect 173486 67448 173492 67500
rect 173544 67488 173550 67500
rect 182318 67488 182324 67500
rect 173544 67460 182324 67488
rect 173544 67448 173550 67460
rect 182318 67448 182324 67460
rect 182376 67448 182382 67500
rect 133006 66904 133012 66956
rect 133064 66944 133070 66956
rect 139630 66944 139636 66956
rect 133064 66916 139636 66944
rect 133064 66904 133070 66916
rect 139630 66904 139636 66916
rect 139688 66904 139694 66956
rect 136686 66768 136692 66820
rect 136744 66808 136750 66820
rect 139722 66808 139728 66820
rect 136744 66780 139728 66808
rect 136744 66768 136750 66780
rect 139722 66768 139728 66780
rect 139780 66768 139786 66820
rect 173854 66700 173860 66752
rect 173912 66740 173918 66752
rect 181398 66740 181404 66752
rect 173912 66712 181404 66740
rect 173912 66700 173918 66712
rect 181398 66700 181404 66712
rect 181456 66700 181462 66752
rect 226294 66700 226300 66752
rect 226352 66740 226358 66752
rect 233470 66740 233476 66752
rect 226352 66712 233476 66740
rect 226352 66700 226358 66712
rect 233470 66700 233476 66712
rect 233528 66700 233534 66752
rect 132178 66632 132184 66684
rect 132236 66672 132242 66684
rect 136778 66672 136784 66684
rect 132236 66644 136784 66672
rect 132236 66632 132242 66644
rect 136778 66632 136784 66644
rect 136836 66632 136842 66684
rect 173578 66632 173584 66684
rect 173636 66672 173642 66684
rect 182318 66672 182324 66684
rect 173636 66644 182324 66672
rect 173636 66632 173642 66644
rect 182318 66632 182324 66644
rect 182376 66632 182382 66684
rect 226018 66632 226024 66684
rect 226076 66672 226082 66684
rect 233562 66672 233568 66684
rect 226076 66644 233568 66672
rect 226076 66632 226082 66644
rect 233562 66632 233568 66644
rect 233620 66632 233626 66684
rect 131350 66564 131356 66616
rect 131408 66604 131414 66616
rect 136502 66604 136508 66616
rect 131408 66576 136508 66604
rect 131408 66564 131414 66576
rect 136502 66564 136508 66576
rect 136560 66564 136566 66616
rect 174038 66564 174044 66616
rect 174096 66604 174102 66616
rect 182226 66604 182232 66616
rect 174096 66576 182232 66604
rect 174096 66564 174102 66576
rect 182226 66564 182232 66576
rect 182284 66564 182290 66616
rect 131350 66156 131356 66208
rect 131408 66196 131414 66208
rect 133006 66196 133012 66208
rect 131408 66168 133012 66196
rect 131408 66156 131414 66168
rect 133006 66156 133012 66168
rect 133064 66156 133070 66208
rect 80198 66088 80204 66140
rect 80256 66128 80262 66140
rect 87190 66128 87196 66140
rect 80256 66100 87196 66128
rect 80256 66088 80262 66100
rect 87190 66088 87196 66100
rect 87248 66088 87254 66140
rect 80106 66020 80112 66072
rect 80164 66060 80170 66072
rect 87282 66060 87288 66072
rect 80164 66032 87288 66060
rect 80164 66020 80170 66032
rect 87282 66020 87288 66032
rect 87340 66020 87346 66072
rect 226386 66020 226392 66072
rect 226444 66060 226450 66072
rect 233470 66060 233476 66072
rect 226444 66032 233476 66060
rect 226444 66020 226450 66032
rect 233470 66020 233476 66032
rect 233528 66020 233534 66072
rect 80198 65340 80204 65392
rect 80256 65380 80262 65392
rect 87190 65380 87196 65392
rect 80256 65352 87196 65380
rect 80256 65340 80262 65352
rect 87190 65340 87196 65352
rect 87248 65340 87254 65392
rect 131810 65340 131816 65392
rect 131868 65380 131874 65392
rect 139630 65380 139636 65392
rect 131868 65352 139636 65380
rect 131868 65340 131874 65352
rect 139630 65340 139636 65352
rect 139688 65340 139694 65392
rect 173486 65340 173492 65392
rect 173544 65380 173550 65392
rect 182318 65380 182324 65392
rect 173544 65352 182324 65380
rect 173544 65340 173550 65352
rect 182318 65340 182324 65352
rect 182376 65340 182382 65392
rect 226294 65340 226300 65392
rect 226352 65380 226358 65392
rect 233470 65380 233476 65392
rect 226352 65352 233476 65380
rect 226352 65340 226358 65352
rect 233470 65340 233476 65352
rect 233528 65340 233534 65392
rect 131442 65272 131448 65324
rect 131500 65312 131506 65324
rect 139722 65312 139728 65324
rect 131500 65284 139728 65312
rect 131500 65272 131506 65284
rect 139722 65272 139728 65284
rect 139780 65272 139786 65324
rect 173762 65272 173768 65324
rect 173820 65312 173826 65324
rect 181398 65312 181404 65324
rect 173820 65284 181404 65312
rect 173820 65272 173826 65284
rect 181398 65272 181404 65284
rect 181456 65272 181462 65324
rect 131350 65204 131356 65256
rect 131408 65244 131414 65256
rect 136686 65244 136692 65256
rect 131408 65216 136692 65244
rect 131408 65204 131414 65216
rect 136686 65204 136692 65216
rect 136744 65204 136750 65256
rect 80106 64728 80112 64780
rect 80164 64768 80170 64780
rect 87190 64768 87196 64780
rect 80164 64740 87196 64768
rect 80164 64728 80170 64740
rect 87190 64728 87196 64740
rect 87248 64728 87254 64780
rect 226294 64728 226300 64780
rect 226352 64768 226358 64780
rect 233562 64768 233568 64780
rect 226352 64740 233568 64768
rect 226352 64728 226358 64740
rect 233562 64728 233568 64740
rect 233620 64728 233626 64780
rect 80198 64660 80204 64712
rect 80256 64700 80262 64712
rect 87282 64700 87288 64712
rect 80256 64672 87288 64700
rect 80256 64660 80262 64672
rect 87282 64660 87288 64672
rect 87340 64660 87346 64712
rect 226386 64660 226392 64712
rect 226444 64700 226450 64712
rect 233470 64700 233476 64712
rect 226444 64672 233476 64700
rect 226444 64660 226450 64672
rect 233470 64660 233476 64672
rect 233528 64660 233534 64712
rect 80198 63980 80204 64032
rect 80256 64020 80262 64032
rect 87650 64020 87656 64032
rect 80256 63992 87656 64020
rect 80256 63980 80262 63992
rect 87650 63980 87656 63992
rect 87708 63980 87714 64032
rect 131350 63980 131356 64032
rect 131408 64020 131414 64032
rect 139630 64020 139636 64032
rect 131408 63992 139636 64020
rect 131408 63980 131414 63992
rect 139630 63980 139636 63992
rect 139688 63980 139694 64032
rect 173854 63980 173860 64032
rect 173912 64020 173918 64032
rect 181030 64020 181036 64032
rect 173912 63992 181036 64020
rect 173912 63980 173918 63992
rect 181030 63980 181036 63992
rect 181088 63980 181094 64032
rect 131810 63912 131816 63964
rect 131868 63952 131874 63964
rect 139722 63952 139728 63964
rect 131868 63924 139728 63952
rect 131868 63912 131874 63924
rect 139722 63912 139728 63924
rect 139780 63912 139786 63964
rect 173946 63912 173952 63964
rect 174004 63952 174010 63964
rect 181122 63952 181128 63964
rect 174004 63924 181128 63952
rect 174004 63912 174010 63924
rect 181122 63912 181128 63924
rect 181180 63912 181186 63964
rect 174038 63844 174044 63896
rect 174096 63884 174102 63896
rect 181306 63884 181312 63896
rect 174096 63856 181312 63884
rect 174096 63844 174102 63856
rect 181306 63844 181312 63856
rect 181364 63844 181370 63896
rect 226294 63436 226300 63488
rect 226352 63476 226358 63488
rect 233654 63476 233660 63488
rect 226352 63448 233660 63476
rect 226352 63436 226358 63448
rect 233654 63436 233660 63448
rect 233712 63436 233718 63488
rect 131994 63368 132000 63420
rect 132052 63408 132058 63420
rect 139630 63408 139636 63420
rect 132052 63380 139636 63408
rect 132052 63368 132058 63380
rect 139630 63368 139636 63380
rect 139688 63368 139694 63420
rect 226386 63368 226392 63420
rect 226444 63408 226450 63420
rect 233470 63408 233476 63420
rect 226444 63380 233476 63408
rect 226444 63368 226450 63380
rect 233470 63368 233476 63380
rect 233528 63368 233534 63420
rect 80198 63300 80204 63352
rect 80256 63340 80262 63352
rect 87190 63340 87196 63352
rect 80256 63312 87196 63340
rect 80256 63300 80262 63312
rect 87190 63300 87196 63312
rect 87248 63300 87254 63352
rect 131350 63300 131356 63352
rect 131408 63340 131414 63352
rect 139722 63340 139728 63352
rect 131408 63312 139728 63340
rect 131408 63300 131414 63312
rect 139722 63300 139728 63312
rect 139780 63300 139786 63352
rect 226294 63300 226300 63352
rect 226352 63340 226358 63352
rect 233562 63340 233568 63352
rect 226352 63312 233568 63340
rect 226352 63300 226358 63312
rect 233562 63300 233568 63312
rect 233620 63300 233626 63352
rect 226294 62620 226300 62672
rect 226352 62660 226358 62672
rect 233470 62660 233476 62672
rect 226352 62632 233476 62660
rect 226352 62620 226358 62632
rect 233470 62620 233476 62632
rect 233528 62620 233534 62672
rect 80198 62552 80204 62604
rect 80256 62592 80262 62604
rect 87282 62592 87288 62604
rect 80256 62564 87288 62592
rect 80256 62552 80262 62564
rect 87282 62552 87288 62564
rect 87340 62552 87346 62604
rect 173762 62552 173768 62604
rect 173820 62592 173826 62604
rect 182318 62592 182324 62604
rect 173820 62564 182324 62592
rect 173820 62552 173826 62564
rect 182318 62552 182324 62564
rect 182376 62552 182382 62604
rect 80106 62484 80112 62536
rect 80164 62524 80170 62536
rect 87190 62524 87196 62536
rect 80164 62496 87196 62524
rect 80164 62484 80170 62496
rect 87190 62484 87196 62496
rect 87248 62484 87254 62536
rect 173302 62484 173308 62536
rect 173360 62524 173366 62536
rect 181398 62524 181404 62536
rect 173360 62496 181404 62524
rect 173360 62484 173366 62496
rect 181398 62484 181404 62496
rect 181456 62484 181462 62536
rect 131442 61940 131448 61992
rect 131500 61980 131506 61992
rect 139722 61980 139728 61992
rect 131500 61952 139728 61980
rect 131500 61940 131506 61952
rect 139722 61940 139728 61952
rect 139780 61940 139786 61992
rect 131350 61872 131356 61924
rect 131408 61912 131414 61924
rect 139630 61912 139636 61924
rect 131408 61884 139636 61912
rect 131408 61872 131414 61884
rect 139630 61872 139636 61884
rect 139688 61872 139694 61924
rect 226386 61872 226392 61924
rect 226444 61912 226450 61924
rect 233470 61912 233476 61924
rect 226444 61884 233476 61912
rect 226444 61872 226450 61884
rect 233470 61872 233476 61884
rect 233528 61872 233534 61924
rect 226202 61328 226208 61380
rect 226260 61368 226266 61380
rect 233470 61368 233476 61380
rect 226260 61340 233476 61368
rect 226260 61328 226266 61340
rect 233470 61328 233476 61340
rect 233528 61328 233534 61380
rect 131350 61260 131356 61312
rect 131408 61300 131414 61312
rect 131408 61272 137284 61300
rect 131408 61260 131414 61272
rect 80198 61192 80204 61244
rect 80256 61232 80262 61244
rect 87282 61232 87288 61244
rect 80256 61204 87288 61232
rect 80256 61192 80262 61204
rect 87282 61192 87288 61204
rect 87340 61192 87346 61244
rect 137256 61232 137284 61272
rect 226294 61260 226300 61312
rect 226352 61300 226358 61312
rect 233562 61300 233568 61312
rect 226352 61272 233568 61300
rect 226352 61260 226358 61272
rect 233562 61260 233568 61272
rect 233620 61260 233626 61312
rect 139630 61232 139636 61244
rect 137256 61204 139636 61232
rect 139630 61192 139636 61204
rect 139688 61192 139694 61244
rect 173670 61192 173676 61244
rect 173728 61232 173734 61244
rect 182226 61232 182232 61244
rect 173728 61204 182232 61232
rect 173728 61192 173734 61204
rect 182226 61192 182232 61204
rect 182284 61192 182290 61244
rect 80106 61124 80112 61176
rect 80164 61164 80170 61176
rect 87190 61164 87196 61176
rect 80164 61136 87196 61164
rect 80164 61124 80170 61136
rect 87190 61124 87196 61136
rect 87248 61124 87254 61176
rect 174038 61124 174044 61176
rect 174096 61164 174102 61176
rect 182134 61164 182140 61176
rect 174096 61136 182140 61164
rect 174096 61124 174102 61136
rect 182134 61124 182140 61136
rect 182192 61124 182198 61176
rect 173946 61056 173952 61108
rect 174004 61096 174010 61108
rect 182042 61096 182048 61108
rect 174004 61068 182048 61096
rect 174004 61056 174010 61068
rect 182042 61056 182048 61068
rect 182100 61056 182106 61108
rect 131350 60580 131356 60632
rect 131408 60620 131414 60632
rect 139722 60620 139728 60632
rect 131408 60592 139728 60620
rect 131408 60580 131414 60592
rect 139722 60580 139728 60592
rect 139780 60580 139786 60632
rect 131442 60512 131448 60564
rect 131500 60552 131506 60564
rect 139630 60552 139636 60564
rect 131500 60524 139636 60552
rect 131500 60512 131506 60524
rect 139630 60512 139636 60524
rect 139688 60512 139694 60564
rect 79094 60308 79100 60360
rect 79152 60348 79158 60360
rect 87006 60348 87012 60360
rect 79152 60320 87012 60348
rect 79152 60308 79158 60320
rect 87006 60308 87012 60320
rect 87064 60308 87070 60360
rect 226386 60104 226392 60156
rect 226444 60144 226450 60156
rect 233746 60144 233752 60156
rect 226444 60116 233752 60144
rect 226444 60104 226450 60116
rect 233746 60104 233752 60116
rect 233804 60104 233810 60156
rect 226294 60036 226300 60088
rect 226352 60076 226358 60088
rect 233838 60076 233844 60088
rect 226352 60048 233844 60076
rect 226352 60036 226358 60048
rect 233838 60036 233844 60048
rect 233896 60036 233902 60088
rect 131810 59968 131816 60020
rect 131868 60008 131874 60020
rect 137238 60008 137244 60020
rect 131868 59980 137244 60008
rect 131868 59968 131874 59980
rect 137238 59968 137244 59980
rect 137296 59968 137302 60020
rect 176890 59968 176896 60020
rect 176948 60008 176954 60020
rect 182226 60008 182232 60020
rect 176948 59980 182232 60008
rect 176948 59968 176954 59980
rect 182226 59968 182232 59980
rect 182284 59968 182290 60020
rect 225742 59968 225748 60020
rect 225800 60008 225806 60020
rect 233470 60008 233476 60020
rect 225800 59980 233476 60008
rect 225800 59968 225806 59980
rect 233470 59968 233476 59980
rect 233528 59968 233534 60020
rect 131350 59900 131356 59952
rect 131408 59940 131414 59952
rect 131408 59912 137560 59940
rect 131408 59900 131414 59912
rect 80106 59832 80112 59884
rect 80164 59872 80170 59884
rect 87190 59872 87196 59884
rect 80164 59844 87196 59872
rect 80164 59832 80170 59844
rect 87190 59832 87196 59844
rect 87248 59832 87254 59884
rect 137532 59872 137560 59912
rect 176982 59900 176988 59952
rect 177040 59940 177046 59952
rect 182318 59940 182324 59952
rect 177040 59912 182324 59940
rect 177040 59900 177046 59912
rect 182318 59900 182324 59912
rect 182376 59900 182382 59952
rect 225926 59900 225932 59952
rect 225984 59940 225990 59952
rect 233562 59940 233568 59952
rect 225984 59912 233568 59940
rect 225984 59900 225990 59912
rect 233562 59900 233568 59912
rect 233620 59900 233626 59952
rect 139630 59872 139636 59884
rect 137532 59844 139636 59872
rect 139630 59832 139636 59844
rect 139688 59832 139694 59884
rect 173854 59832 173860 59884
rect 173912 59872 173918 59884
rect 181950 59872 181956 59884
rect 173912 59844 181956 59872
rect 173912 59832 173918 59844
rect 181950 59832 181956 59844
rect 182008 59832 182014 59884
rect 80198 59764 80204 59816
rect 80256 59804 80262 59816
rect 87098 59804 87104 59816
rect 80256 59776 87104 59804
rect 80256 59764 80262 59776
rect 87098 59764 87104 59776
rect 87156 59764 87162 59816
rect 173670 59764 173676 59816
rect 173728 59804 173734 59816
rect 181858 59804 181864 59816
rect 173728 59776 181864 59804
rect 173728 59764 173734 59776
rect 181858 59764 181864 59776
rect 181916 59764 181922 59816
rect 174038 59696 174044 59748
rect 174096 59736 174102 59748
rect 181766 59736 181772 59748
rect 174096 59708 181772 59736
rect 174096 59696 174102 59708
rect 181766 59696 181772 59708
rect 181824 59696 181830 59748
rect 137238 59220 137244 59272
rect 137296 59260 137302 59272
rect 139722 59260 139728 59272
rect 137296 59232 139728 59260
rect 137296 59220 137302 59232
rect 139722 59220 139728 59232
rect 139780 59220 139786 59272
rect 135769 58787 135827 58793
rect 135769 58753 135781 58787
rect 135815 58784 135827 58787
rect 139814 58784 139820 58796
rect 135815 58756 139820 58784
rect 135815 58753 135827 58756
rect 135769 58747 135827 58753
rect 139814 58744 139820 58756
rect 139872 58744 139878 58796
rect 131534 58676 131540 58728
rect 131592 58716 131598 58728
rect 131592 58688 137560 58716
rect 131592 58676 131598 58688
rect 131442 58608 131448 58660
rect 131500 58648 131506 58660
rect 131500 58620 137468 58648
rect 131500 58608 131506 58620
rect 80014 58540 80020 58592
rect 80072 58580 80078 58592
rect 87190 58580 87196 58592
rect 80072 58552 87196 58580
rect 80072 58540 80078 58552
rect 87190 58540 87196 58552
rect 87248 58540 87254 58592
rect 131350 58540 131356 58592
rect 131408 58580 131414 58592
rect 135769 58583 135827 58589
rect 135769 58580 135781 58583
rect 131408 58552 135781 58580
rect 131408 58540 131414 58552
rect 135769 58549 135781 58552
rect 135815 58549 135827 58583
rect 135769 58543 135827 58549
rect 80106 58472 80112 58524
rect 80164 58512 80170 58524
rect 87006 58512 87012 58524
rect 80164 58484 87012 58512
rect 80164 58472 80170 58484
rect 87006 58472 87012 58484
rect 87064 58472 87070 58524
rect 80198 58404 80204 58456
rect 80256 58444 80262 58456
rect 86914 58444 86920 58456
rect 80256 58416 86920 58444
rect 80256 58404 80262 58416
rect 86914 58404 86920 58416
rect 86972 58404 86978 58456
rect 137440 58444 137468 58620
rect 137532 58512 137560 58688
rect 226202 58676 226208 58728
rect 226260 58716 226266 58728
rect 233470 58716 233476 58728
rect 226260 58688 233476 58716
rect 226260 58676 226266 58688
rect 233470 58676 233476 58688
rect 233528 58676 233534 58728
rect 226386 58608 226392 58660
rect 226444 58648 226450 58660
rect 233562 58648 233568 58660
rect 226444 58620 233568 58648
rect 226444 58608 226450 58620
rect 233562 58608 233568 58620
rect 233620 58608 233626 58660
rect 226294 58540 226300 58592
rect 226352 58580 226358 58592
rect 233654 58580 233660 58592
rect 226352 58552 233660 58580
rect 226352 58540 226358 58552
rect 233654 58540 233660 58552
rect 233712 58540 233718 58592
rect 139630 58512 139636 58524
rect 137532 58484 139636 58512
rect 139630 58472 139636 58484
rect 139688 58472 139694 58524
rect 173762 58472 173768 58524
rect 173820 58512 173826 58524
rect 182134 58512 182140 58524
rect 173820 58484 182140 58512
rect 173820 58472 173826 58484
rect 182134 58472 182140 58484
rect 182192 58472 182198 58524
rect 139722 58444 139728 58456
rect 137440 58416 139728 58444
rect 139722 58404 139728 58416
rect 139780 58404 139786 58456
rect 174038 58404 174044 58456
rect 174096 58444 174102 58456
rect 181674 58444 181680 58456
rect 174096 58416 181680 58444
rect 174096 58404 174102 58416
rect 181674 58404 181680 58416
rect 181732 58404 181738 58456
rect 177994 57656 178000 57708
rect 178052 57696 178058 57708
rect 182318 57696 182324 57708
rect 178052 57668 182324 57696
rect 178052 57656 178058 57668
rect 182318 57656 182324 57668
rect 182376 57656 182382 57708
rect 177626 57520 177632 57572
rect 177684 57560 177690 57572
rect 181674 57560 181680 57572
rect 177684 57532 181680 57560
rect 177684 57520 177690 57532
rect 181674 57520 181680 57532
rect 181732 57520 181738 57572
rect 80198 57316 80204 57368
rect 80256 57356 80262 57368
rect 86822 57356 86828 57368
rect 80256 57328 86828 57356
rect 80256 57316 80262 57328
rect 86822 57316 86828 57328
rect 86880 57316 86886 57368
rect 131350 57316 131356 57368
rect 131408 57356 131414 57368
rect 136226 57356 136232 57368
rect 131408 57328 136232 57356
rect 131408 57316 131414 57328
rect 136226 57316 136232 57328
rect 136284 57316 136290 57368
rect 139906 57356 139912 57368
rect 137440 57328 139912 57356
rect 131534 57248 131540 57300
rect 131592 57288 131598 57300
rect 137330 57288 137336 57300
rect 131592 57260 137336 57288
rect 131592 57248 131598 57260
rect 137330 57248 137336 57260
rect 137388 57248 137394 57300
rect 131442 57180 131448 57232
rect 131500 57220 131506 57232
rect 137440 57220 137468 57328
rect 139906 57316 139912 57328
rect 139964 57316 139970 57368
rect 225742 57316 225748 57368
rect 225800 57356 225806 57368
rect 228042 57356 228048 57368
rect 225800 57328 228048 57356
rect 225800 57316 225806 57328
rect 228042 57316 228048 57328
rect 228100 57316 228106 57368
rect 177718 57248 177724 57300
rect 177776 57288 177782 57300
rect 181582 57288 181588 57300
rect 177776 57260 181588 57288
rect 177776 57248 177782 57260
rect 181582 57248 181588 57260
rect 181640 57248 181646 57300
rect 225834 57248 225840 57300
rect 225892 57288 225898 57300
rect 228594 57288 228600 57300
rect 225892 57260 228600 57288
rect 225892 57248 225898 57260
rect 228594 57248 228600 57260
rect 228652 57248 228658 57300
rect 131500 57192 137468 57220
rect 131500 57180 131506 57192
rect 226478 57180 226484 57232
rect 226536 57220 226542 57232
rect 228686 57220 228692 57232
rect 226536 57192 228692 57220
rect 226536 57180 226542 57192
rect 228686 57180 228692 57192
rect 228744 57180 228750 57232
rect 131626 57112 131632 57164
rect 131684 57152 131690 57164
rect 139722 57152 139728 57164
rect 131684 57124 139728 57152
rect 131684 57112 131690 57124
rect 139722 57112 139728 57124
rect 139780 57112 139786 57164
rect 225926 57112 225932 57164
rect 225984 57152 225990 57164
rect 227950 57152 227956 57164
rect 225984 57124 227956 57152
rect 225984 57112 225990 57124
rect 227950 57112 227956 57124
rect 228008 57112 228014 57164
rect 80106 57044 80112 57096
rect 80164 57084 80170 57096
rect 87282 57084 87288 57096
rect 80164 57056 87288 57084
rect 80164 57044 80170 57056
rect 87282 57044 87288 57056
rect 87340 57044 87346 57096
rect 172934 57044 172940 57096
rect 172992 57084 172998 57096
rect 180938 57084 180944 57096
rect 172992 57056 180944 57084
rect 172992 57044 172998 57056
rect 180938 57044 180944 57056
rect 180996 57044 181002 57096
rect 80198 56976 80204 57028
rect 80256 57016 80262 57028
rect 87374 57016 87380 57028
rect 80256 56988 87380 57016
rect 80256 56976 80262 56988
rect 87374 56976 87380 56988
rect 87432 56976 87438 57028
rect 174038 56976 174044 57028
rect 174096 57016 174102 57028
rect 176890 57016 176896 57028
rect 174096 56988 176896 57016
rect 174096 56976 174102 56988
rect 176890 56976 176896 56988
rect 176948 56976 176954 57028
rect 174038 56772 174044 56824
rect 174096 56812 174102 56824
rect 176982 56812 176988 56824
rect 174096 56784 176988 56812
rect 174096 56772 174102 56784
rect 176982 56772 176988 56784
rect 177040 56772 177046 56824
rect 137330 56568 137336 56620
rect 137388 56608 137394 56620
rect 139630 56608 139636 56620
rect 137388 56580 139636 56608
rect 137388 56568 137394 56580
rect 139630 56568 139636 56580
rect 139688 56568 139694 56620
rect 226294 56160 226300 56212
rect 226352 56200 226358 56212
rect 229422 56200 229428 56212
rect 226352 56172 229428 56200
rect 226352 56160 226358 56172
rect 229422 56160 229428 56172
rect 229480 56160 229486 56212
rect 131442 55888 131448 55940
rect 131500 55928 131506 55940
rect 138066 55928 138072 55940
rect 131500 55900 138072 55928
rect 131500 55888 131506 55900
rect 138066 55888 138072 55900
rect 138124 55888 138130 55940
rect 226294 55888 226300 55940
rect 226352 55928 226358 55940
rect 229330 55928 229336 55940
rect 226352 55900 229336 55928
rect 226352 55888 226358 55900
rect 229330 55888 229336 55900
rect 229388 55888 229394 55940
rect 131350 55820 131356 55872
rect 131408 55860 131414 55872
rect 139446 55860 139452 55872
rect 131408 55832 139452 55860
rect 131408 55820 131414 55832
rect 139446 55820 139452 55832
rect 139504 55820 139510 55872
rect 131534 55752 131540 55804
rect 131592 55792 131598 55804
rect 139538 55792 139544 55804
rect 131592 55764 139544 55792
rect 131592 55752 131598 55764
rect 139538 55752 139544 55764
rect 139596 55752 139602 55804
rect 177350 55752 177356 55804
rect 177408 55792 177414 55804
rect 182318 55792 182324 55804
rect 177408 55764 182324 55792
rect 177408 55752 177414 55764
rect 182318 55752 182324 55764
rect 182376 55752 182382 55804
rect 225926 55752 225932 55804
rect 225984 55792 225990 55804
rect 229606 55792 229612 55804
rect 225984 55764 229612 55792
rect 225984 55752 225990 55764
rect 229606 55752 229612 55764
rect 229664 55752 229670 55804
rect 80106 55684 80112 55736
rect 80164 55724 80170 55736
rect 87098 55724 87104 55736
rect 80164 55696 87104 55724
rect 80164 55684 80170 55696
rect 87098 55684 87104 55696
rect 87156 55684 87162 55736
rect 173302 55684 173308 55736
rect 173360 55724 173366 55736
rect 182226 55724 182232 55736
rect 173360 55696 182232 55724
rect 173360 55684 173366 55696
rect 182226 55684 182232 55696
rect 182284 55684 182290 55736
rect 227950 55684 227956 55736
rect 228008 55724 228014 55736
rect 233562 55724 233568 55736
rect 228008 55696 233568 55724
rect 228008 55684 228014 55696
rect 233562 55684 233568 55696
rect 233620 55684 233626 55736
rect 173762 55616 173768 55668
rect 173820 55656 173826 55668
rect 182042 55656 182048 55668
rect 173820 55628 182048 55656
rect 173820 55616 173826 55628
rect 182042 55616 182048 55628
rect 182100 55616 182106 55668
rect 228042 55616 228048 55668
rect 228100 55656 228106 55668
rect 233470 55656 233476 55668
rect 228100 55628 233476 55656
rect 228100 55616 228106 55628
rect 233470 55616 233476 55628
rect 233528 55616 233534 55668
rect 80198 55412 80204 55464
rect 80256 55452 80262 55464
rect 87006 55452 87012 55464
rect 80256 55424 87012 55452
rect 80256 55412 80262 55424
rect 87006 55412 87012 55424
rect 87064 55412 87070 55464
rect 226294 54664 226300 54716
rect 226352 54704 226358 54716
rect 229514 54704 229520 54716
rect 226352 54676 229520 54704
rect 226352 54664 226358 54676
rect 229514 54664 229520 54676
rect 229572 54664 229578 54716
rect 79738 54528 79744 54580
rect 79796 54568 79802 54580
rect 87282 54568 87288 54580
rect 79796 54540 87288 54568
rect 79796 54528 79802 54540
rect 87282 54528 87288 54540
rect 87340 54528 87346 54580
rect 131350 54528 131356 54580
rect 131408 54568 131414 54580
rect 136778 54568 136784 54580
rect 131408 54540 136784 54568
rect 131408 54528 131414 54540
rect 136778 54528 136784 54540
rect 136836 54528 136842 54580
rect 79462 54460 79468 54512
rect 79520 54500 79526 54512
rect 87190 54500 87196 54512
rect 79520 54472 87196 54500
rect 79520 54460 79526 54472
rect 87190 54460 87196 54472
rect 87248 54460 87254 54512
rect 131442 54460 131448 54512
rect 131500 54500 131506 54512
rect 139906 54500 139912 54512
rect 131500 54472 139912 54500
rect 131500 54460 131506 54472
rect 139906 54460 139912 54472
rect 139964 54460 139970 54512
rect 175234 54460 175240 54512
rect 175292 54500 175298 54512
rect 181674 54500 181680 54512
rect 175292 54472 181680 54500
rect 175292 54460 175298 54472
rect 181674 54460 181680 54472
rect 181732 54460 181738 54512
rect 225742 54460 225748 54512
rect 225800 54500 225806 54512
rect 230894 54500 230900 54512
rect 225800 54472 230900 54500
rect 225800 54460 225806 54472
rect 230894 54460 230900 54472
rect 230952 54460 230958 54512
rect 85902 54392 85908 54444
rect 85960 54432 85966 54444
rect 87282 54432 87288 54444
rect 85960 54404 87288 54432
rect 85960 54392 85966 54404
rect 87282 54392 87288 54404
rect 87340 54392 87346 54444
rect 131534 54392 131540 54444
rect 131592 54432 131598 54444
rect 139630 54432 139636 54444
rect 131592 54404 139636 54432
rect 131592 54392 131598 54404
rect 139630 54392 139636 54404
rect 139688 54392 139694 54444
rect 175326 54392 175332 54444
rect 175384 54432 175390 54444
rect 181582 54432 181588 54444
rect 175384 54404 181588 54432
rect 175384 54392 175390 54404
rect 181582 54392 181588 54404
rect 181640 54392 181646 54444
rect 226386 54392 226392 54444
rect 226444 54432 226450 54444
rect 230710 54432 230716 54444
rect 226444 54404 230716 54432
rect 226444 54392 226450 54404
rect 230710 54392 230716 54404
rect 230768 54392 230774 54444
rect 174038 54324 174044 54376
rect 174096 54364 174102 54376
rect 177994 54364 178000 54376
rect 174096 54336 178000 54364
rect 174096 54324 174102 54336
rect 177994 54324 178000 54336
rect 178052 54324 178058 54376
rect 228594 54324 228600 54376
rect 228652 54364 228658 54376
rect 233470 54364 233476 54376
rect 228652 54336 233476 54364
rect 228652 54324 228658 54336
rect 233470 54324 233476 54336
rect 233528 54324 233534 54376
rect 228686 54256 228692 54308
rect 228744 54296 228750 54308
rect 233562 54296 233568 54308
rect 228744 54268 233568 54296
rect 228744 54256 228750 54268
rect 233562 54256 233568 54268
rect 233620 54256 233626 54308
rect 80198 54188 80204 54240
rect 80256 54228 80262 54240
rect 86730 54228 86736 54240
rect 80256 54200 86736 54228
rect 80256 54188 80262 54200
rect 86730 54188 86736 54200
rect 86788 54188 86794 54240
rect 136226 54188 136232 54240
rect 136284 54228 136290 54240
rect 139722 54228 139728 54240
rect 136284 54200 139728 54228
rect 136284 54188 136290 54200
rect 139722 54188 139728 54200
rect 139780 54188 139786 54240
rect 226294 54188 226300 54240
rect 226352 54228 226358 54240
rect 231722 54228 231728 54240
rect 226352 54200 231728 54228
rect 226352 54188 226358 54200
rect 231722 54188 231728 54200
rect 231780 54188 231786 54240
rect 138066 53916 138072 53968
rect 138124 53956 138130 53968
rect 139998 53956 140004 53968
rect 138124 53928 140004 53956
rect 138124 53916 138130 53928
rect 139998 53916 140004 53928
rect 140056 53916 140062 53968
rect 174038 53780 174044 53832
rect 174096 53820 174102 53832
rect 177626 53820 177632 53832
rect 174096 53792 177632 53820
rect 174096 53780 174102 53792
rect 177626 53780 177632 53792
rect 177684 53780 177690 53832
rect 173486 53712 173492 53764
rect 173544 53752 173550 53764
rect 177718 53752 177724 53764
rect 173544 53724 177724 53752
rect 173544 53712 173550 53724
rect 177718 53712 177724 53724
rect 177776 53712 177782 53764
rect 80198 53304 80204 53356
rect 80256 53344 80262 53356
rect 86546 53344 86552 53356
rect 80256 53316 86552 53344
rect 80256 53304 80262 53316
rect 86546 53304 86552 53316
rect 86604 53304 86610 53356
rect 131442 53032 131448 53084
rect 131500 53072 131506 53084
rect 139722 53072 139728 53084
rect 131500 53044 139728 53072
rect 131500 53032 131506 53044
rect 139722 53032 139728 53044
rect 139780 53032 139786 53084
rect 80014 52964 80020 53016
rect 80072 53004 80078 53016
rect 87190 53004 87196 53016
rect 80072 52976 87196 53004
rect 80072 52964 80078 52976
rect 87190 52964 87196 52976
rect 87248 52964 87254 53016
rect 131350 52964 131356 53016
rect 131408 53004 131414 53016
rect 139814 53004 139820 53016
rect 131408 52976 139820 53004
rect 131408 52964 131414 52976
rect 139814 52964 139820 52976
rect 139872 52964 139878 53016
rect 176890 52964 176896 53016
rect 176948 53004 176954 53016
rect 182318 53004 182324 53016
rect 176948 52976 182324 53004
rect 176948 52964 176954 52976
rect 182318 52964 182324 52976
rect 182376 52964 182382 53016
rect 225834 52964 225840 53016
rect 225892 53004 225898 53016
rect 233562 53004 233568 53016
rect 225892 52976 233568 53004
rect 225892 52964 225898 52976
rect 233562 52964 233568 52976
rect 233620 52964 233626 53016
rect 80106 52896 80112 52948
rect 80164 52936 80170 52948
rect 88386 52936 88392 52948
rect 80164 52908 88392 52936
rect 80164 52896 80170 52908
rect 88386 52896 88392 52908
rect 88444 52896 88450 52948
rect 172842 52896 172848 52948
rect 172900 52936 172906 52948
rect 181214 52936 181220 52948
rect 172900 52908 181220 52936
rect 172900 52896 172906 52908
rect 181214 52896 181220 52908
rect 181272 52896 181278 52948
rect 229606 52896 229612 52948
rect 229664 52936 229670 52948
rect 233470 52936 233476 52948
rect 229664 52908 233476 52936
rect 229664 52896 229670 52908
rect 233470 52896 233476 52908
rect 233528 52896 233534 52948
rect 80198 52828 80204 52880
rect 80256 52868 80262 52880
rect 88202 52868 88208 52880
rect 80256 52840 88208 52868
rect 80256 52828 80262 52840
rect 88202 52828 88208 52840
rect 88260 52828 88266 52880
rect 174038 52828 174044 52880
rect 174096 52868 174102 52880
rect 181306 52868 181312 52880
rect 174096 52840 181312 52868
rect 174096 52828 174102 52840
rect 181306 52828 181312 52840
rect 181364 52828 181370 52880
rect 229422 52828 229428 52880
rect 229480 52868 229486 52880
rect 233654 52868 233660 52880
rect 229480 52840 233660 52868
rect 229480 52828 229486 52840
rect 233654 52828 233660 52840
rect 233712 52828 233718 52880
rect 229330 52760 229336 52812
rect 229388 52800 229394 52812
rect 233470 52800 233476 52812
rect 229388 52772 233476 52800
rect 229388 52760 229394 52772
rect 233470 52760 233476 52772
rect 233528 52760 233534 52812
rect 173946 52692 173952 52744
rect 174004 52732 174010 52744
rect 180294 52732 180300 52744
rect 174004 52704 180300 52732
rect 174004 52692 174010 52704
rect 180294 52692 180300 52704
rect 180352 52692 180358 52744
rect 80198 51536 80204 51588
rect 80256 51576 80262 51588
rect 87926 51576 87932 51588
rect 80256 51548 87932 51576
rect 80256 51536 80262 51548
rect 87926 51536 87932 51548
rect 87984 51536 87990 51588
rect 173946 51536 173952 51588
rect 174004 51576 174010 51588
rect 181122 51576 181128 51588
rect 174004 51548 181128 51576
rect 174004 51536 174010 51548
rect 181122 51536 181128 51548
rect 181180 51536 181186 51588
rect 198786 51536 198792 51588
rect 198844 51576 198850 51588
rect 198844 51548 230848 51576
rect 198844 51536 198850 51548
rect 230820 51508 230848 51548
rect 230894 51536 230900 51588
rect 230952 51576 230958 51588
rect 233470 51576 233476 51588
rect 230952 51548 233476 51576
rect 230952 51536 230958 51548
rect 233470 51536 233476 51548
rect 233528 51536 233534 51588
rect 234114 51508 234120 51520
rect 230820 51480 234120 51508
rect 234114 51468 234120 51480
rect 234172 51468 234178 51520
rect 230710 51400 230716 51452
rect 230768 51440 230774 51452
rect 233654 51440 233660 51452
rect 230768 51412 233660 51440
rect 230768 51400 230774 51412
rect 233654 51400 233660 51412
rect 233712 51400 233718 51452
rect 172934 51196 172940 51248
rect 172992 51236 172998 51248
rect 177350 51236 177356 51248
rect 172992 51208 177356 51236
rect 172992 51196 172998 51208
rect 177350 51196 177356 51208
rect 177408 51196 177414 51248
rect 125186 50924 125192 50976
rect 125244 50964 125250 50976
rect 127026 50964 127032 50976
rect 125244 50936 127032 50964
rect 125244 50924 125250 50936
rect 127026 50924 127032 50936
rect 127084 50964 127090 50976
rect 134754 50964 134760 50976
rect 127084 50936 134760 50964
rect 127084 50924 127090 50936
rect 134754 50924 134760 50936
rect 134812 50924 134818 50976
rect 115158 50856 115164 50908
rect 115216 50896 115222 50908
rect 128590 50896 128596 50908
rect 115216 50868 128596 50896
rect 115216 50856 115222 50868
rect 128590 50856 128596 50868
rect 128648 50856 128654 50908
rect 208814 50856 208820 50908
rect 208872 50896 208878 50908
rect 222430 50896 222436 50908
rect 208872 50868 222436 50896
rect 208872 50856 208878 50868
rect 222430 50856 222436 50868
rect 222488 50856 222494 50908
rect 93998 50652 94004 50704
rect 94056 50692 94062 50704
rect 94550 50692 94556 50704
rect 94056 50664 94556 50692
rect 94056 50652 94062 50664
rect 94550 50652 94556 50664
rect 94608 50652 94614 50704
rect 218842 50380 218848 50432
rect 218900 50420 218906 50432
rect 220958 50420 220964 50432
rect 218900 50392 220964 50420
rect 218900 50380 218906 50392
rect 220958 50380 220964 50392
rect 221016 50380 221022 50432
rect 187838 50244 187844 50296
rect 187896 50284 187902 50296
rect 188850 50284 188856 50296
rect 187896 50256 188856 50284
rect 187896 50244 187902 50256
rect 188850 50244 188856 50256
rect 188908 50244 188914 50296
rect 136778 50176 136784 50228
rect 136836 50216 136842 50228
rect 139630 50216 139636 50228
rect 136836 50188 139636 50216
rect 136836 50176 136842 50188
rect 139630 50176 139636 50188
rect 139688 50176 139694 50228
rect 231722 50176 231728 50228
rect 231780 50216 231786 50228
rect 233470 50216 233476 50228
rect 231780 50188 233476 50216
rect 231780 50176 231786 50188
rect 233470 50176 233476 50188
rect 233528 50176 233534 50228
rect 173302 50108 173308 50160
rect 173360 50148 173366 50160
rect 175234 50148 175240 50160
rect 173360 50120 175240 50148
rect 173360 50108 173366 50120
rect 175234 50108 175240 50120
rect 175292 50108 175298 50160
rect 229514 50108 229520 50160
rect 229572 50148 229578 50160
rect 233654 50148 233660 50160
rect 229572 50120 233660 50148
rect 229572 50108 229578 50120
rect 233654 50108 233660 50120
rect 233712 50108 233718 50160
rect 172750 50040 172756 50092
rect 172808 50080 172814 50092
rect 175326 50080 175332 50092
rect 172808 50052 175332 50080
rect 172808 50040 172814 50052
rect 175326 50040 175332 50052
rect 175384 50040 175390 50092
rect 80198 49224 80204 49276
rect 80256 49264 80262 49276
rect 87098 49264 87104 49276
rect 80256 49236 87104 49264
rect 80256 49224 80262 49236
rect 87098 49224 87104 49236
rect 87156 49224 87162 49276
rect 173118 49156 173124 49208
rect 173176 49196 173182 49208
rect 176890 49196 176896 49208
rect 173176 49168 176896 49196
rect 173176 49156 173182 49168
rect 176890 49156 176896 49168
rect 176948 49156 176954 49208
rect 80106 48884 80112 48936
rect 80164 48924 80170 48936
rect 85902 48924 85908 48936
rect 80164 48896 85908 48924
rect 80164 48884 80170 48896
rect 85902 48884 85908 48896
rect 85960 48884 85966 48936
rect 173302 48612 173308 48664
rect 173360 48652 173366 48664
rect 180938 48652 180944 48664
rect 173360 48624 180944 48652
rect 173360 48612 173366 48624
rect 180938 48612 180944 48624
rect 180996 48612 181002 48664
rect 99518 47456 99524 47508
rect 99576 47496 99582 47508
rect 139630 47496 139636 47508
rect 99576 47468 139636 47496
rect 99576 47456 99582 47468
rect 139630 47456 139636 47468
rect 139688 47456 139694 47508
rect 193358 47456 193364 47508
rect 193416 47496 193422 47508
rect 233470 47496 233476 47508
rect 193416 47468 233476 47496
rect 193416 47456 193422 47468
rect 233470 47456 233476 47468
rect 233528 47456 233534 47508
rect 220958 47388 220964 47440
rect 221016 47428 221022 47440
rect 228134 47428 228140 47440
rect 221016 47400 228140 47428
rect 221016 47388 221022 47400
rect 228134 47388 228140 47400
rect 228192 47428 228198 47440
rect 260426 47428 260432 47440
rect 228192 47400 260432 47428
rect 228192 47388 228198 47400
rect 260426 47388 260432 47400
rect 260484 47388 260490 47440
rect 62902 46028 62908 46080
rect 62960 46068 62966 46080
rect 63638 46068 63644 46080
rect 62960 46040 63644 46068
rect 62960 46028 62966 46040
rect 63638 46028 63644 46040
rect 63696 46028 63702 46080
rect 276066 46028 276072 46080
rect 276124 46068 276130 46080
rect 300170 46068 300176 46080
rect 276124 46040 300176 46068
rect 276124 46028 276130 46040
rect 300170 46028 300176 46040
rect 300228 46028 300234 46080
rect 260426 45348 260432 45400
rect 260484 45388 260490 45400
rect 284530 45388 284536 45400
rect 260484 45360 284536 45388
rect 260484 45348 260490 45360
rect 284530 45348 284536 45360
rect 284588 45348 284594 45400
rect 93078 37732 93084 37784
rect 93136 37772 93142 37784
rect 93998 37772 94004 37784
rect 93136 37744 94004 37772
rect 93136 37732 93142 37744
rect 93998 37732 94004 37744
rect 94056 37732 94062 37784
rect 98782 37732 98788 37784
rect 98840 37772 98846 37784
rect 99518 37772 99524 37784
rect 98840 37744 99524 37772
rect 98840 37732 98846 37744
rect 99518 37732 99524 37744
rect 99576 37732 99582 37784
rect 192438 37732 192444 37784
rect 192496 37772 192502 37784
rect 193358 37772 193364 37784
rect 192496 37744 193364 37772
rect 192496 37732 192502 37744
rect 193358 37732 193364 37744
rect 193416 37732 193422 37784
rect 186734 37392 186740 37444
rect 186792 37432 186798 37444
rect 187838 37432 187844 37444
rect 186792 37404 187844 37432
rect 186792 37392 186798 37404
rect 187838 37392 187844 37404
rect 187896 37392 187902 37444
rect 79554 37188 79560 37240
rect 79612 37228 79618 37240
rect 103842 37228 103848 37240
rect 79612 37200 103848 37228
rect 79612 37188 79618 37200
rect 103842 37188 103848 37200
rect 103900 37188 103906 37240
rect 173394 37188 173400 37240
rect 173452 37228 173458 37240
rect 198142 37228 198148 37240
rect 173452 37200 198148 37228
rect 173452 37188 173458 37200
rect 198142 37188 198148 37200
rect 198200 37188 198206 37240
rect 13498 37120 13504 37172
rect 13556 37160 13562 37172
rect 120954 37160 120960 37172
rect 13556 37132 120960 37160
rect 13556 37120 13562 37132
rect 120954 37120 120960 37132
rect 121012 37120 121018 37172
rect 140918 37120 140924 37172
rect 140976 37160 140982 37172
rect 203846 37160 203852 37172
rect 140976 37132 203852 37160
rect 140976 37120 140982 37132
rect 203846 37120 203852 37132
rect 203904 37120 203910 37172
rect 209550 37120 209556 37172
rect 209608 37160 209614 37172
rect 292626 37160 292632 37172
rect 209608 37132 292632 37160
rect 209608 37120 209614 37132
rect 292626 37120 292632 37132
rect 292684 37120 292690 37172
rect 63638 37052 63644 37104
rect 63696 37092 63702 37104
rect 109546 37092 109552 37104
rect 63696 37064 109552 37092
rect 63696 37052 63702 37064
rect 109546 37052 109552 37064
rect 109604 37052 109610 37104
rect 115802 37052 115808 37104
rect 115860 37092 115866 37104
rect 292534 37092 292540 37104
rect 115860 37064 292540 37092
rect 115860 37052 115866 37064
rect 292534 37052 292540 37064
rect 292592 37052 292598 37104
rect 128866 28008 128872 28060
rect 128924 28048 128930 28060
rect 129510 28048 129516 28060
rect 128924 28020 129516 28048
rect 128924 28008 128930 28020
rect 129510 28008 129516 28020
rect 129568 28008 129574 28060
rect 222798 28008 222804 28060
rect 222856 28048 222862 28060
rect 223534 28048 223540 28060
rect 222856 28020 223540 28048
rect 222856 28008 222862 28020
rect 223534 28008 223540 28020
rect 223592 28008 223598 28060
rect 13314 25356 13320 25408
rect 13372 25396 13378 25408
rect 85074 25396 85080 25408
rect 13372 25368 85080 25396
rect 13372 25356 13378 25368
rect 85074 25356 85080 25368
rect 85132 25356 85138 25408
rect 76518 20868 76524 20920
rect 76576 20908 76582 20920
rect 299802 20908 299808 20920
rect 76576 20880 299808 20908
rect 76576 20868 76582 20880
rect 299802 20868 299808 20880
rect 299860 20868 299866 20920
rect 13590 17060 13596 17112
rect 13648 17100 13654 17112
rect 109546 17100 109552 17112
rect 13648 17072 109552 17100
rect 13648 17060 13654 17072
rect 109546 17060 109552 17072
rect 109604 17060 109610 17112
rect 203846 17060 203852 17112
rect 203904 17100 203910 17112
rect 265854 17100 265860 17112
rect 203904 17072 265860 17100
rect 203904 17060 203910 17072
rect 265854 17060 265860 17072
rect 265912 17060 265918 17112
rect 38154 12436 38160 12488
rect 38212 12476 38218 12488
rect 138434 12476 138440 12488
rect 38212 12448 138440 12476
rect 38212 12436 38218 12448
rect 138434 12436 138440 12448
rect 138492 12436 138498 12488
rect 28218 12368 28224 12420
rect 28276 12408 28282 12420
rect 133374 12408 133380 12420
rect 28276 12380 133380 12408
rect 28276 12368 28282 12380
rect 133374 12368 133380 12380
rect 133432 12368 133438 12420
rect 88478 12300 88484 12352
rect 88536 12340 88542 12352
rect 248742 12340 248748 12352
rect 88536 12312 248748 12340
rect 88536 12300 88542 12312
rect 248742 12300 248748 12312
rect 248800 12300 248806 12352
rect 64926 12232 64932 12284
rect 64984 12272 64990 12284
rect 264658 12272 264664 12284
rect 64984 12244 264664 12272
rect 64984 12232 64990 12244
rect 264658 12232 264664 12244
rect 264716 12232 264722 12284
rect 175234 9376 175240 9428
rect 175292 9416 175298 9428
rect 175418 9416 175424 9428
rect 175292 9388 175424 9416
rect 175292 9376 175298 9388
rect 175418 9376 175424 9388
rect 175476 9376 175482 9428
rect 284530 9376 284536 9428
rect 284588 9416 284594 9428
rect 285450 9416 285456 9428
rect 284588 9388 285456 9416
rect 284588 9376 284594 9388
rect 285450 9376 285456 9388
rect 285508 9376 285514 9428
<< via1 >>
rect 34664 299396 34716 299448
rect 211948 299396 212000 299448
rect 248748 299396 248800 299448
rect 267240 299396 267292 299448
rect 101732 299328 101784 299380
rect 292540 299328 292592 299380
rect 34572 299260 34624 299312
rect 285456 299260 285508 299312
rect 28224 298648 28276 298700
rect 29144 298648 29196 298700
rect 138440 298648 138492 298700
rect 139544 298648 139596 298700
rect 65024 295112 65076 295164
rect 96212 295112 96264 295164
rect 139544 295112 139596 295164
rect 203852 295112 203904 295164
rect 123536 294636 123588 294688
rect 264756 294636 264808 294688
rect 13412 294568 13464 294620
rect 190512 294568 190564 294620
rect 217192 294568 217244 294620
rect 265860 294568 265912 294620
rect 110196 294500 110248 294552
rect 292632 294500 292684 294552
rect 13228 286204 13280 286256
rect 20220 286204 20272 286256
rect 175240 276659 175292 276668
rect 175240 276625 175249 276659
rect 175249 276625 175283 276659
rect 175283 276625 175292 276659
rect 175240 276616 175292 276625
rect 79560 274440 79612 274492
rect 114796 274440 114848 274492
rect 173400 274440 173452 274492
rect 208820 274440 208872 274492
rect 218848 274440 218900 274492
rect 225288 274440 225340 274492
rect 175240 272375 175292 272384
rect 175240 272341 175249 272375
rect 175249 272341 175283 272375
rect 175283 272341 175292 272375
rect 175240 272332 175292 272341
rect 175240 269612 175292 269664
rect 265860 266824 265912 266876
rect 300084 266824 300136 266876
rect 78916 264036 78968 264088
rect 124456 264036 124508 264088
rect 125744 264036 125796 264088
rect 143040 264036 143092 264088
rect 225196 264036 225248 264088
rect 198884 263968 198936 264020
rect 233476 263968 233528 264020
rect 125744 263356 125796 263408
rect 132736 263356 132788 263408
rect 139636 263356 139688 263408
rect 105044 262676 105096 262728
rect 139636 262676 139688 262728
rect 47084 262608 47136 262660
rect 131356 262608 131408 262660
rect 175332 262651 175384 262660
rect 175332 262617 175341 262651
rect 175341 262617 175375 262651
rect 175375 262617 175384 262651
rect 175332 262608 175384 262617
rect 80112 261452 80164 261504
rect 87196 261452 87248 261504
rect 173584 261452 173636 261504
rect 181956 261452 182008 261504
rect 80204 261384 80256 261436
rect 87288 261384 87340 261436
rect 173676 261384 173728 261436
rect 181772 261384 181824 261436
rect 95384 260636 95436 260688
rect 109552 260636 109604 260688
rect 189224 260636 189276 260688
rect 203852 260636 203904 260688
rect 80112 260160 80164 260212
rect 85172 260160 85224 260212
rect 80204 260092 80256 260144
rect 85080 260092 85132 260144
rect 172848 260092 172900 260144
rect 179012 260092 179064 260144
rect 173584 260024 173636 260076
rect 179104 260024 179156 260076
rect 229980 260024 230032 260076
rect 233476 260024 233528 260076
rect 175332 259999 175384 260008
rect 175332 259965 175341 259999
rect 175341 259965 175375 259999
rect 175375 259965 175384 259999
rect 175332 259956 175384 259965
rect 173400 259344 173452 259396
rect 175700 259344 175752 259396
rect 80204 258664 80256 258716
rect 84436 258664 84488 258716
rect 173584 258664 173636 258716
rect 178920 258664 178972 258716
rect 79836 258596 79888 258648
rect 82412 258596 82464 258648
rect 88484 258528 88536 258580
rect 129516 258528 129568 258580
rect 182324 258528 182376 258580
rect 223540 258528 223592 258580
rect 173308 257984 173360 258036
rect 175608 257984 175660 258036
rect 229428 257712 229480 257764
rect 233568 257712 233620 257764
rect 80020 257644 80072 257696
rect 82320 257644 82372 257696
rect 229520 257508 229572 257560
rect 233476 257508 233528 257560
rect 173584 257304 173636 257356
rect 175516 257304 175568 257356
rect 80204 257236 80256 257288
rect 81676 257236 81728 257288
rect 131356 257236 131408 257288
rect 132736 257236 132788 257288
rect 134208 257236 134260 257288
rect 229612 257236 229664 257288
rect 233476 257236 233528 257288
rect 82412 257168 82464 257220
rect 87196 257168 87248 257220
rect 131540 257168 131592 257220
rect 140556 257168 140608 257220
rect 179012 257168 179064 257220
rect 182324 257168 182376 257220
rect 226208 257168 226260 257220
rect 234304 257168 234356 257220
rect 131356 257100 131408 257152
rect 140280 257100 140332 257152
rect 179104 257100 179156 257152
rect 182232 257100 182284 257152
rect 226300 257100 226352 257152
rect 234672 257100 234724 257152
rect 131448 257032 131500 257084
rect 140372 257032 140424 257084
rect 175700 257032 175752 257084
rect 182048 257032 182100 257084
rect 225380 257032 225432 257084
rect 234120 257032 234172 257084
rect 85172 256964 85224 257016
rect 87288 256964 87340 257016
rect 85080 256760 85132 256812
rect 87564 256760 87616 256812
rect 173124 256420 173176 256472
rect 175792 256420 175844 256472
rect 173308 256080 173360 256132
rect 175700 256080 175752 256132
rect 80112 255944 80164 255996
rect 82136 255944 82188 255996
rect 80204 255876 80256 255928
rect 81768 255876 81820 255928
rect 230164 255876 230216 255928
rect 233476 255876 233528 255928
rect 82320 255808 82372 255860
rect 87196 255808 87248 255860
rect 131540 255808 131592 255860
rect 139820 255808 139872 255860
rect 175608 255808 175660 255860
rect 181864 255808 181916 255860
rect 225564 255808 225616 255860
rect 234764 255808 234816 255860
rect 81676 255740 81728 255792
rect 87288 255740 87340 255792
rect 131632 255740 131684 255792
rect 139636 255740 139688 255792
rect 175516 255740 175568 255792
rect 182232 255740 182284 255792
rect 226392 255740 226444 255792
rect 233844 255740 233896 255792
rect 84436 255672 84488 255724
rect 87380 255672 87432 255724
rect 131448 255672 131500 255724
rect 139912 255672 139964 255724
rect 178920 255672 178972 255724
rect 182324 255672 182376 255724
rect 226300 255672 226352 255724
rect 229980 255672 230032 255724
rect 131356 255604 131408 255656
rect 140096 255604 140148 255656
rect 225932 255604 225984 255656
rect 229428 255604 229480 255656
rect 80112 254584 80164 254636
rect 80204 254448 80256 254500
rect 84988 254448 85040 254500
rect 173216 254516 173268 254568
rect 173492 254448 173544 254500
rect 87380 254380 87432 254432
rect 131540 254380 131592 254432
rect 139728 254380 139780 254432
rect 81768 254312 81820 254364
rect 87288 254312 87340 254364
rect 131356 254312 131408 254364
rect 140004 254312 140056 254364
rect 182048 254380 182100 254432
rect 225932 254380 225984 254432
rect 230164 254380 230216 254432
rect 182140 254312 182192 254364
rect 131448 254244 131500 254296
rect 139636 254244 139688 254296
rect 175792 254244 175844 254296
rect 182232 254244 182284 254296
rect 82136 254176 82188 254228
rect 87196 254176 87248 254228
rect 175700 254176 175752 254228
rect 182324 254176 182376 254228
rect 226300 254108 226352 254160
rect 229520 254108 229572 254160
rect 226300 253972 226352 254024
rect 229612 253972 229664 254024
rect 84988 253768 85040 253820
rect 87196 253768 87248 253820
rect 80112 253224 80164 253276
rect 80204 253088 80256 253140
rect 173216 253156 173268 253208
rect 173492 253088 173544 253140
rect 87196 253020 87248 253072
rect 131448 253020 131500 253072
rect 139820 253020 139872 253072
rect 87288 252952 87340 253004
rect 131540 252952 131592 253004
rect 139636 252952 139688 253004
rect 230624 253088 230676 253140
rect 233660 253088 233712 253140
rect 182324 253020 182376 253072
rect 226300 253020 226352 253072
rect 233936 253020 233988 253072
rect 181404 252952 181456 253004
rect 226392 252952 226444 253004
rect 233568 252952 233620 253004
rect 131356 252884 131408 252936
rect 139912 252884 139964 252936
rect 226300 252884 226352 252936
rect 233752 252884 233804 252936
rect 225656 252816 225708 252868
rect 233476 252816 233528 252868
rect 80204 252340 80256 252392
rect 87196 252340 87248 252392
rect 131356 252340 131408 252392
rect 140556 252340 140608 252392
rect 173584 252340 173636 252392
rect 182324 252340 182376 252392
rect 80204 251728 80256 251780
rect 173492 251728 173544 251780
rect 131356 251660 131408 251712
rect 140188 251660 140240 251712
rect 181772 251660 181824 251712
rect 225380 251660 225432 251712
rect 233568 251660 233620 251712
rect 87196 251592 87248 251644
rect 226392 251592 226444 251644
rect 233476 251592 233528 251644
rect 226300 251524 226352 251576
rect 230624 251524 230676 251576
rect 80204 251048 80256 251100
rect 87196 251048 87248 251100
rect 131356 251048 131408 251100
rect 140648 251048 140700 251100
rect 173492 251048 173544 251100
rect 182324 251048 182376 251100
rect 80112 250980 80164 251032
rect 87288 250980 87340 251032
rect 131448 250980 131500 251032
rect 140556 250980 140608 251032
rect 173584 250980 173636 251032
rect 182232 250980 182284 251032
rect 175424 250300 175476 250352
rect 131356 250232 131408 250284
rect 140556 250232 140608 250284
rect 226300 250232 226352 250284
rect 233568 250232 233620 250284
rect 225932 250164 225984 250216
rect 233476 250164 233528 250216
rect 80112 249620 80164 249672
rect 87196 249620 87248 249672
rect 131816 249620 131868 249672
rect 140464 249620 140516 249672
rect 173584 249620 173636 249672
rect 182324 249620 182376 249672
rect 225564 249620 225616 249672
rect 233568 249620 233620 249672
rect 80204 249552 80256 249604
rect 87288 249552 87340 249604
rect 131356 249552 131408 249604
rect 140004 249552 140056 249604
rect 173676 249552 173728 249604
rect 182232 249552 182284 249604
rect 226300 249552 226352 249604
rect 233476 249552 233528 249604
rect 131356 248940 131408 248992
rect 79284 248872 79336 248924
rect 87196 248872 87248 248924
rect 140372 248872 140424 248924
rect 173216 248872 173268 248924
rect 181588 248872 181640 248924
rect 80204 248804 80256 248856
rect 87380 248804 87432 248856
rect 173584 248804 173636 248856
rect 182324 248804 182376 248856
rect 226300 248260 226352 248312
rect 233568 248260 233620 248312
rect 131356 248192 131408 248244
rect 140372 248192 140424 248244
rect 226392 248192 226444 248244
rect 233476 248192 233528 248244
rect 85908 247716 85960 247768
rect 88024 247716 88076 247768
rect 131816 247716 131868 247768
rect 137060 247716 137112 247768
rect 132552 247648 132604 247700
rect 137520 247648 137572 247700
rect 226300 247648 226352 247700
rect 234396 247648 234448 247700
rect 86092 247580 86144 247632
rect 87196 247580 87248 247632
rect 131448 247580 131500 247632
rect 79284 247512 79336 247564
rect 88392 247512 88444 247564
rect 226392 247580 226444 247632
rect 234488 247580 234540 247632
rect 140372 247512 140424 247564
rect 173216 247512 173268 247564
rect 181128 247512 181180 247564
rect 80204 247444 80256 247496
rect 88300 247444 88352 247496
rect 173584 247444 173636 247496
rect 181036 247444 181088 247496
rect 137520 247240 137572 247292
rect 140648 247240 140700 247292
rect 80020 246356 80072 246408
rect 87196 246356 87248 246408
rect 131448 246356 131500 246408
rect 137244 246356 137296 246408
rect 173952 246356 174004 246408
rect 182324 246356 182376 246408
rect 226300 246356 226352 246408
rect 233660 246356 233712 246408
rect 132184 246288 132236 246340
rect 140648 246288 140700 246340
rect 226392 246288 226444 246340
rect 233568 246288 233620 246340
rect 131356 246220 131408 246272
rect 140188 246220 140240 246272
rect 225656 246220 225708 246272
rect 233476 246220 233528 246272
rect 79284 246152 79336 246204
rect 86092 246152 86144 246204
rect 137060 246084 137112 246136
rect 140556 246084 140608 246136
rect 173584 246084 173636 246136
rect 180852 246084 180904 246136
rect 137244 245948 137296 246000
rect 140372 245948 140424 246000
rect 80204 245880 80256 245932
rect 85908 245880 85960 245932
rect 173492 245676 173544 245728
rect 180944 245676 180996 245728
rect 225564 245200 225616 245252
rect 227956 245200 228008 245252
rect 131816 244996 131868 245048
rect 135956 244996 136008 245048
rect 131356 244928 131408 244980
rect 135864 244928 135916 244980
rect 226208 244928 226260 244980
rect 228048 244928 228100 244980
rect 132000 244860 132052 244912
rect 139636 244860 139688 244912
rect 226392 244860 226444 244912
rect 228140 244860 228192 244912
rect 131448 244792 131500 244844
rect 139728 244792 139780 244844
rect 226300 244792 226352 244844
rect 233476 244792 233528 244844
rect 80112 244724 80164 244776
rect 87104 244724 87156 244776
rect 173584 244724 173636 244776
rect 180760 244724 180812 244776
rect 80204 244656 80256 244708
rect 87012 244656 87064 244708
rect 172848 244656 172900 244708
rect 180668 244656 180720 244708
rect 131356 243636 131408 243688
rect 136784 243636 136836 243688
rect 131448 243568 131500 243620
rect 136692 243568 136744 243620
rect 175424 243568 175476 243620
rect 225748 243568 225800 243620
rect 233660 243568 233712 243620
rect 79928 243500 79980 243552
rect 87196 243500 87248 243552
rect 131540 243500 131592 243552
rect 139360 243500 139412 243552
rect 173860 243500 173912 243552
rect 181220 243500 181272 243552
rect 226208 243500 226260 243552
rect 233844 243500 233896 243552
rect 80112 243432 80164 243484
rect 87288 243432 87340 243484
rect 131632 243432 131684 243484
rect 139544 243432 139596 243484
rect 173492 243432 173544 243484
rect 182324 243432 182376 243484
rect 226300 243432 226352 243484
rect 233752 243432 233804 243484
rect 80204 243364 80256 243416
rect 86920 243364 86972 243416
rect 175332 243407 175384 243416
rect 175332 243373 175341 243407
rect 175341 243373 175375 243407
rect 175375 243373 175384 243407
rect 175332 243364 175384 243373
rect 228048 243364 228100 243416
rect 233476 243364 233528 243416
rect 227956 243296 228008 243348
rect 233568 243296 233620 243348
rect 173584 243160 173636 243212
rect 180852 243160 180904 243212
rect 80204 242752 80256 242804
rect 86828 242752 86880 242804
rect 172848 242752 172900 242804
rect 180944 242752 180996 242804
rect 79284 242208 79336 242260
rect 87196 242208 87248 242260
rect 131356 242208 131408 242260
rect 136140 242208 136192 242260
rect 173768 242208 173820 242260
rect 182324 242208 182376 242260
rect 226024 242208 226076 242260
rect 228692 242208 228744 242260
rect 131448 242140 131500 242192
rect 136232 242140 136284 242192
rect 226300 242140 226352 242192
rect 131540 242072 131592 242124
rect 139452 242072 139504 242124
rect 226392 242072 226444 242124
rect 228600 242072 228652 242124
rect 233568 242072 233620 242124
rect 79100 242004 79152 242056
rect 87564 242004 87616 242056
rect 135864 242004 135916 242056
rect 140556 242004 140608 242056
rect 173584 242004 173636 242056
rect 182232 242004 182284 242056
rect 228140 242004 228192 242056
rect 233476 242004 233528 242056
rect 264756 242004 264808 242056
rect 300176 242004 300228 242056
rect 80204 241936 80256 241988
rect 87656 241936 87708 241988
rect 135956 241936 136008 241988
rect 140188 241936 140240 241988
rect 173676 241936 173728 241988
rect 182048 241936 182100 241988
rect 178920 240712 178972 240764
rect 181588 240712 181640 240764
rect 85080 240644 85132 240696
rect 87380 240644 87432 240696
rect 131356 240644 131408 240696
rect 139268 240644 139320 240696
rect 226024 240644 226076 240696
rect 234120 240644 234172 240696
rect 109920 240440 109972 240492
rect 141016 240440 141068 240492
rect 203116 239760 203168 239812
rect 203852 239760 203904 239812
rect 80204 239216 80256 239268
rect 87472 239216 87524 239268
rect 136784 239216 136836 239268
rect 140556 239216 140608 239268
rect 173676 239216 173728 239268
rect 182140 239216 182192 239268
rect 226576 239216 226628 239268
rect 233476 239216 233528 239268
rect 136692 239148 136744 239200
rect 140648 239148 140700 239200
rect 80204 237856 80256 237908
rect 86552 237856 86604 237908
rect 228692 237856 228744 237908
rect 233476 237856 233528 237908
rect 136232 237788 136284 237840
rect 140556 237788 140608 237840
rect 228600 237788 228652 237840
rect 233568 237788 233620 237840
rect 136140 237516 136192 237568
rect 140280 237516 140332 237568
rect 173584 237380 173636 237432
rect 180392 237380 180444 237432
rect 80204 237312 80256 237364
rect 86460 237312 86512 237364
rect 173400 236904 173452 236956
rect 180300 236904 180352 236956
rect 173584 236496 173636 236548
rect 178920 236496 178972 236548
rect 80204 235272 80256 235324
rect 85080 235272 85132 235324
rect 151780 233708 151832 233760
rect 163188 233708 163240 233760
rect 249116 233708 249168 233760
rect 259236 233708 259288 233760
rect 60884 233640 60936 233692
rect 60148 233572 60200 233624
rect 154908 233640 154960 233692
rect 167880 233640 167932 233692
rect 249300 233640 249352 233692
rect 57940 233504 57992 233556
rect 66220 233504 66272 233556
rect 60608 233436 60660 233488
rect 71648 233572 71700 233624
rect 154632 233572 154684 233624
rect 247736 233572 247788 233624
rect 259788 233640 259840 233692
rect 138164 233504 138216 233556
rect 142856 233504 142908 233556
rect 153160 233504 153212 233556
rect 72384 233436 72436 233488
rect 137980 233436 138032 233488
rect 143960 233436 144012 233488
rect 61252 233368 61304 233420
rect 74408 233368 74460 233420
rect 137888 233368 137940 233420
rect 144604 233368 144656 233420
rect 153252 233368 153304 233420
rect 159508 233504 159560 233556
rect 162084 233504 162136 233556
rect 248656 233504 248708 233556
rect 255832 233504 255884 233556
rect 261996 233504 262048 233556
rect 166684 233436 166736 233488
rect 248932 233436 248984 233488
rect 261444 233436 261496 233488
rect 57664 233232 57716 233284
rect 65484 233232 65536 233284
rect 154540 233300 154592 233352
rect 156104 233300 156156 233352
rect 73028 233232 73080 233284
rect 138072 233232 138124 233284
rect 143776 233232 143828 233284
rect 153712 233232 153764 233284
rect 164936 233368 164988 233420
rect 249024 233368 249076 233420
rect 255556 233368 255608 233420
rect 166132 233300 166184 233352
rect 165948 233232 166000 233284
rect 247000 233232 247052 233284
rect 249576 233232 249628 233284
rect 61712 233164 61764 233216
rect 62080 233164 62132 233216
rect 62264 233164 62316 233216
rect 75788 233164 75840 233216
rect 137796 233164 137848 233216
rect 145156 233164 145208 233216
rect 151596 233164 151648 233216
rect 156196 233164 156248 233216
rect 53248 233096 53300 233148
rect 62356 233096 62408 233148
rect 62448 233096 62500 233148
rect 76432 233096 76484 233148
rect 155276 233096 155328 233148
rect 168616 233164 168668 233216
rect 231820 233164 231872 233216
rect 239180 233164 239232 233216
rect 245344 233164 245396 233216
rect 249392 233164 249444 233216
rect 249484 233164 249536 233216
rect 256384 233232 256436 233284
rect 258960 233232 259012 233284
rect 250312 233164 250364 233216
rect 263100 233164 263152 233216
rect 38160 233028 38212 233080
rect 49200 233028 49252 233080
rect 62080 233028 62132 233080
rect 75052 233028 75104 233080
rect 137612 233028 137664 233080
rect 145708 233028 145760 233080
rect 150492 233028 150544 233080
rect 154816 233028 154868 233080
rect 167328 233096 167380 233148
rect 248472 233096 248524 233148
rect 261076 233096 261128 233148
rect 56008 232960 56060 233012
rect 66036 232960 66088 233012
rect 154724 232960 154776 233012
rect 161808 233028 161860 233080
rect 231728 233028 231780 233080
rect 239640 233028 239692 233080
rect 245804 233028 245856 233080
rect 249668 233028 249720 233080
rect 249852 233028 249904 233080
rect 262548 233028 262600 233080
rect 63644 232892 63696 232944
rect 152792 232892 152844 232944
rect 155184 232892 155236 232944
rect 56652 232824 56704 232876
rect 66404 232824 66456 232876
rect 150584 232824 150636 232876
rect 242492 232960 242544 233012
rect 247644 232960 247696 233012
rect 258316 232960 258368 233012
rect 158036 232892 158088 232944
rect 161164 232892 161216 232944
rect 243596 232892 243648 232944
rect 248288 232892 248340 232944
rect 256936 232892 256988 232944
rect 159784 232824 159836 232876
rect 162636 232824 162688 232876
rect 244148 232824 244200 232876
rect 247552 232824 247604 232876
rect 59320 232756 59372 232808
rect 58032 232688 58084 232740
rect 61344 232688 61396 232740
rect 61528 232688 61580 232740
rect 68244 232688 68296 232740
rect 60792 232620 60844 232672
rect 61620 232620 61672 232672
rect 67600 232620 67652 232672
rect 149848 232756 149900 232808
rect 151872 232756 151924 232808
rect 151964 232756 152016 232808
rect 156288 232756 156340 232808
rect 156840 232756 156892 232808
rect 160060 232756 160112 232808
rect 246724 232756 246776 232808
rect 248012 232756 248064 232808
rect 254176 232824 254228 232876
rect 248564 232756 248616 232808
rect 254728 232756 254780 232808
rect 153344 232688 153396 232740
rect 158220 232688 158272 232740
rect 158588 232688 158640 232740
rect 160980 232688 161032 232740
rect 169076 232688 169128 232740
rect 247184 232688 247236 232740
rect 258684 232688 258736 232740
rect 71004 232620 71056 232672
rect 153988 232620 154040 232672
rect 155000 232620 155052 232672
rect 155092 232620 155144 232672
rect 158312 232620 158364 232672
rect 159048 232620 159100 232672
rect 161072 232620 161124 232672
rect 231636 232620 231688 232672
rect 238536 232620 238588 232672
rect 244424 232620 244476 232672
rect 247368 232620 247420 232672
rect 248104 232620 248156 232672
rect 249944 232620 249996 232672
rect 252060 232620 252112 232672
rect 257028 232620 257080 232672
rect 57296 232552 57348 232604
rect 61436 232552 61488 232604
rect 61804 232552 61856 232604
rect 63460 232552 63512 232604
rect 67968 232552 68020 232604
rect 70268 232552 70320 232604
rect 157484 232552 157536 232604
rect 159876 232552 159928 232604
rect 231544 232552 231596 232604
rect 237984 232552 238036 232604
rect 245804 232552 245856 232604
rect 253072 232552 253124 232604
rect 62172 232484 62224 232536
rect 66864 232484 66916 232536
rect 67876 232484 67928 232536
rect 69624 232484 69676 232536
rect 151044 232484 151096 232536
rect 153436 232484 153488 232536
rect 156380 232484 156432 232536
rect 159140 232484 159192 232536
rect 231452 232484 231504 232536
rect 237616 232484 237668 232536
rect 243044 232484 243096 232536
rect 247000 232484 247052 232536
rect 248196 232484 248248 232536
rect 260340 232484 260392 232536
rect 60056 232416 60108 232468
rect 61160 232416 61212 232468
rect 61988 232416 62040 232468
rect 68980 232416 69032 232468
rect 158404 232416 158456 232468
rect 159692 232416 159744 232468
rect 162360 232416 162412 232468
rect 163832 232416 163884 232468
rect 231360 232416 231412 232468
rect 236880 232416 236932 232468
rect 241572 232416 241624 232468
rect 245436 232416 245488 232468
rect 246448 232416 246500 232468
rect 251416 232416 251468 232468
rect 256200 232416 256252 232468
rect 257488 232416 257540 232468
rect 155736 231464 155788 231516
rect 126480 229628 126532 229680
rect 159600 229628 159652 229680
rect 220504 229628 220556 229680
rect 254728 229628 254780 229680
rect 137704 228200 137756 228252
rect 146812 228200 146864 228252
rect 232004 228200 232056 228252
rect 240744 228200 240796 228252
rect 156104 226840 156156 226892
rect 56192 225412 56244 225464
rect 57664 225412 57716 225464
rect 58676 225412 58728 225464
rect 59504 225412 59556 225464
rect 231912 225480 231964 225532
rect 234120 225480 234172 225532
rect 55272 225344 55324 225396
rect 51868 225276 51920 225328
rect 64288 225412 64340 225464
rect 151412 225412 151464 225464
rect 159692 225412 159744 225464
rect 161164 225412 161216 225464
rect 163556 225412 163608 225464
rect 244424 225412 244476 225464
rect 248564 225412 248616 225464
rect 250036 225412 250088 225464
rect 254728 225412 254780 225464
rect 258684 225412 258736 225464
rect 64012 225344 64064 225396
rect 149848 225344 149900 225396
rect 160336 225344 160388 225396
rect 160980 225344 161032 225396
rect 163924 225344 163976 225396
rect 244056 225344 244108 225396
rect 248012 225344 248064 225396
rect 248288 225344 248340 225396
rect 252060 225344 252112 225396
rect 252704 225344 252756 225396
rect 258316 225344 258368 225396
rect 65944 225276 65996 225328
rect 156196 225276 156248 225328
rect 159232 225276 159284 225328
rect 159784 225276 159836 225328
rect 163096 225276 163148 225328
rect 175332 225276 175384 225328
rect 281868 225276 281920 225328
rect 55824 225208 55876 225260
rect 59688 225208 59740 225260
rect 60976 225208 61028 225260
rect 54628 225140 54680 225192
rect 52512 225072 52564 225124
rect 56560 225140 56612 225192
rect 57940 225140 57992 225192
rect 58124 225140 58176 225192
rect 61988 225140 62040 225192
rect 62816 225208 62868 225260
rect 70268 225208 70320 225260
rect 154816 225208 154868 225260
rect 158404 225208 158456 225260
rect 245436 225208 245488 225260
rect 250864 225208 250916 225260
rect 251324 225208 251376 225260
rect 67876 225140 67928 225192
rect 150216 225140 150268 225192
rect 160428 225140 160480 225192
rect 247000 225140 247052 225192
rect 251692 225140 251744 225192
rect 257580 225140 257632 225192
rect 51224 225004 51276 225056
rect 51132 224868 51184 224920
rect 29144 224800 29196 224852
rect 31628 224800 31680 224852
rect 49844 224732 49896 224784
rect 59412 225072 59464 225124
rect 58584 224936 58636 224988
rect 61896 225072 61948 225124
rect 69532 225072 69584 225124
rect 148652 225072 148704 225124
rect 157300 225072 157352 225124
rect 157668 225072 157720 225124
rect 63644 225004 63696 225056
rect 69072 225004 69124 225056
rect 149480 225004 149532 225056
rect 158588 225004 158640 225056
rect 159600 225072 159652 225124
rect 164660 225072 164712 225124
rect 247644 225072 247696 225124
rect 251324 225072 251376 225124
rect 251416 225072 251468 225124
rect 253992 225072 254044 225124
rect 160888 225004 160940 225056
rect 161072 225004 161124 225056
rect 164292 225004 164344 225056
rect 245620 225004 245672 225056
rect 249484 225004 249536 225056
rect 251048 225004 251100 225056
rect 68336 224936 68388 224988
rect 156288 224936 156340 224988
rect 159600 224936 159652 224988
rect 159876 224936 159928 224988
rect 162728 224936 162780 224988
rect 243320 224936 243372 224988
rect 253164 224936 253216 224988
rect 257120 224936 257172 224988
rect 61160 224868 61212 224920
rect 61712 224868 61764 224920
rect 69900 224868 69952 224920
rect 151044 224868 151096 224920
rect 159508 224868 159560 224920
rect 243688 224868 243740 224920
rect 253624 224868 253676 224920
rect 256752 224868 256804 224920
rect 64380 224800 64432 224852
rect 152608 224800 152660 224852
rect 164568 224800 164620 224852
rect 247552 224800 247604 224852
rect 252428 224800 252480 224852
rect 256016 224800 256068 224852
rect 63368 224732 63420 224784
rect 149112 224732 149164 224784
rect 156380 224732 156432 224784
rect 156472 224732 156524 224784
rect 170180 224732 170232 224784
rect 247276 224732 247328 224784
rect 250680 224732 250732 224784
rect 263836 224732 263888 224784
rect 267240 224732 267292 224784
rect 289872 224732 289924 224784
rect 57296 224664 57348 224716
rect 62172 224664 62224 224716
rect 62356 224664 62408 224716
rect 64840 224664 64892 224716
rect 149204 224664 149256 224716
rect 247552 224664 247604 224716
rect 249116 224664 249168 224716
rect 249208 224664 249260 224716
rect 53984 224596 54036 224648
rect 65208 224596 65260 224648
rect 147824 224596 147876 224648
rect 156840 224596 156892 224648
rect 158220 224596 158272 224648
rect 160428 224596 160480 224648
rect 244884 224596 244936 224648
rect 249024 224596 249076 224648
rect 249760 224596 249812 224648
rect 256384 224664 256436 224716
rect 57756 224528 57808 224580
rect 61528 224528 61580 224580
rect 68704 224528 68756 224580
rect 158312 224528 158364 224580
rect 161532 224528 161584 224580
rect 245252 224528 245304 224580
rect 248656 224528 248708 224580
rect 249668 224528 249720 224580
rect 253624 224528 253676 224580
rect 254452 224528 254504 224580
rect 57388 224460 57440 224512
rect 61620 224460 61672 224512
rect 61712 224460 61764 224512
rect 67140 224460 67192 224512
rect 151872 224460 151924 224512
rect 158036 224460 158088 224512
rect 249392 224460 249444 224512
rect 253256 224460 253308 224512
rect 62816 224392 62868 224444
rect 62908 224392 62960 224444
rect 67968 224392 68020 224444
rect 155184 224392 155236 224444
rect 159968 224392 160020 224444
rect 246448 224392 246500 224444
rect 256200 224392 256252 224444
rect 55088 224324 55140 224376
rect 55732 224256 55784 224308
rect 65576 224324 65628 224376
rect 153436 224324 153488 224376
rect 158864 224324 158916 224376
rect 249944 224324 249996 224376
rect 255188 224324 255240 224376
rect 61804 224256 61856 224308
rect 61896 224256 61948 224308
rect 67508 224256 67560 224308
rect 152148 224256 152200 224308
rect 162268 224256 162320 224308
rect 249576 224256 249628 224308
rect 254820 224256 254872 224308
rect 58952 224188 59004 224240
rect 61160 224188 61212 224240
rect 38252 224120 38304 224172
rect 59504 224052 59556 224104
rect 67968 224120 68020 224172
rect 155000 224188 155052 224240
rect 160796 224188 160848 224240
rect 248380 224188 248432 224240
rect 70636 224120 70688 224172
rect 155828 224120 155880 224172
rect 161992 224120 162044 224172
rect 255556 224120 255608 224172
rect 137704 224052 137756 224104
rect 146720 224052 146772 224104
rect 155920 224052 155972 224104
rect 162360 224052 162412 224104
rect 232004 224052 232056 224104
rect 240376 224052 240428 224104
rect 247368 224052 247420 224104
rect 252796 224052 252848 224104
rect 63736 223984 63788 224036
rect 63276 223644 63328 223696
rect 257028 223032 257080 223084
rect 257902 223032 257954 223084
rect 148744 221332 148796 221384
rect 165120 221332 165172 221384
rect 231084 221332 231136 221384
rect 239364 221332 239416 221384
rect 12952 219972 13004 220024
rect 18840 219972 18892 220024
rect 230992 218816 231044 218868
rect 232740 218816 232792 218868
rect 231728 218680 231780 218732
rect 240928 218680 240980 218732
rect 137428 218612 137480 218664
rect 145616 218612 145668 218664
rect 292816 217116 292868 217168
rect 300176 217116 300228 217168
rect 232004 215960 232056 216012
rect 238260 215960 238312 216012
rect 137336 215824 137388 215876
rect 145616 215824 145668 215876
rect 231820 215824 231872 215876
rect 240468 215824 240520 215876
rect 165120 215756 165172 215808
rect 175516 215756 175568 215808
rect 137152 213104 137204 213156
rect 145616 213104 145668 213156
rect 231912 213104 231964 213156
rect 240928 213104 240980 213156
rect 262364 212832 262416 212884
rect 265216 212832 265268 212884
rect 232004 212288 232056 212340
rect 236880 212288 236932 212340
rect 137244 211676 137296 211728
rect 145616 211676 145668 211728
rect 231636 211676 231688 211728
rect 240928 211676 240980 211728
rect 232004 209228 232056 209280
rect 235500 209228 235552 209280
rect 137060 208956 137112 209008
rect 145616 208956 145668 209008
rect 231544 208956 231596 209008
rect 240468 208956 240520 209008
rect 258960 208888 259012 208940
rect 274876 208888 274928 208940
rect 232004 206440 232056 206492
rect 234212 206440 234264 206492
rect 232004 206168 232056 206220
rect 240652 206168 240704 206220
rect 136968 204808 137020 204860
rect 145616 204808 145668 204860
rect 231452 204808 231504 204860
rect 240928 204808 240980 204860
rect 143040 202020 143092 202072
rect 145524 202020 145576 202072
rect 231268 202020 231320 202072
rect 240376 202020 240428 202072
rect 231728 199300 231780 199352
rect 240468 199300 240520 199352
rect 140280 197872 140332 197924
rect 145616 197872 145668 197924
rect 231820 197872 231872 197924
rect 240928 197872 240980 197924
rect 263744 196512 263796 196564
rect 274876 196512 274928 196564
rect 140372 195152 140424 195204
rect 145616 195152 145668 195204
rect 234304 195152 234356 195204
rect 240928 195152 240980 195204
rect 137428 195084 137480 195136
rect 145800 195084 145852 195136
rect 236972 192432 237024 192484
rect 240468 192432 240520 192484
rect 143132 192364 143184 192416
rect 145800 192364 145852 192416
rect 167880 192364 167932 192416
rect 175516 192364 175568 192416
rect 262364 192364 262416 192416
rect 275520 192364 275572 192416
rect 137428 191072 137480 191124
rect 143040 191072 143092 191124
rect 74040 190936 74092 190988
rect 81676 190936 81728 190988
rect 137060 189644 137112 189696
rect 145156 189644 145208 189696
rect 230808 189644 230860 189696
rect 240652 189644 240704 189696
rect 137428 189372 137480 189424
rect 144420 189372 144472 189424
rect 292816 188896 292868 188948
rect 293552 188896 293604 188948
rect 47084 188216 47136 188268
rect 51316 188216 51368 188268
rect 137336 188216 137388 188268
rect 145616 188216 145668 188268
rect 231268 188216 231320 188268
rect 240744 188216 240796 188268
rect 137428 188148 137480 188200
rect 140280 188148 140332 188200
rect 38804 186788 38856 186840
rect 47084 186788 47136 186840
rect 137428 186788 137480 186840
rect 140372 186788 140424 186840
rect 231820 186788 231872 186840
rect 234304 186788 234356 186840
rect 237616 185496 237668 185548
rect 240928 185496 240980 185548
rect 231820 185428 231872 185480
rect 236972 185428 237024 185480
rect 137428 184204 137480 184256
rect 143132 184204 143184 184256
rect 63828 181348 63880 181400
rect 18840 181280 18892 181332
rect 23716 181280 23768 181332
rect 31628 181280 31680 181332
rect 55824 181280 55876 181332
rect 63736 181280 63788 181332
rect 150676 181280 150728 181332
rect 151688 181280 151740 181332
rect 153068 181280 153120 181332
rect 156288 181280 156340 181332
rect 157484 181280 157536 181332
rect 158404 181280 158456 181332
rect 244424 181280 244476 181332
rect 245436 181280 245488 181332
rect 62080 181212 62132 181264
rect 69808 181212 69860 181264
rect 149204 181212 149256 181264
rect 160704 181212 160756 181264
rect 243320 181212 243372 181264
rect 245160 181212 245212 181264
rect 245712 181212 245764 181264
rect 249576 181280 249628 181332
rect 249944 181280 249996 181332
rect 250496 181348 250548 181400
rect 253440 181280 253492 181332
rect 253624 181280 253676 181332
rect 255188 181280 255240 181332
rect 249300 181212 249352 181264
rect 250772 181212 250824 181264
rect 250864 181212 250916 181264
rect 253716 181212 253768 181264
rect 59872 181144 59924 181196
rect 69900 181144 69952 181196
rect 145156 181144 145208 181196
rect 157208 181144 157260 181196
rect 243044 181144 243096 181196
rect 251416 181144 251468 181196
rect 20220 181076 20272 181128
rect 59044 181076 59096 181128
rect 69348 181076 69400 181128
rect 152240 181076 152292 181128
rect 245712 181076 245764 181128
rect 248932 181076 248984 181128
rect 250680 181076 250732 181128
rect 251324 181076 251376 181128
rect 257212 181076 257264 181128
rect 55456 181008 55508 181060
rect 69256 181008 69308 181060
rect 147732 181008 147784 181060
rect 159508 181008 159560 181060
rect 245344 181008 245396 181060
rect 249760 181008 249812 181060
rect 252428 181008 252480 181060
rect 53984 180940 54036 180992
rect 65484 180940 65536 180992
rect 147824 180940 147876 180992
rect 160244 180940 160296 180992
rect 242952 180940 243004 180992
rect 251600 180940 251652 180992
rect 58676 180872 58728 180924
rect 67048 180872 67100 180924
rect 149480 180872 149532 180924
rect 153160 180872 153212 180924
rect 153252 180872 153304 180924
rect 231636 180872 231688 180924
rect 237616 180872 237668 180924
rect 242860 180872 242912 180924
rect 251968 180872 252020 180924
rect 252060 180872 252112 180924
rect 254820 180872 254872 180924
rect 56652 180804 56704 180856
rect 65116 180804 65168 180856
rect 147640 180804 147692 180856
rect 159876 180804 159928 180856
rect 244884 180804 244936 180856
rect 254176 180804 254228 180856
rect 63460 180736 63512 180788
rect 146444 180736 146496 180788
rect 159048 180736 159100 180788
rect 163096 180736 163148 180788
rect 247184 180736 247236 180788
rect 251140 180736 251192 180788
rect 257580 180736 257632 180788
rect 49844 180668 49896 180720
rect 51132 180600 51184 180652
rect 58216 180668 58268 180720
rect 63552 180668 63604 180720
rect 70636 180668 70688 180720
rect 144880 180668 144932 180720
rect 158312 180668 158364 180720
rect 246908 180668 246960 180720
rect 56284 180600 56336 180652
rect 65208 180600 65260 180652
rect 144972 180600 145024 180652
rect 157852 180600 157904 180652
rect 158220 180600 158272 180652
rect 164660 180600 164712 180652
rect 242400 180600 242452 180652
rect 251048 180600 251100 180652
rect 63092 180532 63144 180584
rect 65760 180532 65812 180584
rect 153436 180532 153488 180584
rect 163832 180532 163884 180584
rect 245804 180532 245856 180584
rect 253164 180600 253216 180652
rect 261076 180600 261128 180652
rect 251232 180532 251284 180584
rect 258316 180532 258368 180584
rect 52512 180464 52564 180516
rect 64288 180464 64340 180516
rect 150308 180464 150360 180516
rect 152976 180464 153028 180516
rect 155460 180464 155512 180516
rect 156104 180464 156156 180516
rect 162452 180464 162504 180516
rect 243688 180464 243740 180516
rect 245252 180464 245304 180516
rect 246080 180464 246132 180516
rect 249208 180464 249260 180516
rect 249300 180464 249352 180516
rect 252796 180464 252848 180516
rect 52604 180396 52656 180448
rect 64656 180396 64708 180448
rect 151780 180396 151832 180448
rect 162636 180396 162688 180448
rect 247184 180396 247236 180448
rect 254360 180396 254412 180448
rect 57020 180328 57072 180380
rect 60608 180328 60660 180380
rect 63092 180328 63144 180380
rect 68612 180328 68664 180380
rect 146352 180328 146404 180380
rect 70268 180260 70320 180312
rect 152056 180260 152108 180312
rect 153896 180328 153948 180380
rect 163740 180328 163792 180380
rect 249852 180328 249904 180380
rect 256384 180328 256436 180380
rect 158680 180260 158732 180312
rect 253716 180260 253768 180312
rect 55088 180192 55140 180244
rect 60148 180192 60200 180244
rect 60424 180192 60476 180244
rect 66680 180192 66732 180244
rect 157116 180192 157168 180244
rect 162360 180192 162412 180244
rect 247736 180192 247788 180244
rect 249576 180192 249628 180244
rect 253532 180192 253584 180244
rect 60056 180124 60108 180176
rect 63000 180124 63052 180176
rect 68244 180124 68296 180176
rect 149112 180124 149164 180176
rect 152884 180124 152936 180176
rect 57572 180056 57624 180108
rect 65024 180056 65076 180108
rect 149848 180056 149900 180108
rect 152792 180056 152844 180108
rect 57480 179988 57532 180040
rect 60240 179988 60292 180040
rect 63736 179988 63788 180040
rect 64472 179988 64524 180040
rect 69440 179988 69492 180040
rect 137428 179988 137480 180040
rect 144788 179988 144840 180040
rect 151044 179988 151096 180040
rect 156840 180124 156892 180176
rect 248840 180124 248892 180176
rect 163464 180056 163516 180108
rect 244148 180056 244200 180108
rect 245344 180056 245396 180108
rect 246540 180056 246592 180108
rect 248932 180056 248984 180108
rect 153252 179988 153304 180040
rect 157024 179988 157076 180040
rect 164292 179988 164344 180040
rect 248104 179988 248156 180040
rect 249392 179988 249444 180040
rect 57848 179920 57900 179972
rect 61068 179920 61120 179972
rect 61804 179920 61856 179972
rect 61896 179920 61948 179972
rect 62264 179920 62316 179972
rect 62632 179920 62684 179972
rect 63644 179920 63696 179972
rect 60516 179784 60568 179836
rect 62264 179784 62316 179836
rect 64380 179920 64432 179972
rect 69072 179920 69124 179972
rect 143684 179920 143736 179972
rect 153344 179920 153396 179972
rect 137428 179852 137480 179904
rect 145800 179852 145852 179904
rect 163556 179920 163608 179972
rect 248380 179920 248432 179972
rect 249024 179920 249076 179972
rect 257028 180124 257080 180176
rect 250588 180056 250640 180108
rect 250956 180056 251008 180108
rect 252704 180056 252756 180108
rect 258408 180056 258460 180108
rect 256936 179988 256988 180040
rect 257120 179920 257172 179972
rect 231636 179852 231688 179904
rect 239640 179852 239692 179904
rect 88208 177948 88260 178000
rect 86828 177880 86880 177932
rect 87104 177744 87156 177796
rect 90876 177880 90928 177932
rect 88484 177744 88536 177796
rect 91244 177744 91296 177796
rect 249576 176248 249628 176300
rect 249576 176044 249628 176096
rect 85540 175772 85592 175824
rect 179564 175772 179616 175824
rect 188948 175772 189000 175824
rect 198240 175772 198292 175824
rect 228692 175772 228744 175824
rect 261168 175772 261220 175824
rect 94924 175704 94976 175756
rect 104216 175704 104268 175756
rect 132736 175704 132788 175756
rect 226760 175704 226812 175756
rect 115164 175636 115216 175688
rect 173400 175636 173452 175688
rect 203852 175636 203904 175688
rect 211948 175636 212000 175688
rect 79744 175568 79796 175620
rect 109828 175568 109880 175620
rect 111116 175568 111168 175620
rect 140280 175568 140332 175620
rect 173860 175568 173912 175620
rect 206520 175568 206572 175620
rect 228140 175568 228192 175620
rect 228692 175568 228744 175620
rect 79560 175500 79612 175552
rect 112496 175500 112548 175552
rect 173676 175500 173728 175552
rect 209188 175500 209240 175552
rect 213236 175500 213288 175552
rect 51224 175432 51276 175484
rect 65576 175432 65628 175484
rect 65852 175432 65904 175484
rect 79652 175432 79704 175484
rect 152700 175432 152752 175484
rect 152976 175432 153028 175484
rect 173492 175432 173544 175484
rect 232832 175432 232884 175484
rect 79836 175364 79888 175416
rect 117924 175364 117976 175416
rect 173768 175364 173820 175416
rect 214616 175364 214668 175416
rect 215996 175364 216048 175416
rect 224460 175364 224512 175416
rect 79928 175296 79980 175348
rect 123260 175296 123312 175348
rect 173584 175296 173636 175348
rect 217284 175296 217336 175348
rect 80204 175228 80256 175280
rect 126020 175228 126072 175280
rect 176160 175228 176212 175280
rect 220044 175228 220096 175280
rect 221332 175228 221384 175280
rect 264848 175228 264900 175280
rect 80020 175160 80072 175212
rect 128688 175160 128740 175212
rect 174780 175160 174832 175212
rect 222712 175160 222764 175212
rect 65116 175092 65168 175144
rect 65852 175092 65904 175144
rect 80112 175092 80164 175144
rect 120592 175092 120644 175144
rect 121972 175092 122024 175144
rect 170640 175092 170692 175144
rect 190328 175092 190380 175144
rect 199620 175092 199672 175144
rect 202472 175092 202524 175144
rect 264756 175092 264808 175144
rect 92256 175024 92308 175076
rect 97500 175024 97552 175076
rect 93636 174956 93688 175008
rect 98880 174956 98932 175008
rect 89588 174888 89640 174940
rect 95476 174888 95528 174940
rect 96304 174820 96356 174872
rect 105688 175024 105740 175076
rect 256936 175024 256988 175076
rect 257580 175024 257632 175076
rect 186280 174752 186332 174804
rect 191340 174752 191392 174804
rect 187660 174616 187712 174668
rect 192720 174616 192772 174668
rect 97684 174412 97736 174464
rect 98144 174412 98196 174464
rect 98972 174412 99024 174464
rect 99524 174412 99576 174464
rect 100352 174412 100404 174464
rect 100904 174412 100956 174464
rect 101732 174412 101784 174464
rect 102284 174412 102336 174464
rect 103020 174412 103072 174464
rect 103664 174412 103716 174464
rect 104400 174412 104452 174464
rect 105044 174412 105096 174464
rect 105780 174412 105832 174464
rect 106424 174412 106476 174464
rect 107068 174412 107120 174464
rect 107804 174412 107856 174464
rect 116544 174412 116596 174464
rect 117464 174412 117516 174464
rect 119212 174412 119264 174464
rect 120224 174412 120276 174464
rect 124640 174412 124692 174464
rect 125744 174412 125796 174464
rect 134116 174412 134168 174464
rect 134760 174412 134812 174464
rect 171376 174412 171428 174464
rect 183612 174412 183664 174464
rect 189316 174412 189368 174464
rect 197044 174412 197096 174464
rect 197504 174412 197556 174464
rect 198424 174412 198476 174464
rect 198884 174412 198936 174464
rect 199804 174412 199856 174464
rect 200264 174412 200316 174464
rect 201092 174412 201144 174464
rect 201644 174412 201696 174464
rect 205140 174412 205192 174464
rect 205784 174412 205836 174464
rect 210568 174412 210620 174464
rect 211304 174412 211356 174464
rect 243044 173120 243096 173172
rect 151412 173052 151464 173104
rect 60792 172984 60844 173036
rect 64472 172984 64524 173036
rect 65944 172984 65996 173036
rect 68980 172984 69032 173036
rect 69900 172984 69952 173036
rect 71648 172984 71700 173036
rect 144604 172984 144656 173036
rect 144972 172984 145024 173036
rect 145708 172984 145760 173036
rect 146352 172984 146404 173036
rect 148468 172984 148520 173036
rect 149204 172984 149256 173036
rect 151320 172984 151372 173036
rect 151780 172984 151832 173036
rect 161808 172984 161860 173036
rect 162452 172984 162504 173036
rect 163188 172984 163240 173036
rect 163832 172984 163884 173036
rect 164660 172984 164712 173036
rect 231360 172984 231412 173036
rect 236788 172984 236840 173036
rect 236880 172984 236932 173036
rect 238352 172984 238404 173036
rect 242308 172984 242360 173036
rect 242860 172984 242912 173036
rect 243044 172984 243096 173036
rect 246724 172984 246776 173036
rect 247184 172984 247236 173036
rect 248840 172984 248892 173036
rect 249852 172984 249904 173036
rect 250588 172984 250640 173036
rect 251324 172984 251376 173036
rect 252152 172984 252204 173036
rect 252704 172984 252756 173036
rect 253716 172984 253768 173036
rect 254268 172984 254320 173036
rect 59412 172916 59464 172968
rect 63092 172916 63144 172968
rect 143868 172916 143920 172968
rect 145064 172916 145116 172968
rect 58676 172848 58728 172900
rect 63000 172848 63052 172900
rect 150124 172848 150176 172900
rect 162360 172916 162412 172968
rect 163464 172916 163516 172968
rect 163740 172916 163792 172968
rect 165212 172916 165264 172968
rect 235500 172916 235552 172968
rect 237800 172916 237852 172968
rect 245344 172916 245396 172968
rect 253164 172916 253216 172968
rect 253532 172916 253584 172968
rect 254820 172916 254872 172968
rect 152424 172848 152476 172900
rect 152976 172848 153028 172900
rect 156840 172848 156892 172900
rect 161256 172848 161308 172900
rect 161900 172848 161952 172900
rect 234212 172848 234264 172900
rect 237248 172848 237300 172900
rect 245436 172848 245488 172900
rect 60516 172780 60568 172832
rect 68244 172780 68296 172832
rect 150584 172780 150636 172832
rect 162268 172780 162320 172832
rect 245252 172780 245304 172832
rect 252796 172780 252848 172832
rect 253440 172848 253492 172900
rect 255556 172848 255608 172900
rect 253808 172780 253860 172832
rect 57296 172712 57348 172764
rect 67416 172712 67468 172764
rect 151688 172712 151740 172764
rect 153344 172712 153396 172764
rect 157024 172712 157076 172764
rect 248380 172712 248432 172764
rect 255924 172712 255976 172764
rect 58032 172644 58084 172696
rect 67876 172644 67928 172696
rect 138072 172644 138124 172696
rect 154816 172644 154868 172696
rect 248564 172644 248616 172696
rect 256292 172644 256344 172696
rect 54628 172576 54680 172628
rect 65576 172576 65628 172628
rect 138164 172576 138216 172628
rect 154172 172576 154224 172628
rect 156104 172576 156156 172628
rect 167420 172576 167472 172628
rect 245068 172576 245120 172628
rect 245804 172576 245856 172628
rect 249576 172576 249628 172628
rect 258316 172576 258368 172628
rect 50488 172508 50540 172560
rect 51224 172508 51276 172560
rect 61988 172508 62040 172560
rect 74408 172508 74460 172560
rect 137888 172508 137940 172560
rect 155644 172508 155696 172560
rect 155828 172508 155880 172560
rect 167972 172508 168024 172560
rect 250772 172508 250824 172560
rect 260340 172508 260392 172560
rect 137796 172440 137848 172492
rect 156196 172440 156248 172492
rect 157484 172440 157536 172492
rect 168616 172440 168668 172492
rect 241572 172440 241624 172492
rect 242400 172440 242452 172492
rect 249392 172440 249444 172492
rect 258684 172440 258736 172492
rect 61804 172372 61856 172424
rect 73672 172372 73724 172424
rect 137980 172372 138032 172424
rect 155092 172372 155144 172424
rect 155736 172372 155788 172424
rect 167236 172372 167288 172424
rect 250680 172372 250732 172424
rect 259788 172372 259840 172424
rect 38160 172304 38212 172356
rect 49200 172304 49252 172356
rect 63644 172304 63696 172356
rect 76432 172304 76484 172356
rect 137612 172304 137664 172356
rect 156840 172304 156892 172356
rect 157392 172304 157444 172356
rect 169076 172304 169128 172356
rect 249208 172304 249260 172356
rect 255924 172304 255976 172356
rect 259236 172304 259288 172356
rect 60332 172236 60384 172288
rect 60240 172168 60292 172220
rect 63644 172168 63696 172220
rect 65116 172236 65168 172288
rect 66220 172236 66272 172288
rect 151872 172236 151924 172288
rect 162544 172236 162596 172288
rect 67600 172168 67652 172220
rect 149020 172168 149072 172220
rect 154080 172168 154132 172220
rect 158220 172168 158272 172220
rect 248932 172168 248984 172220
rect 256476 172168 256528 172220
rect 55272 172032 55324 172084
rect 65116 172100 65168 172152
rect 160704 172100 160756 172152
rect 245160 172100 245212 172152
rect 252244 172100 252296 172152
rect 60608 172032 60660 172084
rect 66864 172032 66916 172084
rect 152884 172032 152936 172084
rect 159048 172032 159100 172084
rect 247828 172032 247880 172084
rect 253624 172032 253676 172084
rect 56008 171964 56060 172016
rect 60424 171964 60476 172016
rect 161072 171964 161124 172016
rect 232740 171964 232792 172016
rect 239272 171964 239324 172016
rect 247092 171964 247144 172016
rect 252060 171964 252112 172016
rect 146536 171896 146588 171948
rect 147732 171896 147784 171948
rect 152792 171896 152844 171948
rect 158496 171896 158548 171948
rect 234120 171896 234172 171948
rect 240560 171896 240612 171948
rect 245620 171896 245672 171948
rect 250864 171896 250916 171948
rect 152700 171828 152752 171880
rect 160336 171828 160388 171880
rect 243964 171828 244016 171880
rect 249668 171828 249720 171880
rect 56652 171760 56704 171812
rect 60056 171760 60108 171812
rect 152608 171760 152660 171812
rect 159600 171760 159652 171812
rect 244424 171760 244476 171812
rect 249300 171760 249352 171812
rect 53248 171692 53300 171744
rect 57572 171692 57624 171744
rect 64380 171692 64432 171744
rect 149572 171692 149624 171744
rect 161440 171692 161492 171744
rect 238260 171692 238312 171744
rect 238996 171692 239048 171744
rect 249024 171692 249076 171744
rect 60056 171624 60108 171676
rect 120224 170196 120276 170248
rect 170732 170196 170784 170248
rect 211304 170196 211356 170248
rect 233476 170196 233528 170248
rect 125744 170128 125796 170180
rect 139636 170128 139688 170180
rect 239364 169992 239416 170044
rect 240008 169992 240060 170044
rect 117464 168836 117516 168888
rect 139636 168836 139688 168888
rect 205784 168836 205836 168888
rect 233476 168836 233528 168888
rect 236696 168836 236748 168888
rect 292632 168836 292684 168888
rect 228692 168156 228744 168208
rect 228876 168156 228928 168208
rect 174044 167816 174096 167868
rect 177540 167816 177592 167868
rect 173308 167680 173360 167732
rect 180300 167680 180352 167732
rect 265860 167544 265912 167596
rect 300176 167544 300228 167596
rect 98144 167272 98196 167324
rect 109460 167272 109512 167324
rect 191984 167272 192036 167324
rect 203760 167272 203812 167324
rect 100904 167204 100956 167256
rect 114152 167204 114204 167256
rect 194744 167204 194796 167256
rect 208452 167204 208504 167256
rect 99524 167136 99576 167188
rect 112036 167136 112088 167188
rect 193364 167136 193416 167188
rect 206152 167136 206204 167188
rect 102284 167068 102336 167120
rect 116544 167068 116596 167120
rect 196124 167068 196176 167120
rect 210844 167068 210896 167120
rect 105044 167000 105096 167052
rect 121236 167000 121288 167052
rect 197504 167000 197556 167052
rect 213236 167000 213288 167052
rect 103664 166932 103716 166984
rect 118936 166932 118988 166984
rect 184992 166932 185044 166984
rect 191984 166932 192036 166984
rect 198884 166932 198936 166984
rect 215536 166932 215588 166984
rect 106424 166864 106476 166916
rect 123628 166864 123680 166916
rect 182232 166864 182284 166916
rect 187292 166864 187344 166916
rect 200264 166864 200316 166916
rect 217928 166864 217980 166916
rect 87104 166796 87156 166848
rect 90692 166796 90744 166848
rect 91244 166796 91296 166848
rect 97684 166796 97736 166848
rect 98880 166796 98932 166848
rect 102376 166796 102428 166848
rect 104400 166796 104452 166848
rect 105136 166796 105188 166848
rect 107804 166796 107856 166848
rect 125928 166796 125980 166848
rect 180852 166796 180904 166848
rect 184992 166796 185044 166848
rect 198240 166796 198292 166848
rect 199068 166796 199120 166848
rect 201644 166796 201696 166848
rect 220228 166796 220280 166848
rect 192720 166660 192772 166712
rect 196676 166660 196728 166712
rect 199620 166660 199672 166712
rect 201460 166660 201512 166712
rect 97500 166592 97552 166644
rect 100076 166592 100128 166644
rect 173124 166592 173176 166644
rect 178920 166592 178972 166644
rect 191340 166524 191392 166576
rect 194376 166524 194428 166576
rect 231820 166524 231872 166576
rect 233476 166524 233528 166576
rect 88484 166456 88536 166508
rect 92992 166456 93044 166508
rect 105780 166456 105832 166508
rect 107160 166456 107212 166508
rect 135036 166252 135088 166304
rect 139728 166252 139780 166304
rect 76708 166184 76760 166236
rect 128688 166184 128740 166236
rect 132092 166184 132144 166236
rect 139636 166184 139688 166236
rect 170732 166184 170784 166236
rect 222620 166184 222672 166236
rect 230900 166184 230952 166236
rect 233476 166184 233528 166236
rect 80204 164756 80256 164808
rect 174044 164756 174096 164808
rect 181588 164756 181640 164808
rect 87196 164688 87248 164740
rect 225932 164688 225984 164740
rect 233660 164688 233712 164740
rect 80204 163872 80256 163924
rect 85448 163872 85500 163924
rect 131908 163532 131960 163584
rect 140556 163532 140608 163584
rect 177908 163532 177960 163584
rect 181772 163532 181824 163584
rect 80204 163464 80256 163516
rect 132276 163464 132328 163516
rect 140648 163464 140700 163516
rect 132368 163396 132420 163448
rect 140372 163396 140424 163448
rect 174044 163396 174096 163448
rect 181772 163396 181824 163448
rect 87196 163328 87248 163380
rect 226392 163328 226444 163380
rect 231820 163328 231872 163380
rect 85448 163260 85500 163312
rect 87288 163260 87340 163312
rect 226484 163260 226536 163312
rect 230900 163260 230952 163312
rect 225564 163192 225616 163244
rect 233568 163192 233620 163244
rect 225932 162988 225984 163040
rect 233476 162988 233528 163040
rect 172940 162784 172992 162836
rect 179104 162784 179156 162836
rect 80112 162716 80164 162768
rect 87196 162716 87248 162768
rect 80204 162648 80256 162700
rect 87288 162648 87340 162700
rect 132644 162308 132696 162360
rect 139728 162308 139780 162360
rect 172940 162240 172992 162292
rect 179012 162240 179064 162292
rect 132644 162172 132696 162224
rect 139912 162172 139964 162224
rect 132460 162104 132512 162156
rect 135312 162104 135364 162156
rect 136232 162104 136284 162156
rect 140464 162104 140516 162156
rect 132552 162036 132604 162088
rect 134116 162036 134168 162088
rect 136324 162036 136376 162088
rect 140556 162036 140608 162088
rect 179656 162036 179708 162088
rect 182324 162036 182376 162088
rect 229336 162036 229388 162088
rect 233476 162036 233528 162088
rect 226484 161628 226536 161680
rect 233752 161628 233804 161680
rect 226484 161492 226536 161544
rect 233844 161492 233896 161544
rect 80204 161424 80256 161476
rect 87196 161424 87248 161476
rect 80112 161356 80164 161408
rect 87380 161356 87432 161408
rect 80020 161288 80072 161340
rect 87288 161288 87340 161340
rect 225932 161152 225984 161204
rect 233568 161152 233620 161204
rect 181036 160948 181088 161000
rect 181864 160948 181916 161000
rect 132644 160880 132696 160932
rect 140004 160880 140056 160932
rect 173952 160880 174004 160932
rect 181956 160880 182008 160932
rect 136416 160812 136468 160864
rect 139820 160812 139872 160864
rect 174044 160812 174096 160864
rect 181036 160812 181088 160864
rect 173124 160744 173176 160796
rect 173952 160744 174004 160796
rect 174872 160744 174924 160796
rect 182324 160744 182376 160796
rect 132552 160676 132604 160728
rect 140096 160676 140148 160728
rect 180116 160676 180168 160728
rect 182140 160676 182192 160728
rect 136508 160608 136560 160660
rect 140464 160608 140516 160660
rect 175424 160608 175476 160660
rect 181404 160608 181456 160660
rect 226484 160540 226536 160592
rect 229336 160540 229388 160592
rect 225932 160472 225984 160524
rect 233476 160472 233528 160524
rect 173032 160379 173084 160388
rect 173032 160345 173041 160379
rect 173041 160345 173075 160379
rect 173075 160345 173084 160379
rect 173032 160336 173084 160345
rect 225564 160268 225616 160320
rect 233660 160268 233712 160320
rect 80112 159928 80164 159980
rect 87196 159928 87248 159980
rect 173308 159928 173360 159980
rect 180484 159928 180536 159980
rect 80204 159860 80256 159912
rect 87288 159860 87340 159912
rect 226484 159724 226536 159776
rect 233568 159724 233620 159776
rect 172756 159588 172808 159640
rect 180668 159588 180720 159640
rect 173216 159520 173268 159572
rect 174044 159520 174096 159572
rect 132644 159452 132696 159504
rect 140924 159452 140976 159504
rect 176068 159452 176120 159504
rect 181404 159452 181456 159504
rect 132460 159384 132512 159436
rect 139268 159384 139320 159436
rect 174044 159384 174096 159436
rect 180392 159384 180444 159436
rect 132552 159316 132604 159368
rect 140740 159316 140792 159368
rect 176896 159316 176948 159368
rect 181312 159316 181364 159368
rect 132644 159248 132696 159300
rect 134944 159248 134996 159300
rect 176988 159248 177040 159300
rect 181036 159248 181088 159300
rect 80204 159180 80256 159232
rect 87196 159180 87248 159232
rect 226484 158908 226536 158960
rect 233476 158908 233528 158960
rect 225564 158636 225616 158688
rect 233568 158636 233620 158688
rect 80204 158500 80256 158552
rect 87288 158500 87340 158552
rect 226392 158228 226444 158280
rect 233476 158228 233528 158280
rect 173308 158160 173360 158212
rect 176344 158160 176396 158212
rect 132552 158092 132604 158144
rect 140648 158092 140700 158144
rect 132644 158024 132696 158076
rect 140556 158024 140608 158076
rect 135220 157956 135272 158008
rect 140372 157956 140424 158008
rect 80112 157820 80164 157872
rect 87196 157820 87248 157872
rect 80204 157752 80256 157804
rect 87288 157752 87340 157804
rect 132368 157888 132420 157940
rect 132460 157888 132512 157940
rect 136140 157888 136192 157940
rect 173124 157888 173176 157940
rect 176252 157888 176304 157940
rect 178276 157888 178328 157940
rect 181496 157888 181548 157940
rect 79468 157684 79520 157736
rect 87380 157684 87432 157736
rect 132276 157684 132328 157736
rect 226300 157684 226352 157736
rect 233476 157684 233528 157736
rect 173124 157616 173176 157668
rect 180944 157616 180996 157668
rect 173216 157548 173268 157600
rect 177908 157548 177960 157600
rect 226484 157412 226536 157464
rect 233476 157412 233528 157464
rect 131540 157140 131592 157192
rect 140832 157140 140884 157192
rect 173216 157140 173268 157192
rect 132552 157072 132604 157124
rect 137520 157072 137572 157124
rect 172940 157072 172992 157124
rect 177632 157072 177684 157124
rect 138808 156936 138860 156988
rect 140188 156936 140240 156988
rect 226484 156936 226536 156988
rect 233476 156936 233528 156988
rect 132644 156732 132696 156784
rect 140464 156732 140516 156784
rect 139728 156664 139780 156716
rect 140096 156664 140148 156716
rect 132552 156596 132604 156648
rect 138900 156596 138952 156648
rect 132644 156528 132696 156580
rect 140372 156528 140424 156580
rect 225380 156528 225432 156580
rect 233476 156528 233528 156580
rect 131908 156460 131960 156512
rect 132552 156460 132604 156512
rect 180208 156460 180260 156512
rect 182048 156460 182100 156512
rect 80112 156392 80164 156444
rect 87196 156392 87248 156444
rect 177540 156392 177592 156444
rect 181036 156392 181088 156444
rect 80204 156324 80256 156376
rect 87288 156324 87340 156376
rect 174044 156324 174096 156376
rect 181128 156324 181180 156376
rect 173952 156188 174004 156240
rect 181220 156188 181272 156240
rect 226484 155984 226536 156036
rect 233476 155984 233528 156036
rect 226484 155576 226536 155628
rect 233568 155576 233620 155628
rect 225564 155304 225616 155356
rect 233476 155304 233528 155356
rect 131816 155100 131868 155152
rect 134852 155100 134904 155152
rect 135128 155100 135180 155152
rect 139728 155100 139780 155152
rect 80112 155032 80164 155084
rect 87380 155032 87432 155084
rect 131356 155032 131408 155084
rect 135036 155032 135088 155084
rect 135312 155032 135364 155084
rect 139636 155032 139688 155084
rect 172940 155032 172992 155084
rect 175424 155032 175476 155084
rect 178920 155032 178972 155084
rect 181220 155032 181272 155084
rect 80020 154964 80072 155016
rect 87196 154964 87248 155016
rect 131448 154964 131500 155016
rect 134116 154964 134168 155016
rect 139728 154964 139780 155016
rect 173952 154964 174004 155016
rect 179656 154964 179708 155016
rect 173032 154896 173084 154948
rect 181036 154964 181088 155016
rect 131356 154828 131408 154880
rect 138992 154828 139044 154880
rect 174044 154828 174096 154880
rect 181128 154828 181180 154880
rect 139084 154760 139136 154812
rect 80204 154556 80256 154608
rect 87104 154556 87156 154608
rect 225748 154488 225800 154540
rect 233568 154488 233620 154540
rect 173124 154420 173176 154472
rect 174872 154420 174924 154472
rect 225840 154080 225892 154132
rect 233660 154080 233712 154132
rect 79928 153876 79980 153928
rect 87196 153876 87248 153928
rect 226116 153808 226168 153860
rect 233476 153808 233528 153860
rect 226484 153740 226536 153792
rect 233752 153740 233804 153792
rect 173216 153604 173268 153656
rect 181220 153604 181272 153656
rect 173308 153536 173360 153588
rect 181036 153536 181088 153588
rect 172848 153468 172900 153520
rect 173308 153400 173360 153452
rect 176068 153400 176120 153452
rect 181128 153400 181180 153452
rect 226116 153400 226168 153452
rect 233568 153400 233620 153452
rect 174044 153332 174096 153384
rect 180116 153332 180168 153384
rect 80204 153196 80256 153248
rect 87012 153196 87064 153248
rect 80204 152924 80256 152976
rect 86920 152924 86972 152976
rect 225380 152584 225432 152636
rect 233844 152584 233896 152636
rect 85816 152448 85868 152500
rect 87932 152448 87984 152500
rect 85908 152380 85960 152432
rect 87564 152380 87616 152432
rect 225748 152380 225800 152432
rect 233476 152380 233528 152432
rect 80112 152312 80164 152364
rect 87104 152312 87156 152364
rect 131540 152312 131592 152364
rect 136508 152312 136560 152364
rect 179104 152312 179156 152364
rect 181036 152312 181088 152364
rect 131356 152244 131408 152296
rect 136232 152244 136284 152296
rect 174044 152244 174096 152296
rect 176896 152244 176948 152296
rect 179012 152244 179064 152296
rect 181128 152244 181180 152296
rect 131448 152176 131500 152228
rect 136416 152176 136468 152228
rect 131356 152108 131408 152160
rect 136324 152108 136376 152160
rect 173308 151836 173360 151888
rect 176988 151836 177040 151888
rect 225932 151700 225984 151752
rect 227956 151700 228008 151752
rect 80204 151496 80256 151548
rect 86828 151496 86880 151548
rect 173952 151428 174004 151480
rect 178276 151428 178328 151480
rect 225380 151360 225432 151412
rect 229244 151360 229296 151412
rect 79376 151088 79428 151140
rect 87288 151088 87340 151140
rect 226484 151088 226536 151140
rect 228048 151088 228100 151140
rect 79744 151020 79796 151072
rect 87380 151020 87432 151072
rect 79284 150952 79336 151004
rect 87196 150952 87248 151004
rect 226116 150952 226168 151004
rect 229152 150952 229204 151004
rect 133380 150884 133432 150936
rect 139636 150884 139688 150936
rect 131356 150816 131408 150868
rect 139360 150816 139412 150868
rect 172940 150816 172992 150868
rect 182324 150816 182376 150868
rect 174044 150748 174096 150800
rect 182140 150748 182192 150800
rect 131448 150680 131500 150732
rect 139452 150680 139504 150732
rect 131356 150476 131408 150528
rect 135220 150476 135272 150528
rect 80112 150340 80164 150392
rect 85908 150340 85960 150392
rect 80204 150136 80256 150188
rect 85816 150136 85868 150188
rect 225564 150068 225616 150120
rect 230624 150068 230676 150120
rect 80020 149728 80072 149780
rect 87380 149728 87432 149780
rect 79928 149660 79980 149712
rect 87288 149660 87340 149712
rect 79836 149592 79888 149644
rect 87196 149592 87248 149644
rect 225748 149592 225800 149644
rect 230348 149592 230400 149644
rect 80204 149524 80256 149576
rect 87748 149524 87800 149576
rect 131632 149524 131684 149576
rect 139544 149524 139596 149576
rect 176252 149524 176304 149576
rect 182324 149524 182376 149576
rect 227956 149524 228008 149576
rect 233476 149524 233528 149576
rect 80112 149456 80164 149508
rect 88116 149456 88168 149508
rect 131540 149456 131592 149508
rect 139820 149456 139872 149508
rect 173308 149456 173360 149508
rect 173860 149456 173912 149508
rect 176344 149456 176396 149508
rect 181772 149456 181824 149508
rect 229152 149456 229204 149508
rect 233568 149456 233620 149508
rect 131448 149388 131500 149440
rect 139176 149388 139228 149440
rect 174044 149388 174096 149440
rect 180760 149388 180812 149440
rect 131356 149320 131408 149372
rect 138808 149320 138860 149372
rect 173860 149320 173912 149372
rect 180208 149320 180260 149372
rect 225380 149048 225432 149100
rect 233752 149048 233804 149100
rect 132276 148844 132328 148896
rect 139636 148844 139688 148896
rect 174044 148844 174096 148896
rect 180944 148844 180996 148896
rect 226484 148640 226536 148692
rect 233936 148640 233988 148692
rect 225564 148300 225616 148352
rect 233660 148300 233712 148352
rect 226484 148232 226536 148284
rect 233844 148232 233896 148284
rect 134944 148164 134996 148216
rect 139728 148164 139780 148216
rect 229244 148164 229296 148216
rect 233476 148164 233528 148216
rect 131356 148096 131408 148148
rect 135128 148096 135180 148148
rect 228048 148096 228100 148148
rect 233568 148096 233620 148148
rect 177632 148028 177684 148080
rect 182324 148028 182376 148080
rect 172756 147824 172808 147876
rect 180852 147824 180904 147876
rect 174044 147756 174096 147808
rect 180576 147756 180628 147808
rect 225564 147348 225616 147400
rect 232004 147348 232056 147400
rect 136140 146736 136192 146788
rect 139728 146736 139780 146788
rect 174044 146668 174096 146720
rect 181956 146668 182008 146720
rect 230624 146668 230676 146720
rect 233476 146668 233528 146720
rect 172756 146328 172808 146380
rect 174780 146328 174832 146380
rect 230348 146328 230400 146380
rect 233476 146328 233528 146380
rect 228324 145963 228376 145972
rect 228324 145929 228333 145963
rect 228333 145929 228367 145963
rect 228367 145929 228376 145963
rect 228324 145920 228376 145929
rect 80204 145376 80256 145428
rect 87472 145376 87524 145428
rect 137520 145376 137572 145428
rect 139912 145376 139964 145428
rect 173676 145376 173728 145428
rect 176160 145376 176212 145428
rect 203852 145376 203904 145428
rect 226576 145308 226628 145360
rect 233476 145308 233528 145360
rect 228324 145283 228376 145292
rect 228324 145249 228333 145283
rect 228333 145249 228367 145283
rect 228367 145249 228376 145283
rect 228324 145240 228376 145249
rect 170824 144696 170876 144748
rect 171376 144696 171428 144748
rect 80020 144016 80072 144068
rect 87196 144016 87248 144068
rect 109552 144016 109604 144068
rect 134760 144016 134812 144068
rect 134852 144016 134904 144068
rect 139728 144016 139780 144068
rect 296220 144016 296272 144068
rect 300176 144016 300228 144068
rect 80204 143948 80256 144000
rect 87564 143948 87616 144000
rect 80112 143880 80164 143932
rect 87288 143880 87340 143932
rect 80204 142656 80256 142708
rect 87380 142656 87432 142708
rect 232004 142656 232056 142708
rect 233476 142656 233528 142708
rect 169996 141704 170048 141756
rect 170640 141704 170692 141756
rect 168432 141636 168484 141688
rect 170732 141636 170784 141688
rect 56744 139868 56796 139920
rect 60056 139868 60108 139920
rect 56468 139800 56520 139852
rect 60976 139800 61028 139852
rect 65116 139868 65168 139920
rect 132000 139868 132052 139920
rect 168984 139868 169036 139920
rect 224460 139868 224512 139920
rect 67140 139800 67192 139852
rect 140280 139800 140332 139852
rect 169444 139800 169496 139852
rect 59964 139732 60016 139784
rect 71832 139732 71884 139784
rect 149388 139732 149440 139784
rect 157852 139732 157904 139784
rect 57112 139664 57164 139716
rect 61712 139664 61764 139716
rect 63828 139664 63880 139716
rect 150492 139664 150544 139716
rect 59872 139596 59924 139648
rect 71096 139596 71148 139648
rect 155276 139664 155328 139716
rect 165764 139664 165816 139716
rect 242768 139664 242820 139716
rect 159232 139596 159284 139648
rect 54444 139528 54496 139580
rect 57572 139528 57624 139580
rect 59688 139528 59740 139580
rect 60516 139528 60568 139580
rect 61160 139528 61212 139580
rect 61988 139528 62040 139580
rect 62448 139528 62500 139580
rect 65760 139528 65812 139580
rect 67232 139528 67284 139580
rect 70452 139528 70504 139580
rect 73764 139528 73816 139580
rect 155000 139528 155052 139580
rect 166316 139528 166368 139580
rect 243044 139528 243096 139580
rect 250772 139800 250824 139852
rect 263836 139868 263888 139920
rect 254176 139800 254228 139852
rect 247644 139732 247696 139784
rect 250864 139732 250916 139784
rect 254452 139732 254504 139784
rect 249668 139664 249720 139716
rect 244884 139596 244936 139648
rect 249392 139596 249444 139648
rect 250036 139596 250088 139648
rect 251968 139596 252020 139648
rect 255556 139596 255608 139648
rect 260432 139596 260484 139648
rect 245804 139528 245856 139580
rect 249116 139528 249168 139580
rect 249208 139528 249260 139580
rect 250680 139528 250732 139580
rect 251876 139528 251928 139580
rect 252704 139528 252756 139580
rect 58492 139460 58544 139512
rect 60608 139460 60660 139512
rect 60700 139460 60752 139512
rect 72476 139460 72528 139512
rect 149112 139460 149164 139512
rect 157576 139460 157628 139512
rect 160520 139460 160572 139512
rect 242216 139460 242268 139512
rect 247920 139460 247972 139512
rect 59136 139392 59188 139444
rect 60424 139392 60476 139444
rect 59044 139324 59096 139376
rect 63184 139392 63236 139444
rect 63644 139392 63696 139444
rect 75788 139392 75840 139444
rect 153252 139392 153304 139444
rect 60792 139324 60844 139376
rect 73120 139324 73172 139376
rect 137980 139324 138032 139376
rect 145156 139324 145208 139376
rect 155184 139324 155236 139376
rect 155920 139324 155972 139376
rect 166868 139392 166920 139444
rect 251048 139460 251100 139512
rect 251324 139460 251376 139512
rect 261444 139460 261496 139512
rect 163648 139324 163700 139376
rect 245344 139324 245396 139376
rect 250128 139392 250180 139444
rect 253440 139392 253492 139444
rect 259880 139392 259932 139444
rect 249760 139324 249812 139376
rect 252152 139324 252204 139376
rect 258776 139324 258828 139376
rect 55180 139256 55232 139308
rect 57480 139256 57532 139308
rect 59780 139256 59832 139308
rect 60884 139256 60936 139308
rect 61344 139256 61396 139308
rect 74500 139256 74552 139308
rect 138992 139256 139044 139308
rect 146260 139256 146312 139308
rect 38252 139188 38304 139240
rect 49200 139188 49252 139240
rect 53156 139188 53208 139240
rect 61804 139188 61856 139240
rect 60148 139120 60200 139172
rect 66496 139188 66548 139240
rect 67140 139188 67192 139240
rect 69808 139188 69860 139240
rect 75144 139188 75196 139240
rect 137888 139188 137940 139240
rect 145708 139188 145760 139240
rect 60240 139052 60292 139104
rect 61252 139052 61304 139104
rect 65484 139052 65536 139104
rect 149940 139052 149992 139104
rect 158864 139256 158916 139308
rect 163096 139256 163148 139308
rect 231820 139256 231872 139308
rect 238996 139256 239048 139308
rect 245436 139256 245488 139308
rect 249300 139256 249352 139308
rect 154172 139188 154224 139240
rect 155552 139188 155604 139240
rect 155828 139188 155880 139240
rect 167328 139188 167380 139240
rect 231728 139188 231780 139240
rect 239456 139188 239508 139240
rect 245712 139188 245764 139240
rect 250496 139256 250548 139308
rect 259328 139256 259380 139308
rect 249576 139188 249628 139240
rect 256936 139188 256988 139240
rect 155368 139120 155420 139172
rect 159416 139120 159468 139172
rect 248932 139120 248984 139172
rect 255004 139120 255056 139172
rect 154724 139052 154776 139104
rect 155460 139052 155512 139104
rect 155736 139052 155788 139104
rect 159968 139052 160020 139104
rect 249852 139052 249904 139104
rect 261168 139188 261220 139240
rect 55824 138984 55876 139036
rect 58860 138984 58912 139036
rect 59504 138984 59556 139036
rect 61436 138984 61488 139036
rect 152700 138984 152752 139036
rect 60332 138916 60384 138968
rect 61528 138916 61580 138968
rect 64472 138916 64524 138968
rect 153620 138916 153672 138968
rect 154724 138916 154776 138968
rect 156012 138984 156064 139036
rect 156748 138984 156800 139036
rect 165212 138984 165264 139036
rect 246540 138984 246592 139036
rect 249484 138984 249536 139036
rect 250220 138984 250272 139036
rect 252888 138984 252940 139036
rect 156932 138916 156984 138968
rect 164752 138916 164804 138968
rect 243872 138916 243924 138968
rect 249024 138916 249076 138968
rect 57848 138848 57900 138900
rect 61896 138848 61948 138900
rect 69164 138848 69216 138900
rect 151044 138848 151096 138900
rect 157576 138848 157628 138900
rect 158404 138848 158456 138900
rect 161072 138848 161124 138900
rect 231360 138848 231412 138900
rect 237248 138848 237300 138900
rect 245620 138848 245672 138900
rect 249208 138848 249260 138900
rect 256108 138848 256160 138900
rect 67784 138780 67836 138832
rect 137796 138780 137848 138832
rect 144696 138780 144748 138832
rect 151504 138780 151556 138832
rect 158220 138780 158272 138832
rect 158312 138780 158364 138832
rect 161532 138780 161584 138832
rect 68428 138712 68480 138764
rect 137704 138712 137756 138764
rect 144144 138712 144196 138764
rect 147824 138712 147876 138764
rect 154264 138712 154316 138764
rect 155644 138712 155696 138764
rect 158956 138712 159008 138764
rect 161072 138712 161124 138764
rect 164200 138780 164252 138832
rect 231636 138780 231688 138832
rect 238352 138780 238404 138832
rect 248380 138780 248432 138832
rect 254820 138780 254872 138832
rect 258316 138780 258368 138832
rect 163740 138712 163792 138764
rect 167880 138712 167932 138764
rect 231544 138712 231596 138764
rect 237800 138712 237852 138764
rect 250404 138712 250456 138764
rect 66680 138644 66732 138696
rect 137612 138644 137664 138696
rect 143592 138644 143644 138696
rect 147272 138644 147324 138696
rect 154080 138644 154132 138696
rect 60976 138576 61028 138628
rect 63000 138576 63052 138628
rect 62264 138508 62316 138560
rect 137520 138576 137572 138628
rect 142764 138576 142816 138628
rect 148376 138576 148428 138628
rect 149020 138576 149072 138628
rect 152056 138576 152108 138628
rect 153160 138576 153212 138628
rect 156288 138644 156340 138696
rect 157484 138644 157536 138696
rect 157576 138644 157628 138696
rect 158496 138644 158548 138696
rect 160980 138644 161032 138696
rect 162636 138644 162688 138696
rect 231452 138644 231504 138696
rect 236788 138644 236840 138696
rect 244424 138644 244476 138696
rect 246540 138644 246592 138696
rect 247092 138644 247144 138696
rect 253440 138644 253492 138696
rect 254912 138644 254964 138696
rect 257764 138644 257816 138696
rect 152884 138508 152936 138560
rect 156840 138576 156892 138628
rect 157300 138576 157352 138628
rect 161164 138576 161216 138628
rect 162084 138576 162136 138628
rect 167880 138576 167932 138628
rect 170824 138576 170876 138628
rect 232924 138576 232976 138628
rect 240008 138576 240060 138628
rect 245804 138576 245856 138628
rect 255004 138576 255056 138628
rect 257212 138576 257264 138628
rect 261996 138576 262048 138628
rect 263192 138576 263244 138628
rect 263744 138576 263796 138628
rect 126480 135788 126532 135840
rect 159600 135788 159652 135840
rect 220504 135788 220556 135840
rect 255464 135788 255516 135840
rect 136876 132932 136928 132984
rect 146812 132932 146864 132984
rect 231912 132932 231964 132984
rect 240560 132932 240612 132984
rect 250036 131708 250088 131760
rect 148928 131640 148980 131692
rect 149204 131640 149256 131692
rect 56192 131572 56244 131624
rect 56744 131572 56796 131624
rect 57388 131572 57440 131624
rect 60056 131572 60108 131624
rect 60424 131572 60476 131624
rect 68336 131572 68388 131624
rect 150216 131572 150268 131624
rect 155368 131572 155420 131624
rect 155460 131572 155512 131624
rect 157300 131572 157352 131624
rect 163924 131572 163976 131624
rect 244884 131572 244936 131624
rect 245344 131572 245396 131624
rect 248012 131572 248064 131624
rect 248564 131572 248616 131624
rect 250496 131572 250548 131624
rect 55088 131504 55140 131556
rect 59044 131504 59096 131556
rect 57572 131436 57624 131488
rect 65576 131504 65628 131556
rect 149848 131504 149900 131556
rect 155644 131504 155696 131556
rect 157392 131504 157444 131556
rect 164292 131504 164344 131556
rect 243320 131504 243372 131556
rect 249484 131504 249536 131556
rect 254268 131572 254320 131624
rect 255464 131572 255516 131624
rect 258408 131572 258460 131624
rect 255004 131504 255056 131556
rect 59688 131436 59740 131488
rect 60424 131436 60476 131488
rect 57480 131368 57532 131420
rect 60516 131368 60568 131420
rect 53984 131300 54036 131352
rect 65208 131436 65260 131488
rect 153160 131436 153212 131488
rect 160428 131436 160480 131488
rect 250036 131436 250088 131488
rect 61528 131368 61580 131420
rect 61620 131368 61672 131420
rect 64380 131300 64432 131352
rect 60884 131232 60936 131284
rect 63368 131232 63420 131284
rect 67232 131368 67284 131420
rect 151044 131368 151096 131420
rect 152700 131368 152752 131420
rect 152976 131368 153028 131420
rect 157484 131368 157536 131420
rect 163556 131368 163608 131420
rect 248472 131368 248524 131420
rect 255648 131436 255700 131488
rect 252060 131368 252112 131420
rect 252704 131368 252756 131420
rect 258316 131368 258368 131420
rect 154724 131300 154776 131352
rect 161532 131300 161584 131352
rect 248012 131300 248064 131352
rect 254820 131300 254872 131352
rect 52420 131164 52472 131216
rect 59320 131164 59372 131216
rect 149480 131164 149532 131216
rect 157668 131232 157720 131284
rect 160980 131232 161032 131284
rect 175424 131232 175476 131284
rect 281868 131232 281920 131284
rect 152608 131164 152660 131216
rect 156472 131164 156524 131216
rect 163740 131164 163792 131216
rect 249392 131164 249444 131216
rect 252980 131164 253032 131216
rect 51040 131096 51092 131148
rect 57020 131096 57072 131148
rect 60332 131096 60384 131148
rect 60424 131096 60476 131148
rect 69072 131096 69124 131148
rect 149204 131096 149256 131148
rect 158036 131096 158088 131148
rect 159600 131096 159652 131148
rect 164660 131096 164712 131148
rect 246540 131096 246592 131148
rect 249944 131096 249996 131148
rect 256936 131096 256988 131148
rect 63276 131028 63328 131080
rect 153712 131028 153764 131080
rect 51224 130960 51276 131012
rect 58768 130960 58820 131012
rect 58860 130960 58912 131012
rect 60608 130960 60660 131012
rect 67968 130960 68020 131012
rect 149020 130960 149072 131012
rect 157668 130960 157720 131012
rect 162360 131028 162412 131080
rect 249024 131028 249076 131080
rect 252244 131028 252296 131080
rect 161072 130960 161124 131012
rect 250312 130960 250364 131012
rect 257212 130960 257264 131012
rect 49844 130892 49896 130944
rect 62816 130892 62868 130944
rect 52604 130824 52656 130876
rect 64012 130892 64064 130944
rect 65760 130892 65812 130944
rect 70268 130892 70320 130944
rect 63000 130824 63052 130876
rect 66772 130824 66824 130876
rect 151412 130824 151464 130876
rect 56560 130756 56612 130808
rect 61252 130756 61304 130808
rect 61988 130756 62040 130808
rect 69532 130756 69584 130808
rect 151780 130756 151832 130808
rect 158312 130892 158364 130944
rect 241664 130892 241716 130944
rect 250588 130892 250640 130944
rect 252888 130892 252940 130944
rect 158404 130824 158456 130876
rect 247184 130824 247236 130876
rect 253716 130824 253768 130876
rect 155552 130756 155604 130808
rect 160796 130756 160848 130808
rect 243688 130756 243740 130808
rect 58124 130688 58176 130740
rect 60148 130688 60200 130740
rect 58584 130620 58636 130672
rect 59504 130620 59556 130672
rect 61712 130688 61764 130740
rect 61896 130688 61948 130740
rect 67508 130688 67560 130740
rect 153068 130688 153120 130740
rect 55456 130552 55508 130604
rect 62172 130620 62224 130672
rect 69900 130620 69952 130672
rect 60976 130552 61028 130604
rect 68704 130552 68756 130604
rect 150584 130552 150636 130604
rect 155736 130620 155788 130672
rect 155920 130688 155972 130740
rect 156104 130620 156156 130672
rect 154264 130552 154316 130604
rect 157300 130552 157352 130604
rect 161164 130620 161216 130672
rect 244056 130688 244108 130740
rect 250220 130756 250272 130808
rect 250680 130756 250732 130808
rect 245252 130688 245304 130740
rect 245712 130688 245764 130740
rect 246816 130688 246868 130740
rect 249576 130688 249628 130740
rect 162728 130620 162780 130672
rect 250312 130688 250364 130740
rect 251324 130688 251376 130740
rect 163096 130552 163148 130604
rect 244332 130552 244384 130604
rect 246448 130552 246500 130604
rect 249208 130552 249260 130604
rect 58952 130484 59004 130536
rect 67140 130484 67192 130536
rect 154172 130484 154224 130536
rect 156932 130484 156984 130536
rect 161992 130484 162044 130536
rect 249116 130484 249168 130536
rect 251232 130620 251284 130672
rect 255556 130688 255608 130740
rect 250772 130552 250824 130604
rect 251784 130552 251836 130604
rect 256108 130620 256160 130672
rect 257672 130552 257724 130604
rect 250864 130484 250916 130536
rect 254912 130484 254964 130536
rect 57756 130416 57808 130468
rect 60240 130416 60292 130468
rect 55824 130348 55876 130400
rect 61344 130348 61396 130400
rect 61712 130348 61764 130400
rect 61896 130416 61948 130468
rect 64840 130416 64892 130468
rect 62448 130348 62500 130400
rect 63644 130348 63696 130400
rect 66404 130416 66456 130468
rect 154080 130416 154132 130468
rect 156564 130416 156616 130468
rect 13780 130280 13832 130332
rect 31904 130280 31956 130332
rect 38344 130280 38396 130332
rect 65944 130348 65996 130400
rect 70636 130348 70688 130400
rect 154540 130348 154592 130400
rect 156840 130348 156892 130400
rect 152148 130280 152200 130332
rect 136876 130212 136928 130264
rect 138992 130212 139044 130264
rect 154908 130280 154960 130332
rect 155276 130280 155328 130332
rect 155736 130280 155788 130332
rect 156012 130280 156064 130332
rect 161164 130416 161216 130468
rect 247552 130416 247604 130468
rect 254820 130416 254872 130468
rect 158220 130348 158272 130400
rect 159968 130348 160020 130400
rect 247920 130348 247972 130400
rect 250956 130348 251008 130400
rect 251048 130348 251100 130400
rect 251416 130348 251468 130400
rect 252152 130348 252204 130400
rect 256476 130348 256528 130400
rect 158496 130280 158548 130332
rect 159600 130280 159652 130332
rect 249300 130280 249352 130332
rect 253348 130280 253400 130332
rect 253440 130280 253492 130332
rect 254544 130280 254596 130332
rect 232004 130212 232056 130264
rect 232924 130212 232976 130264
rect 136876 127492 136928 127544
rect 145340 127492 145392 127544
rect 228508 127560 228560 127612
rect 230716 127492 230768 127544
rect 239640 127492 239692 127544
rect 228416 127424 228468 127476
rect 148744 126608 148796 126660
rect 165120 126608 165172 126660
rect 231636 124976 231688 125028
rect 238260 124976 238312 125028
rect 138164 124840 138216 124892
rect 144420 124840 144472 124892
rect 137888 124772 137940 124824
rect 145616 124772 145668 124824
rect 231912 124772 231964 124824
rect 240928 124772 240980 124824
rect 228416 124747 228468 124756
rect 228416 124713 228425 124747
rect 228425 124713 228459 124747
rect 228459 124713 228468 124747
rect 228416 124704 228468 124713
rect 47820 122188 47872 122240
rect 51316 122188 51368 122240
rect 138164 122052 138216 122104
rect 143040 122052 143092 122104
rect 231636 122052 231688 122104
rect 236880 122052 236932 122104
rect 137980 121984 138032 122036
rect 145616 121984 145668 122036
rect 232004 121984 232056 122036
rect 240928 121984 240980 122036
rect 165120 121916 165172 121968
rect 175516 121916 175568 121968
rect 228508 120488 228560 120540
rect 138072 119264 138124 119316
rect 145616 119264 145668 119316
rect 231912 119264 231964 119316
rect 240928 119264 240980 119316
rect 231636 118448 231688 118500
rect 235500 118448 235552 118500
rect 138164 117904 138216 117956
rect 141660 117904 141712 117956
rect 137796 117836 137848 117888
rect 145616 117836 145668 117888
rect 231636 117836 231688 117888
rect 240928 117836 240980 117888
rect 292816 117836 292868 117888
rect 300176 117836 300228 117888
rect 137336 115184 137388 115236
rect 140280 115184 140332 115236
rect 231268 115184 231320 115236
rect 234120 115184 234172 115236
rect 137704 115116 137756 115168
rect 145616 115116 145668 115168
rect 231544 115116 231596 115168
rect 240928 115116 240980 115168
rect 263744 115048 263796 115100
rect 274876 115048 274928 115100
rect 138164 112532 138216 112584
rect 138992 112532 139044 112584
rect 292816 112507 292868 112516
rect 292816 112473 292825 112507
rect 292825 112473 292859 112507
rect 292859 112473 292868 112507
rect 292816 112464 292868 112473
rect 137428 112328 137480 112380
rect 145616 112328 145668 112380
rect 231268 112328 231320 112380
rect 240744 112328 240796 112380
rect 292816 111920 292868 111972
rect 293552 111920 293604 111972
rect 138164 110968 138216 111020
rect 145616 110968 145668 111020
rect 232004 110968 232056 111020
rect 240928 110968 240980 111020
rect 292816 110263 292868 110272
rect 292816 110229 292825 110263
rect 292825 110229 292859 110263
rect 292859 110229 292868 110263
rect 292816 110220 292868 110229
rect 231544 109540 231596 109592
rect 232832 109540 232884 109592
rect 47084 109472 47136 109524
rect 51316 109472 51368 109524
rect 137336 108180 137388 108232
rect 145616 108180 145668 108232
rect 228508 108180 228560 108232
rect 231452 108180 231504 108232
rect 240836 108180 240888 108232
rect 228508 108044 228560 108096
rect 140372 105460 140424 105512
rect 145616 105460 145668 105512
rect 231728 105460 231780 105512
rect 240928 105460 240980 105512
rect 143132 103080 143184 103132
rect 145432 103080 145484 103132
rect 236972 102672 237024 102724
rect 240744 102672 240796 102724
rect 265124 102672 265176 102724
rect 274876 102672 274928 102724
rect 140464 101312 140516 101364
rect 145616 101312 145668 101364
rect 234212 101312 234264 101364
rect 240376 101312 240428 101364
rect 140556 98524 140608 98576
rect 145616 98524 145668 98576
rect 167880 98524 167932 98576
rect 175516 98524 175568 98576
rect 234304 98524 234356 98576
rect 240836 98524 240888 98576
rect 262364 98524 262416 98576
rect 272760 98524 272812 98576
rect 74040 97096 74092 97148
rect 81676 97096 81728 97148
rect 238352 95804 238404 95856
rect 240928 95804 240980 95856
rect 138164 95736 138216 95788
rect 140372 95736 140424 95788
rect 228508 95779 228560 95788
rect 228508 95745 228517 95779
rect 228517 95745 228551 95779
rect 228551 95745 228560 95779
rect 228508 95736 228560 95745
rect 45796 94376 45848 94428
rect 51316 94376 51368 94428
rect 143776 94376 143828 94428
rect 146352 94376 146404 94428
rect 237616 94376 237668 94428
rect 240928 94376 240980 94428
rect 292816 94376 292868 94428
rect 299716 94376 299768 94428
rect 272760 94308 272812 94360
rect 274876 94308 274928 94360
rect 231820 94172 231872 94224
rect 236972 94172 237024 94224
rect 138164 93832 138216 93884
rect 143132 93832 143184 93884
rect 38804 92948 38856 93000
rect 45796 92948 45848 93000
rect 231452 92948 231504 93000
rect 234212 92948 234264 93000
rect 137796 92676 137848 92728
rect 140464 92676 140516 92728
rect 143684 91656 143736 91708
rect 145248 91656 145300 91708
rect 236328 91656 236380 91708
rect 240928 91656 240980 91708
rect 137612 91588 137664 91640
rect 140556 91588 140608 91640
rect 231452 91588 231504 91640
rect 234304 91588 234356 91640
rect 228508 90883 228560 90892
rect 228508 90849 228517 90883
rect 228517 90849 228551 90883
rect 228551 90849 228560 90883
rect 228508 90840 228560 90849
rect 231636 90024 231688 90076
rect 238352 90024 238404 90076
rect 138164 89140 138216 89192
rect 144604 89140 144656 89192
rect 155276 88936 155328 88988
rect 155552 88936 155604 88988
rect 143500 88868 143552 88920
rect 145248 88868 145300 88920
rect 236236 88868 236288 88920
rect 240928 88868 240980 88920
rect 137612 88800 137664 88852
rect 143776 88800 143828 88852
rect 231636 88460 231688 88512
rect 237616 88460 237668 88512
rect 292540 88120 292592 88172
rect 292724 88120 292776 88172
rect 23900 87440 23952 87492
rect 31904 87440 31956 87492
rect 34572 87440 34624 87492
rect 55088 87440 55140 87492
rect 56100 87440 56152 87492
rect 58676 87440 58728 87492
rect 65484 87440 65536 87492
rect 154172 87440 154224 87492
rect 157392 87440 157444 87492
rect 160704 87440 160756 87492
rect 160980 87440 161032 87492
rect 162268 87440 162320 87492
rect 254360 87440 254412 87492
rect 59872 87372 59924 87424
rect 70728 87372 70780 87424
rect 152700 87372 152752 87424
rect 158404 87372 158456 87424
rect 159600 87372 159652 87424
rect 161072 87372 161124 87424
rect 249944 87372 249996 87424
rect 256936 87372 256988 87424
rect 34664 87304 34716 87356
rect 58216 87304 58268 87356
rect 67140 87304 67192 87356
rect 153068 87304 153120 87356
rect 158220 87304 158272 87356
rect 246080 87304 246132 87356
rect 255740 87304 255792 87356
rect 53984 87236 54036 87288
rect 60240 87236 60292 87288
rect 70820 87236 70872 87288
rect 152700 87236 152752 87288
rect 157484 87236 157536 87288
rect 161072 87236 161124 87288
rect 161900 87236 161952 87288
rect 246540 87236 246592 87288
rect 256936 87236 256988 87288
rect 67232 87168 67284 87220
rect 150308 87168 150360 87220
rect 159324 87168 159376 87220
rect 246908 87168 246960 87220
rect 257028 87168 257080 87220
rect 63828 87100 63880 87152
rect 154080 87100 154132 87152
rect 157484 87100 157536 87152
rect 158312 87100 158364 87152
rect 248104 87100 248156 87152
rect 256292 87100 256344 87152
rect 52604 87032 52656 87084
rect 64656 87032 64708 87084
rect 149848 87032 149900 87084
rect 158956 87032 159008 87084
rect 247736 87032 247788 87084
rect 256476 87032 256528 87084
rect 51224 86964 51276 87016
rect 63460 86964 63512 87016
rect 151320 86964 151372 87016
rect 157116 86964 157168 87016
rect 159048 86964 159100 87016
rect 247184 86964 247236 87016
rect 251048 86964 251100 87016
rect 257212 86964 257264 87016
rect 52512 86896 52564 86948
rect 64288 86896 64340 86948
rect 152240 86896 152292 86948
rect 157852 86896 157904 86948
rect 247000 86896 247052 86948
rect 251324 86896 251376 86948
rect 257580 86896 257632 86948
rect 49844 86828 49896 86880
rect 63092 86828 63144 86880
rect 63644 86828 63696 86880
rect 70636 86828 70688 86880
rect 149112 86828 149164 86880
rect 157760 86828 157812 86880
rect 158864 86828 158916 86880
rect 164660 86828 164712 86880
rect 245712 86828 245764 86880
rect 256200 86828 256252 86880
rect 51132 86760 51184 86812
rect 59044 86760 59096 86812
rect 66772 86760 66824 86812
rect 156012 86760 156064 86812
rect 158680 86760 158732 86812
rect 245344 86760 245396 86812
rect 256108 86760 256160 86812
rect 57480 86692 57532 86744
rect 61804 86692 61856 86744
rect 153344 86692 153396 86744
rect 155644 86692 155696 86744
rect 159508 86692 159560 86744
rect 245160 86692 245212 86744
rect 251140 86692 251192 86744
rect 254268 86692 254320 86744
rect 61344 86624 61396 86676
rect 69808 86624 69860 86676
rect 150584 86624 150636 86676
rect 60884 86556 60936 86608
rect 69440 86556 69492 86608
rect 150676 86556 150728 86608
rect 155368 86556 155420 86608
rect 57020 86488 57072 86540
rect 61712 86488 61764 86540
rect 61988 86488 62040 86540
rect 69900 86488 69952 86540
rect 155184 86488 155236 86540
rect 156104 86624 156156 86676
rect 162636 86624 162688 86676
rect 247920 86624 247972 86676
rect 251600 86624 251652 86676
rect 252704 86624 252756 86676
rect 258316 86624 258368 86676
rect 155920 86556 155972 86608
rect 163096 86556 163148 86608
rect 247828 86556 247880 86608
rect 251508 86556 251560 86608
rect 59412 86420 59464 86472
rect 67324 86420 67376 86472
rect 151044 86420 151096 86472
rect 155552 86420 155604 86472
rect 156656 86488 156708 86540
rect 159784 86488 159836 86540
rect 244884 86488 244936 86540
rect 249484 86488 249536 86540
rect 250956 86488 251008 86540
rect 251232 86488 251284 86540
rect 57848 86352 57900 86404
rect 61620 86352 61672 86404
rect 61896 86352 61948 86404
rect 65852 86352 65904 86404
rect 153436 86352 153488 86404
rect 156656 86352 156708 86404
rect 55824 86284 55876 86336
rect 60516 86284 60568 86336
rect 61068 86284 61120 86336
rect 61988 86284 62040 86336
rect 62264 86284 62316 86336
rect 70268 86284 70320 86336
rect 151504 86284 151556 86336
rect 155460 86284 155512 86336
rect 157392 86420 157444 86472
rect 163832 86420 163884 86472
rect 248932 86420 248984 86472
rect 251416 86420 251468 86472
rect 157484 86352 157536 86404
rect 164292 86352 164344 86404
rect 249392 86352 249444 86404
rect 252428 86352 252480 86404
rect 163464 86284 163516 86336
rect 243320 86284 243372 86336
rect 248380 86284 248432 86336
rect 249116 86284 249168 86336
rect 249852 86284 249904 86336
rect 250680 86284 250732 86336
rect 253624 86284 253676 86336
rect 55456 86216 55508 86268
rect 60332 86216 60384 86268
rect 64380 86216 64432 86268
rect 67416 86216 67468 86268
rect 154264 86216 154316 86268
rect 157024 86216 157076 86268
rect 157116 86216 157168 86268
rect 159876 86216 159928 86268
rect 244424 86216 244476 86268
rect 248288 86216 248340 86268
rect 249576 86216 249628 86268
rect 251968 86216 252020 86268
rect 252612 86216 252664 86268
rect 258408 86216 258460 86268
rect 56284 86148 56336 86200
rect 60424 86148 60476 86200
rect 61988 86148 62040 86200
rect 65024 86148 65076 86200
rect 65760 86148 65812 86200
rect 67048 86148 67100 86200
rect 154632 86148 154684 86200
rect 156932 86148 156984 86200
rect 157208 86148 157260 86200
rect 160244 86148 160296 86200
rect 243688 86148 243740 86200
rect 248012 86148 248064 86200
rect 249300 86148 249352 86200
rect 249852 86148 249904 86200
rect 56652 86080 56704 86132
rect 60240 86080 60292 86132
rect 62632 86080 62684 86132
rect 63552 86080 63604 86132
rect 65852 86080 65904 86132
rect 66680 86080 66732 86132
rect 66772 86080 66824 86132
rect 67416 86080 67468 86132
rect 67508 86080 67560 86132
rect 69072 86080 69124 86132
rect 149480 86080 149532 86132
rect 150492 86080 150544 86132
rect 153896 86080 153948 86132
rect 154724 86080 154776 86132
rect 155092 86080 155144 86132
rect 155828 86080 155880 86132
rect 156288 86080 156340 86132
rect 157300 86080 157352 86132
rect 158312 86080 158364 86132
rect 159692 86080 159744 86132
rect 161440 86080 161492 86132
rect 244148 86080 244200 86132
rect 248196 86080 248248 86132
rect 252796 86148 252848 86200
rect 253440 86148 253492 86200
rect 255188 86148 255240 86200
rect 250772 86080 250824 86132
rect 253164 86080 253216 86132
rect 253532 86080 253584 86132
rect 254820 86080 254872 86132
rect 255556 86080 255608 86132
rect 256384 86080 256436 86132
rect 231636 86012 231688 86064
rect 236328 86012 236380 86064
rect 249300 86012 249352 86064
rect 256016 85876 256068 85928
rect 256200 85876 256252 85928
rect 256292 85604 256344 85656
rect 256568 85604 256620 85656
rect 136876 85196 136928 85248
rect 143684 85196 143736 85248
rect 136876 84652 136928 84704
rect 143500 84652 143552 84704
rect 231636 84652 231688 84704
rect 236236 84652 236288 84704
rect 155552 84244 155604 84296
rect 160428 84244 160480 84296
rect 92256 83972 92308 84024
rect 89588 83904 89640 83956
rect 90876 83904 90928 83956
rect 67876 83836 67928 83888
rect 68244 83836 68296 83888
rect 86828 83879 86880 83888
rect 86828 83845 86837 83879
rect 86837 83845 86871 83879
rect 86871 83845 86880 83879
rect 86828 83836 86880 83845
rect 88208 83836 88260 83888
rect 93636 83879 93688 83888
rect 93636 83845 93645 83879
rect 93645 83845 93679 83879
rect 93679 83845 93688 83879
rect 93636 83836 93688 83845
rect 94924 83879 94976 83888
rect 94924 83845 94933 83879
rect 94933 83845 94967 83879
rect 94967 83845 94976 83879
rect 94924 83836 94976 83845
rect 116544 83904 116596 83956
rect 120592 83947 120644 83956
rect 120592 83913 120601 83947
rect 120601 83913 120635 83947
rect 120635 83913 120644 83947
rect 120592 83904 120644 83913
rect 124640 83904 124692 83956
rect 127308 83904 127360 83956
rect 134852 83904 134904 83956
rect 96304 83836 96356 83888
rect 97684 83836 97736 83888
rect 91980 83768 92032 83820
rect 96120 83768 96172 83820
rect 98972 83836 99024 83888
rect 100352 83836 100404 83888
rect 101732 83836 101784 83888
rect 103020 83836 103072 83888
rect 104400 83836 104452 83888
rect 105780 83836 105832 83888
rect 107068 83836 107120 83888
rect 108448 83836 108500 83888
rect 109828 83879 109880 83888
rect 109828 83845 109837 83879
rect 109837 83845 109871 83879
rect 109871 83845 109880 83879
rect 109828 83836 109880 83845
rect 111116 83836 111168 83888
rect 112496 83879 112548 83888
rect 112496 83845 112505 83879
rect 112505 83845 112539 83879
rect 112539 83845 112548 83879
rect 112496 83836 112548 83845
rect 113876 83836 113928 83888
rect 115164 83879 115216 83888
rect 99524 83768 99576 83820
rect 100904 83768 100956 83820
rect 102284 83768 102336 83820
rect 103664 83768 103716 83820
rect 105044 83768 105096 83820
rect 106424 83768 106476 83820
rect 107804 83768 107856 83820
rect 112956 83768 113008 83820
rect 115164 83845 115173 83879
rect 115173 83845 115207 83879
rect 115207 83845 115216 83879
rect 115164 83836 115216 83845
rect 96396 83700 96448 83752
rect 97776 83700 97828 83752
rect 113968 83700 114020 83752
rect 117924 83879 117976 83888
rect 117924 83845 117933 83879
rect 117933 83845 117967 83879
rect 117967 83845 117976 83879
rect 117924 83836 117976 83845
rect 119212 83836 119264 83888
rect 121972 83836 122024 83888
rect 123260 83879 123312 83888
rect 123260 83845 123269 83879
rect 123269 83845 123303 83879
rect 123303 83845 123312 83879
rect 123260 83836 123312 83845
rect 126020 83879 126072 83888
rect 126020 83845 126029 83879
rect 126029 83845 126063 83879
rect 126063 83845 126072 83879
rect 126020 83836 126072 83845
rect 128688 83879 128740 83888
rect 128688 83845 128697 83879
rect 128697 83845 128731 83879
rect 128731 83845 128740 83879
rect 128688 83836 128740 83845
rect 132736 83836 132788 83888
rect 300360 84244 300412 84296
rect 250496 83836 250548 83888
rect 251140 83836 251192 83888
rect 125560 83768 125612 83820
rect 133380 83768 133432 83820
rect 182140 83768 182192 83820
rect 116636 83700 116688 83752
rect 119304 83700 119356 83752
rect 85080 81932 85132 81984
rect 179564 81932 179616 81984
rect 186280 81932 186332 81984
rect 194100 81932 194152 81984
rect 203852 81932 203904 81984
rect 99616 81864 99668 81916
rect 133380 81864 133432 81916
rect 226760 81864 226812 81916
rect 89220 81796 89272 81848
rect 79560 81728 79612 81780
rect 79744 81660 79796 81712
rect 174044 81728 174096 81780
rect 197044 81728 197096 81780
rect 197504 81728 197556 81780
rect 198424 81728 198476 81780
rect 198884 81728 198936 81780
rect 199804 81728 199856 81780
rect 200264 81728 200316 81780
rect 201092 81728 201144 81780
rect 201644 81728 201696 81780
rect 173768 81660 173820 81712
rect 209188 81660 209240 81712
rect 79836 81592 79888 81644
rect 173492 81592 173544 81644
rect 211948 81592 212000 81644
rect 79652 81524 79704 81576
rect 173860 81524 173912 81576
rect 214616 81524 214668 81576
rect 79928 81456 79980 81508
rect 173676 81456 173728 81508
rect 217284 81456 217336 81508
rect 80020 81388 80072 81440
rect 173952 81388 174004 81440
rect 220044 81388 220096 81440
rect 221332 81388 221384 81440
rect 264848 81388 264900 81440
rect 80112 81320 80164 81372
rect 173308 81320 173360 81372
rect 222712 81320 222764 81372
rect 80204 81252 80256 81304
rect 173584 81252 173636 81304
rect 206520 81252 206572 81304
rect 207900 81252 207952 81304
rect 264756 81252 264808 81304
rect 99616 81184 99668 81236
rect 100260 81184 100312 81236
rect 187660 81184 187712 81236
rect 195572 81184 195624 81236
rect 101732 81116 101784 81168
rect 188948 81116 189000 81168
rect 195480 81116 195532 81168
rect 101640 80708 101692 80760
rect 182232 80640 182284 80692
rect 185820 80640 185872 80692
rect 180852 80572 180904 80624
rect 183060 80572 183112 80624
rect 184900 80572 184952 80624
rect 191340 80572 191392 80624
rect 134760 80504 134812 80556
rect 167236 80504 167288 80556
rect 111208 80139 111260 80148
rect 111208 80105 111217 80139
rect 111217 80105 111251 80139
rect 111251 80105 111260 80139
rect 111208 80096 111260 80105
rect 124732 80139 124784 80148
rect 124732 80105 124741 80139
rect 124741 80105 124775 80139
rect 124775 80105 124784 80139
rect 124732 80096 124784 80105
rect 167236 79756 167288 79808
rect 170180 79756 170232 79808
rect 155736 79416 155788 79468
rect 145340 79348 145392 79400
rect 145984 79348 146036 79400
rect 257028 79348 257080 79400
rect 257488 79348 257540 79400
rect 155368 79280 155420 79332
rect 155644 79212 155696 79264
rect 50488 79144 50540 79196
rect 51224 79144 51276 79196
rect 51776 79144 51828 79196
rect 52512 79144 52564 79196
rect 56468 79144 56520 79196
rect 54444 79008 54496 79060
rect 61896 79008 61948 79060
rect 62448 79144 62500 79196
rect 63644 79144 63696 79196
rect 138992 79144 139044 79196
rect 143224 79144 143276 79196
rect 158404 79144 158456 79196
rect 162636 79144 162688 79196
rect 231360 79144 231412 79196
rect 237616 79144 237668 79196
rect 238260 79144 238312 79196
rect 239732 79144 239784 79196
rect 241572 79144 241624 79196
rect 245160 79144 245212 79196
rect 246448 79144 246500 79196
rect 247000 79144 247052 79196
rect 249760 79144 249812 79196
rect 255556 79144 255608 79196
rect 256384 79144 256436 79196
rect 258684 79144 258736 79196
rect 264296 79144 264348 79196
rect 265124 79144 265176 79196
rect 137520 79076 137572 79128
rect 142764 79076 142816 79128
rect 65760 79008 65812 79060
rect 141660 79008 141712 79060
rect 144328 79076 144380 79128
rect 158312 79076 158364 79128
rect 162084 79076 162136 79128
rect 242492 79076 242544 79128
rect 247828 79076 247880 79128
rect 249208 79076 249260 79128
rect 255832 79076 255884 79128
rect 256292 79076 256344 79128
rect 143040 79008 143092 79060
rect 145248 79008 145300 79060
rect 153988 79008 154040 79060
rect 159784 79008 159836 79060
rect 167972 79008 168024 79060
rect 236880 79008 236932 79060
rect 239180 79008 239232 79060
rect 244424 79008 244476 79060
rect 249300 79008 249352 79060
rect 255740 79008 255792 79060
rect 256384 79008 256436 79060
rect 256568 79076 256620 79128
rect 259236 79076 259288 79128
rect 260340 79008 260392 79060
rect 60516 78940 60568 78992
rect 64472 78940 64524 78992
rect 140280 78940 140332 78992
rect 143776 78940 143828 78992
rect 151412 78940 151464 78992
rect 157116 78940 157168 78992
rect 158220 78940 158272 78992
rect 163188 78940 163240 78992
rect 246908 78940 246960 78992
rect 247184 78940 247236 78992
rect 248104 78940 248156 78992
rect 253440 78940 253492 78992
rect 256200 78940 256252 78992
rect 256568 78940 256620 78992
rect 59136 78872 59188 78924
rect 61712 78804 61764 78856
rect 66496 78804 66548 78856
rect 67140 78872 67192 78924
rect 68428 78872 68480 78924
rect 157024 78872 157076 78924
rect 164752 78872 164804 78924
rect 232740 78872 232792 78924
rect 240744 78872 240796 78924
rect 244148 78872 244200 78924
rect 249392 78872 249444 78924
rect 68060 78804 68112 78856
rect 69900 78804 69952 78856
rect 73120 78804 73172 78856
rect 156932 78804 156984 78856
rect 165304 78804 165356 78856
rect 61804 78736 61856 78788
rect 67140 78736 67192 78788
rect 147640 78736 147692 78788
rect 151320 78736 151372 78788
rect 154724 78736 154776 78788
rect 164568 78736 164620 78788
rect 243044 78736 243096 78788
rect 247920 78736 247972 78788
rect 255648 78736 255700 78788
rect 61620 78668 61672 78720
rect 67784 78668 67836 78720
rect 166408 78668 166460 78720
rect 247000 78668 247052 78720
rect 253532 78668 253584 78720
rect 61988 78600 62040 78652
rect 68244 78600 68296 78652
rect 151964 78600 152016 78652
rect 161716 78600 161768 78652
rect 243596 78600 243648 78652
rect 249576 78600 249628 78652
rect 251232 78600 251284 78652
rect 263100 78600 263152 78652
rect 55180 78532 55232 78584
rect 38252 78464 38304 78516
rect 49200 78464 49252 78516
rect 53156 78464 53208 78516
rect 60332 78532 60384 78584
rect 63828 78532 63880 78584
rect 151780 78532 151832 78584
rect 157208 78532 157260 78584
rect 157300 78532 157352 78584
rect 167420 78532 167472 78584
rect 248472 78532 248524 78584
rect 249484 78532 249536 78584
rect 254728 78532 254780 78584
rect 63552 78464 63604 78516
rect 75788 78464 75840 78516
rect 138900 78464 138952 78516
rect 146536 78464 146588 78516
rect 150492 78464 150544 78516
rect 60424 78396 60476 78448
rect 65116 78396 65168 78448
rect 67968 78396 68020 78448
rect 156656 78464 156708 78516
rect 163740 78464 163792 78516
rect 234120 78464 234172 78516
rect 237984 78464 238036 78516
rect 251140 78464 251192 78516
rect 262548 78464 262600 78516
rect 264480 78464 264532 78516
rect 295576 78464 295628 78516
rect 158312 78396 158364 78448
rect 161072 78396 161124 78448
rect 248288 78396 248340 78448
rect 254176 78396 254228 78448
rect 67416 78328 67468 78380
rect 69808 78328 69860 78380
rect 144420 78328 144472 78380
rect 145432 78328 145484 78380
rect 150492 78328 150544 78380
rect 155736 78328 155788 78380
rect 155828 78328 155880 78380
rect 165856 78328 165908 78380
rect 235500 78328 235552 78380
rect 238536 78328 238588 78380
rect 248012 78328 248064 78380
rect 253072 78328 253124 78380
rect 149756 78260 149808 78312
rect 155368 78260 155420 78312
rect 155644 78260 155696 78312
rect 160336 78260 160388 78312
rect 248196 78260 248248 78312
rect 253624 78260 253676 78312
rect 58492 78192 58544 78244
rect 60424 78192 60476 78244
rect 65208 78192 65260 78244
rect 67232 78192 67284 78244
rect 69164 78192 69216 78244
rect 148744 78192 148796 78244
rect 154080 78192 154132 78244
rect 157668 78192 157720 78244
rect 158864 78192 158916 78244
rect 245344 78192 245396 78244
rect 250772 78192 250824 78244
rect 55824 78124 55876 78176
rect 65852 78124 65904 78176
rect 149204 78124 149256 78176
rect 154172 78124 154224 78176
rect 155092 78124 155144 78176
rect 156104 78124 156156 78176
rect 245804 78124 245856 78176
rect 250680 78124 250732 78176
rect 57848 78056 57900 78108
rect 65760 78056 65812 78108
rect 67324 78056 67376 78108
rect 70452 78056 70504 78108
rect 153160 78056 153212 78108
rect 232832 78056 232884 78108
rect 236880 78056 236932 78108
rect 239640 78056 239692 78108
rect 240376 78056 240428 78108
rect 248380 78056 248432 78108
rect 252796 78124 252848 78176
rect 252060 78056 252112 78108
rect 252704 78056 252756 78108
rect 59780 77988 59832 78040
rect 67508 77988 67560 78040
rect 153068 77988 153120 78040
rect 159692 77988 159744 78040
rect 56100 77920 56152 77972
rect 63184 77920 63236 77972
rect 148192 77920 148244 77972
rect 152700 77920 152752 77972
rect 154632 77920 154684 77972
rect 160888 77920 160940 77972
rect 57112 77852 57164 77904
rect 64380 77852 64432 77904
rect 150400 77852 150452 77904
rect 150584 77852 150636 77904
rect 152516 77852 152568 77904
rect 153344 77852 153396 77904
rect 155184 77852 155236 77904
rect 156012 77852 156064 77904
rect 156840 77852 156892 77904
rect 157392 77852 157444 77904
rect 159600 77852 159652 77904
rect 155460 77784 155512 77836
rect 160980 77784 161032 77836
rect 89772 77691 89824 77700
rect 89772 77657 89781 77691
rect 89781 77657 89815 77691
rect 89815 77657 89824 77691
rect 89772 77648 89824 77657
rect 124732 76356 124784 76408
rect 169996 76356 170048 76408
rect 218664 76356 218716 76408
rect 233476 76356 233528 76408
rect 119304 76288 119356 76340
rect 139636 76288 139688 76340
rect 111208 74996 111260 75048
rect 170732 74996 170784 75048
rect 205140 74996 205192 75048
rect 233660 74996 233712 75048
rect 113968 74928 114020 74980
rect 170824 74928 170876 74980
rect 213236 74928 213288 74980
rect 233568 74928 233620 74980
rect 116636 74860 116688 74912
rect 170640 74860 170692 74912
rect 215996 74860 216048 74912
rect 233476 74860 233528 74912
rect 138072 73704 138124 73756
rect 139636 73704 139688 73756
rect 100260 73636 100312 73688
rect 100996 73636 101048 73688
rect 183704 73636 183756 73688
rect 190144 73636 190196 73688
rect 190604 73636 190656 73688
rect 96396 73500 96448 73552
rect 108264 73500 108316 73552
rect 202656 73500 202708 73552
rect 97776 73432 97828 73484
rect 110748 73432 110800 73484
rect 191984 73432 192036 73484
rect 205140 73432 205192 73484
rect 100904 73364 100956 73416
rect 115716 73364 115768 73416
rect 193364 73364 193416 73416
rect 207624 73364 207676 73416
rect 99524 73296 99576 73348
rect 113416 73296 113468 73348
rect 194744 73296 194796 73348
rect 210108 73296 210160 73348
rect 102284 73228 102336 73280
rect 118292 73228 118344 73280
rect 196124 73228 196176 73280
rect 212684 73228 212736 73280
rect 103664 73160 103716 73212
rect 120776 73160 120828 73212
rect 197504 73160 197556 73212
rect 215168 73160 215220 73212
rect 105044 73092 105096 73144
rect 123260 73092 123312 73144
rect 198884 73092 198936 73144
rect 217652 73092 217704 73144
rect 106424 73024 106476 73076
rect 125836 73024 125888 73076
rect 200264 73024 200316 73076
rect 220136 73024 220188 73076
rect 107804 72956 107856 73008
rect 128596 72956 128648 73008
rect 201644 72956 201696 73008
rect 222620 72956 222672 73008
rect 89772 72888 89824 72940
rect 95752 72888 95804 72940
rect 96120 72888 96172 72940
rect 98236 72888 98288 72940
rect 101640 72684 101692 72736
rect 105780 72684 105832 72736
rect 91980 72616 92032 72668
rect 93268 72616 93320 72668
rect 101732 72616 101784 72668
rect 103204 72616 103256 72668
rect 136508 72412 136560 72464
rect 139728 72412 139780 72464
rect 195480 72412 195532 72464
rect 200172 72412 200224 72464
rect 89220 72344 89272 72396
rect 90784 72344 90836 72396
rect 136784 72344 136836 72396
rect 139636 72344 139688 72396
rect 183060 72344 183112 72396
rect 184716 72344 184768 72396
rect 185820 72344 185872 72396
rect 187660 72344 187712 72396
rect 191340 72344 191392 72396
rect 192628 72344 192680 72396
rect 194100 72344 194152 72396
rect 195112 72344 195164 72396
rect 195572 72344 195624 72396
rect 197504 72344 197556 72396
rect 230624 72344 230676 72396
rect 233476 72344 233528 72396
rect 80204 70916 80256 70968
rect 84436 70916 84488 70968
rect 135956 70916 136008 70968
rect 139636 70916 139688 70968
rect 131356 70848 131408 70900
rect 138072 70848 138124 70900
rect 226024 70848 226076 70900
rect 230624 70848 230676 70900
rect 276164 70848 276216 70900
rect 300176 70848 300228 70900
rect 84436 70236 84488 70288
rect 87196 70236 87248 70288
rect 136416 69692 136468 69744
rect 139820 69692 139872 69744
rect 229888 69692 229940 69744
rect 233660 69692 233712 69744
rect 79468 69624 79520 69676
rect 80204 69556 80256 69608
rect 136600 69624 136652 69676
rect 139728 69624 139780 69676
rect 136692 69556 136744 69608
rect 139636 69556 139688 69608
rect 87196 69488 87248 69540
rect 131540 69488 131592 69540
rect 135956 69488 136008 69540
rect 173308 69488 173360 69540
rect 181772 69488 181824 69540
rect 226024 69488 226076 69540
rect 233568 69488 233620 69540
rect 87288 69420 87340 69472
rect 131356 69420 131408 69472
rect 136508 69420 136560 69472
rect 225748 69420 225800 69472
rect 233476 69420 233528 69472
rect 131448 69352 131500 69404
rect 136784 69352 136836 69404
rect 80204 68808 80256 68860
rect 87196 68808 87248 68860
rect 172848 68808 172900 68860
rect 182324 68808 182376 68860
rect 226300 68740 226352 68792
rect 229888 68740 229940 68792
rect 80112 68264 80164 68316
rect 80204 68196 80256 68248
rect 136508 68264 136560 68316
rect 139728 68264 139780 68316
rect 136784 68196 136836 68248
rect 139636 68196 139688 68248
rect 87196 68128 87248 68180
rect 132000 68128 132052 68180
rect 139912 68128 139964 68180
rect 174044 68128 174096 68180
rect 181772 68128 181824 68180
rect 225472 68128 225524 68180
rect 233568 68128 233620 68180
rect 87288 68060 87340 68112
rect 132552 68060 132604 68112
rect 136416 68060 136468 68112
rect 173952 68060 174004 68112
rect 181588 68060 181640 68112
rect 225564 68060 225616 68112
rect 233660 68060 233712 68112
rect 131816 67992 131868 68044
rect 136600 67992 136652 68044
rect 225840 67992 225892 68044
rect 233476 67992 233528 68044
rect 131356 67924 131408 67976
rect 136692 67924 136744 67976
rect 226300 67924 226352 67976
rect 233752 67924 233804 67976
rect 80204 67516 80256 67568
rect 87196 67516 87248 67568
rect 80112 67448 80164 67500
rect 87288 67448 87340 67500
rect 173492 67448 173544 67500
rect 182324 67448 182376 67500
rect 133012 66904 133064 66956
rect 139636 66904 139688 66956
rect 136692 66768 136744 66820
rect 139728 66768 139780 66820
rect 173860 66700 173912 66752
rect 181404 66700 181456 66752
rect 226300 66700 226352 66752
rect 233476 66700 233528 66752
rect 132184 66632 132236 66684
rect 136784 66632 136836 66684
rect 173584 66632 173636 66684
rect 182324 66632 182376 66684
rect 226024 66632 226076 66684
rect 233568 66632 233620 66684
rect 131356 66564 131408 66616
rect 136508 66564 136560 66616
rect 174044 66564 174096 66616
rect 182232 66564 182284 66616
rect 131356 66156 131408 66208
rect 133012 66156 133064 66208
rect 80204 66088 80256 66140
rect 87196 66088 87248 66140
rect 80112 66020 80164 66072
rect 87288 66020 87340 66072
rect 226392 66020 226444 66072
rect 233476 66020 233528 66072
rect 80204 65340 80256 65392
rect 87196 65340 87248 65392
rect 131816 65340 131868 65392
rect 139636 65340 139688 65392
rect 173492 65340 173544 65392
rect 182324 65340 182376 65392
rect 226300 65340 226352 65392
rect 233476 65340 233528 65392
rect 131448 65272 131500 65324
rect 139728 65272 139780 65324
rect 173768 65272 173820 65324
rect 181404 65272 181456 65324
rect 131356 65204 131408 65256
rect 136692 65204 136744 65256
rect 80112 64728 80164 64780
rect 87196 64728 87248 64780
rect 226300 64728 226352 64780
rect 233568 64728 233620 64780
rect 80204 64660 80256 64712
rect 87288 64660 87340 64712
rect 226392 64660 226444 64712
rect 233476 64660 233528 64712
rect 80204 63980 80256 64032
rect 87656 63980 87708 64032
rect 131356 63980 131408 64032
rect 139636 63980 139688 64032
rect 173860 63980 173912 64032
rect 181036 63980 181088 64032
rect 131816 63912 131868 63964
rect 139728 63912 139780 63964
rect 173952 63912 174004 63964
rect 181128 63912 181180 63964
rect 174044 63844 174096 63896
rect 181312 63844 181364 63896
rect 226300 63436 226352 63488
rect 233660 63436 233712 63488
rect 132000 63368 132052 63420
rect 139636 63368 139688 63420
rect 226392 63368 226444 63420
rect 233476 63368 233528 63420
rect 80204 63300 80256 63352
rect 87196 63300 87248 63352
rect 131356 63300 131408 63352
rect 139728 63300 139780 63352
rect 226300 63300 226352 63352
rect 233568 63300 233620 63352
rect 226300 62620 226352 62672
rect 233476 62620 233528 62672
rect 80204 62552 80256 62604
rect 87288 62552 87340 62604
rect 173768 62552 173820 62604
rect 182324 62552 182376 62604
rect 80112 62484 80164 62536
rect 87196 62484 87248 62536
rect 173308 62484 173360 62536
rect 181404 62484 181456 62536
rect 131448 61940 131500 61992
rect 139728 61940 139780 61992
rect 131356 61872 131408 61924
rect 139636 61872 139688 61924
rect 226392 61872 226444 61924
rect 233476 61872 233528 61924
rect 226208 61328 226260 61380
rect 233476 61328 233528 61380
rect 131356 61260 131408 61312
rect 80204 61192 80256 61244
rect 87288 61192 87340 61244
rect 226300 61260 226352 61312
rect 233568 61260 233620 61312
rect 139636 61192 139688 61244
rect 173676 61192 173728 61244
rect 182232 61192 182284 61244
rect 80112 61124 80164 61176
rect 87196 61124 87248 61176
rect 174044 61124 174096 61176
rect 182140 61124 182192 61176
rect 173952 61056 174004 61108
rect 182048 61056 182100 61108
rect 131356 60580 131408 60632
rect 139728 60580 139780 60632
rect 131448 60512 131500 60564
rect 139636 60512 139688 60564
rect 79100 60308 79152 60360
rect 87012 60308 87064 60360
rect 226392 60104 226444 60156
rect 233752 60104 233804 60156
rect 226300 60036 226352 60088
rect 233844 60036 233896 60088
rect 131816 59968 131868 60020
rect 137244 59968 137296 60020
rect 176896 59968 176948 60020
rect 182232 59968 182284 60020
rect 225748 59968 225800 60020
rect 233476 59968 233528 60020
rect 131356 59900 131408 59952
rect 80112 59832 80164 59884
rect 87196 59832 87248 59884
rect 176988 59900 177040 59952
rect 182324 59900 182376 59952
rect 225932 59900 225984 59952
rect 233568 59900 233620 59952
rect 139636 59832 139688 59884
rect 173860 59832 173912 59884
rect 181956 59832 182008 59884
rect 80204 59764 80256 59816
rect 87104 59764 87156 59816
rect 173676 59764 173728 59816
rect 181864 59764 181916 59816
rect 174044 59696 174096 59748
rect 181772 59696 181824 59748
rect 137244 59220 137296 59272
rect 139728 59220 139780 59272
rect 139820 58744 139872 58796
rect 131540 58676 131592 58728
rect 131448 58608 131500 58660
rect 80020 58540 80072 58592
rect 87196 58540 87248 58592
rect 131356 58540 131408 58592
rect 80112 58472 80164 58524
rect 87012 58472 87064 58524
rect 80204 58404 80256 58456
rect 86920 58404 86972 58456
rect 226208 58676 226260 58728
rect 233476 58676 233528 58728
rect 226392 58608 226444 58660
rect 233568 58608 233620 58660
rect 226300 58540 226352 58592
rect 233660 58540 233712 58592
rect 139636 58472 139688 58524
rect 173768 58472 173820 58524
rect 182140 58472 182192 58524
rect 139728 58404 139780 58456
rect 174044 58404 174096 58456
rect 181680 58404 181732 58456
rect 178000 57656 178052 57708
rect 182324 57656 182376 57708
rect 177632 57520 177684 57572
rect 181680 57520 181732 57572
rect 80204 57316 80256 57368
rect 86828 57316 86880 57368
rect 131356 57316 131408 57368
rect 136232 57316 136284 57368
rect 131540 57248 131592 57300
rect 137336 57248 137388 57300
rect 131448 57180 131500 57232
rect 139912 57316 139964 57368
rect 225748 57316 225800 57368
rect 228048 57316 228100 57368
rect 177724 57248 177776 57300
rect 181588 57248 181640 57300
rect 225840 57248 225892 57300
rect 228600 57248 228652 57300
rect 226484 57180 226536 57232
rect 228692 57180 228744 57232
rect 131632 57112 131684 57164
rect 139728 57112 139780 57164
rect 225932 57112 225984 57164
rect 227956 57112 228008 57164
rect 80112 57044 80164 57096
rect 87288 57044 87340 57096
rect 172940 57044 172992 57096
rect 180944 57044 180996 57096
rect 80204 56976 80256 57028
rect 87380 56976 87432 57028
rect 174044 56976 174096 57028
rect 176896 56976 176948 57028
rect 174044 56772 174096 56824
rect 176988 56772 177040 56824
rect 137336 56568 137388 56620
rect 139636 56568 139688 56620
rect 226300 56160 226352 56212
rect 229428 56160 229480 56212
rect 131448 55888 131500 55940
rect 138072 55888 138124 55940
rect 226300 55888 226352 55940
rect 229336 55888 229388 55940
rect 131356 55820 131408 55872
rect 139452 55820 139504 55872
rect 131540 55752 131592 55804
rect 139544 55752 139596 55804
rect 177356 55752 177408 55804
rect 182324 55752 182376 55804
rect 225932 55752 225984 55804
rect 229612 55752 229664 55804
rect 80112 55684 80164 55736
rect 87104 55684 87156 55736
rect 173308 55684 173360 55736
rect 182232 55684 182284 55736
rect 227956 55684 228008 55736
rect 233568 55684 233620 55736
rect 173768 55616 173820 55668
rect 182048 55616 182100 55668
rect 228048 55616 228100 55668
rect 233476 55616 233528 55668
rect 80204 55412 80256 55464
rect 87012 55412 87064 55464
rect 226300 54664 226352 54716
rect 229520 54664 229572 54716
rect 79744 54528 79796 54580
rect 87288 54528 87340 54580
rect 131356 54528 131408 54580
rect 136784 54528 136836 54580
rect 79468 54460 79520 54512
rect 87196 54460 87248 54512
rect 131448 54460 131500 54512
rect 139912 54460 139964 54512
rect 175240 54460 175292 54512
rect 181680 54460 181732 54512
rect 225748 54460 225800 54512
rect 230900 54460 230952 54512
rect 85908 54392 85960 54444
rect 87288 54392 87340 54444
rect 131540 54392 131592 54444
rect 139636 54392 139688 54444
rect 175332 54392 175384 54444
rect 181588 54392 181640 54444
rect 226392 54392 226444 54444
rect 230716 54392 230768 54444
rect 174044 54324 174096 54376
rect 178000 54324 178052 54376
rect 228600 54324 228652 54376
rect 233476 54324 233528 54376
rect 228692 54256 228744 54308
rect 233568 54256 233620 54308
rect 80204 54188 80256 54240
rect 86736 54188 86788 54240
rect 136232 54188 136284 54240
rect 139728 54188 139780 54240
rect 226300 54188 226352 54240
rect 231728 54188 231780 54240
rect 138072 53916 138124 53968
rect 140004 53916 140056 53968
rect 174044 53780 174096 53832
rect 177632 53780 177684 53832
rect 173492 53712 173544 53764
rect 177724 53712 177776 53764
rect 80204 53304 80256 53356
rect 86552 53304 86604 53356
rect 131448 53032 131500 53084
rect 139728 53032 139780 53084
rect 80020 52964 80072 53016
rect 87196 52964 87248 53016
rect 131356 52964 131408 53016
rect 139820 52964 139872 53016
rect 176896 52964 176948 53016
rect 182324 52964 182376 53016
rect 225840 52964 225892 53016
rect 233568 52964 233620 53016
rect 80112 52896 80164 52948
rect 88392 52896 88444 52948
rect 172848 52896 172900 52948
rect 181220 52896 181272 52948
rect 229612 52896 229664 52948
rect 233476 52896 233528 52948
rect 80204 52828 80256 52880
rect 88208 52828 88260 52880
rect 174044 52828 174096 52880
rect 181312 52828 181364 52880
rect 229428 52828 229480 52880
rect 233660 52828 233712 52880
rect 229336 52760 229388 52812
rect 233476 52760 233528 52812
rect 173952 52692 174004 52744
rect 180300 52692 180352 52744
rect 80204 51536 80256 51588
rect 87932 51536 87984 51588
rect 173952 51536 174004 51588
rect 181128 51536 181180 51588
rect 198792 51536 198844 51588
rect 230900 51536 230952 51588
rect 233476 51536 233528 51588
rect 234120 51468 234172 51520
rect 230716 51400 230768 51452
rect 233660 51400 233712 51452
rect 172940 51196 172992 51248
rect 177356 51196 177408 51248
rect 125192 50924 125244 50976
rect 127032 50924 127084 50976
rect 134760 50924 134812 50976
rect 115164 50856 115216 50908
rect 128596 50856 128648 50908
rect 208820 50856 208872 50908
rect 222436 50856 222488 50908
rect 94004 50652 94056 50704
rect 94556 50652 94608 50704
rect 218848 50380 218900 50432
rect 220964 50380 221016 50432
rect 187844 50244 187896 50296
rect 188856 50244 188908 50296
rect 136784 50176 136836 50228
rect 139636 50176 139688 50228
rect 231728 50176 231780 50228
rect 233476 50176 233528 50228
rect 173308 50108 173360 50160
rect 175240 50108 175292 50160
rect 229520 50108 229572 50160
rect 233660 50108 233712 50160
rect 172756 50040 172808 50092
rect 175332 50040 175384 50092
rect 80204 49224 80256 49276
rect 87104 49224 87156 49276
rect 173124 49156 173176 49208
rect 176896 49156 176948 49208
rect 80112 48884 80164 48936
rect 85908 48884 85960 48936
rect 173308 48612 173360 48664
rect 180944 48612 180996 48664
rect 99524 47456 99576 47508
rect 139636 47456 139688 47508
rect 193364 47456 193416 47508
rect 233476 47456 233528 47508
rect 220964 47388 221016 47440
rect 228140 47388 228192 47440
rect 260432 47388 260484 47440
rect 62908 46028 62960 46080
rect 63644 46028 63696 46080
rect 276072 46028 276124 46080
rect 300176 46028 300228 46080
rect 260432 45348 260484 45400
rect 284536 45348 284588 45400
rect 93084 37732 93136 37784
rect 94004 37732 94056 37784
rect 98788 37732 98840 37784
rect 99524 37732 99576 37784
rect 192444 37732 192496 37784
rect 193364 37732 193416 37784
rect 186740 37392 186792 37444
rect 187844 37392 187896 37444
rect 79560 37188 79612 37240
rect 103848 37188 103900 37240
rect 173400 37188 173452 37240
rect 198148 37188 198200 37240
rect 13504 37120 13556 37172
rect 120960 37120 121012 37172
rect 140924 37120 140976 37172
rect 203852 37120 203904 37172
rect 209556 37120 209608 37172
rect 292632 37120 292684 37172
rect 63644 37052 63696 37104
rect 109552 37052 109604 37104
rect 115808 37052 115860 37104
rect 292540 37052 292592 37104
rect 128872 28008 128924 28060
rect 129516 28008 129568 28060
rect 222804 28008 222856 28060
rect 223540 28008 223592 28060
rect 13320 25356 13372 25408
rect 85080 25356 85132 25408
rect 76524 20868 76576 20920
rect 299808 20868 299860 20920
rect 13596 17060 13648 17112
rect 109552 17060 109604 17112
rect 203852 17060 203904 17112
rect 265860 17060 265912 17112
rect 38160 12436 38212 12488
rect 138440 12436 138492 12488
rect 28224 12368 28276 12420
rect 133380 12368 133432 12420
rect 88484 12300 88536 12352
rect 248748 12300 248800 12352
rect 64932 12232 64984 12284
rect 264664 12232 264716 12284
rect 175240 9376 175292 9428
rect 175424 9376 175476 9428
rect 284536 9376 284588 9428
rect 285456 9376 285508 9428
<< metal2 >>
rect 28222 302344 28278 302824
rect 64930 302344 64986 302824
rect 101730 302344 101786 302824
rect 138438 302344 138494 302824
rect 175238 302344 175294 302824
rect 211946 302344 212002 302824
rect 248746 302344 248802 302824
rect 285454 302344 285510 302824
rect 28236 298706 28264 302344
rect 64944 302258 64972 302344
rect 64944 302230 65064 302258
rect 34664 299448 34716 299454
rect 34664 299390 34716 299396
rect 34572 299312 34624 299318
rect 34572 299254 34624 299260
rect 28224 298700 28276 298706
rect 28224 298642 28276 298648
rect 29144 298700 29196 298706
rect 29144 298642 29196 298648
rect 13412 294620 13464 294626
rect 13412 294562 13464 294568
rect 13318 287856 13374 287865
rect 13318 287791 13374 287800
rect 13226 286496 13282 286505
rect 13226 286431 13282 286440
rect 13240 286262 13268 286431
rect 13228 286256 13280 286262
rect 13228 286198 13280 286204
rect 12950 221216 13006 221225
rect 12950 221151 13006 221160
rect 12964 220030 12992 221151
rect 12952 220024 13004 220030
rect 12952 219966 13004 219972
rect 13332 57889 13360 287791
rect 13424 123169 13452 294562
rect 20220 286256 20272 286262
rect 20220 286198 20272 286204
rect 13686 253856 13742 253865
rect 13686 253791 13742 253800
rect 13502 188576 13558 188585
rect 13502 188511 13558 188520
rect 13410 123160 13466 123169
rect 13410 123095 13466 123104
rect 13318 57880 13374 57889
rect 13318 57815 13374 57824
rect 13516 37178 13544 188511
rect 13594 155800 13650 155809
rect 13594 155735 13650 155744
rect 13504 37172 13556 37178
rect 13504 37114 13556 37120
rect 13320 25408 13372 25414
rect 13320 25350 13372 25356
rect 13332 25249 13360 25350
rect 13318 25240 13374 25249
rect 13318 25175 13374 25184
rect 13608 17118 13636 155735
rect 13700 131601 13728 253791
rect 18840 220024 18892 220030
rect 18840 219966 18892 219972
rect 18852 181338 18880 219966
rect 18840 181332 18892 181338
rect 18840 181274 18892 181280
rect 20232 181134 20260 286198
rect 29156 224858 29184 298642
rect 29144 224852 29196 224858
rect 29144 224794 29196 224800
rect 31628 224852 31680 224858
rect 31628 224794 31680 224800
rect 24174 224208 24230 224217
rect 24174 224143 24230 224152
rect 24188 222698 24216 224143
rect 31640 222834 31668 224794
rect 31640 222806 31930 222834
rect 23926 222670 24216 222698
rect 23728 182822 23926 182850
rect 31640 182822 31930 182850
rect 23728 181338 23756 182822
rect 31640 181338 31668 182822
rect 23716 181332 23768 181338
rect 23716 181274 23768 181280
rect 31628 181332 31680 181338
rect 31628 181274 31680 181280
rect 20220 181128 20272 181134
rect 20220 181070 20272 181076
rect 13686 131592 13742 131601
rect 13686 131527 13742 131536
rect 23898 130368 23954 130377
rect 13780 130332 13832 130338
rect 23898 130303 23954 130312
rect 31904 130332 31956 130338
rect 13780 130274 13832 130280
rect 13792 90529 13820 130274
rect 23912 128708 23940 130303
rect 31904 130274 31956 130280
rect 31916 128708 31944 130274
rect 13778 90520 13834 90529
rect 13778 90455 13834 90464
rect 23912 87498 23940 88860
rect 31916 87498 31944 88860
rect 34584 87498 34612 299254
rect 23900 87492 23952 87498
rect 23900 87434 23952 87440
rect 31904 87492 31956 87498
rect 31904 87434 31956 87440
rect 34572 87492 34624 87498
rect 34572 87434 34624 87440
rect 34676 87362 34704 299390
rect 65036 295170 65064 302230
rect 101744 299386 101772 302344
rect 101732 299380 101784 299386
rect 101732 299322 101784 299328
rect 138452 298706 138480 302344
rect 175252 302258 175280 302344
rect 175252 302230 175464 302258
rect 138440 298700 138492 298706
rect 138440 298642 138492 298648
rect 139544 298700 139596 298706
rect 139544 298642 139596 298648
rect 139556 295170 139584 298642
rect 65024 295164 65076 295170
rect 65024 295106 65076 295112
rect 96212 295164 96264 295170
rect 96212 295106 96264 295112
rect 139544 295164 139596 295170
rect 139544 295106 139596 295112
rect 96224 292738 96252 295106
rect 123536 294688 123588 294694
rect 123536 294630 123588 294636
rect 110196 294552 110248 294558
rect 110196 294494 110248 294500
rect 110208 292738 110236 294494
rect 123548 292738 123576 294630
rect 96224 292710 96560 292738
rect 109900 292710 110236 292738
rect 123240 292710 123576 292738
rect 175436 286210 175464 302230
rect 211960 299454 211988 302344
rect 248760 299454 248788 302344
rect 211948 299448 212000 299454
rect 211948 299390 212000 299396
rect 248748 299448 248800 299454
rect 248748 299390 248800 299396
rect 267240 299448 267292 299454
rect 267240 299390 267292 299396
rect 203852 295164 203904 295170
rect 203852 295106 203904 295112
rect 190512 294620 190564 294626
rect 190512 294562 190564 294568
rect 190524 292724 190552 294562
rect 203864 292724 203892 295106
rect 264756 294688 264808 294694
rect 264756 294630 264808 294636
rect 217192 294620 217244 294626
rect 217192 294562 217244 294568
rect 217204 292724 217232 294562
rect 175252 286182 175464 286210
rect 88482 284864 88538 284873
rect 88482 284799 88538 284808
rect 79560 274492 79612 274498
rect 79560 274434 79612 274440
rect 62906 265552 62962 265561
rect 62906 265487 62962 265496
rect 62920 263756 62948 265487
rect 78916 264088 78968 264094
rect 78916 264030 78968 264036
rect 78928 263793 78956 264030
rect 78914 263784 78970 263793
rect 78914 263719 78970 263728
rect 79572 263385 79600 274434
rect 79558 263376 79614 263385
rect 79558 263311 79614 263320
rect 47084 262660 47136 262666
rect 47084 262602 47136 262608
rect 47096 249921 47124 262602
rect 80110 262152 80166 262161
rect 80110 262087 80166 262096
rect 80124 261510 80152 262087
rect 80112 261504 80164 261510
rect 87196 261504 87248 261510
rect 80112 261446 80164 261452
rect 80202 261472 80258 261481
rect 87196 261446 87248 261452
rect 80202 261407 80204 261416
rect 80256 261407 80258 261416
rect 80204 261378 80256 261384
rect 80110 260792 80166 260801
rect 80110 260727 80166 260736
rect 80124 260218 80152 260727
rect 80112 260212 80164 260218
rect 80112 260154 80164 260160
rect 85172 260212 85224 260218
rect 85172 260154 85224 260160
rect 80204 260144 80256 260150
rect 80202 260112 80204 260121
rect 85080 260144 85132 260150
rect 80256 260112 80258 260121
rect 85080 260086 85132 260092
rect 80202 260047 80258 260056
rect 79834 259432 79890 259441
rect 79834 259367 79890 259376
rect 79848 258654 79876 259367
rect 80202 258752 80258 258761
rect 80202 258687 80204 258696
rect 80256 258687 80258 258696
rect 84436 258716 84488 258722
rect 80204 258658 80256 258664
rect 84436 258658 84488 258664
rect 79836 258648 79888 258654
rect 79836 258590 79888 258596
rect 82412 258648 82464 258654
rect 82412 258590 82464 258596
rect 80018 258072 80074 258081
rect 80018 258007 80074 258016
rect 80032 257702 80060 258007
rect 80020 257696 80072 257702
rect 80020 257638 80072 257644
rect 82320 257696 82372 257702
rect 82320 257638 82372 257644
rect 80202 257392 80258 257401
rect 80202 257327 80258 257336
rect 80216 257294 80244 257327
rect 80204 257288 80256 257294
rect 80204 257230 80256 257236
rect 81676 257288 81728 257294
rect 81676 257230 81728 257236
rect 80110 256848 80166 256857
rect 80110 256783 80166 256792
rect 80124 256002 80152 256783
rect 80202 256168 80258 256177
rect 80202 256103 80258 256112
rect 80112 255996 80164 256002
rect 80112 255938 80164 255944
rect 80216 255934 80244 256103
rect 80204 255928 80256 255934
rect 80204 255870 80256 255876
rect 81688 255798 81716 257230
rect 82136 255996 82188 256002
rect 82136 255938 82188 255944
rect 81768 255928 81820 255934
rect 81768 255870 81820 255876
rect 81676 255792 81728 255798
rect 81676 255734 81728 255740
rect 80110 255488 80166 255497
rect 80110 255423 80166 255432
rect 80124 254642 80152 255423
rect 80202 254808 80258 254817
rect 80202 254743 80258 254752
rect 80112 254636 80164 254642
rect 80112 254578 80164 254584
rect 80216 254506 80244 254743
rect 80204 254500 80256 254506
rect 80204 254442 80256 254448
rect 81780 254370 81808 255870
rect 81768 254364 81820 254370
rect 81768 254306 81820 254312
rect 82148 254234 82176 255938
rect 82332 255866 82360 257638
rect 82424 257226 82452 258590
rect 82412 257220 82464 257226
rect 82412 257162 82464 257168
rect 82320 255860 82372 255866
rect 82320 255802 82372 255808
rect 84448 255730 84476 258658
rect 85092 256818 85120 260086
rect 85184 257022 85212 260154
rect 87208 258353 87236 261446
rect 87288 261436 87340 261442
rect 87288 261378 87340 261384
rect 87194 258344 87250 258353
rect 87194 258279 87250 258288
rect 87300 257537 87328 261378
rect 88496 258586 88524 284799
rect 131354 280784 131410 280793
rect 131354 280719 131410 280728
rect 94904 276934 95424 276962
rect 104840 276934 105084 276962
rect 95396 260694 95424 276934
rect 105056 262734 105084 276934
rect 114854 276690 114882 276948
rect 114808 276662 114882 276690
rect 124468 276934 124896 276962
rect 114808 274498 114836 276662
rect 114796 274492 114848 274498
rect 114796 274434 114848 274440
rect 124468 264094 124496 276934
rect 124456 264088 124508 264094
rect 124456 264030 124508 264036
rect 125744 264088 125796 264094
rect 125744 264030 125796 264036
rect 125756 263414 125784 264030
rect 125744 263408 125796 263414
rect 125744 263350 125796 263356
rect 105044 262728 105096 262734
rect 105044 262670 105096 262676
rect 131368 262666 131396 280719
rect 175252 276674 175280 286182
rect 182322 284864 182378 284873
rect 182322 284799 182378 284808
rect 175240 276668 175292 276674
rect 175240 276610 175292 276616
rect 173400 274492 173452 274498
rect 173400 274434 173452 274440
rect 143040 264088 143092 264094
rect 143040 264030 143092 264036
rect 139634 263512 139690 263521
rect 139634 263447 139690 263456
rect 139648 263414 139676 263447
rect 132736 263408 132788 263414
rect 132736 263350 132788 263356
rect 139636 263408 139688 263414
rect 139636 263350 139688 263356
rect 131356 262660 131408 262666
rect 131356 262602 131408 262608
rect 95384 260688 95436 260694
rect 95384 260630 95436 260636
rect 109552 260688 109604 260694
rect 109552 260630 109604 260636
rect 88484 258580 88536 258586
rect 88484 258522 88536 258528
rect 109564 257786 109592 260630
rect 129516 258580 129568 258586
rect 129516 258522 129568 258528
rect 109564 257758 109900 257786
rect 129528 257537 129556 258522
rect 131354 257664 131410 257673
rect 131354 257599 131410 257608
rect 87286 257528 87342 257537
rect 87286 257463 87342 257472
rect 129514 257528 129570 257537
rect 129514 257463 129570 257472
rect 131368 257294 131396 257599
rect 132748 257294 132776 263350
rect 143052 263249 143080 264030
rect 143038 263240 143094 263249
rect 143038 263175 143094 263184
rect 173412 262841 173440 274434
rect 175240 272384 175292 272390
rect 175240 272326 175292 272332
rect 175252 269670 175280 272326
rect 175240 269664 175292 269670
rect 175240 269606 175292 269612
rect 173398 262832 173454 262841
rect 173398 262767 173454 262776
rect 139636 262728 139688 262734
rect 139634 262696 139636 262705
rect 139688 262696 139690 262705
rect 139634 262631 139690 262640
rect 175332 262660 175384 262666
rect 175332 262602 175384 262608
rect 173674 262152 173730 262161
rect 173674 262087 173730 262096
rect 173584 261504 173636 261510
rect 140278 261472 140334 261481
rect 140278 261407 140334 261416
rect 173582 261472 173584 261481
rect 173636 261472 173638 261481
rect 173688 261442 173716 262087
rect 173582 261407 173638 261416
rect 173676 261436 173728 261442
rect 140094 259568 140150 259577
rect 140094 259503 140150 259512
rect 139910 258888 139966 258897
rect 139910 258823 139966 258832
rect 139818 258208 139874 258217
rect 139818 258143 139874 258152
rect 139634 257664 139690 257673
rect 139634 257599 139690 257608
rect 131356 257288 131408 257294
rect 131356 257230 131408 257236
rect 132736 257288 132788 257294
rect 132736 257230 132788 257236
rect 134208 257288 134260 257294
rect 134208 257230 134260 257236
rect 87196 257220 87248 257226
rect 87196 257162 87248 257168
rect 131540 257220 131592 257226
rect 131540 257162 131592 257168
rect 85172 257016 85224 257022
rect 85172 256958 85224 256964
rect 85080 256812 85132 256818
rect 85080 256754 85132 256760
rect 87208 256313 87236 257162
rect 131356 257152 131408 257158
rect 131356 257094 131408 257100
rect 87288 257016 87340 257022
rect 87288 256958 87340 256964
rect 87300 256857 87328 256958
rect 131368 256857 131396 257094
rect 131448 257084 131500 257090
rect 131448 257026 131500 257032
rect 87286 256848 87342 256857
rect 131354 256848 131410 256857
rect 87286 256783 87342 256792
rect 87564 256812 87616 256818
rect 131354 256783 131410 256792
rect 87564 256754 87616 256760
rect 87576 256721 87604 256754
rect 131460 256721 131488 257026
rect 87562 256712 87618 256721
rect 87562 256647 87618 256656
rect 131446 256712 131502 256721
rect 131446 256647 131502 256656
rect 131552 256313 131580 257162
rect 87194 256304 87250 256313
rect 87194 256239 87250 256248
rect 131538 256304 131594 256313
rect 131538 256239 131594 256248
rect 87196 255860 87248 255866
rect 87196 255802 87248 255808
rect 131540 255860 131592 255866
rect 131540 255802 131592 255808
rect 84436 255724 84488 255730
rect 84436 255666 84488 255672
rect 87208 255497 87236 255802
rect 87288 255792 87340 255798
rect 87288 255734 87340 255740
rect 131354 255760 131410 255769
rect 87194 255488 87250 255497
rect 87194 255423 87250 255432
rect 87300 255089 87328 255734
rect 87380 255724 87432 255730
rect 131354 255695 131410 255704
rect 131448 255724 131500 255730
rect 87380 255666 87432 255672
rect 87392 255633 87420 255666
rect 131368 255662 131396 255695
rect 131448 255666 131500 255672
rect 131356 255656 131408 255662
rect 87378 255624 87434 255633
rect 131356 255598 131408 255604
rect 87378 255559 87434 255568
rect 131460 255361 131488 255666
rect 131446 255352 131502 255361
rect 131446 255287 131502 255296
rect 131552 255225 131580 255802
rect 131632 255792 131684 255798
rect 131632 255734 131684 255740
rect 131538 255216 131594 255225
rect 131538 255151 131594 255160
rect 87286 255080 87342 255089
rect 87286 255015 87342 255024
rect 131644 254817 131672 255734
rect 131630 254808 131686 254817
rect 131630 254743 131686 254752
rect 84988 254500 85040 254506
rect 84988 254442 85040 254448
rect 82136 254228 82188 254234
rect 82136 254170 82188 254176
rect 80110 254128 80166 254137
rect 80110 254063 80166 254072
rect 80124 253282 80152 254063
rect 85000 253826 85028 254442
rect 87380 254432 87432 254438
rect 87194 254400 87250 254409
rect 87380 254374 87432 254380
rect 131540 254432 131592 254438
rect 131540 254374 131592 254380
rect 87194 254335 87250 254344
rect 87288 254364 87340 254370
rect 87208 254234 87236 254335
rect 87288 254306 87340 254312
rect 87300 254273 87328 254306
rect 87286 254264 87342 254273
rect 87196 254228 87248 254234
rect 87286 254199 87342 254208
rect 87196 254170 87248 254176
rect 87392 253865 87420 254374
rect 131356 254364 131408 254370
rect 131356 254306 131408 254312
rect 131368 254137 131396 254306
rect 131448 254296 131500 254302
rect 131448 254238 131500 254244
rect 131354 254128 131410 254137
rect 131354 254063 131410 254072
rect 87378 253856 87434 253865
rect 84988 253820 85040 253826
rect 84988 253762 85040 253768
rect 87196 253820 87248 253826
rect 87378 253791 87434 253800
rect 87196 253762 87248 253768
rect 87208 253457 87236 253762
rect 131460 253729 131488 254238
rect 131552 253865 131580 254374
rect 131538 253856 131594 253865
rect 131538 253791 131594 253800
rect 131446 253720 131502 253729
rect 131446 253655 131502 253664
rect 80202 253448 80258 253457
rect 80202 253383 80258 253392
rect 87194 253448 87250 253457
rect 87194 253383 87250 253392
rect 80112 253276 80164 253282
rect 80112 253218 80164 253224
rect 80216 253146 80244 253383
rect 80204 253140 80256 253146
rect 80204 253082 80256 253088
rect 87196 253072 87248 253078
rect 87194 253040 87196 253049
rect 131448 253072 131500 253078
rect 87248 253040 87250 253049
rect 131354 253040 131410 253049
rect 87194 252975 87250 252984
rect 87288 253004 87340 253010
rect 131448 253014 131500 253020
rect 131354 252975 131410 252984
rect 87288 252946 87340 252952
rect 80202 252768 80258 252777
rect 80202 252703 80258 252712
rect 80216 252398 80244 252703
rect 87300 252641 87328 252946
rect 131368 252942 131396 252975
rect 131356 252936 131408 252942
rect 131460 252913 131488 253014
rect 131540 253004 131592 253010
rect 131540 252946 131592 252952
rect 131356 252878 131408 252884
rect 131446 252904 131502 252913
rect 131446 252839 131502 252848
rect 87286 252632 87342 252641
rect 87286 252567 87342 252576
rect 131552 252505 131580 252946
rect 131538 252496 131594 252505
rect 131538 252431 131594 252440
rect 80204 252392 80256 252398
rect 80204 252334 80256 252340
rect 87196 252392 87248 252398
rect 87196 252334 87248 252340
rect 131356 252392 131408 252398
rect 131356 252334 131408 252340
rect 87208 252233 87236 252334
rect 87194 252224 87250 252233
rect 87194 252159 87250 252168
rect 80202 252088 80258 252097
rect 80202 252023 80258 252032
rect 80216 251786 80244 252023
rect 131368 251961 131396 252334
rect 131354 251952 131410 251961
rect 131354 251887 131410 251896
rect 80204 251780 80256 251786
rect 80204 251722 80256 251728
rect 131356 251712 131408 251718
rect 131356 251654 131408 251660
rect 87196 251644 87248 251650
rect 87196 251586 87248 251592
rect 87208 251553 87236 251586
rect 131368 251553 131396 251654
rect 87194 251544 87250 251553
rect 87194 251479 87250 251488
rect 131354 251544 131410 251553
rect 131354 251479 131410 251488
rect 80202 251408 80258 251417
rect 80202 251343 80258 251352
rect 80216 251106 80244 251343
rect 87194 251136 87250 251145
rect 80204 251100 80256 251106
rect 87194 251071 87196 251080
rect 80204 251042 80256 251048
rect 87248 251071 87250 251080
rect 131354 251136 131410 251145
rect 131354 251071 131356 251080
rect 87196 251042 87248 251048
rect 131408 251071 131410 251080
rect 131356 251042 131408 251048
rect 80112 251032 80164 251038
rect 87288 251032 87340 251038
rect 80112 250974 80164 250980
rect 87286 251000 87288 251009
rect 131448 251032 131500 251038
rect 87340 251000 87342 251009
rect 80124 250737 80152 250974
rect 131448 250974 131500 250980
rect 87286 250935 87342 250944
rect 131460 250737 131488 250974
rect 80110 250728 80166 250737
rect 80110 250663 80166 250672
rect 131446 250728 131502 250737
rect 131446 250663 131502 250672
rect 87194 250320 87250 250329
rect 87194 250255 87250 250264
rect 131354 250320 131410 250329
rect 131354 250255 131356 250264
rect 80110 250184 80166 250193
rect 80110 250119 80166 250128
rect 47082 249912 47138 249921
rect 47082 249847 47138 249856
rect 80124 249678 80152 250119
rect 87208 249678 87236 250255
rect 131408 250255 131410 250264
rect 131356 250226 131408 250232
rect 87286 250048 87342 250057
rect 87286 249983 87342 249992
rect 131354 250048 131410 250057
rect 131354 249983 131410 249992
rect 80112 249672 80164 249678
rect 80112 249614 80164 249620
rect 87196 249672 87248 249678
rect 87196 249614 87248 249620
rect 87300 249610 87328 249983
rect 87378 249640 87434 249649
rect 80204 249604 80256 249610
rect 80204 249546 80256 249552
rect 87288 249604 87340 249610
rect 131368 249610 131396 249983
rect 131816 249672 131868 249678
rect 131814 249640 131816 249649
rect 131868 249640 131870 249649
rect 87378 249575 87434 249584
rect 131356 249604 131408 249610
rect 87288 249546 87340 249552
rect 80216 249513 80244 249546
rect 80202 249504 80258 249513
rect 80202 249439 80258 249448
rect 87194 249232 87250 249241
rect 87194 249167 87250 249176
rect 87208 248930 87236 249167
rect 79284 248924 79336 248930
rect 79284 248866 79336 248872
rect 87196 248924 87248 248930
rect 87196 248866 87248 248872
rect 79296 248561 79324 248866
rect 87392 248862 87420 249575
rect 131814 249575 131870 249584
rect 131356 249546 131408 249552
rect 131354 249232 131410 249241
rect 131354 249167 131410 249176
rect 131368 248998 131396 249167
rect 131356 248992 131408 248998
rect 131356 248934 131408 248940
rect 80204 248856 80256 248862
rect 80202 248824 80204 248833
rect 87380 248856 87432 248862
rect 80256 248824 80258 248833
rect 87380 248798 87432 248804
rect 88298 248824 88354 248833
rect 80202 248759 80258 248768
rect 88298 248759 88354 248768
rect 131354 248824 131410 248833
rect 131354 248759 131410 248768
rect 79282 248552 79338 248561
rect 79282 248487 79338 248496
rect 88022 248008 88078 248017
rect 88022 247943 88078 247952
rect 88036 247774 88064 247943
rect 85908 247768 85960 247774
rect 85908 247710 85960 247716
rect 88024 247768 88076 247774
rect 88024 247710 88076 247716
rect 79284 247564 79336 247570
rect 79284 247506 79336 247512
rect 79296 247201 79324 247506
rect 80204 247496 80256 247502
rect 80202 247464 80204 247473
rect 80256 247464 80258 247473
rect 80202 247399 80258 247408
rect 79282 247192 79338 247201
rect 79282 247127 79338 247136
rect 80020 246408 80072 246414
rect 80020 246350 80072 246356
rect 79284 246204 79336 246210
rect 79284 246146 79336 246152
rect 79296 245841 79324 246146
rect 79282 245832 79338 245841
rect 79282 245767 79338 245776
rect 79928 243552 79980 243558
rect 79928 243494 79980 243500
rect 79284 242260 79336 242266
rect 79284 242202 79336 242208
rect 79100 242056 79152 242062
rect 79100 241998 79152 242004
rect 79112 241353 79140 241998
rect 79098 241344 79154 241353
rect 79098 241279 79154 241288
rect 79296 238633 79324 242202
rect 79940 239993 79968 243494
rect 80032 243393 80060 246350
rect 80202 246104 80258 246113
rect 80202 246039 80258 246048
rect 80216 245938 80244 246039
rect 85920 245938 85948 247710
rect 86092 247632 86144 247638
rect 87196 247632 87248 247638
rect 86092 247574 86144 247580
rect 87194 247600 87196 247609
rect 87248 247600 87250 247609
rect 86104 246210 86132 247574
rect 87194 247535 87250 247544
rect 88312 247502 88340 248759
rect 88390 248416 88446 248425
rect 88390 248351 88446 248360
rect 88404 247570 88432 248351
rect 131368 248250 131396 248759
rect 131446 248416 131502 248425
rect 131446 248351 131502 248360
rect 131356 248244 131408 248250
rect 131356 248186 131408 248192
rect 131460 247638 131488 248351
rect 132550 248008 132606 248017
rect 132550 247943 132606 247952
rect 131816 247768 131868 247774
rect 131814 247736 131816 247745
rect 131868 247736 131870 247745
rect 132564 247706 132592 247943
rect 131814 247671 131870 247680
rect 132552 247700 132604 247706
rect 132552 247642 132604 247648
rect 131448 247632 131500 247638
rect 131448 247574 131500 247580
rect 88392 247564 88444 247570
rect 88392 247506 88444 247512
rect 88300 247496 88352 247502
rect 88300 247438 88352 247444
rect 131446 247328 131502 247337
rect 131446 247263 131502 247272
rect 87010 247192 87066 247201
rect 87010 247127 87066 247136
rect 86092 246204 86144 246210
rect 86092 246146 86144 246152
rect 86918 245968 86974 245977
rect 80204 245932 80256 245938
rect 80204 245874 80256 245880
rect 85908 245932 85960 245938
rect 86918 245903 86974 245912
rect 85908 245874 85960 245880
rect 86826 245560 86882 245569
rect 86826 245495 86882 245504
rect 80112 244776 80164 244782
rect 80112 244718 80164 244724
rect 80202 244744 80258 244753
rect 80124 244481 80152 244718
rect 80202 244679 80204 244688
rect 80256 244679 80258 244688
rect 80204 244650 80256 244656
rect 80110 244472 80166 244481
rect 80110 244407 80166 244416
rect 80112 243484 80164 243490
rect 80112 243426 80164 243432
rect 80018 243384 80074 243393
rect 80018 243319 80074 243328
rect 80124 240673 80152 243426
rect 80204 243416 80256 243422
rect 80204 243358 80256 243364
rect 80216 243121 80244 243358
rect 80202 243112 80258 243121
rect 80202 243047 80258 243056
rect 86840 242810 86868 245495
rect 86932 243422 86960 245903
rect 87024 244714 87052 247127
rect 87102 246784 87158 246793
rect 87102 246719 87158 246728
rect 87116 244782 87144 246719
rect 131354 246512 131410 246521
rect 131354 246447 131410 246456
rect 87196 246408 87248 246414
rect 87194 246376 87196 246385
rect 87248 246376 87250 246385
rect 87194 246311 87250 246320
rect 131368 246278 131396 246447
rect 131460 246414 131488 247263
rect 132182 246920 132238 246929
rect 132182 246855 132238 246864
rect 131448 246408 131500 246414
rect 131448 246350 131500 246356
rect 132196 246346 132224 246855
rect 132184 246340 132236 246346
rect 132184 246282 132236 246288
rect 131356 246272 131408 246278
rect 131356 246214 131408 246220
rect 131998 246104 132054 246113
rect 131998 246039 132054 246048
rect 131446 245832 131502 245841
rect 131446 245767 131502 245776
rect 131354 245424 131410 245433
rect 131354 245359 131410 245368
rect 87654 245152 87710 245161
rect 87654 245087 87710 245096
rect 87104 244776 87156 244782
rect 87104 244718 87156 244724
rect 87562 244744 87618 244753
rect 87012 244708 87064 244714
rect 87562 244679 87618 244688
rect 87012 244650 87064 244656
rect 87286 244336 87342 244345
rect 87286 244271 87342 244280
rect 87194 243928 87250 243937
rect 87194 243863 87250 243872
rect 87208 243558 87236 243863
rect 87196 243552 87248 243558
rect 87196 243494 87248 243500
rect 87300 243490 87328 244271
rect 87470 243520 87526 243529
rect 87288 243484 87340 243490
rect 87470 243455 87526 243464
rect 87288 243426 87340 243432
rect 86920 243416 86972 243422
rect 86920 243358 86972 243364
rect 87194 243112 87250 243121
rect 87194 243047 87250 243056
rect 80204 242804 80256 242810
rect 80204 242746 80256 242752
rect 86828 242804 86880 242810
rect 86828 242746 86880 242752
rect 80216 242441 80244 242746
rect 86550 242704 86606 242713
rect 86550 242639 86606 242648
rect 80202 242432 80258 242441
rect 80202 242367 80258 242376
rect 86458 242296 86514 242305
rect 86458 242231 86514 242240
rect 80204 241988 80256 241994
rect 80204 241930 80256 241936
rect 80216 241761 80244 241930
rect 80202 241752 80258 241761
rect 80202 241687 80258 241696
rect 85080 240696 85132 240702
rect 80110 240664 80166 240673
rect 85080 240638 85132 240644
rect 80110 240599 80166 240608
rect 79926 239984 79982 239993
rect 79926 239919 79982 239928
rect 80204 239268 80256 239274
rect 80204 239210 80256 239216
rect 80216 239041 80244 239210
rect 80202 239032 80258 239041
rect 80202 238967 80258 238976
rect 79282 238624 79338 238633
rect 79282 238559 79338 238568
rect 80204 237908 80256 237914
rect 80204 237850 80256 237856
rect 80216 237681 80244 237850
rect 80202 237672 80258 237681
rect 80202 237607 80258 237616
rect 80204 237364 80256 237370
rect 80204 237306 80256 237312
rect 80216 237001 80244 237306
rect 80202 236992 80258 237001
rect 80202 236927 80258 236936
rect 80202 236176 80258 236185
rect 80202 236111 80258 236120
rect 64300 235998 64866 236026
rect 49212 233086 49240 235876
rect 38160 233080 38212 233086
rect 38160 233022 38212 233028
rect 49200 233080 49252 233086
rect 49200 233022 49252 233028
rect 38172 203409 38200 233022
rect 49856 224790 49884 235876
rect 50514 235862 51172 235890
rect 51144 224926 51172 235862
rect 51236 225062 51264 235876
rect 51880 225334 51908 235876
rect 52524 235862 52630 235890
rect 51868 225328 51920 225334
rect 51868 225270 51920 225276
rect 52524 225130 52552 235862
rect 53260 233154 53288 235876
rect 53918 235862 54024 235890
rect 53248 233148 53300 233154
rect 53248 233090 53300 233096
rect 52512 225124 52564 225130
rect 52512 225066 52564 225072
rect 51224 225056 51276 225062
rect 51224 224998 51276 225004
rect 51132 224920 51184 224926
rect 51132 224862 51184 224868
rect 49844 224784 49896 224790
rect 49844 224726 49896 224732
rect 53996 224654 54024 235862
rect 54640 225198 54668 235876
rect 55284 225402 55312 235876
rect 56020 233018 56048 235876
rect 56008 233012 56060 233018
rect 56008 232954 56060 232960
rect 56664 232882 56692 235876
rect 56652 232876 56704 232882
rect 56652 232818 56704 232824
rect 57308 232610 57336 235876
rect 57940 233556 57992 233562
rect 57940 233498 57992 233504
rect 57664 233284 57716 233290
rect 57664 233226 57716 233232
rect 57296 232604 57348 232610
rect 57296 232546 57348 232552
rect 57676 225470 57704 233226
rect 56192 225464 56244 225470
rect 56192 225406 56244 225412
rect 57664 225464 57716 225470
rect 57664 225406 57716 225412
rect 55272 225396 55324 225402
rect 55272 225338 55324 225344
rect 55824 225260 55876 225266
rect 55824 225202 55876 225208
rect 54628 225192 54680 225198
rect 54628 225134 54680 225140
rect 53984 224648 54036 224654
rect 53984 224590 54036 224596
rect 55088 224376 55140 224382
rect 55088 224318 55140 224324
rect 38252 224172 38304 224178
rect 38252 224114 38304 224120
rect 38264 211297 38292 224114
rect 55100 222820 55128 224318
rect 55732 224308 55784 224314
rect 55732 224250 55784 224256
rect 55744 222834 55772 224250
rect 55482 222806 55772 222834
rect 55836 222820 55864 225202
rect 56204 222820 56232 225406
rect 57952 225198 57980 233498
rect 58044 232746 58072 235876
rect 58032 232740 58084 232746
rect 58032 232682 58084 232688
rect 58688 225470 58716 235876
rect 59320 232808 59372 232814
rect 59320 232750 59372 232756
rect 58676 225464 58728 225470
rect 58676 225406 58728 225412
rect 56560 225192 56612 225198
rect 56560 225134 56612 225140
rect 57940 225192 57992 225198
rect 57940 225134 57992 225140
rect 58124 225192 58176 225198
rect 58124 225134 58176 225140
rect 56572 222820 56600 225134
rect 57296 224716 57348 224722
rect 57296 224658 57348 224664
rect 57308 222834 57336 224658
rect 57756 224580 57808 224586
rect 57756 224522 57808 224528
rect 57388 224512 57440 224518
rect 57388 224454 57440 224460
rect 57046 222806 57336 222834
rect 57400 222820 57428 224454
rect 57768 222820 57796 224522
rect 58136 222820 58164 225134
rect 58584 224988 58636 224994
rect 58584 224930 58636 224936
rect 58596 222820 58624 224930
rect 58952 224240 59004 224246
rect 58952 224182 59004 224188
rect 58964 222820 58992 224182
rect 59332 222820 59360 232750
rect 59424 225130 59452 235876
rect 60068 232474 60096 235876
rect 60148 233624 60200 233630
rect 60148 233566 60200 233572
rect 60056 232468 60108 232474
rect 60056 232410 60108 232416
rect 59504 225464 59556 225470
rect 59504 225406 59556 225412
rect 59412 225124 59464 225130
rect 59412 225066 59464 225072
rect 59516 224110 59544 225406
rect 59688 225260 59740 225266
rect 59688 225202 59740 225208
rect 59504 224104 59556 224110
rect 59504 224046 59556 224052
rect 59700 222820 59728 225202
rect 60160 222820 60188 233566
rect 60608 233488 60660 233494
rect 60608 233430 60660 233436
rect 60620 225146 60648 233430
rect 60698 233048 60754 233057
rect 60698 232983 60754 232992
rect 60712 225282 60740 232983
rect 60804 232678 60832 235876
rect 61462 235862 62028 235890
rect 60884 233692 60936 233698
rect 60884 233634 60936 233640
rect 60792 232672 60844 232678
rect 60792 232614 60844 232620
rect 60896 225418 60924 233634
rect 61252 233420 61304 233426
rect 61252 233362 61304 233368
rect 61160 232468 61212 232474
rect 61160 232410 61212 232416
rect 60896 225390 61016 225418
rect 60712 225254 60924 225282
rect 60988 225266 61016 225390
rect 60620 225118 60740 225146
rect 60712 222834 60740 225118
rect 60542 222806 60740 222834
rect 60896 222820 60924 225254
rect 60976 225260 61028 225266
rect 60976 225202 61028 225208
rect 61172 224926 61200 232410
rect 61160 224920 61212 224926
rect 61160 224862 61212 224868
rect 61158 224344 61214 224353
rect 61158 224279 61214 224288
rect 61172 224246 61200 224279
rect 61160 224240 61212 224246
rect 61160 224182 61212 224188
rect 61264 222820 61292 233362
rect 61712 233216 61764 233222
rect 61712 233158 61764 233164
rect 61344 232740 61396 232746
rect 61344 232682 61396 232688
rect 61528 232740 61580 232746
rect 61528 232682 61580 232688
rect 61356 224194 61384 232682
rect 61436 232604 61488 232610
rect 61436 232546 61488 232552
rect 61448 224330 61476 232546
rect 61540 224586 61568 232682
rect 61620 232672 61672 232678
rect 61620 232614 61672 232620
rect 61528 224580 61580 224586
rect 61528 224522 61580 224528
rect 61632 224518 61660 232614
rect 61724 224926 61752 233158
rect 62000 232626 62028 235862
rect 62092 233222 62120 235876
rect 62080 233216 62132 233222
rect 62080 233158 62132 233164
rect 62264 233216 62316 233222
rect 62264 233158 62316 233164
rect 62080 233080 62132 233086
rect 62080 233022 62132 233028
rect 61804 232604 61856 232610
rect 61804 232546 61856 232552
rect 61908 232598 62028 232626
rect 61712 224920 61764 224926
rect 61712 224862 61764 224868
rect 61620 224512 61672 224518
rect 61620 224454 61672 224460
rect 61712 224512 61764 224518
rect 61712 224454 61764 224460
rect 61724 224330 61752 224454
rect 61448 224302 61752 224330
rect 61816 224314 61844 232546
rect 61908 225130 61936 232598
rect 61988 232468 62040 232474
rect 61988 232410 62040 232416
rect 62000 225198 62028 232410
rect 61988 225192 62040 225198
rect 61988 225134 62040 225140
rect 61896 225124 61948 225130
rect 61896 225066 61948 225072
rect 61804 224308 61856 224314
rect 61804 224250 61856 224256
rect 61896 224308 61948 224314
rect 61896 224250 61948 224256
rect 61908 224194 61936 224250
rect 61356 224166 61936 224194
rect 62092 223242 62120 233022
rect 62172 232536 62224 232542
rect 62172 232478 62224 232484
rect 62184 224722 62212 232478
rect 62172 224716 62224 224722
rect 62172 224658 62224 224664
rect 62000 223214 62120 223242
rect 62000 222834 62028 223214
rect 62276 222834 62304 233158
rect 62356 233148 62408 233154
rect 62356 233090 62408 233096
rect 62448 233148 62500 233154
rect 62448 233090 62500 233096
rect 62368 224722 62396 233090
rect 62356 224716 62408 224722
rect 62356 224658 62408 224664
rect 61738 222806 62028 222834
rect 62106 222806 62304 222834
rect 62460 222820 62488 233090
rect 62828 225266 62856 235876
rect 63472 232610 63500 235876
rect 63748 235862 64222 235890
rect 63644 232944 63696 232950
rect 63644 232886 63696 232892
rect 63460 232604 63512 232610
rect 63460 232546 63512 232552
rect 62816 225260 62868 225266
rect 62816 225202 62868 225208
rect 63656 225062 63684 232886
rect 63644 225056 63696 225062
rect 63644 224998 63696 225004
rect 63368 224784 63420 224790
rect 63368 224726 63420 224732
rect 62816 224444 62868 224450
rect 62816 224386 62868 224392
rect 62908 224444 62960 224450
rect 62908 224386 62960 224392
rect 62828 222820 62856 224386
rect 62920 224353 62948 224386
rect 62906 224344 62962 224353
rect 62906 224279 62962 224288
rect 63276 223696 63328 223702
rect 63276 223638 63328 223644
rect 63288 222820 63316 223638
rect 63380 222698 63408 224726
rect 63748 224042 63776 235862
rect 64300 225470 64328 235998
rect 65496 233290 65524 235876
rect 66232 233562 66260 235876
rect 66220 233556 66272 233562
rect 66220 233498 66272 233504
rect 65484 233284 65536 233290
rect 65484 233226 65536 233232
rect 66036 233012 66088 233018
rect 66036 232954 66088 232960
rect 64288 225464 64340 225470
rect 64288 225406 64340 225412
rect 64012 225396 64064 225402
rect 64012 225338 64064 225344
rect 63736 224036 63788 224042
rect 63736 223978 63788 223984
rect 64024 222820 64052 225338
rect 65944 225328 65996 225334
rect 65944 225270 65996 225276
rect 64380 224852 64432 224858
rect 64380 224794 64432 224800
rect 64392 222820 64420 224794
rect 64840 224716 64892 224722
rect 64840 224658 64892 224664
rect 64852 222820 64880 224658
rect 65208 224648 65260 224654
rect 65208 224590 65260 224596
rect 65220 222820 65248 224590
rect 65576 224376 65628 224382
rect 65576 224318 65628 224324
rect 65588 222820 65616 224318
rect 65956 222820 65984 225270
rect 66048 222698 66076 232954
rect 66404 232876 66456 232882
rect 66404 232818 66456 232824
rect 66416 225418 66444 232818
rect 66876 232542 66904 235876
rect 67612 232678 67640 235876
rect 68256 232746 68284 235876
rect 68244 232740 68296 232746
rect 68244 232682 68296 232688
rect 67600 232672 67652 232678
rect 67600 232614 67652 232620
rect 67968 232604 68020 232610
rect 67968 232546 68020 232552
rect 66864 232536 66916 232542
rect 66864 232478 66916 232484
rect 67876 232536 67928 232542
rect 67876 232478 67928 232484
rect 66416 225390 66812 225418
rect 66784 222820 66812 225390
rect 67888 225198 67916 232478
rect 67876 225192 67928 225198
rect 67876 225134 67928 225140
rect 67140 224512 67192 224518
rect 67140 224454 67192 224460
rect 67152 222820 67180 224454
rect 67980 224450 68008 232546
rect 68992 232474 69020 235876
rect 69636 232542 69664 235876
rect 70280 232610 70308 235876
rect 71016 232678 71044 235876
rect 71660 233630 71688 235876
rect 71648 233624 71700 233630
rect 71648 233566 71700 233572
rect 72396 233494 72424 235876
rect 72384 233488 72436 233494
rect 72384 233430 72436 233436
rect 73040 233290 73068 235876
rect 73028 233284 73080 233290
rect 73028 233226 73080 233232
rect 73684 233057 73712 235876
rect 74420 233426 74448 235876
rect 74408 233420 74460 233426
rect 74408 233362 74460 233368
rect 75064 233086 75092 235876
rect 75800 233222 75828 235876
rect 75788 233216 75840 233222
rect 75788 233158 75840 233164
rect 76444 233154 76472 235876
rect 80216 235330 80244 236111
rect 85092 235330 85120 240638
rect 86472 237370 86500 242231
rect 86564 237914 86592 242639
rect 87208 242266 87236 243047
rect 87196 242260 87248 242266
rect 87196 242202 87248 242208
rect 87378 242024 87434 242033
rect 87378 241959 87434 241968
rect 87392 240702 87420 241959
rect 87380 240696 87432 240702
rect 87380 240638 87432 240644
rect 87484 239274 87512 243455
rect 87576 242062 87604 244679
rect 87564 242056 87616 242062
rect 87564 241998 87616 242004
rect 87668 241994 87696 245087
rect 131368 244986 131396 245359
rect 131356 244980 131408 244986
rect 131356 244922 131408 244928
rect 131460 244850 131488 245767
rect 131816 245048 131868 245054
rect 131814 245016 131816 245025
rect 131868 245016 131870 245025
rect 131814 244951 131870 244960
rect 132012 244918 132040 246039
rect 132000 244912 132052 244918
rect 132000 244854 132052 244860
rect 131448 244844 131500 244850
rect 131448 244786 131500 244792
rect 131630 244608 131686 244617
rect 131630 244543 131686 244552
rect 131538 244200 131594 244209
rect 131538 244135 131594 244144
rect 131354 243928 131410 243937
rect 131354 243863 131410 243872
rect 131368 243694 131396 243863
rect 131356 243688 131408 243694
rect 131356 243630 131408 243636
rect 131448 243620 131500 243626
rect 131448 243562 131500 243568
rect 131460 243529 131488 243562
rect 131552 243558 131580 244135
rect 131540 243552 131592 243558
rect 131446 243520 131502 243529
rect 131540 243494 131592 243500
rect 131644 243490 131672 244543
rect 131446 243455 131502 243464
rect 131632 243484 131684 243490
rect 131632 243426 131684 243432
rect 131538 243112 131594 243121
rect 131538 243047 131594 243056
rect 131446 242704 131502 242713
rect 131446 242639 131502 242648
rect 131354 242296 131410 242305
rect 131354 242231 131356 242240
rect 131408 242231 131410 242240
rect 131356 242202 131408 242208
rect 131460 242198 131488 242639
rect 131448 242192 131500 242198
rect 131448 242134 131500 242140
rect 131552 242130 131580 243047
rect 131540 242124 131592 242130
rect 131540 242066 131592 242072
rect 131354 242024 131410 242033
rect 87656 241988 87708 241994
rect 131354 241959 131410 241968
rect 87656 241930 87708 241936
rect 109886 241602 109914 241860
rect 109886 241574 109960 241602
rect 109932 240498 109960 241574
rect 131368 240702 131396 241959
rect 131356 240696 131408 240702
rect 131356 240638 131408 240644
rect 109920 240492 109972 240498
rect 109920 240434 109972 240440
rect 87472 239268 87524 239274
rect 87472 239210 87524 239216
rect 86552 237908 86604 237914
rect 86552 237850 86604 237856
rect 86460 237364 86512 237370
rect 86460 237306 86512 237312
rect 80204 235324 80256 235330
rect 80204 235266 80256 235272
rect 85080 235324 85132 235330
rect 85080 235266 85132 235272
rect 76432 233148 76484 233154
rect 76432 233090 76484 233096
rect 75052 233080 75104 233086
rect 73670 233048 73726 233057
rect 75052 233022 75104 233028
rect 73670 232983 73726 232992
rect 71004 232672 71056 232678
rect 71004 232614 71056 232620
rect 70268 232604 70320 232610
rect 70268 232546 70320 232552
rect 69624 232536 69676 232542
rect 69624 232478 69676 232484
rect 68980 232468 69032 232474
rect 68980 232410 69032 232416
rect 126480 229680 126532 229686
rect 126480 229622 126532 229628
rect 126492 227716 126520 229622
rect 70268 225260 70320 225266
rect 70268 225202 70320 225208
rect 69532 225124 69584 225130
rect 69532 225066 69584 225072
rect 69072 225056 69124 225062
rect 69072 224998 69124 225004
rect 68336 224988 68388 224994
rect 68336 224930 68388 224936
rect 67968 224444 68020 224450
rect 67968 224386 68020 224392
rect 67508 224308 67560 224314
rect 67508 224250 67560 224256
rect 67520 222820 67548 224250
rect 67968 224172 68020 224178
rect 67968 224114 68020 224120
rect 67980 222820 68008 224114
rect 68348 222820 68376 224930
rect 68704 224580 68756 224586
rect 68704 224522 68756 224528
rect 68716 222820 68744 224522
rect 69084 222820 69112 224998
rect 69544 222820 69572 225066
rect 69900 224920 69952 224926
rect 69900 224862 69952 224868
rect 69912 222820 69940 224862
rect 70280 222820 70308 225202
rect 70636 224172 70688 224178
rect 70636 224114 70688 224120
rect 70648 222820 70676 224114
rect 63380 222670 63670 222698
rect 66048 222670 66430 222698
rect 51958 216184 52014 216193
rect 51958 216119 52014 216128
rect 38250 211288 38306 211297
rect 38250 211223 38306 211232
rect 38158 203400 38214 203409
rect 38158 203335 38214 203344
rect 51972 202185 52000 216119
rect 134220 211818 134248 257230
rect 139648 255798 139676 257599
rect 139726 256304 139782 256313
rect 139726 256239 139782 256248
rect 139636 255792 139688 255798
rect 139636 255734 139688 255740
rect 139634 255624 139690 255633
rect 139634 255559 139690 255568
rect 139648 254302 139676 255559
rect 139740 254438 139768 256239
rect 139832 255866 139860 258143
rect 139820 255860 139872 255866
rect 139820 255802 139872 255808
rect 139924 255730 139952 258823
rect 140002 256984 140058 256993
rect 140002 256919 140058 256928
rect 139912 255724 139964 255730
rect 139912 255666 139964 255672
rect 139910 254944 139966 254953
rect 139910 254879 139966 254888
rect 139728 254432 139780 254438
rect 139728 254374 139780 254380
rect 139818 254400 139874 254409
rect 139818 254335 139874 254344
rect 139636 254296 139688 254302
rect 139636 254238 139688 254244
rect 139634 253720 139690 253729
rect 139634 253655 139690 253664
rect 139648 253010 139676 253655
rect 139832 253078 139860 254335
rect 139820 253072 139872 253078
rect 139820 253014 139872 253020
rect 139636 253004 139688 253010
rect 139636 252946 139688 252952
rect 139924 252942 139952 254879
rect 140016 254370 140044 256919
rect 140108 255662 140136 259503
rect 140292 257158 140320 261407
rect 173676 261378 173728 261384
rect 140370 260928 140426 260937
rect 140370 260863 140426 260872
rect 140280 257152 140332 257158
rect 140280 257094 140332 257100
rect 140384 257090 140412 260863
rect 172846 260792 172902 260801
rect 172846 260727 172902 260736
rect 140554 260248 140610 260257
rect 140554 260183 140610 260192
rect 140568 257226 140596 260183
rect 172860 260150 172888 260727
rect 172848 260144 172900 260150
rect 172848 260086 172900 260092
rect 173582 260112 173638 260121
rect 173582 260047 173584 260056
rect 173636 260047 173638 260056
rect 173584 260018 173636 260024
rect 175344 260014 175372 262602
rect 181956 261504 182008 261510
rect 181956 261446 182008 261452
rect 181772 261436 181824 261442
rect 181772 261378 181824 261384
rect 179012 260144 179064 260150
rect 179012 260086 179064 260092
rect 175332 260008 175384 260014
rect 175332 259950 175384 259956
rect 173398 259432 173454 259441
rect 173398 259367 173400 259376
rect 173452 259367 173454 259376
rect 175700 259396 175752 259402
rect 173400 259338 173452 259344
rect 175700 259338 175752 259344
rect 173582 258752 173638 258761
rect 173582 258687 173584 258696
rect 173636 258687 173638 258696
rect 173584 258658 173636 258664
rect 173306 258072 173362 258081
rect 173306 258007 173308 258016
rect 173360 258007 173362 258016
rect 175608 258036 175660 258042
rect 173308 257978 173360 257984
rect 175608 257978 175660 257984
rect 173582 257392 173638 257401
rect 173582 257327 173584 257336
rect 173636 257327 173638 257336
rect 175516 257356 175568 257362
rect 173584 257298 173636 257304
rect 175516 257298 175568 257304
rect 140556 257220 140608 257226
rect 140556 257162 140608 257168
rect 140372 257084 140424 257090
rect 140372 257026 140424 257032
rect 173122 256848 173178 256857
rect 173122 256783 173178 256792
rect 173136 256478 173164 256783
rect 173124 256472 173176 256478
rect 173124 256414 173176 256420
rect 173306 256168 173362 256177
rect 173306 256103 173308 256112
rect 173360 256103 173362 256112
rect 173308 256074 173360 256080
rect 175528 255798 175556 257298
rect 175620 255866 175648 257978
rect 175712 257090 175740 259338
rect 178920 258716 178972 258722
rect 178920 258658 178972 258664
rect 175700 257084 175752 257090
rect 175700 257026 175752 257032
rect 175792 256472 175844 256478
rect 175792 256414 175844 256420
rect 175700 256132 175752 256138
rect 175700 256074 175752 256080
rect 175608 255860 175660 255866
rect 175608 255802 175660 255808
rect 175516 255792 175568 255798
rect 175516 255734 175568 255740
rect 140096 255656 140148 255662
rect 140096 255598 140148 255604
rect 173214 255488 173270 255497
rect 173214 255423 173270 255432
rect 173228 254574 173256 255423
rect 173490 254808 173546 254817
rect 173490 254743 173546 254752
rect 173216 254568 173268 254574
rect 173216 254510 173268 254516
rect 173504 254506 173532 254743
rect 173492 254500 173544 254506
rect 173492 254442 173544 254448
rect 140004 254364 140056 254370
rect 140004 254306 140056 254312
rect 175712 254234 175740 256074
rect 175804 254302 175832 256414
rect 178932 255730 178960 258658
rect 179024 257226 179052 260086
rect 179104 260076 179156 260082
rect 179104 260018 179156 260024
rect 179012 257220 179064 257226
rect 179012 257162 179064 257168
rect 179116 257158 179144 260018
rect 181784 258353 181812 261378
rect 181770 258344 181826 258353
rect 181770 258279 181826 258288
rect 181968 257537 181996 261446
rect 182336 258586 182364 284799
rect 225194 280784 225250 280793
rect 225194 280719 225250 280728
rect 188882 276934 189264 276962
rect 189236 260694 189264 276934
rect 198712 276934 198818 276962
rect 198712 276690 198740 276934
rect 198712 276662 198924 276690
rect 198896 264026 198924 276662
rect 208832 274498 208860 276948
rect 218860 274498 218888 276948
rect 208820 274492 208872 274498
rect 208820 274434 208872 274440
rect 218848 274492 218900 274498
rect 218848 274434 218900 274440
rect 225208 264094 225236 280719
rect 225288 274492 225340 274498
rect 225288 274434 225340 274440
rect 225196 264088 225248 264094
rect 225196 264030 225248 264036
rect 198884 264020 198936 264026
rect 198884 263962 198936 263968
rect 189224 260688 189276 260694
rect 189224 260630 189276 260636
rect 203852 260688 203904 260694
rect 203852 260630 203904 260636
rect 182324 258580 182376 258586
rect 182324 258522 182376 258528
rect 203864 257772 203892 260630
rect 223540 258580 223592 258586
rect 223540 258522 223592 258528
rect 223552 257537 223580 258522
rect 225300 257673 225328 274434
rect 233476 264020 233528 264026
rect 233476 263962 233528 263968
rect 233488 263929 233516 263962
rect 233474 263920 233530 263929
rect 233474 263855 233530 263864
rect 234302 262696 234358 262705
rect 234302 262631 234358 262640
rect 234118 262016 234174 262025
rect 234118 261951 234174 261960
rect 233474 260656 233530 260665
rect 233474 260591 233530 260600
rect 233488 260082 233516 260591
rect 229980 260076 230032 260082
rect 229980 260018 230032 260024
rect 233476 260076 233528 260082
rect 233476 260018 233528 260024
rect 229428 257764 229480 257770
rect 229428 257706 229480 257712
rect 225286 257664 225342 257673
rect 225286 257599 225342 257608
rect 181954 257528 182010 257537
rect 181954 257463 182010 257472
rect 223538 257528 223594 257537
rect 223538 257463 223594 257472
rect 182324 257220 182376 257226
rect 182324 257162 182376 257168
rect 226208 257220 226260 257226
rect 226208 257162 226260 257168
rect 179104 257152 179156 257158
rect 179104 257094 179156 257100
rect 182232 257152 182284 257158
rect 182336 257129 182364 257162
rect 182232 257094 182284 257100
rect 182322 257120 182378 257129
rect 182048 257084 182100 257090
rect 182048 257026 182100 257032
rect 182060 256313 182088 257026
rect 182244 256721 182272 257094
rect 182322 257055 182378 257064
rect 225380 257084 225432 257090
rect 225380 257026 225432 257032
rect 182230 256712 182286 256721
rect 182230 256647 182286 256656
rect 225392 256449 225420 257026
rect 226220 256857 226248 257162
rect 226300 257152 226352 257158
rect 226300 257094 226352 257100
rect 226206 256848 226262 256857
rect 226206 256783 226262 256792
rect 225378 256440 225434 256449
rect 225378 256375 225434 256384
rect 182046 256304 182102 256313
rect 182046 256239 182102 256248
rect 226312 256041 226340 257094
rect 226298 256032 226354 256041
rect 226298 255967 226354 255976
rect 181864 255860 181916 255866
rect 181864 255802 181916 255808
rect 225564 255860 225616 255866
rect 225564 255802 225616 255808
rect 178920 255724 178972 255730
rect 178920 255666 178972 255672
rect 181876 255497 181904 255802
rect 182232 255792 182284 255798
rect 182232 255734 182284 255740
rect 181862 255488 181918 255497
rect 181862 255423 181918 255432
rect 182244 255089 182272 255734
rect 182324 255724 182376 255730
rect 182324 255666 182376 255672
rect 182336 255633 182364 255666
rect 182322 255624 182378 255633
rect 182322 255559 182378 255568
rect 182230 255080 182286 255089
rect 182230 255015 182286 255024
rect 225576 254953 225604 255802
rect 226392 255792 226444 255798
rect 226298 255760 226354 255769
rect 226392 255734 226444 255740
rect 226298 255695 226300 255704
rect 226352 255695 226354 255704
rect 226300 255666 226352 255672
rect 225932 255656 225984 255662
rect 225932 255598 225984 255604
rect 225562 254944 225618 254953
rect 225562 254879 225618 254888
rect 225944 254545 225972 255598
rect 226404 255361 226432 255734
rect 229440 255662 229468 257706
rect 229520 257560 229572 257566
rect 229520 257502 229572 257508
rect 229428 255656 229480 255662
rect 229428 255598 229480 255604
rect 226390 255352 226446 255361
rect 226390 255287 226446 255296
rect 225930 254536 225986 254545
rect 225930 254471 225986 254480
rect 182048 254432 182100 254438
rect 225932 254432 225984 254438
rect 182048 254374 182100 254380
rect 182230 254400 182286 254409
rect 175792 254296 175844 254302
rect 175792 254238 175844 254244
rect 175700 254228 175752 254234
rect 175700 254170 175752 254176
rect 173214 254128 173270 254137
rect 173214 254063 173270 254072
rect 173228 253214 173256 254063
rect 182060 253865 182088 254374
rect 182140 254364 182192 254370
rect 225932 254374 225984 254380
rect 182230 254335 182286 254344
rect 182140 254306 182192 254312
rect 182046 253856 182102 253865
rect 182046 253791 182102 253800
rect 182152 253457 182180 254306
rect 182244 254302 182272 254335
rect 182232 254296 182284 254302
rect 182232 254238 182284 254244
rect 182324 254228 182376 254234
rect 182324 254170 182376 254176
rect 182336 254001 182364 254170
rect 182322 253992 182378 254001
rect 182322 253927 182378 253936
rect 225944 253457 225972 254374
rect 229532 254166 229560 257502
rect 229612 257288 229664 257294
rect 229612 257230 229664 257236
rect 226300 254160 226352 254166
rect 226298 254128 226300 254137
rect 229520 254160 229572 254166
rect 226352 254128 226354 254137
rect 229520 254102 229572 254108
rect 226298 254063 226354 254072
rect 229624 254030 229652 257230
rect 229992 255730 230020 260018
rect 233842 259976 233898 259985
rect 233842 259911 233898 259920
rect 233566 258616 233622 258625
rect 233566 258551 233622 258560
rect 233474 257936 233530 257945
rect 233474 257871 233530 257880
rect 233488 257566 233516 257871
rect 233580 257770 233608 258551
rect 233568 257764 233620 257770
rect 233568 257706 233620 257712
rect 233476 257560 233528 257566
rect 233476 257502 233528 257508
rect 233476 257288 233528 257294
rect 233474 257256 233476 257265
rect 233528 257256 233530 257265
rect 233474 257191 233530 257200
rect 233474 256576 233530 256585
rect 233474 256511 233530 256520
rect 233488 255934 233516 256511
rect 230164 255928 230216 255934
rect 230164 255870 230216 255876
rect 233476 255928 233528 255934
rect 233476 255870 233528 255876
rect 229980 255724 230032 255730
rect 229980 255666 230032 255672
rect 230176 254438 230204 255870
rect 233856 255798 233884 259911
rect 234132 257090 234160 261951
rect 234316 257226 234344 262631
rect 234670 261336 234726 261345
rect 234670 261271 234726 261280
rect 234304 257220 234356 257226
rect 234304 257162 234356 257168
rect 234684 257158 234712 261271
rect 234762 259296 234818 259305
rect 234762 259231 234818 259240
rect 234672 257152 234724 257158
rect 234672 257094 234724 257100
rect 234120 257084 234172 257090
rect 234120 257026 234172 257032
rect 233934 255896 233990 255905
rect 234776 255866 234804 259231
rect 233934 255831 233990 255840
rect 234764 255860 234816 255866
rect 233844 255792 233896 255798
rect 233844 255734 233896 255740
rect 233750 255216 233806 255225
rect 233750 255151 233806 255160
rect 233566 254536 233622 254545
rect 233566 254471 233622 254480
rect 230164 254432 230216 254438
rect 230164 254374 230216 254380
rect 226300 254024 226352 254030
rect 226300 253966 226352 253972
rect 229612 254024 229664 254030
rect 229612 253966 229664 253972
rect 226312 253865 226340 253966
rect 226298 253856 226354 253865
rect 226298 253791 226354 253800
rect 233474 253856 233530 253865
rect 233474 253791 233530 253800
rect 173490 253448 173546 253457
rect 173490 253383 173546 253392
rect 182138 253448 182194 253457
rect 182138 253383 182194 253392
rect 225930 253448 225986 253457
rect 225930 253383 225986 253392
rect 173216 253208 173268 253214
rect 173216 253150 173268 253156
rect 173504 253146 173532 253383
rect 173492 253140 173544 253146
rect 173492 253082 173544 253088
rect 230624 253140 230676 253146
rect 230624 253082 230676 253088
rect 182324 253072 182376 253078
rect 140554 253040 140610 253049
rect 182322 253040 182324 253049
rect 226300 253072 226352 253078
rect 182376 253040 182378 253049
rect 140554 252975 140610 252984
rect 181404 253004 181456 253010
rect 139912 252936 139964 252942
rect 139912 252878 139964 252884
rect 140568 252398 140596 252975
rect 182322 252975 182378 252984
rect 226298 253040 226300 253049
rect 226352 253040 226354 253049
rect 226298 252975 226354 252984
rect 226392 253004 226444 253010
rect 181404 252946 181456 252952
rect 226392 252946 226444 252952
rect 173582 252768 173638 252777
rect 173582 252703 173638 252712
rect 173596 252398 173624 252703
rect 181416 252641 181444 252946
rect 226300 252936 226352 252942
rect 226300 252878 226352 252884
rect 225656 252868 225708 252874
rect 225656 252810 225708 252816
rect 181402 252632 181458 252641
rect 181402 252567 181458 252576
rect 140556 252392 140608 252398
rect 140186 252360 140242 252369
rect 140556 252334 140608 252340
rect 173584 252392 173636 252398
rect 173584 252334 173636 252340
rect 182324 252392 182376 252398
rect 182324 252334 182376 252340
rect 140186 252295 140242 252304
rect 140200 251718 140228 252295
rect 173490 252088 173546 252097
rect 173490 252023 173546 252032
rect 173504 251786 173532 252023
rect 182336 251961 182364 252334
rect 225668 251961 225696 252810
rect 226312 252641 226340 252878
rect 226298 252632 226354 252641
rect 226298 252567 226354 252576
rect 226404 252233 226432 252946
rect 226390 252224 226446 252233
rect 226390 252159 226446 252168
rect 182322 251952 182378 251961
rect 182322 251887 182378 251896
rect 225654 251952 225710 251961
rect 225654 251887 225710 251896
rect 173492 251780 173544 251786
rect 173492 251722 173544 251728
rect 140188 251712 140240 251718
rect 181772 251712 181824 251718
rect 140188 251654 140240 251660
rect 140646 251680 140702 251689
rect 181772 251654 181824 251660
rect 225380 251712 225432 251718
rect 225380 251654 225432 251660
rect 140646 251615 140702 251624
rect 140554 251136 140610 251145
rect 140660 251106 140688 251615
rect 181784 251553 181812 251654
rect 181770 251544 181826 251553
rect 181770 251479 181826 251488
rect 173490 251408 173546 251417
rect 173490 251343 173546 251352
rect 173504 251106 173532 251343
rect 225392 251145 225420 251654
rect 226392 251644 226444 251650
rect 226392 251586 226444 251592
rect 226300 251576 226352 251582
rect 226298 251544 226300 251553
rect 226352 251544 226354 251553
rect 226298 251479 226354 251488
rect 182322 251136 182378 251145
rect 140554 251071 140610 251080
rect 140648 251100 140700 251106
rect 140568 251038 140596 251071
rect 140648 251042 140700 251048
rect 173492 251100 173544 251106
rect 182322 251071 182324 251080
rect 173492 251042 173544 251048
rect 182376 251071 182378 251080
rect 225378 251136 225434 251145
rect 225378 251071 225434 251080
rect 182324 251042 182376 251048
rect 140556 251032 140608 251038
rect 140556 250974 140608 250980
rect 173584 251032 173636 251038
rect 182232 251032 182284 251038
rect 173584 250974 173636 250980
rect 182230 251000 182232 251009
rect 182284 251000 182286 251009
rect 173596 250737 173624 250974
rect 182230 250935 182286 250944
rect 226404 250737 226432 251586
rect 230636 251582 230664 253082
rect 233488 252874 233516 253791
rect 233580 253010 233608 254471
rect 233658 253176 233714 253185
rect 233658 253111 233660 253120
rect 233712 253111 233714 253120
rect 233660 253082 233712 253088
rect 233568 253004 233620 253010
rect 233568 252946 233620 252952
rect 233764 252942 233792 255151
rect 233948 253078 233976 255831
rect 234764 255802 234816 255808
rect 233936 253072 233988 253078
rect 233936 253014 233988 253020
rect 233752 252936 233804 252942
rect 233752 252878 233804 252884
rect 233476 252868 233528 252874
rect 233476 252810 233528 252816
rect 233566 252496 233622 252505
rect 233566 252431 233622 252440
rect 233474 251816 233530 251825
rect 233474 251751 233530 251760
rect 233488 251650 233516 251751
rect 233580 251718 233608 252431
rect 233568 251712 233620 251718
rect 233568 251654 233620 251660
rect 233476 251644 233528 251650
rect 233476 251586 233528 251592
rect 230624 251576 230676 251582
rect 230624 251518 230676 251524
rect 233566 251136 233622 251145
rect 233566 251071 233622 251080
rect 173582 250728 173638 250737
rect 173582 250663 173638 250672
rect 226390 250728 226446 250737
rect 226390 250663 226446 250672
rect 140554 250456 140610 250465
rect 140554 250391 140610 250400
rect 233474 250456 233530 250465
rect 233474 250391 233530 250400
rect 140568 250290 140596 250391
rect 175424 250352 175476 250358
rect 175424 250294 175476 250300
rect 182230 250320 182286 250329
rect 140556 250284 140608 250290
rect 140556 250226 140608 250232
rect 173674 250184 173730 250193
rect 173674 250119 173730 250128
rect 140002 249776 140058 249785
rect 140002 249711 140058 249720
rect 140016 249610 140044 249711
rect 140464 249672 140516 249678
rect 140462 249640 140464 249649
rect 173584 249672 173636 249678
rect 140516 249640 140518 249649
rect 140004 249604 140056 249610
rect 173584 249614 173636 249620
rect 140462 249575 140518 249584
rect 140004 249546 140056 249552
rect 173596 249513 173624 249614
rect 173688 249610 173716 250119
rect 173676 249604 173728 249610
rect 173676 249546 173728 249552
rect 173582 249504 173638 249513
rect 173582 249439 173638 249448
rect 140372 248924 140424 248930
rect 140372 248866 140424 248872
rect 173216 248924 173268 248930
rect 173216 248866 173268 248872
rect 140384 248833 140412 248866
rect 173228 248833 173256 248866
rect 173584 248856 173636 248862
rect 140370 248824 140426 248833
rect 140370 248759 140426 248768
rect 173214 248824 173270 248833
rect 173584 248798 173636 248804
rect 173214 248759 173270 248768
rect 140372 248244 140424 248250
rect 140372 248186 140424 248192
rect 140384 248153 140412 248186
rect 173596 248153 173624 248798
rect 140370 248144 140426 248153
rect 140370 248079 140426 248088
rect 173582 248144 173638 248153
rect 173582 248079 173638 248088
rect 137060 247768 137112 247774
rect 137060 247710 137112 247716
rect 137072 246142 137100 247710
rect 137520 247700 137572 247706
rect 137520 247642 137572 247648
rect 137532 247298 137560 247642
rect 140372 247564 140424 247570
rect 140372 247506 140424 247512
rect 173216 247564 173268 247570
rect 173216 247506 173268 247512
rect 140384 247473 140412 247506
rect 173228 247473 173256 247506
rect 173584 247496 173636 247502
rect 140370 247464 140426 247473
rect 140370 247399 140426 247408
rect 173214 247464 173270 247473
rect 173584 247438 173636 247444
rect 173214 247399 173270 247408
rect 137520 247292 137572 247298
rect 137520 247234 137572 247240
rect 140648 247292 140700 247298
rect 140648 247234 140700 247240
rect 140660 247065 140688 247234
rect 140646 247056 140702 247065
rect 140646 246991 140702 247000
rect 173596 246793 173624 247438
rect 173582 246784 173638 246793
rect 173582 246719 173638 246728
rect 137244 246408 137296 246414
rect 137244 246350 137296 246356
rect 173952 246408 174004 246414
rect 173952 246350 174004 246356
rect 137060 246136 137112 246142
rect 137060 246078 137112 246084
rect 137256 246006 137284 246350
rect 140648 246340 140700 246346
rect 140648 246282 140700 246288
rect 140188 246272 140240 246278
rect 140188 246214 140240 246220
rect 137244 246000 137296 246006
rect 137244 245942 137296 245948
rect 135956 245048 136008 245054
rect 135956 244990 136008 244996
rect 135864 244980 135916 244986
rect 135864 244922 135916 244928
rect 135876 242062 135904 244922
rect 135864 242056 135916 242062
rect 135864 241998 135916 242004
rect 135968 241994 135996 244990
rect 139636 244912 139688 244918
rect 139636 244854 139688 244860
rect 136784 243688 136836 243694
rect 136784 243630 136836 243636
rect 136692 243620 136744 243626
rect 136692 243562 136744 243568
rect 136140 242260 136192 242266
rect 136140 242202 136192 242208
rect 135956 241988 136008 241994
rect 135956 241930 136008 241936
rect 136152 237574 136180 242202
rect 136232 242192 136284 242198
rect 136232 242134 136284 242140
rect 136244 237846 136272 242134
rect 136704 239206 136732 243562
rect 136796 239274 136824 243630
rect 139360 243552 139412 243558
rect 139360 243494 139412 243500
rect 139268 240696 139320 240702
rect 139268 240638 139320 240644
rect 136784 239268 136836 239274
rect 136784 239210 136836 239216
rect 136692 239200 136744 239206
rect 136692 239142 136744 239148
rect 136232 237840 136284 237846
rect 136232 237782 136284 237788
rect 136140 237568 136192 237574
rect 136140 237510 136192 237516
rect 139280 236457 139308 240638
rect 139372 240401 139400 243494
rect 139544 243484 139596 243490
rect 139544 243426 139596 243432
rect 139452 242124 139504 242130
rect 139452 242066 139504 242072
rect 139358 240392 139414 240401
rect 139358 240327 139414 240336
rect 139464 238633 139492 242066
rect 139556 240673 139584 243426
rect 139648 243257 139676 244854
rect 139728 244844 139780 244850
rect 139728 244786 139780 244792
rect 139634 243248 139690 243257
rect 139634 243183 139690 243192
rect 139740 243121 139768 244786
rect 140200 244481 140228 246214
rect 140556 246136 140608 246142
rect 140554 246104 140556 246113
rect 140608 246104 140610 246113
rect 140554 246039 140610 246048
rect 140372 246000 140424 246006
rect 140372 245942 140424 245948
rect 140384 245569 140412 245942
rect 140370 245560 140426 245569
rect 140370 245495 140426 245504
rect 140660 244617 140688 246282
rect 173584 246136 173636 246142
rect 173582 246104 173584 246113
rect 173636 246104 173638 246113
rect 173582 246039 173638 246048
rect 173492 245728 173544 245734
rect 173492 245670 173544 245676
rect 173504 245433 173532 245670
rect 173490 245424 173546 245433
rect 173490 245359 173546 245368
rect 173584 244776 173636 244782
rect 173582 244744 173584 244753
rect 173636 244744 173638 244753
rect 172848 244708 172900 244714
rect 173582 244679 173638 244688
rect 172848 244650 172900 244656
rect 140646 244608 140702 244617
rect 140646 244543 140702 244552
rect 140186 244472 140242 244481
rect 140186 244407 140242 244416
rect 172860 244073 172888 244650
rect 172846 244064 172902 244073
rect 172846 243999 172902 244008
rect 173860 243552 173912 243558
rect 173860 243494 173912 243500
rect 173492 243484 173544 243490
rect 173492 243426 173544 243432
rect 139726 243112 139782 243121
rect 139726 243047 139782 243056
rect 172848 242804 172900 242810
rect 172848 242746 172900 242752
rect 172860 242169 172888 242746
rect 172846 242160 172902 242169
rect 172846 242095 172902 242104
rect 140556 242056 140608 242062
rect 140554 242024 140556 242033
rect 140608 242024 140610 242033
rect 140188 241988 140240 241994
rect 140554 241959 140610 241968
rect 140188 241930 140240 241936
rect 140200 241897 140228 241930
rect 140186 241888 140242 241897
rect 140186 241823 140242 241832
rect 139542 240664 139598 240673
rect 139542 240599 139598 240608
rect 141014 240528 141070 240537
rect 141014 240463 141016 240472
rect 141068 240463 141070 240472
rect 141016 240434 141068 240440
rect 173504 240129 173532 243426
rect 173584 243212 173636 243218
rect 173584 243154 173636 243160
rect 173596 242849 173624 243154
rect 173582 242840 173638 242849
rect 173582 242775 173638 242784
rect 173768 242260 173820 242266
rect 173768 242202 173820 242208
rect 173584 242056 173636 242062
rect 173584 241998 173636 242004
rect 173596 241489 173624 241998
rect 173676 241988 173728 241994
rect 173676 241930 173728 241936
rect 173582 241480 173638 241489
rect 173582 241415 173638 241424
rect 173688 240809 173716 241930
rect 173674 240800 173730 240809
rect 173674 240735 173730 240744
rect 173490 240120 173546 240129
rect 173490 240055 173546 240064
rect 140554 239304 140610 239313
rect 140554 239239 140556 239248
rect 140608 239239 140610 239248
rect 173676 239268 173728 239274
rect 140556 239210 140608 239216
rect 173676 239210 173728 239216
rect 140648 239200 140700 239206
rect 140646 239168 140648 239177
rect 140700 239168 140702 239177
rect 140646 239103 140702 239112
rect 173688 238769 173716 239210
rect 173674 238760 173730 238769
rect 173674 238695 173730 238704
rect 139450 238624 139506 238633
rect 139450 238559 139506 238568
rect 173780 238089 173808 242202
rect 173872 239449 173900 243494
rect 173964 243393 173992 246350
rect 175436 243626 175464 250294
rect 182230 250255 182286 250264
rect 226298 250320 226354 250329
rect 226298 250255 226300 250264
rect 181586 249640 181642 249649
rect 182244 249610 182272 250255
rect 226352 250255 226354 250264
rect 226300 250226 226352 250232
rect 233488 250222 233516 250391
rect 233580 250290 233608 251071
rect 233568 250284 233620 250290
rect 233568 250226 233620 250232
rect 225932 250216 225984 250222
rect 225932 250158 225984 250164
rect 233476 250216 233528 250222
rect 233476 250158 233528 250164
rect 225944 250057 225972 250158
rect 182322 250048 182378 250057
rect 182322 249983 182378 249992
rect 225930 250048 225986 250057
rect 225930 249983 225986 249992
rect 182336 249678 182364 249983
rect 233474 249776 233530 249785
rect 233474 249711 233530 249720
rect 182324 249672 182376 249678
rect 182324 249614 182376 249620
rect 225564 249672 225616 249678
rect 225564 249614 225616 249620
rect 226298 249640 226354 249649
rect 181586 249575 181642 249584
rect 182232 249604 182284 249610
rect 181600 248930 181628 249575
rect 182232 249546 182284 249552
rect 225576 249241 225604 249614
rect 233488 249610 233516 249711
rect 233568 249672 233620 249678
rect 233566 249640 233568 249649
rect 233620 249640 233622 249649
rect 226298 249575 226300 249584
rect 226352 249575 226354 249584
rect 233476 249604 233528 249610
rect 226300 249546 226352 249552
rect 233566 249575 233622 249584
rect 233476 249546 233528 249552
rect 182322 249232 182378 249241
rect 182322 249167 182378 249176
rect 225562 249232 225618 249241
rect 225562 249167 225618 249176
rect 181588 248924 181640 248930
rect 181588 248866 181640 248872
rect 182336 248862 182364 249167
rect 182324 248856 182376 248862
rect 181126 248824 181182 248833
rect 182324 248798 182376 248804
rect 226390 248824 226446 248833
rect 181126 248759 181182 248768
rect 226390 248759 226446 248768
rect 181034 248416 181090 248425
rect 181034 248351 181090 248360
rect 180850 248008 180906 248017
rect 180850 247943 180906 247952
rect 180758 247192 180814 247201
rect 180758 247127 180814 247136
rect 180666 246784 180722 246793
rect 180666 246719 180722 246728
rect 180680 244714 180708 246719
rect 180772 244782 180800 247127
rect 180864 246142 180892 247943
rect 180942 247600 180998 247609
rect 180942 247535 180998 247544
rect 180852 246136 180904 246142
rect 180852 246078 180904 246084
rect 180850 245968 180906 245977
rect 180850 245903 180906 245912
rect 180760 244776 180812 244782
rect 180760 244718 180812 244724
rect 180668 244708 180720 244714
rect 180668 244650 180720 244656
rect 175424 243620 175476 243626
rect 175424 243562 175476 243568
rect 175332 243416 175384 243422
rect 173950 243384 174006 243393
rect 175332 243358 175384 243364
rect 173950 243319 174006 243328
rect 173858 239440 173914 239449
rect 173858 239375 173914 239384
rect 173766 238080 173822 238089
rect 173766 238015 173822 238024
rect 140556 237840 140608 237846
rect 140556 237782 140608 237788
rect 140280 237568 140332 237574
rect 140280 237510 140332 237516
rect 140292 237273 140320 237510
rect 140568 237409 140596 237782
rect 173584 237432 173636 237438
rect 140554 237400 140610 237409
rect 140554 237335 140610 237344
rect 173582 237400 173584 237409
rect 173636 237400 173638 237409
rect 173582 237335 173638 237344
rect 140278 237264 140334 237273
rect 140278 237199 140334 237208
rect 173400 236956 173452 236962
rect 173400 236898 173452 236904
rect 173412 236729 173440 236898
rect 173398 236720 173454 236729
rect 173398 236655 173454 236664
rect 173584 236548 173636 236554
rect 173584 236490 173636 236496
rect 139266 236448 139322 236457
rect 139266 236383 139322 236392
rect 173596 236185 173624 236490
rect 173582 236176 173638 236185
rect 173582 236111 173638 236120
rect 142868 235862 143204 235890
rect 143756 235862 143816 235890
rect 142868 233562 142896 235862
rect 138164 233556 138216 233562
rect 138164 233498 138216 233504
rect 142856 233556 142908 233562
rect 142856 233498 142908 233504
rect 137980 233488 138032 233494
rect 137980 233430 138032 233436
rect 137888 233420 137940 233426
rect 137888 233362 137940 233368
rect 137796 233216 137848 233222
rect 137796 233158 137848 233164
rect 137612 233080 137664 233086
rect 137612 233022 137664 233028
rect 137518 225568 137574 225577
rect 137518 225503 137574 225512
rect 137428 218664 137480 218670
rect 137428 218606 137480 218612
rect 137336 215876 137388 215882
rect 137336 215818 137388 215824
rect 137152 213156 137204 213162
rect 137152 213098 137204 213104
rect 134574 211832 134630 211841
rect 134220 211790 134574 211818
rect 74038 202856 74094 202865
rect 74038 202791 74094 202800
rect 51958 202176 52014 202185
rect 51958 202111 52014 202120
rect 38158 194696 38214 194705
rect 38158 194631 38214 194640
rect 38172 172362 38200 194631
rect 74052 190994 74080 202791
rect 74040 190988 74092 190994
rect 74040 190930 74092 190936
rect 81676 190988 81728 190994
rect 81676 190930 81728 190936
rect 81688 190489 81716 190930
rect 81674 190480 81730 190489
rect 81674 190415 81730 190424
rect 51314 189528 51370 189537
rect 51314 189463 51370 189472
rect 51328 188274 51356 189463
rect 47084 188268 47136 188274
rect 47084 188210 47136 188216
rect 51316 188268 51368 188274
rect 51316 188210 51368 188216
rect 47096 186846 47124 188210
rect 38804 186840 38856 186846
rect 38802 186808 38804 186817
rect 47084 186840 47136 186846
rect 38856 186808 38858 186817
rect 47084 186782 47136 186788
rect 38802 186743 38858 186752
rect 53984 180992 54036 180998
rect 53984 180934 54036 180940
rect 49844 180720 49896 180726
rect 49844 180662 49896 180668
rect 38160 172356 38212 172362
rect 38160 172298 38212 172304
rect 49200 172356 49252 172362
rect 49200 172298 49252 172304
rect 49212 169780 49240 172298
rect 49856 169780 49884 180662
rect 51132 180652 51184 180658
rect 51132 180594 51184 180600
rect 50488 172560 50540 172566
rect 50488 172502 50540 172508
rect 50500 169780 50528 172502
rect 51144 169794 51172 180594
rect 52512 180516 52564 180522
rect 52512 180458 52564 180464
rect 51224 175484 51276 175490
rect 51224 175426 51276 175432
rect 51236 172566 51264 175426
rect 51224 172560 51276 172566
rect 51224 172502 51276 172508
rect 51144 169766 51250 169794
rect 52524 169658 52552 180458
rect 52604 180448 52656 180454
rect 52604 180390 52656 180396
rect 52616 169780 52644 180390
rect 53248 171744 53300 171750
rect 53248 171686 53300 171692
rect 53260 169780 53288 171686
rect 53996 169794 54024 180934
rect 55100 180250 55128 182836
rect 55468 181066 55496 182836
rect 55836 181338 55864 182836
rect 55824 181332 55876 181338
rect 55824 181274 55876 181280
rect 55456 181060 55508 181066
rect 55456 181002 55508 181008
rect 56296 180658 56324 182836
rect 56664 180862 56692 182836
rect 56652 180856 56704 180862
rect 56652 180798 56704 180804
rect 56284 180652 56336 180658
rect 56284 180594 56336 180600
rect 57032 180386 57060 182836
rect 57020 180380 57072 180386
rect 57020 180322 57072 180328
rect 55088 180244 55140 180250
rect 55088 180186 55140 180192
rect 57492 180046 57520 182836
rect 57572 180108 57624 180114
rect 57572 180050 57624 180056
rect 57480 180040 57532 180046
rect 57480 179982 57532 179988
rect 57296 172764 57348 172770
rect 57296 172706 57348 172712
rect 54628 172628 54680 172634
rect 54628 172570 54680 172576
rect 53918 169766 54024 169794
rect 54640 169780 54668 172570
rect 55272 172084 55324 172090
rect 55272 172026 55324 172032
rect 55284 169780 55312 172026
rect 56008 172016 56060 172022
rect 56008 171958 56060 171964
rect 56020 169780 56048 171958
rect 56652 171812 56704 171818
rect 56652 171754 56704 171760
rect 56664 169780 56692 171754
rect 57308 169780 57336 172706
rect 57584 171750 57612 180050
rect 57860 179978 57888 182836
rect 58228 180726 58256 182836
rect 58688 180930 58716 182836
rect 59056 181134 59084 182836
rect 59438 182822 59544 182850
rect 59044 181128 59096 181134
rect 59044 181070 59096 181076
rect 58676 180924 58728 180930
rect 58676 180866 58728 180872
rect 58216 180720 58268 180726
rect 58216 180662 58268 180668
rect 57848 179972 57900 179978
rect 57848 179914 57900 179920
rect 59412 172968 59464 172974
rect 59412 172910 59464 172916
rect 58676 172900 58728 172906
rect 58676 172842 58728 172848
rect 58032 172696 58084 172702
rect 58032 172638 58084 172644
rect 57572 171744 57624 171750
rect 57572 171686 57624 171692
rect 58044 169780 58072 172638
rect 58688 169780 58716 172842
rect 59424 169780 59452 172910
rect 59516 172673 59544 182822
rect 59884 181202 59912 182836
rect 60266 182822 60556 182850
rect 60634 182822 60924 182850
rect 59872 181196 59924 181202
rect 59872 181138 59924 181144
rect 60528 180538 60556 182822
rect 60528 180510 60740 180538
rect 60608 180380 60660 180386
rect 60608 180322 60660 180328
rect 60148 180244 60200 180250
rect 60148 180186 60200 180192
rect 60424 180244 60476 180250
rect 60424 180186 60476 180192
rect 60056 180176 60108 180182
rect 60056 180118 60108 180124
rect 59502 172664 59558 172673
rect 59502 172599 59558 172608
rect 60068 171818 60096 180118
rect 60160 178906 60188 180186
rect 60240 180040 60292 180046
rect 60240 179982 60292 179988
rect 60252 179042 60280 179982
rect 60252 179014 60372 179042
rect 60160 178878 60280 178906
rect 60252 172226 60280 178878
rect 60344 172294 60372 179014
rect 60332 172288 60384 172294
rect 60332 172230 60384 172236
rect 60240 172220 60292 172226
rect 60240 172162 60292 172168
rect 60436 172022 60464 180186
rect 60516 179836 60568 179842
rect 60516 179778 60568 179784
rect 60528 172838 60556 179778
rect 60516 172832 60568 172838
rect 60516 172774 60568 172780
rect 60620 172090 60648 180322
rect 60712 172537 60740 180510
rect 60792 173036 60844 173042
rect 60792 172978 60844 172984
rect 60698 172528 60754 172537
rect 60698 172463 60754 172472
rect 60608 172084 60660 172090
rect 60608 172026 60660 172032
rect 60424 172016 60476 172022
rect 60424 171958 60476 171964
rect 60056 171812 60108 171818
rect 60056 171754 60108 171760
rect 60056 171676 60108 171682
rect 60056 171618 60108 171624
rect 60068 169780 60096 171618
rect 60804 169780 60832 172978
rect 60896 172809 60924 182822
rect 61080 179978 61108 182836
rect 61462 182822 61752 182850
rect 61830 182822 62212 182850
rect 61724 180130 61752 182822
rect 62080 181264 62132 181270
rect 62080 181206 62132 181212
rect 61724 180102 62028 180130
rect 61068 179972 61120 179978
rect 61068 179914 61120 179920
rect 61804 179972 61856 179978
rect 61804 179914 61856 179920
rect 61896 179972 61948 179978
rect 61896 179914 61948 179920
rect 60882 172800 60938 172809
rect 60882 172735 60938 172744
rect 61816 172430 61844 179914
rect 61804 172424 61856 172430
rect 61908 172401 61936 179914
rect 62000 172566 62028 180102
rect 61988 172560 62040 172566
rect 61988 172502 62040 172508
rect 61804 172366 61856 172372
rect 61894 172392 61950 172401
rect 61894 172327 61950 172336
rect 62092 170202 62120 181206
rect 62184 172265 62212 182822
rect 62276 179978 62304 182836
rect 62644 179978 62672 182836
rect 63104 180590 63132 182836
rect 63472 180794 63500 182836
rect 63840 181406 63868 182836
rect 63828 181400 63880 181406
rect 63828 181342 63880 181348
rect 63736 181332 63788 181338
rect 63736 181274 63788 181280
rect 63460 180788 63512 180794
rect 63460 180730 63512 180736
rect 63552 180720 63604 180726
rect 63552 180662 63604 180668
rect 63092 180584 63144 180590
rect 63092 180526 63144 180532
rect 63092 180380 63144 180386
rect 63092 180322 63144 180328
rect 63000 180176 63052 180182
rect 63000 180118 63052 180124
rect 62264 179972 62316 179978
rect 62264 179914 62316 179920
rect 62632 179972 62684 179978
rect 62632 179914 62684 179920
rect 62264 179836 62316 179842
rect 62264 179778 62316 179784
rect 62170 172256 62226 172265
rect 62170 172191 62226 172200
rect 61908 170174 62120 170202
rect 61908 169658 61936 170174
rect 62276 169794 62304 179778
rect 63012 172906 63040 180118
rect 63104 172974 63132 180322
rect 63092 172968 63144 172974
rect 63092 172910 63144 172916
rect 63000 172900 63052 172906
rect 63000 172842 63052 172848
rect 63564 169930 63592 180662
rect 63748 180130 63776 181274
rect 64300 180522 64328 182836
rect 64288 180516 64340 180522
rect 64288 180458 64340 180464
rect 64668 180454 64696 182836
rect 64656 180448 64708 180454
rect 64656 180390 64708 180396
rect 63748 180102 63868 180130
rect 65036 180114 65064 182836
rect 65496 180998 65524 182836
rect 65484 180992 65536 180998
rect 65484 180934 65536 180940
rect 65116 180856 65168 180862
rect 65116 180798 65168 180804
rect 63736 180040 63788 180046
rect 63736 179982 63788 179988
rect 63644 179972 63696 179978
rect 63644 179914 63696 179920
rect 63656 172362 63684 179914
rect 63644 172356 63696 172362
rect 63644 172298 63696 172304
rect 63644 172220 63696 172226
rect 63644 172162 63696 172168
rect 62106 169766 62304 169794
rect 63380 169902 63592 169930
rect 63380 169658 63408 169902
rect 63656 169794 63684 172162
rect 63486 169766 63684 169794
rect 63748 169794 63776 179982
rect 63840 171562 63868 180102
rect 65024 180108 65076 180114
rect 65024 180050 65076 180056
rect 64472 180040 64524 180046
rect 64472 179982 64524 179988
rect 64380 179972 64432 179978
rect 64380 179914 64432 179920
rect 64392 171750 64420 179914
rect 64484 173042 64512 179982
rect 65128 175150 65156 180798
rect 65208 180652 65260 180658
rect 65208 180594 65260 180600
rect 65116 175144 65168 175150
rect 65116 175086 65168 175092
rect 64472 173036 64524 173042
rect 64472 172978 64524 172984
rect 65116 172288 65168 172294
rect 65116 172230 65168 172236
rect 65128 172158 65156 172230
rect 65116 172152 65168 172158
rect 65116 172094 65168 172100
rect 64380 171744 64432 171750
rect 64380 171686 64432 171692
rect 63840 171534 64512 171562
rect 64484 169794 64512 171534
rect 65220 169794 65248 180594
rect 65760 180584 65812 180590
rect 65760 180526 65812 180532
rect 65576 175484 65628 175490
rect 65576 175426 65628 175432
rect 65588 172634 65616 175426
rect 65772 175370 65800 180526
rect 65864 175490 65892 182836
rect 65852 175484 65904 175490
rect 65852 175426 65904 175432
rect 65772 175342 65984 175370
rect 65852 175144 65904 175150
rect 65852 175086 65904 175092
rect 65576 172628 65628 172634
rect 65576 172570 65628 172576
rect 65864 169794 65892 175086
rect 65956 173042 65984 175342
rect 65944 173036 65996 173042
rect 65944 172978 65996 172984
rect 66232 172294 66260 182836
rect 66692 180250 66720 182836
rect 67060 180930 67088 182836
rect 67048 180924 67100 180930
rect 67048 180866 67100 180872
rect 66680 180244 66732 180250
rect 66680 180186 66732 180192
rect 67428 172770 67456 182836
rect 67416 172764 67468 172770
rect 67416 172706 67468 172712
rect 67888 172702 67916 182836
rect 68256 180182 68284 182836
rect 68624 180386 68652 182836
rect 68612 180380 68664 180386
rect 68612 180322 68664 180328
rect 68244 180176 68296 180182
rect 68244 180118 68296 180124
rect 69084 179978 69112 182836
rect 69348 181128 69400 181134
rect 69348 181070 69400 181076
rect 69256 181060 69308 181066
rect 69256 181002 69308 181008
rect 69072 179972 69124 179978
rect 69072 179914 69124 179920
rect 68980 173036 69032 173042
rect 68980 172978 69032 172984
rect 68244 172832 68296 172838
rect 68244 172774 68296 172780
rect 67876 172696 67928 172702
rect 67876 172638 67928 172644
rect 66220 172288 66272 172294
rect 66220 172230 66272 172236
rect 67600 172220 67652 172226
rect 67600 172162 67652 172168
rect 66864 172084 66916 172090
rect 66864 172026 66916 172032
rect 63748 169766 64222 169794
rect 64484 169766 64866 169794
rect 65220 169766 65510 169794
rect 65864 169766 66246 169794
rect 66876 169780 66904 172026
rect 67612 169780 67640 172162
rect 68256 169780 68284 172774
rect 68992 169780 69020 172978
rect 69268 169794 69296 181002
rect 69360 169930 69388 181070
rect 69452 180046 69480 182836
rect 69820 181270 69848 182836
rect 69808 181264 69860 181270
rect 69808 181206 69860 181212
rect 69900 181196 69952 181202
rect 69900 181138 69952 181144
rect 69440 180040 69492 180046
rect 69440 179982 69492 179988
rect 69912 173042 69940 181138
rect 70280 180318 70308 182836
rect 70648 180726 70676 182836
rect 70636 180720 70688 180726
rect 70636 180662 70688 180668
rect 70268 180312 70320 180318
rect 70268 180254 70320 180260
rect 88208 178000 88260 178006
rect 134220 177954 134248 211790
rect 134574 211767 134630 211776
rect 137060 209008 137112 209014
rect 137060 208950 137112 208956
rect 136968 204860 137020 204866
rect 136968 204802 137020 204808
rect 136980 192665 137008 204802
rect 137072 195793 137100 208950
rect 137164 198921 137192 213098
rect 137244 211728 137296 211734
rect 137244 211670 137296 211676
rect 137150 198912 137206 198921
rect 137150 198847 137206 198856
rect 137256 197425 137284 211670
rect 137348 200553 137376 215818
rect 137440 202049 137468 218606
rect 137426 202040 137482 202049
rect 137426 201975 137482 201984
rect 137334 200544 137390 200553
rect 137334 200479 137390 200488
rect 137242 197416 137298 197425
rect 137242 197351 137298 197360
rect 137058 195784 137114 195793
rect 137058 195719 137114 195728
rect 137428 195136 137480 195142
rect 137428 195078 137480 195084
rect 137440 194297 137468 195078
rect 137426 194288 137482 194297
rect 137426 194223 137482 194232
rect 136966 192656 137022 192665
rect 136966 192591 137022 192600
rect 137426 191160 137482 191169
rect 137426 191095 137428 191104
rect 137480 191095 137482 191104
rect 137428 191066 137480 191072
rect 137060 189696 137112 189702
rect 137060 189638 137112 189644
rect 137072 183281 137100 189638
rect 137426 189528 137482 189537
rect 137426 189463 137482 189472
rect 137440 189430 137468 189463
rect 137428 189424 137480 189430
rect 137428 189366 137480 189372
rect 137336 188268 137388 188274
rect 137336 188210 137388 188216
rect 137058 183272 137114 183281
rect 137058 183207 137114 183216
rect 137348 181785 137376 188210
rect 137428 188200 137480 188206
rect 137428 188142 137480 188148
rect 137440 188041 137468 188142
rect 137426 188032 137482 188041
rect 137426 187967 137482 187976
rect 137428 186840 137480 186846
rect 137428 186782 137480 186788
rect 137440 186409 137468 186782
rect 137426 186400 137482 186409
rect 137426 186335 137482 186344
rect 137426 184632 137482 184641
rect 137426 184567 137482 184576
rect 137440 184262 137468 184567
rect 137428 184256 137480 184262
rect 137428 184198 137480 184204
rect 137334 181776 137390 181785
rect 137334 181711 137390 181720
rect 137426 180144 137482 180153
rect 137426 180079 137482 180088
rect 137440 180046 137468 180079
rect 137428 180040 137480 180046
rect 137428 179982 137480 179988
rect 137428 179904 137480 179910
rect 137428 179846 137480 179852
rect 137440 178657 137468 179846
rect 137426 178648 137482 178657
rect 137426 178583 137482 178592
rect 88208 177942 88260 177948
rect 88220 177940 88248 177942
rect 134142 177940 134248 177954
rect 85552 175830 85580 177940
rect 86840 177938 86868 177940
rect 86828 177932 86880 177938
rect 86828 177874 86880 177880
rect 87104 177796 87156 177802
rect 87104 177738 87156 177744
rect 88484 177796 88536 177802
rect 88484 177738 88536 177744
rect 85540 175824 85592 175830
rect 85540 175766 85592 175772
rect 79744 175620 79796 175626
rect 79744 175562 79796 175568
rect 79560 175552 79612 175558
rect 79560 175494 79612 175500
rect 69900 173036 69952 173042
rect 69900 172978 69952 172984
rect 71648 173036 71700 173042
rect 71648 172978 71700 172984
rect 71002 172664 71058 172673
rect 71002 172599 71058 172608
rect 69360 169902 69756 169930
rect 69268 169766 69650 169794
rect 51894 169630 52552 169658
rect 61462 169630 61936 169658
rect 62842 169630 63408 169658
rect 69728 169658 69756 169902
rect 71016 169780 71044 172599
rect 71660 169780 71688 172978
rect 73026 172800 73082 172809
rect 73026 172735 73082 172744
rect 72382 172528 72438 172537
rect 72382 172463 72438 172472
rect 72396 169780 72424 172463
rect 73040 169780 73068 172735
rect 74408 172560 74460 172566
rect 74408 172502 74460 172508
rect 73672 172424 73724 172430
rect 73672 172366 73724 172372
rect 73684 169780 73712 172366
rect 74420 169780 74448 172502
rect 75786 172392 75842 172401
rect 75786 172327 75842 172336
rect 76432 172356 76484 172362
rect 75050 172256 75106 172265
rect 75050 172191 75106 172200
rect 75064 169780 75092 172191
rect 75800 169780 75828 172327
rect 76432 172298 76484 172304
rect 76444 169780 76472 172298
rect 69728 169630 70294 169658
rect 76536 166242 76748 166258
rect 76536 166236 76760 166242
rect 76536 166230 76708 166236
rect 46990 162872 47046 162881
rect 46990 162807 47046 162816
rect 47004 144113 47032 162807
rect 76536 160546 76564 166230
rect 76708 166178 76760 166184
rect 79572 166009 79600 175494
rect 79652 175484 79704 175490
rect 79652 175426 79704 175432
rect 79664 166689 79692 175426
rect 79650 166680 79706 166689
rect 79650 166615 79706 166624
rect 79558 166000 79614 166009
rect 79558 165935 79614 165944
rect 79756 165465 79784 175562
rect 79836 175416 79888 175422
rect 79836 175358 79888 175364
rect 79848 167233 79876 175358
rect 79928 175348 79980 175354
rect 79928 175290 79980 175296
rect 79940 168457 79968 175290
rect 80204 175280 80256 175286
rect 80204 175222 80256 175228
rect 80020 175212 80072 175218
rect 80020 175154 80072 175160
rect 80032 169545 80060 175154
rect 80112 175144 80164 175150
rect 80112 175086 80164 175092
rect 80018 169536 80074 169545
rect 80018 169471 80074 169480
rect 79926 168448 79982 168457
rect 79926 168383 79982 168392
rect 80124 167777 80152 175086
rect 80216 169001 80244 175222
rect 85552 174713 85580 175766
rect 85538 174704 85594 174713
rect 85538 174639 85594 174648
rect 80202 168992 80258 169001
rect 80202 168927 80258 168936
rect 80110 167768 80166 167777
rect 80110 167703 80166 167712
rect 79834 167224 79890 167233
rect 79834 167159 79890 167168
rect 87116 166854 87144 177738
rect 87104 166848 87156 166854
rect 87104 166790 87156 166796
rect 88496 166514 88524 177738
rect 89600 174946 89628 177940
rect 90888 177938 90916 177940
rect 90876 177932 90928 177938
rect 90876 177874 90928 177880
rect 91244 177796 91296 177802
rect 91244 177738 91296 177744
rect 89588 174940 89640 174946
rect 89588 174882 89640 174888
rect 91256 166854 91284 177738
rect 92268 175082 92296 177940
rect 92256 175076 92308 175082
rect 92256 175018 92308 175024
rect 93648 175014 93676 177940
rect 94936 175762 94964 177940
rect 94924 175756 94976 175762
rect 94924 175698 94976 175704
rect 93636 175008 93688 175014
rect 93636 174950 93688 174956
rect 95476 174940 95528 174946
rect 95476 174882 95528 174888
rect 90692 166848 90744 166854
rect 90692 166790 90744 166796
rect 91244 166848 91296 166854
rect 91244 166790 91296 166796
rect 88484 166508 88536 166514
rect 88484 166450 88536 166456
rect 79742 165456 79798 165465
rect 79742 165391 79798 165400
rect 80202 164912 80258 164921
rect 80202 164847 80258 164856
rect 80216 164814 80244 164847
rect 80204 164808 80256 164814
rect 80204 164750 80256 164756
rect 87196 164740 87248 164746
rect 87196 164682 87248 164688
rect 87208 164377 87236 164682
rect 87194 164368 87250 164377
rect 87194 164303 87250 164312
rect 80202 164096 80258 164105
rect 80202 164031 80258 164040
rect 80216 163930 80244 164031
rect 80204 163924 80256 163930
rect 80204 163866 80256 163872
rect 85448 163924 85500 163930
rect 85448 163866 85500 163872
rect 80202 163688 80258 163697
rect 80202 163623 80258 163632
rect 80216 163522 80244 163623
rect 80204 163516 80256 163522
rect 80204 163458 80256 163464
rect 85460 163318 85488 163866
rect 90704 163810 90732 166790
rect 92992 166508 93044 166514
rect 92992 166450 93044 166456
rect 93004 163810 93032 166450
rect 95488 163810 95516 174882
rect 96316 174878 96344 177940
rect 97500 175076 97552 175082
rect 97500 175018 97552 175024
rect 96304 174872 96356 174878
rect 96304 174814 96356 174820
rect 97512 166650 97540 175018
rect 97696 174470 97724 177940
rect 98880 175008 98932 175014
rect 98880 174950 98932 174956
rect 97684 174464 97736 174470
rect 97684 174406 97736 174412
rect 98144 174464 98196 174470
rect 98144 174406 98196 174412
rect 98156 167330 98184 174406
rect 98144 167324 98196 167330
rect 98144 167266 98196 167272
rect 98892 166854 98920 174950
rect 98984 174470 99012 177940
rect 100364 174470 100392 177940
rect 101744 174470 101772 177940
rect 103032 174470 103060 177940
rect 104216 175756 104268 175762
rect 104216 175698 104268 175704
rect 98972 174464 99024 174470
rect 98972 174406 99024 174412
rect 99524 174464 99576 174470
rect 99524 174406 99576 174412
rect 100352 174464 100404 174470
rect 100352 174406 100404 174412
rect 100904 174464 100956 174470
rect 100904 174406 100956 174412
rect 101732 174464 101784 174470
rect 101732 174406 101784 174412
rect 102284 174464 102336 174470
rect 102284 174406 102336 174412
rect 103020 174464 103072 174470
rect 103020 174406 103072 174412
rect 103664 174464 103716 174470
rect 103664 174406 103716 174412
rect 99536 167194 99564 174406
rect 100916 167262 100944 174406
rect 100904 167256 100956 167262
rect 100904 167198 100956 167204
rect 99524 167188 99576 167194
rect 99524 167130 99576 167136
rect 102296 167126 102324 174406
rect 102284 167120 102336 167126
rect 102284 167062 102336 167068
rect 103676 166990 103704 174406
rect 104228 174282 104256 175698
rect 104412 174470 104440 177940
rect 105688 175076 105740 175082
rect 105688 175018 105740 175024
rect 104400 174464 104452 174470
rect 104400 174406 104452 174412
rect 105044 174464 105096 174470
rect 105044 174406 105096 174412
rect 104228 174254 104440 174282
rect 103664 166984 103716 166990
rect 103664 166926 103716 166932
rect 104412 166854 104440 174254
rect 105056 167058 105084 174406
rect 105700 174282 105728 175018
rect 105792 174470 105820 177940
rect 107080 174470 107108 177940
rect 105780 174464 105832 174470
rect 105780 174406 105832 174412
rect 106424 174464 106476 174470
rect 106424 174406 106476 174412
rect 107068 174464 107120 174470
rect 107068 174406 107120 174412
rect 107804 174464 107856 174470
rect 107804 174406 107856 174412
rect 105700 174254 105820 174282
rect 105044 167052 105096 167058
rect 105044 166994 105096 167000
rect 97684 166848 97736 166854
rect 97684 166790 97736 166796
rect 98880 166848 98932 166854
rect 98880 166790 98932 166796
rect 102376 166848 102428 166854
rect 102376 166790 102428 166796
rect 104400 166848 104452 166854
rect 104400 166790 104452 166796
rect 105136 166848 105188 166854
rect 105136 166790 105188 166796
rect 97500 166644 97552 166650
rect 97500 166586 97552 166592
rect 97696 163810 97724 166790
rect 100076 166644 100128 166650
rect 100076 166586 100128 166592
rect 100088 163810 100116 166586
rect 102388 163810 102416 166790
rect 105148 163810 105176 166790
rect 105792 166514 105820 174254
rect 106436 166922 106464 174406
rect 106424 166916 106476 166922
rect 106424 166858 106476 166864
rect 107816 166854 107844 174406
rect 108460 172265 108488 177940
rect 109840 175626 109868 177940
rect 111128 175626 111156 177940
rect 109828 175620 109880 175626
rect 109828 175562 109880 175568
rect 111116 175620 111168 175626
rect 111116 175562 111168 175568
rect 112508 175558 112536 177940
rect 112496 175552 112548 175558
rect 112496 175494 112548 175500
rect 113888 172401 113916 177940
rect 115176 175694 115204 177940
rect 115164 175688 115216 175694
rect 115164 175630 115216 175636
rect 116556 174470 116584 177940
rect 117936 175422 117964 177940
rect 117924 175416 117976 175422
rect 117924 175358 117976 175364
rect 119224 174470 119252 177940
rect 120604 175150 120632 177940
rect 121984 175150 122012 177940
rect 123272 175354 123300 177940
rect 123260 175348 123312 175354
rect 123260 175290 123312 175296
rect 120592 175144 120644 175150
rect 120592 175086 120644 175092
rect 121972 175144 122024 175150
rect 121972 175086 122024 175092
rect 124652 174470 124680 177940
rect 126032 175286 126060 177940
rect 126020 175280 126072 175286
rect 126020 175222 126072 175228
rect 127320 174577 127348 177940
rect 128700 175218 128728 177940
rect 132748 175762 132776 177940
rect 134128 177926 134248 177940
rect 132736 175756 132788 175762
rect 132736 175698 132788 175704
rect 128688 175212 128740 175218
rect 128688 175154 128740 175160
rect 132748 174713 132776 175698
rect 132734 174704 132790 174713
rect 132734 174639 132790 174648
rect 127306 174568 127362 174577
rect 127306 174503 127362 174512
rect 134128 174470 134156 177926
rect 116544 174464 116596 174470
rect 116544 174406 116596 174412
rect 117464 174464 117516 174470
rect 117464 174406 117516 174412
rect 119212 174464 119264 174470
rect 119212 174406 119264 174412
rect 120224 174464 120276 174470
rect 120224 174406 120276 174412
rect 124640 174464 124692 174470
rect 124640 174406 124692 174412
rect 125744 174464 125796 174470
rect 125744 174406 125796 174412
rect 134116 174464 134168 174470
rect 134116 174406 134168 174412
rect 134760 174464 134812 174470
rect 134760 174406 134812 174412
rect 113874 172392 113930 172401
rect 113874 172327 113930 172336
rect 108446 172256 108502 172265
rect 108446 172191 108502 172200
rect 117476 168894 117504 174406
rect 120236 170254 120264 174406
rect 120224 170248 120276 170254
rect 120224 170190 120276 170196
rect 125756 170186 125784 174406
rect 125744 170180 125796 170186
rect 125744 170122 125796 170128
rect 117464 168888 117516 168894
rect 117464 168830 117516 168836
rect 109460 167324 109512 167330
rect 109460 167266 109512 167272
rect 107804 166848 107856 166854
rect 107804 166790 107856 166796
rect 105780 166508 105832 166514
rect 105780 166450 105832 166456
rect 107160 166508 107212 166514
rect 107160 166450 107212 166456
rect 90704 163782 91040 163810
rect 93004 163782 93340 163810
rect 95488 163782 95732 163810
rect 97696 163782 98032 163810
rect 100088 163782 100424 163810
rect 102388 163782 102724 163810
rect 105116 163782 105176 163810
rect 107172 163810 107200 166450
rect 109472 163810 109500 167266
rect 114152 167256 114204 167262
rect 114152 167198 114204 167204
rect 112036 167188 112088 167194
rect 112036 167130 112088 167136
rect 112048 163810 112076 167130
rect 114164 163810 114192 167198
rect 116544 167120 116596 167126
rect 116544 167062 116596 167068
rect 116556 163810 116584 167062
rect 121236 167052 121288 167058
rect 121236 166994 121288 167000
rect 118936 166984 118988 166990
rect 118936 166926 118988 166932
rect 118948 163810 118976 166926
rect 121248 163810 121276 166994
rect 123628 166916 123680 166922
rect 123628 166858 123680 166864
rect 123640 163810 123668 166858
rect 125928 166848 125980 166854
rect 125928 166790 125980 166796
rect 125940 163810 125968 166790
rect 128688 166236 128740 166242
rect 128688 166178 128740 166184
rect 132092 166236 132144 166242
rect 132092 166178 132144 166184
rect 128700 163810 128728 166178
rect 107172 163782 107508 163810
rect 109472 163782 109808 163810
rect 112048 163782 112200 163810
rect 114164 163782 114500 163810
rect 116556 163782 116892 163810
rect 118948 163782 119284 163810
rect 121248 163782 121584 163810
rect 123640 163782 123976 163810
rect 125940 163782 126276 163810
rect 128668 163782 128728 163810
rect 131998 163688 132054 163697
rect 131998 163623 132054 163632
rect 131908 163584 131960 163590
rect 131908 163526 131960 163532
rect 87196 163380 87248 163386
rect 87196 163322 87248 163328
rect 85448 163312 85500 163318
rect 85448 163254 85500 163260
rect 80110 163144 80166 163153
rect 80110 163079 80166 163088
rect 80124 162774 80152 163079
rect 87208 162881 87236 163322
rect 87288 163312 87340 163318
rect 87286 163280 87288 163289
rect 87340 163280 87342 163289
rect 87286 163215 87342 163224
rect 87194 162872 87250 162881
rect 87194 162807 87250 162816
rect 80112 162768 80164 162774
rect 80112 162710 80164 162716
rect 87196 162768 87248 162774
rect 87196 162710 87248 162716
rect 80204 162700 80256 162706
rect 80204 162642 80256 162648
rect 80216 162609 80244 162642
rect 80202 162600 80258 162609
rect 80202 162535 80258 162544
rect 87208 162473 87236 162710
rect 87288 162700 87340 162706
rect 87288 162642 87340 162648
rect 87194 162464 87250 162473
rect 87194 162399 87250 162408
rect 87300 162065 87328 162642
rect 87286 162056 87342 162065
rect 87286 161991 87342 162000
rect 80018 161648 80074 161657
rect 80018 161583 80074 161592
rect 87286 161648 87342 161657
rect 87286 161583 87342 161592
rect 80032 161346 80060 161583
rect 80204 161476 80256 161482
rect 80204 161418 80256 161424
rect 87196 161476 87248 161482
rect 87196 161418 87248 161424
rect 80112 161408 80164 161414
rect 80216 161385 80244 161418
rect 80112 161350 80164 161356
rect 80202 161376 80258 161385
rect 80020 161340 80072 161346
rect 80020 161282 80072 161288
rect 80124 160841 80152 161350
rect 80202 161311 80258 161320
rect 87208 161249 87236 161418
rect 87300 161346 87328 161583
rect 87380 161408 87432 161414
rect 87380 161350 87432 161356
rect 87288 161340 87340 161346
rect 87288 161282 87340 161288
rect 87194 161240 87250 161249
rect 87194 161175 87250 161184
rect 87392 160841 87420 161350
rect 80110 160832 80166 160841
rect 80110 160767 80166 160776
rect 87378 160832 87434 160841
rect 87378 160767 87434 160776
rect 76536 160518 76656 160546
rect 47082 148864 47138 148873
rect 47082 148799 47138 148808
rect 46990 144104 47046 144113
rect 46990 144039 47046 144048
rect 38252 139240 38304 139246
rect 38252 139182 38304 139188
rect 38158 124792 38214 124801
rect 38158 124727 38214 124736
rect 34664 87356 34716 87362
rect 34664 87298 34716 87304
rect 13596 17112 13648 17118
rect 13596 17054 13648 17060
rect 38172 12494 38200 124727
rect 38264 109433 38292 139182
rect 38344 130332 38396 130338
rect 38344 130274 38396 130280
rect 38356 117457 38384 130274
rect 38342 117448 38398 117457
rect 38342 117383 38398 117392
rect 47096 109530 47124 148799
rect 76628 142050 76656 160518
rect 87286 160424 87342 160433
rect 87286 160359 87342 160368
rect 80202 160288 80258 160297
rect 80202 160223 80258 160232
rect 80112 159980 80164 159986
rect 80112 159922 80164 159928
rect 80124 159617 80152 159922
rect 80216 159918 80244 160223
rect 87194 160016 87250 160025
rect 87194 159951 87196 159960
rect 87248 159951 87250 159960
rect 87196 159922 87248 159928
rect 87300 159918 87328 160359
rect 80204 159912 80256 159918
rect 80204 159854 80256 159860
rect 87288 159912 87340 159918
rect 87288 159854 87340 159860
rect 80110 159608 80166 159617
rect 80110 159543 80166 159552
rect 87194 159608 87250 159617
rect 87194 159543 87250 159552
rect 87208 159238 87236 159543
rect 80204 159232 80256 159238
rect 80204 159174 80256 159180
rect 87196 159232 87248 159238
rect 87196 159174 87248 159180
rect 87286 159200 87342 159209
rect 80216 159073 80244 159174
rect 87286 159135 87342 159144
rect 80202 159064 80258 159073
rect 80202 158999 80258 159008
rect 87300 158558 87328 159135
rect 87378 158792 87434 158801
rect 87378 158727 87434 158736
rect 80204 158552 80256 158558
rect 80202 158520 80204 158529
rect 87288 158552 87340 158558
rect 80256 158520 80258 158529
rect 87288 158494 87340 158500
rect 80202 158455 80258 158464
rect 87286 158384 87342 158393
rect 87286 158319 87342 158328
rect 87194 157976 87250 157985
rect 87194 157911 87250 157920
rect 87208 157878 87236 157911
rect 80112 157872 80164 157878
rect 79466 157840 79522 157849
rect 80112 157814 80164 157820
rect 87196 157872 87248 157878
rect 87196 157814 87248 157820
rect 79466 157775 79522 157784
rect 79480 157742 79508 157775
rect 79468 157736 79520 157742
rect 79468 157678 79520 157684
rect 80124 156761 80152 157814
rect 87300 157810 87328 158319
rect 80204 157804 80256 157810
rect 80204 157746 80256 157752
rect 87288 157804 87340 157810
rect 87288 157746 87340 157752
rect 80216 157305 80244 157746
rect 87392 157742 87420 158727
rect 87380 157736 87432 157742
rect 87380 157678 87432 157684
rect 87286 157568 87342 157577
rect 87286 157503 87342 157512
rect 80202 157296 80258 157305
rect 80202 157231 80258 157240
rect 87194 157160 87250 157169
rect 87194 157095 87250 157104
rect 80110 156752 80166 156761
rect 80110 156687 80166 156696
rect 87102 156752 87158 156761
rect 87102 156687 87158 156696
rect 80112 156444 80164 156450
rect 80112 156386 80164 156392
rect 80124 155537 80152 156386
rect 80204 156376 80256 156382
rect 80204 156318 80256 156324
rect 80216 156217 80244 156318
rect 80202 156208 80258 156217
rect 80202 156143 80258 156152
rect 87010 155664 87066 155673
rect 87010 155599 87066 155608
rect 80110 155528 80166 155537
rect 80110 155463 80166 155472
rect 86918 155256 86974 155265
rect 86918 155191 86974 155200
rect 80112 155084 80164 155090
rect 80112 155026 80164 155032
rect 80020 155016 80072 155022
rect 80020 154958 80072 154964
rect 79928 153928 79980 153934
rect 79928 153870 79980 153876
rect 79940 151298 79968 153870
rect 80032 153769 80060 154958
rect 80124 154449 80152 155026
rect 80202 154984 80258 154993
rect 80202 154919 80258 154928
rect 80216 154614 80244 154919
rect 86826 154848 86882 154857
rect 86826 154783 86882 154792
rect 80204 154608 80256 154614
rect 80204 154550 80256 154556
rect 80110 154440 80166 154449
rect 80110 154375 80166 154384
rect 80018 153760 80074 153769
rect 80018 153695 80074 153704
rect 80204 153248 80256 153254
rect 80202 153216 80204 153225
rect 80256 153216 80258 153225
rect 80202 153151 80258 153160
rect 80204 152976 80256 152982
rect 80204 152918 80256 152924
rect 80216 152681 80244 152918
rect 80202 152672 80258 152681
rect 80202 152607 80258 152616
rect 85816 152500 85868 152506
rect 85816 152442 85868 152448
rect 80112 152364 80164 152370
rect 80112 152306 80164 152312
rect 80124 151457 80152 152306
rect 80202 151720 80258 151729
rect 80202 151655 80258 151664
rect 80216 151554 80244 151655
rect 80204 151548 80256 151554
rect 80204 151490 80256 151496
rect 80110 151448 80166 151457
rect 80110 151383 80166 151392
rect 79940 151270 80152 151298
rect 79376 151140 79428 151146
rect 79376 151082 79428 151088
rect 79284 151004 79336 151010
rect 79284 150946 79336 150952
rect 79296 146833 79324 150946
rect 79388 147377 79416 151082
rect 79744 151072 79796 151078
rect 79744 151014 79796 151020
rect 79756 147921 79784 151014
rect 80124 150913 80152 151270
rect 80110 150904 80166 150913
rect 80110 150839 80166 150848
rect 80112 150392 80164 150398
rect 80112 150334 80164 150340
rect 80202 150360 80258 150369
rect 80020 149780 80072 149786
rect 80020 149722 80072 149728
rect 79928 149712 79980 149718
rect 79928 149654 79980 149660
rect 79836 149644 79888 149650
rect 79836 149586 79888 149592
rect 79742 147912 79798 147921
rect 79742 147847 79798 147856
rect 79374 147368 79430 147377
rect 79374 147303 79430 147312
rect 79282 146824 79338 146833
rect 79282 146759 79338 146768
rect 79848 145065 79876 149586
rect 79940 145609 79968 149654
rect 80032 146289 80060 149722
rect 80124 149689 80152 150334
rect 80202 150295 80258 150304
rect 80216 150194 80244 150295
rect 85828 150194 85856 152442
rect 85908 152432 85960 152438
rect 85908 152374 85960 152380
rect 85920 150398 85948 152374
rect 86840 151554 86868 154783
rect 86932 152982 86960 155191
rect 87024 153254 87052 155599
rect 87116 154614 87144 156687
rect 87208 156450 87236 157095
rect 87196 156444 87248 156450
rect 87196 156386 87248 156392
rect 87300 156382 87328 157503
rect 131540 157192 131592 157198
rect 131540 157134 131592 157140
rect 87288 156376 87340 156382
rect 87288 156318 87340 156324
rect 87378 156344 87434 156353
rect 87378 156279 87434 156288
rect 87194 156072 87250 156081
rect 87194 156007 87250 156016
rect 87208 155022 87236 156007
rect 87392 155090 87420 156279
rect 131552 155401 131580 157134
rect 131920 156518 131948 163526
rect 131908 156512 131960 156518
rect 131908 156454 131960 156460
rect 131814 156208 131870 156217
rect 131814 156143 131870 156152
rect 131538 155392 131594 155401
rect 131538 155327 131594 155336
rect 131828 155158 131856 156143
rect 131816 155152 131868 155158
rect 131816 155094 131868 155100
rect 87380 155084 87432 155090
rect 87380 155026 87432 155032
rect 131356 155084 131408 155090
rect 131356 155026 131408 155032
rect 87196 155016 87248 155022
rect 131368 154993 131396 155026
rect 131448 155016 131500 155022
rect 87196 154958 87248 154964
rect 131354 154984 131410 154993
rect 131448 154958 131500 154964
rect 131354 154919 131410 154928
rect 131356 154880 131408 154886
rect 131356 154822 131408 154828
rect 87104 154608 87156 154614
rect 87104 154550 87156 154556
rect 87102 154440 87158 154449
rect 87102 154375 87158 154384
rect 87012 153248 87064 153254
rect 87012 153190 87064 153196
rect 86920 152976 86972 152982
rect 86920 152918 86972 152924
rect 87116 152370 87144 154375
rect 87194 154032 87250 154041
rect 87194 153967 87250 153976
rect 87208 153934 87236 153967
rect 87196 153928 87248 153934
rect 131368 153905 131396 154822
rect 131460 154313 131488 154958
rect 131446 154304 131502 154313
rect 131446 154239 131502 154248
rect 87196 153870 87248 153876
rect 131354 153896 131410 153905
rect 131354 153831 131410 153840
rect 87930 153624 87986 153633
rect 87930 153559 87986 153568
rect 87562 153216 87618 153225
rect 87562 153151 87618 153160
rect 87576 152438 87604 153151
rect 87746 152808 87802 152817
rect 87746 152743 87802 152752
rect 87564 152432 87616 152438
rect 87564 152374 87616 152380
rect 87104 152364 87156 152370
rect 87104 152306 87156 152312
rect 87378 151992 87434 152001
rect 87378 151927 87434 151936
rect 87286 151584 87342 151593
rect 86828 151548 86880 151554
rect 87286 151519 87342 151528
rect 86828 151490 86880 151496
rect 87194 151176 87250 151185
rect 87300 151146 87328 151519
rect 87194 151111 87250 151120
rect 87288 151140 87340 151146
rect 87208 151010 87236 151111
rect 87288 151082 87340 151088
rect 87392 151078 87420 151927
rect 87380 151072 87432 151078
rect 87380 151014 87432 151020
rect 87196 151004 87248 151010
rect 87196 150946 87248 150952
rect 87378 150768 87434 150777
rect 87378 150703 87434 150712
rect 85908 150392 85960 150398
rect 85908 150334 85960 150340
rect 87286 150360 87342 150369
rect 87286 150295 87342 150304
rect 80204 150188 80256 150194
rect 80204 150130 80256 150136
rect 85816 150188 85868 150194
rect 85816 150130 85868 150136
rect 87194 149952 87250 149961
rect 87194 149887 87250 149896
rect 80110 149680 80166 149689
rect 87208 149650 87236 149887
rect 87300 149718 87328 150295
rect 87392 149786 87420 150703
rect 87380 149780 87432 149786
rect 87380 149722 87432 149728
rect 87288 149712 87340 149718
rect 87288 149654 87340 149660
rect 80110 149615 80166 149624
rect 87196 149644 87248 149650
rect 87196 149586 87248 149592
rect 87760 149582 87788 152743
rect 87944 152506 87972 153559
rect 87932 152500 87984 152506
rect 87932 152442 87984 152448
rect 88114 152400 88170 152409
rect 88114 152335 88170 152344
rect 131540 152364 131592 152370
rect 80204 149576 80256 149582
rect 87748 149576 87800 149582
rect 80204 149518 80256 149524
rect 87470 149544 87526 149553
rect 80112 149508 80164 149514
rect 80112 149450 80164 149456
rect 80124 148601 80152 149450
rect 80216 149145 80244 149518
rect 87748 149518 87800 149524
rect 88128 149514 88156 152335
rect 131540 152306 131592 152312
rect 131356 152296 131408 152302
rect 131354 152264 131356 152273
rect 131408 152264 131410 152273
rect 131354 152199 131410 152208
rect 131448 152228 131500 152234
rect 131448 152170 131500 152176
rect 131356 152160 131408 152166
rect 131356 152102 131408 152108
rect 131368 151865 131396 152102
rect 131354 151856 131410 151865
rect 131354 151791 131410 151800
rect 131460 151457 131488 152170
rect 131446 151448 131502 151457
rect 131446 151383 131502 151392
rect 131552 151185 131580 152306
rect 131538 151176 131594 151185
rect 131538 151111 131594 151120
rect 131356 150868 131408 150874
rect 131356 150810 131408 150816
rect 131368 150777 131396 150810
rect 131354 150768 131410 150777
rect 131354 150703 131410 150712
rect 131448 150732 131500 150738
rect 131448 150674 131500 150680
rect 131356 150528 131408 150534
rect 131356 150470 131408 150476
rect 131368 149961 131396 150470
rect 131460 150369 131488 150674
rect 131446 150360 131502 150369
rect 131446 150295 131502 150304
rect 131354 149952 131410 149961
rect 131354 149887 131410 149896
rect 131632 149576 131684 149582
rect 131446 149544 131502 149553
rect 87470 149479 87526 149488
rect 88116 149508 88168 149514
rect 80202 149136 80258 149145
rect 80202 149071 80258 149080
rect 87194 148728 87250 148737
rect 87194 148663 87250 148672
rect 80110 148592 80166 148601
rect 80110 148527 80166 148536
rect 80018 146280 80074 146289
rect 80018 146215 80074 146224
rect 79926 145600 79982 145609
rect 79926 145535 79982 145544
rect 80204 145428 80256 145434
rect 80204 145370 80256 145376
rect 79834 145056 79890 145065
rect 79834 144991 79890 145000
rect 80216 144521 80244 145370
rect 80202 144512 80258 144521
rect 80202 144447 80258 144456
rect 87208 144074 87236 148663
rect 87286 148320 87342 148329
rect 87286 148255 87342 148264
rect 80020 144068 80072 144074
rect 80020 144010 80072 144016
rect 87196 144068 87248 144074
rect 87196 144010 87248 144016
rect 80032 143297 80060 144010
rect 80204 144000 80256 144006
rect 80204 143942 80256 143948
rect 80112 143932 80164 143938
rect 80112 143874 80164 143880
rect 80018 143288 80074 143297
rect 80018 143223 80074 143232
rect 80124 142753 80152 143874
rect 80216 143841 80244 143942
rect 87300 143938 87328 148255
rect 87378 148048 87434 148057
rect 87378 147983 87434 147992
rect 87288 143932 87340 143938
rect 87288 143874 87340 143880
rect 80202 143832 80258 143841
rect 80202 143767 80258 143776
rect 80110 142744 80166 142753
rect 87392 142714 87420 147983
rect 87484 145434 87512 149479
rect 131632 149518 131684 149524
rect 131446 149479 131502 149488
rect 131540 149508 131592 149514
rect 88116 149450 88168 149456
rect 131460 149446 131488 149479
rect 131540 149450 131592 149456
rect 131448 149440 131500 149446
rect 131448 149382 131500 149388
rect 131356 149372 131408 149378
rect 131356 149314 131408 149320
rect 131368 149145 131396 149314
rect 87562 149136 87618 149145
rect 87562 149071 87618 149080
rect 131354 149136 131410 149145
rect 131354 149071 131410 149080
rect 87472 145428 87524 145434
rect 87472 145370 87524 145376
rect 87576 144006 87604 149071
rect 131552 148329 131580 149450
rect 131644 148737 131672 149518
rect 131630 148728 131686 148737
rect 131630 148663 131686 148672
rect 131538 148320 131594 148329
rect 131538 148255 131594 148264
rect 131356 148148 131408 148154
rect 131356 148090 131408 148096
rect 131368 148057 131396 148090
rect 131354 148048 131410 148057
rect 131354 147983 131410 147992
rect 109564 147870 109900 147898
rect 109564 144074 109592 147870
rect 109552 144068 109604 144074
rect 109552 144010 109604 144016
rect 87564 144000 87616 144006
rect 109564 143977 109592 144010
rect 87564 143942 87616 143948
rect 109550 143968 109606 143977
rect 109550 143903 109606 143912
rect 80110 142679 80166 142688
rect 80204 142708 80256 142714
rect 80204 142650 80256 142656
rect 87380 142708 87432 142714
rect 87380 142650 87432 142656
rect 80216 142209 80244 142650
rect 80202 142200 80258 142209
rect 80202 142135 80258 142144
rect 76458 142022 76656 142050
rect 49212 139246 49240 141900
rect 49200 139240 49252 139246
rect 49200 139182 49252 139188
rect 49856 130950 49884 141900
rect 50514 141886 51080 141914
rect 51158 141886 51264 141914
rect 51802 141886 52460 141914
rect 52538 141886 52644 141914
rect 51052 131154 51080 141886
rect 51040 131148 51092 131154
rect 51040 131090 51092 131096
rect 51236 131018 51264 141886
rect 52432 131222 52460 141886
rect 52420 131216 52472 131222
rect 52420 131158 52472 131164
rect 51224 131012 51276 131018
rect 51224 130954 51276 130960
rect 49844 130944 49896 130950
rect 49844 130886 49896 130892
rect 52616 130882 52644 141886
rect 53168 139246 53196 141900
rect 53826 141886 54024 141914
rect 53156 139240 53208 139246
rect 53156 139182 53208 139188
rect 53996 131358 54024 141886
rect 54456 139586 54484 141900
rect 54444 139580 54496 139586
rect 54444 139522 54496 139528
rect 55192 139314 55220 141900
rect 55180 139308 55232 139314
rect 55180 139250 55232 139256
rect 55836 139042 55864 141900
rect 56480 139858 56508 141900
rect 56744 139920 56796 139926
rect 56744 139862 56796 139868
rect 56468 139852 56520 139858
rect 56468 139794 56520 139800
rect 55824 139036 55876 139042
rect 55824 138978 55876 138984
rect 56756 131630 56784 139862
rect 57124 139722 57152 141900
rect 57112 139716 57164 139722
rect 57112 139658 57164 139664
rect 57572 139580 57624 139586
rect 57572 139522 57624 139528
rect 57480 139308 57532 139314
rect 57480 139250 57532 139256
rect 56192 131624 56244 131630
rect 56192 131566 56244 131572
rect 56744 131624 56796 131630
rect 56744 131566 56796 131572
rect 57388 131624 57440 131630
rect 57388 131566 57440 131572
rect 55088 131556 55140 131562
rect 55088 131498 55140 131504
rect 53984 131352 54036 131358
rect 53984 131294 54036 131300
rect 52604 130876 52656 130882
rect 52604 130818 52656 130824
rect 55100 128708 55128 131498
rect 55456 130604 55508 130610
rect 55456 130546 55508 130552
rect 55468 128708 55496 130546
rect 55824 130400 55876 130406
rect 55824 130342 55876 130348
rect 55836 128708 55864 130342
rect 56204 128708 56232 131566
rect 57020 131148 57072 131154
rect 57020 131090 57072 131096
rect 56560 130808 56612 130814
rect 56560 130750 56612 130756
rect 56572 128708 56600 130750
rect 57032 128708 57060 131090
rect 57400 128708 57428 131566
rect 57492 131426 57520 139250
rect 57584 131494 57612 139522
rect 57860 138906 57888 141900
rect 58504 139518 58532 141900
rect 58492 139512 58544 139518
rect 58492 139454 58544 139460
rect 59148 139450 59176 141900
rect 59688 139580 59740 139586
rect 59688 139522 59740 139528
rect 59136 139444 59188 139450
rect 59136 139386 59188 139392
rect 59044 139376 59096 139382
rect 59044 139318 59096 139324
rect 58860 139036 58912 139042
rect 58860 138978 58912 138984
rect 57848 138900 57900 138906
rect 57848 138842 57900 138848
rect 57572 131488 57624 131494
rect 57572 131430 57624 131436
rect 57480 131420 57532 131426
rect 57480 131362 57532 131368
rect 58766 131184 58822 131193
rect 58766 131119 58822 131128
rect 58780 131018 58808 131119
rect 58872 131018 58900 138978
rect 59056 131562 59084 139318
rect 59504 139036 59556 139042
rect 59504 138978 59556 138984
rect 59044 131556 59096 131562
rect 59044 131498 59096 131504
rect 59320 131216 59372 131222
rect 59320 131158 59372 131164
rect 58768 131012 58820 131018
rect 58768 130954 58820 130960
rect 58860 131012 58912 131018
rect 58860 130954 58912 130960
rect 58124 130740 58176 130746
rect 58124 130682 58176 130688
rect 57756 130468 57808 130474
rect 57756 130410 57808 130416
rect 57768 128708 57796 130410
rect 58136 128708 58164 130682
rect 58584 130672 58636 130678
rect 58584 130614 58636 130620
rect 58596 128708 58624 130614
rect 58952 130536 59004 130542
rect 58952 130478 59004 130484
rect 58964 128708 58992 130478
rect 59332 128708 59360 131158
rect 59516 130678 59544 138978
rect 59700 131494 59728 139522
rect 59792 139314 59820 141900
rect 60056 139920 60108 139926
rect 60056 139862 60108 139868
rect 59964 139784 60016 139790
rect 59964 139726 60016 139732
rect 59872 139648 59924 139654
rect 59872 139590 59924 139596
rect 59780 139308 59832 139314
rect 59780 139250 59832 139256
rect 59688 131488 59740 131494
rect 59688 131430 59740 131436
rect 59504 130672 59556 130678
rect 59504 130614 59556 130620
rect 59884 128722 59912 139590
rect 59714 128694 59912 128722
rect 59976 128722 60004 139726
rect 60068 131630 60096 139862
rect 60528 139586 60556 141900
rect 60976 139852 61028 139858
rect 60976 139794 61028 139800
rect 60516 139580 60568 139586
rect 60516 139522 60568 139528
rect 60608 139512 60660 139518
rect 60608 139454 60660 139460
rect 60700 139512 60752 139518
rect 60700 139454 60752 139460
rect 60424 139444 60476 139450
rect 60424 139386 60476 139392
rect 60148 139172 60200 139178
rect 60148 139114 60200 139120
rect 60056 131624 60108 131630
rect 60056 131566 60108 131572
rect 60160 130746 60188 139114
rect 60240 139104 60292 139110
rect 60240 139046 60292 139052
rect 60148 130740 60200 130746
rect 60148 130682 60200 130688
rect 60252 130474 60280 139046
rect 60332 138968 60384 138974
rect 60332 138910 60384 138916
rect 60344 131154 60372 138910
rect 60436 131630 60464 139386
rect 60424 131624 60476 131630
rect 60424 131566 60476 131572
rect 60424 131488 60476 131494
rect 60424 131430 60476 131436
rect 60514 131456 60570 131465
rect 60436 131154 60464 131430
rect 60514 131391 60516 131400
rect 60568 131391 60570 131400
rect 60516 131362 60568 131368
rect 60332 131148 60384 131154
rect 60332 131090 60384 131096
rect 60424 131148 60476 131154
rect 60424 131090 60476 131096
rect 60620 131018 60648 139454
rect 60608 131012 60660 131018
rect 60608 130954 60660 130960
rect 60240 130468 60292 130474
rect 60240 130410 60292 130416
rect 60712 128722 60740 139454
rect 60792 139376 60844 139382
rect 60792 139318 60844 139324
rect 59976 128694 60174 128722
rect 60542 128694 60740 128722
rect 60804 128722 60832 139318
rect 60884 139308 60936 139314
rect 60884 139250 60936 139256
rect 60896 131986 60924 139250
rect 60988 138634 61016 139794
rect 61172 139586 61200 141900
rect 61830 141886 62212 141914
rect 61712 139716 61764 139722
rect 61712 139658 61764 139664
rect 61160 139580 61212 139586
rect 61160 139522 61212 139528
rect 61344 139308 61396 139314
rect 61344 139250 61396 139256
rect 61252 139104 61304 139110
rect 61252 139046 61304 139052
rect 60976 138628 61028 138634
rect 60976 138570 61028 138576
rect 60896 131958 61016 131986
rect 60884 131284 60936 131290
rect 60884 131226 60936 131232
rect 60896 131193 60924 131226
rect 60882 131184 60938 131193
rect 60882 131119 60938 131128
rect 60988 130610 61016 131958
rect 61264 130814 61292 139046
rect 61252 130808 61304 130814
rect 61252 130750 61304 130756
rect 60976 130604 61028 130610
rect 60976 130546 61028 130552
rect 61356 130406 61384 139250
rect 61436 139036 61488 139042
rect 61436 138978 61488 138984
rect 61344 130400 61396 130406
rect 61344 130342 61396 130348
rect 61448 128722 61476 138978
rect 61528 138968 61580 138974
rect 61528 138910 61580 138916
rect 61540 131426 61568 138910
rect 61618 131456 61674 131465
rect 61528 131420 61580 131426
rect 61618 131391 61620 131400
rect 61528 131362 61580 131368
rect 61672 131391 61674 131400
rect 61620 131362 61672 131368
rect 61724 130746 61752 139658
rect 61988 139580 62040 139586
rect 61988 139522 62040 139528
rect 61804 139240 61856 139246
rect 61804 139182 61856 139188
rect 61712 130740 61764 130746
rect 61712 130682 61764 130688
rect 61816 130490 61844 139182
rect 61896 138900 61948 138906
rect 61896 138842 61948 138848
rect 61908 130746 61936 138842
rect 62000 130814 62028 139522
rect 61988 130808 62040 130814
rect 61988 130750 62040 130756
rect 61896 130740 61948 130746
rect 61896 130682 61948 130688
rect 62184 130678 62212 141886
rect 62460 139586 62488 141900
rect 62448 139580 62500 139586
rect 62448 139522 62500 139528
rect 63196 139450 63224 141900
rect 63840 139722 63868 141900
rect 63828 139716 63880 139722
rect 63828 139658 63880 139664
rect 63184 139444 63236 139450
rect 63184 139386 63236 139392
rect 63644 139444 63696 139450
rect 63644 139386 63696 139392
rect 63000 138628 63052 138634
rect 63000 138570 63052 138576
rect 62264 138560 62316 138566
rect 62264 138502 62316 138508
rect 62172 130672 62224 130678
rect 62172 130614 62224 130620
rect 61816 130474 61936 130490
rect 61816 130468 61948 130474
rect 61816 130462 61896 130468
rect 61896 130410 61948 130416
rect 61712 130400 61764 130406
rect 61712 130342 61764 130348
rect 60804 128694 60910 128722
rect 61278 128694 61476 128722
rect 61724 128708 61752 130342
rect 62276 128722 62304 138502
rect 62816 130944 62868 130950
rect 62816 130886 62868 130892
rect 62448 130400 62500 130406
rect 62448 130342 62500 130348
rect 62106 128694 62304 128722
rect 62460 128708 62488 130342
rect 62828 128708 62856 130886
rect 63012 130882 63040 138570
rect 63368 131284 63420 131290
rect 63368 131226 63420 131232
rect 63276 131080 63328 131086
rect 63276 131022 63328 131028
rect 63000 130876 63052 130882
rect 63000 130818 63052 130824
rect 63288 128708 63316 131022
rect 63380 128722 63408 131226
rect 63656 130406 63684 139386
rect 64484 138974 64512 141900
rect 65128 139926 65156 141900
rect 65496 141886 65786 141914
rect 65116 139920 65168 139926
rect 65116 139862 65168 139868
rect 65496 139110 65524 141886
rect 65760 139580 65812 139586
rect 65760 139522 65812 139528
rect 65484 139104 65536 139110
rect 65484 139046 65536 139052
rect 64472 138968 64524 138974
rect 64472 138910 64524 138916
rect 65576 131556 65628 131562
rect 65576 131498 65628 131504
rect 65208 131488 65260 131494
rect 65208 131430 65260 131436
rect 64380 131352 64432 131358
rect 64380 131294 64432 131300
rect 64012 130944 64064 130950
rect 64012 130886 64064 130892
rect 63644 130400 63696 130406
rect 63644 130342 63696 130348
rect 63380 128694 63670 128722
rect 64024 128708 64052 130886
rect 64392 128708 64420 131294
rect 64840 130468 64892 130474
rect 64840 130410 64892 130416
rect 64852 128708 64880 130410
rect 65220 128708 65248 131430
rect 65588 128708 65616 131498
rect 65772 130950 65800 139522
rect 66508 139246 66536 141900
rect 67152 139858 67180 141900
rect 67140 139852 67192 139858
rect 67140 139794 67192 139800
rect 67232 139580 67284 139586
rect 67232 139522 67284 139528
rect 66496 139240 66548 139246
rect 66496 139182 66548 139188
rect 67140 139240 67192 139246
rect 67140 139182 67192 139188
rect 66680 138696 66732 138702
rect 66680 138638 66732 138644
rect 66692 131034 66720 138638
rect 66692 131006 67088 131034
rect 65760 130944 65812 130950
rect 65760 130886 65812 130892
rect 66772 130876 66824 130882
rect 66772 130818 66824 130824
rect 66404 130468 66456 130474
rect 66404 130410 66456 130416
rect 65944 130400 65996 130406
rect 65944 130342 65996 130348
rect 65956 128708 65984 130342
rect 66416 128708 66444 130410
rect 66784 128708 66812 130818
rect 67060 128722 67088 131006
rect 67152 130542 67180 139182
rect 67244 131426 67272 139522
rect 67796 138838 67824 141900
rect 67784 138832 67836 138838
rect 67784 138774 67836 138780
rect 68440 138770 68468 141900
rect 69176 138906 69204 141900
rect 69820 139246 69848 141900
rect 70464 139586 70492 141900
rect 71108 139654 71136 141900
rect 71844 139790 71872 141900
rect 71832 139784 71884 139790
rect 71832 139726 71884 139732
rect 71096 139648 71148 139654
rect 71096 139590 71148 139596
rect 70452 139580 70504 139586
rect 70452 139522 70504 139528
rect 72488 139518 72516 141900
rect 72476 139512 72528 139518
rect 72476 139454 72528 139460
rect 73132 139382 73160 141900
rect 73776 139586 73804 141900
rect 73764 139580 73816 139586
rect 73764 139522 73816 139528
rect 73120 139376 73172 139382
rect 73120 139318 73172 139324
rect 74512 139314 74540 141900
rect 74500 139308 74552 139314
rect 74500 139250 74552 139256
rect 75156 139246 75184 141900
rect 75800 139450 75828 141900
rect 132012 139926 132040 163623
rect 132104 154585 132132 166178
rect 132276 163516 132328 163522
rect 132276 163458 132328 163464
rect 132288 157826 132316 163458
rect 132368 163448 132420 163454
rect 132368 163390 132420 163396
rect 132380 157946 132408 163390
rect 132458 163280 132514 163289
rect 132458 163215 132514 163224
rect 132472 162162 132500 163215
rect 132550 162872 132606 162881
rect 132550 162807 132606 162816
rect 132460 162156 132512 162162
rect 132460 162098 132512 162104
rect 132564 162094 132592 162807
rect 132642 162464 132698 162473
rect 132642 162399 132698 162408
rect 132656 162366 132684 162399
rect 132644 162360 132696 162366
rect 132644 162302 132696 162308
rect 132644 162224 132696 162230
rect 132644 162166 132696 162172
rect 132552 162088 132604 162094
rect 132656 162065 132684 162166
rect 134116 162088 134168 162094
rect 132552 162030 132604 162036
rect 132642 162056 132698 162065
rect 134116 162030 134168 162036
rect 132642 161991 132698 162000
rect 132642 161648 132698 161657
rect 132642 161583 132698 161592
rect 132550 161240 132606 161249
rect 132550 161175 132606 161184
rect 132564 160734 132592 161175
rect 132656 160938 132684 161583
rect 132644 160932 132696 160938
rect 132644 160874 132696 160880
rect 133378 160832 133434 160841
rect 133378 160767 133434 160776
rect 132552 160728 132604 160734
rect 132552 160670 132604 160676
rect 132458 160560 132514 160569
rect 132458 160495 132514 160504
rect 132472 159442 132500 160495
rect 132642 160152 132698 160161
rect 132642 160087 132698 160096
rect 132550 159744 132606 159753
rect 132550 159679 132606 159688
rect 132460 159436 132512 159442
rect 132460 159378 132512 159384
rect 132564 159374 132592 159679
rect 132656 159510 132684 160087
rect 132644 159504 132696 159510
rect 132644 159446 132696 159452
rect 132552 159368 132604 159374
rect 132552 159310 132604 159316
rect 132642 159336 132698 159345
rect 132642 159271 132644 159280
rect 132696 159271 132698 159280
rect 132644 159242 132696 159248
rect 132550 158928 132606 158937
rect 132550 158863 132606 158872
rect 132458 158520 132514 158529
rect 132458 158455 132514 158464
rect 132472 157946 132500 158455
rect 132564 158150 132592 158863
rect 132552 158144 132604 158150
rect 132552 158086 132604 158092
rect 132642 158112 132698 158121
rect 132642 158047 132644 158056
rect 132696 158047 132698 158056
rect 132644 158018 132696 158024
rect 132368 157940 132420 157946
rect 132368 157882 132420 157888
rect 132460 157940 132512 157946
rect 132460 157882 132512 157888
rect 132288 157798 132500 157826
rect 132276 157736 132328 157742
rect 132276 157678 132328 157684
rect 132288 155922 132316 157678
rect 132196 155894 132316 155922
rect 132090 154576 132146 154585
rect 132090 154511 132146 154520
rect 132196 153497 132224 155894
rect 132274 155800 132330 155809
rect 132274 155735 132330 155744
rect 132182 153488 132238 153497
rect 132182 153423 132238 153432
rect 132288 148902 132316 155735
rect 132472 152681 132500 157798
rect 132550 157704 132606 157713
rect 132550 157639 132606 157648
rect 132564 157130 132592 157639
rect 132642 157432 132698 157441
rect 132642 157367 132698 157376
rect 132552 157124 132604 157130
rect 132552 157066 132604 157072
rect 132550 157024 132606 157033
rect 132550 156959 132606 156968
rect 132564 156654 132592 156959
rect 132656 156790 132684 157367
rect 132644 156784 132696 156790
rect 132644 156726 132696 156732
rect 132552 156648 132604 156654
rect 132552 156590 132604 156596
rect 132642 156616 132698 156625
rect 132642 156551 132644 156560
rect 132696 156551 132698 156560
rect 132644 156522 132696 156528
rect 132552 156512 132604 156518
rect 132552 156454 132604 156460
rect 132564 153089 132592 156454
rect 132550 153080 132606 153089
rect 132550 153015 132606 153024
rect 132458 152672 132514 152681
rect 132458 152607 132514 152616
rect 133392 150942 133420 160767
rect 134128 155022 134156 162030
rect 134116 155016 134168 155022
rect 134116 154958 134168 154964
rect 133380 150936 133432 150942
rect 133380 150878 133432 150884
rect 132276 148896 132328 148902
rect 132276 148838 132328 148844
rect 134772 144074 134800 174406
rect 137532 172537 137560 225503
rect 137624 220817 137652 233022
rect 137704 228252 137756 228258
rect 137704 228194 137756 228200
rect 137716 227073 137744 228194
rect 137702 227064 137758 227073
rect 137702 226999 137758 227008
rect 137704 224104 137756 224110
rect 137704 224046 137756 224052
rect 137716 223945 137744 224046
rect 137702 223936 137758 223945
rect 137702 223871 137758 223880
rect 137702 221760 137758 221769
rect 137702 221695 137758 221704
rect 137610 220808 137666 220817
rect 137610 220743 137666 220752
rect 137610 218904 137666 218913
rect 137610 218839 137666 218848
rect 137518 172528 137574 172537
rect 137518 172463 137574 172472
rect 137624 172362 137652 218839
rect 137716 172673 137744 221695
rect 137808 217689 137836 233158
rect 137794 217680 137850 217689
rect 137794 217615 137850 217624
rect 137794 215912 137850 215921
rect 137794 215847 137850 215856
rect 137702 172664 137758 172673
rect 137702 172599 137758 172608
rect 137808 172498 137836 215847
rect 137900 214561 137928 233362
rect 137886 214552 137942 214561
rect 137886 214487 137942 214496
rect 137886 212376 137942 212385
rect 137886 212311 137942 212320
rect 137900 172566 137928 212311
rect 137992 211433 138020 233430
rect 138072 233284 138124 233290
rect 138072 233226 138124 233232
rect 137978 211424 138034 211433
rect 137978 211359 138034 211368
rect 137978 209384 138034 209393
rect 137978 209319 138034 209328
rect 137888 172560 137940 172566
rect 137888 172502 137940 172508
rect 137796 172492 137848 172498
rect 137796 172434 137848 172440
rect 137992 172430 138020 209319
rect 138084 208305 138112 233226
rect 138070 208296 138126 208305
rect 138070 208231 138126 208240
rect 138070 206256 138126 206265
rect 138070 206191 138126 206200
rect 138084 172702 138112 206191
rect 138176 205177 138204 233498
rect 143788 233290 143816 235862
rect 143972 235862 144308 235890
rect 144616 235862 144952 235890
rect 145168 235862 145504 235890
rect 145720 235862 146056 235890
rect 146700 235862 146760 235890
rect 143972 233494 144000 235862
rect 143960 233488 144012 233494
rect 143960 233430 144012 233436
rect 144616 233426 144644 235862
rect 144604 233420 144656 233426
rect 144604 233362 144656 233368
rect 143776 233284 143828 233290
rect 143776 233226 143828 233232
rect 145168 233222 145196 235862
rect 145156 233216 145208 233222
rect 145156 233158 145208 233164
rect 145720 233086 145748 235862
rect 145708 233080 145760 233086
rect 145708 233022 145760 233028
rect 146732 224110 146760 235862
rect 146824 235862 147252 235890
rect 147804 235862 147864 235890
rect 148448 235862 148692 235890
rect 149000 235862 149244 235890
rect 149552 235862 149888 235890
rect 150196 235862 150532 235890
rect 150748 235862 151084 235890
rect 151300 235862 151636 235890
rect 151944 235862 152004 235890
rect 152496 235862 152832 235890
rect 153048 235862 153384 235890
rect 153692 235862 154028 235890
rect 154244 235862 154580 235890
rect 154796 235862 155132 235890
rect 155440 235862 155868 235890
rect 155992 235862 156052 235890
rect 156544 235862 156880 235890
rect 157188 235862 157524 235890
rect 157740 235862 158076 235890
rect 158292 235862 158628 235890
rect 158936 235862 159088 235890
rect 146824 228258 146852 235862
rect 146812 228252 146864 228258
rect 146812 228194 146864 228200
rect 147836 224654 147864 235862
rect 148664 225130 148692 235862
rect 148652 225124 148704 225130
rect 148652 225066 148704 225072
rect 149112 224784 149164 224790
rect 149112 224726 149164 224732
rect 147824 224648 147876 224654
rect 147824 224590 147876 224596
rect 146720 224104 146772 224110
rect 146720 224046 146772 224052
rect 149124 222820 149152 224726
rect 149216 224722 149244 235862
rect 149860 232814 149888 235862
rect 150504 233086 150532 235862
rect 150492 233080 150544 233086
rect 150492 233022 150544 233028
rect 150584 232876 150636 232882
rect 150584 232818 150636 232824
rect 149848 232808 149900 232814
rect 149848 232750 149900 232756
rect 149848 225396 149900 225402
rect 149848 225338 149900 225344
rect 149480 225056 149532 225062
rect 149480 224998 149532 225004
rect 149204 224716 149256 224722
rect 149204 224658 149256 224664
rect 149492 222820 149520 224998
rect 149860 222820 149888 225338
rect 150216 225192 150268 225198
rect 150216 225134 150268 225140
rect 150228 222820 150256 225134
rect 150596 222820 150624 232818
rect 151056 232542 151084 235862
rect 151608 233222 151636 235862
rect 151780 233760 151832 233766
rect 151780 233702 151832 233708
rect 151596 233216 151648 233222
rect 151596 233158 151648 233164
rect 151044 232536 151096 232542
rect 151044 232478 151096 232484
rect 151412 225464 151464 225470
rect 151412 225406 151464 225412
rect 151044 224920 151096 224926
rect 151044 224862 151096 224868
rect 151056 222820 151084 224862
rect 151424 222820 151452 225406
rect 151792 222820 151820 233702
rect 151976 232814 152004 235862
rect 152804 232950 152832 235862
rect 153160 233556 153212 233562
rect 153160 233498 153212 233504
rect 152792 232944 152844 232950
rect 152792 232886 152844 232892
rect 151872 232808 151924 232814
rect 151872 232750 151924 232756
rect 151964 232808 152016 232814
rect 151964 232750 152016 232756
rect 151884 224518 151912 232750
rect 153172 231017 153200 233498
rect 153252 233420 153304 233426
rect 153252 233362 153304 233368
rect 152974 231008 153030 231017
rect 152974 230943 153030 230952
rect 153158 231008 153214 231017
rect 153158 230943 153214 230952
rect 152608 224852 152660 224858
rect 152608 224794 152660 224800
rect 151872 224512 151924 224518
rect 151872 224454 151924 224460
rect 152148 224308 152200 224314
rect 152148 224250 152200 224256
rect 152160 222820 152188 224250
rect 152620 222820 152648 224794
rect 152988 222820 153016 230943
rect 153264 228682 153292 233362
rect 153356 232746 153384 235862
rect 153712 233284 153764 233290
rect 153712 233226 153764 233232
rect 153344 232740 153396 232746
rect 153344 232682 153396 232688
rect 153436 232536 153488 232542
rect 153436 232478 153488 232484
rect 153264 228654 153384 228682
rect 153356 222820 153384 228654
rect 153448 224382 153476 232478
rect 153436 224376 153488 224382
rect 153436 224318 153488 224324
rect 153724 222820 153752 233226
rect 154000 232678 154028 235862
rect 154552 233358 154580 235862
rect 154908 233692 154960 233698
rect 154908 233634 154960 233640
rect 154632 233624 154684 233630
rect 154632 233566 154684 233572
rect 154540 233352 154592 233358
rect 154540 233294 154592 233300
rect 153988 232672 154040 232678
rect 153988 232614 154040 232620
rect 154644 222970 154672 233566
rect 154816 233080 154868 233086
rect 154816 233022 154868 233028
rect 154724 233012 154776 233018
rect 154724 232954 154776 232960
rect 154460 222942 154672 222970
rect 154460 222698 154488 222942
rect 154736 222698 154764 232954
rect 154828 225266 154856 233022
rect 154816 225260 154868 225266
rect 154816 225202 154868 225208
rect 154920 222820 154948 233634
rect 155104 232678 155132 235862
rect 155276 233148 155328 233154
rect 155276 233090 155328 233096
rect 155184 232944 155236 232950
rect 155184 232886 155236 232892
rect 155000 232672 155052 232678
rect 155000 232614 155052 232620
rect 155092 232672 155144 232678
rect 155092 232614 155144 232620
rect 155012 224246 155040 232614
rect 155196 224450 155224 232886
rect 155184 224444 155236 224450
rect 155184 224386 155236 224392
rect 155000 224240 155052 224246
rect 155000 224182 155052 224188
rect 155288 222820 155316 233090
rect 155736 231516 155788 231522
rect 155736 231458 155788 231464
rect 155748 222820 155776 231458
rect 155840 224178 155868 235862
rect 156024 233170 156052 235862
rect 156104 233352 156156 233358
rect 156104 233294 156156 233300
rect 155932 233142 156052 233170
rect 155828 224172 155880 224178
rect 155828 224114 155880 224120
rect 155932 224110 155960 233142
rect 156010 233048 156066 233057
rect 156010 232983 156066 232992
rect 156024 226778 156052 232983
rect 156116 226898 156144 233294
rect 156196 233216 156248 233222
rect 156196 233158 156248 233164
rect 156104 226892 156156 226898
rect 156104 226834 156156 226840
rect 156024 226750 156144 226778
rect 155920 224104 155972 224110
rect 155920 224046 155972 224052
rect 156116 222820 156144 226750
rect 156208 225334 156236 233158
rect 156852 232814 156880 235862
rect 156288 232808 156340 232814
rect 156288 232750 156340 232756
rect 156840 232808 156892 232814
rect 156840 232750 156892 232756
rect 156196 225328 156248 225334
rect 156196 225270 156248 225276
rect 156300 224994 156328 232750
rect 157496 232610 157524 235862
rect 158048 232950 158076 235862
rect 158036 232944 158088 232950
rect 158036 232886 158088 232892
rect 158600 232746 158628 235862
rect 158220 232740 158272 232746
rect 158220 232682 158272 232688
rect 158588 232740 158640 232746
rect 158588 232682 158640 232688
rect 157484 232604 157536 232610
rect 157484 232546 157536 232552
rect 156380 232536 156432 232542
rect 156380 232478 156432 232484
rect 156288 224988 156340 224994
rect 156288 224930 156340 224936
rect 156392 224790 156420 232478
rect 157300 225124 157352 225130
rect 157300 225066 157352 225072
rect 157668 225124 157720 225130
rect 157668 225066 157720 225072
rect 156380 224784 156432 224790
rect 156380 224726 156432 224732
rect 156472 224784 156524 224790
rect 156472 224726 156524 224732
rect 156484 222820 156512 224726
rect 156840 224648 156892 224654
rect 156840 224590 156892 224596
rect 156852 222820 156880 224590
rect 157312 222820 157340 225066
rect 157680 222820 157708 225066
rect 158232 224654 158260 232682
rect 159060 232678 159088 235862
rect 159152 235862 159488 235890
rect 159704 235862 160040 235890
rect 160348 235862 160684 235890
rect 160900 235862 161236 235890
rect 161788 235862 161848 235890
rect 158312 232672 158364 232678
rect 158312 232614 158364 232620
rect 159048 232672 159100 232678
rect 159048 232614 159100 232620
rect 158220 224648 158272 224654
rect 158220 224590 158272 224596
rect 158324 224586 158352 232614
rect 159152 232542 159180 235862
rect 159508 233556 159560 233562
rect 159508 233498 159560 233504
rect 159140 232536 159192 232542
rect 159140 232478 159192 232484
rect 158404 232468 158456 232474
rect 158404 232410 158456 232416
rect 158416 225418 158444 232410
rect 158416 225390 158628 225418
rect 158404 225260 158456 225266
rect 158404 225202 158456 225208
rect 158312 224580 158364 224586
rect 158312 224522 158364 224528
rect 158036 224512 158088 224518
rect 158036 224454 158088 224460
rect 158048 222820 158076 224454
rect 158416 222820 158444 225202
rect 158600 225062 158628 225390
rect 159232 225328 159284 225334
rect 159232 225270 159284 225276
rect 158588 225056 158640 225062
rect 158588 224998 158640 225004
rect 158864 224376 158916 224382
rect 158864 224318 158916 224324
rect 158876 222820 158904 224318
rect 159244 222820 159272 225270
rect 159520 224926 159548 233498
rect 159704 232474 159732 235862
rect 159784 232876 159836 232882
rect 159784 232818 159836 232824
rect 159692 232468 159744 232474
rect 159692 232410 159744 232416
rect 159796 230586 159824 232818
rect 160060 232808 160112 232814
rect 160060 232750 160112 232756
rect 159876 232604 159928 232610
rect 159876 232546 159928 232552
rect 159704 230558 159824 230586
rect 159600 229680 159652 229686
rect 159600 229622 159652 229628
rect 159612 225130 159640 229622
rect 159704 225470 159732 230558
rect 159888 230450 159916 232546
rect 159796 230422 159916 230450
rect 159692 225464 159744 225470
rect 159692 225406 159744 225412
rect 159796 225334 159824 230422
rect 160072 230314 160100 232750
rect 159888 230286 160100 230314
rect 159784 225328 159836 225334
rect 159784 225270 159836 225276
rect 159600 225124 159652 225130
rect 159600 225066 159652 225072
rect 159888 224994 159916 230286
rect 160348 225402 160376 235862
rect 160900 232082 160928 235862
rect 161820 233086 161848 235862
rect 162096 235862 162432 235890
rect 162648 235862 162984 235890
rect 163200 235862 163536 235890
rect 163844 235862 164180 235890
rect 164580 235862 164732 235890
rect 164948 235862 165284 235890
rect 165928 235862 165988 235890
rect 162096 233562 162124 235862
rect 162084 233556 162136 233562
rect 162084 233498 162136 233504
rect 161808 233080 161860 233086
rect 161808 233022 161860 233028
rect 161164 232944 161216 232950
rect 161164 232886 161216 232892
rect 160980 232740 161032 232746
rect 160980 232682 161032 232688
rect 160440 232054 160928 232082
rect 160336 225396 160388 225402
rect 160336 225338 160388 225344
rect 160440 225198 160468 232054
rect 160992 225402 161020 232682
rect 161072 232672 161124 232678
rect 161072 232614 161124 232620
rect 160980 225396 161032 225402
rect 160980 225338 161032 225344
rect 160428 225192 160480 225198
rect 160428 225134 160480 225140
rect 161084 225062 161112 232614
rect 161176 225470 161204 232886
rect 162648 232882 162676 235862
rect 163200 233766 163228 235862
rect 163188 233760 163240 233766
rect 163188 233702 163240 233708
rect 162636 232876 162688 232882
rect 162636 232818 162688 232824
rect 163844 232474 163872 235862
rect 162360 232468 162412 232474
rect 162360 232410 162412 232416
rect 163832 232468 163884 232474
rect 163832 232410 163884 232416
rect 161164 225464 161216 225470
rect 161164 225406 161216 225412
rect 160888 225056 160940 225062
rect 160888 224998 160940 225004
rect 161072 225056 161124 225062
rect 161072 224998 161124 225004
rect 159600 224988 159652 224994
rect 159600 224930 159652 224936
rect 159876 224988 159928 224994
rect 159876 224930 159928 224936
rect 159508 224920 159560 224926
rect 159508 224862 159560 224868
rect 159612 222820 159640 224930
rect 160428 224648 160480 224654
rect 160428 224590 160480 224596
rect 159968 224444 160020 224450
rect 159968 224386 160020 224392
rect 159980 222820 160008 224386
rect 160440 222820 160468 224590
rect 160796 224240 160848 224246
rect 160796 224182 160848 224188
rect 160808 222820 160836 224182
rect 160900 222834 160928 224998
rect 162372 224874 162400 232410
rect 163556 225464 163608 225470
rect 163556 225406 163608 225412
rect 163096 225328 163148 225334
rect 163096 225270 163148 225276
rect 162728 224988 162780 224994
rect 162728 224930 162780 224936
rect 162280 224846 162400 224874
rect 161532 224580 161584 224586
rect 161532 224522 161584 224528
rect 160900 222806 161190 222834
rect 161544 222820 161572 224522
rect 162280 224314 162308 224846
rect 162268 224308 162320 224314
rect 162268 224250 162320 224256
rect 161992 224172 162044 224178
rect 161992 224114 162044 224120
rect 162004 222820 162032 224114
rect 162360 224104 162412 224110
rect 162360 224046 162412 224052
rect 162372 222820 162400 224046
rect 162740 222820 162768 224930
rect 163108 222820 163136 225270
rect 163568 222820 163596 225406
rect 163924 225396 163976 225402
rect 163924 225338 163976 225344
rect 163936 222820 163964 225338
rect 164292 225056 164344 225062
rect 164292 224998 164344 225004
rect 164304 222820 164332 224998
rect 164580 224858 164608 235862
rect 164948 233426 164976 235862
rect 164936 233420 164988 233426
rect 164936 233362 164988 233368
rect 165960 233290 165988 235862
rect 166144 235862 166480 235890
rect 166696 235862 167032 235890
rect 167340 235862 167676 235890
rect 167892 235862 168228 235890
rect 168628 235862 168780 235890
rect 169088 235862 169424 235890
rect 169976 235862 170036 235890
rect 166144 233358 166172 235862
rect 166696 233494 166724 235862
rect 166684 233488 166736 233494
rect 166684 233430 166736 233436
rect 166132 233352 166184 233358
rect 166132 233294 166184 233300
rect 165948 233284 166000 233290
rect 165948 233226 166000 233232
rect 167340 233154 167368 235862
rect 167892 233698 167920 235862
rect 167880 233692 167932 233698
rect 167880 233634 167932 233640
rect 168628 233222 168656 235862
rect 168616 233216 168668 233222
rect 168616 233158 168668 233164
rect 167328 233148 167380 233154
rect 167328 233090 167380 233096
rect 169088 232746 169116 235862
rect 170008 233057 170036 235862
rect 170192 235862 170528 235890
rect 169994 233048 170050 233057
rect 169994 232983 170050 232992
rect 169076 232740 169128 232746
rect 169076 232682 169128 232688
rect 164660 225124 164712 225130
rect 164660 225066 164712 225072
rect 164568 224852 164620 224858
rect 164568 224794 164620 224800
rect 164672 222820 164700 225066
rect 170192 224790 170220 235862
rect 175344 225334 175372 243358
rect 180864 243218 180892 245903
rect 180956 245734 180984 247535
rect 181048 247502 181076 248351
rect 181140 247570 181168 248759
rect 226298 248416 226354 248425
rect 226298 248351 226354 248360
rect 226312 248318 226340 248351
rect 226300 248312 226352 248318
rect 226300 248254 226352 248260
rect 226404 248250 226432 248759
rect 233474 248416 233530 248425
rect 233474 248351 233530 248360
rect 233488 248250 233516 248351
rect 233568 248312 233620 248318
rect 233566 248280 233568 248289
rect 233620 248280 233622 248289
rect 226392 248244 226444 248250
rect 226392 248186 226444 248192
rect 233476 248244 233528 248250
rect 233566 248215 233622 248224
rect 233476 248186 233528 248192
rect 226390 248008 226446 248017
rect 226390 247943 226446 247952
rect 226298 247736 226354 247745
rect 226298 247671 226300 247680
rect 226352 247671 226354 247680
rect 226300 247642 226352 247648
rect 226404 247638 226432 247943
rect 234396 247700 234448 247706
rect 234396 247642 234448 247648
rect 226392 247632 226444 247638
rect 226392 247574 226444 247580
rect 181128 247564 181180 247570
rect 181128 247506 181180 247512
rect 181036 247496 181088 247502
rect 181036 247438 181088 247444
rect 225654 247328 225710 247337
rect 225654 247263 225710 247272
rect 182324 246408 182376 246414
rect 182322 246376 182324 246385
rect 182376 246376 182378 246385
rect 182322 246311 182378 246320
rect 225668 246278 225696 247263
rect 234408 246929 234436 247642
rect 234488 247632 234540 247638
rect 234488 247574 234540 247580
rect 234500 247337 234528 247574
rect 234486 247328 234542 247337
rect 234486 247263 234542 247272
rect 226390 246920 226446 246929
rect 226390 246855 226446 246864
rect 234394 246920 234450 246929
rect 234394 246855 234450 246864
rect 226298 246512 226354 246521
rect 226298 246447 226354 246456
rect 226312 246414 226340 246447
rect 226300 246408 226352 246414
rect 226300 246350 226352 246356
rect 226404 246346 226432 246855
rect 233660 246408 233712 246414
rect 233660 246350 233712 246356
rect 226392 246340 226444 246346
rect 226392 246282 226444 246288
rect 233568 246340 233620 246346
rect 233568 246282 233620 246288
rect 225656 246272 225708 246278
rect 225656 246214 225708 246220
rect 233476 246272 233528 246278
rect 233476 246214 233528 246220
rect 226298 246104 226354 246113
rect 226298 246039 226354 246048
rect 226206 245832 226262 245841
rect 226206 245767 226262 245776
rect 180944 245728 180996 245734
rect 180944 245670 180996 245676
rect 180942 245560 180998 245569
rect 180942 245495 180998 245504
rect 180852 243212 180904 243218
rect 180852 243154 180904 243160
rect 180956 242810 180984 245495
rect 225562 245424 225618 245433
rect 225562 245359 225618 245368
rect 225576 245258 225604 245359
rect 225564 245252 225616 245258
rect 225564 245194 225616 245200
rect 182230 245152 182286 245161
rect 182230 245087 182286 245096
rect 182046 244744 182102 244753
rect 182046 244679 182102 244688
rect 181218 243928 181274 243937
rect 181218 243863 181274 243872
rect 181232 243558 181260 243863
rect 181220 243552 181272 243558
rect 181220 243494 181272 243500
rect 180944 242804 180996 242810
rect 180944 242746 180996 242752
rect 180390 242704 180446 242713
rect 180390 242639 180446 242648
rect 180298 242296 180354 242305
rect 180298 242231 180354 242240
rect 178920 240764 178972 240770
rect 178920 240706 178972 240712
rect 178932 236554 178960 240706
rect 180312 236962 180340 242231
rect 180404 237438 180432 242639
rect 181586 242024 181642 242033
rect 182060 241994 182088 244679
rect 182138 243520 182194 243529
rect 182138 243455 182194 243464
rect 181586 241959 181642 241968
rect 182048 241988 182100 241994
rect 181600 240770 181628 241959
rect 182048 241930 182100 241936
rect 181588 240764 181640 240770
rect 181588 240706 181640 240712
rect 182152 239274 182180 243455
rect 182244 242062 182272 245087
rect 226220 244986 226248 245767
rect 226208 244980 226260 244986
rect 226208 244922 226260 244928
rect 226312 244850 226340 246039
rect 233488 245977 233516 246214
rect 233474 245968 233530 245977
rect 233474 245903 233530 245912
rect 233580 245569 233608 246282
rect 233566 245560 233622 245569
rect 233566 245495 233622 245504
rect 227956 245252 228008 245258
rect 227956 245194 228008 245200
rect 226390 245016 226446 245025
rect 226390 244951 226446 244960
rect 226404 244918 226432 244951
rect 226392 244912 226444 244918
rect 226392 244854 226444 244860
rect 226300 244844 226352 244850
rect 226300 244786 226352 244792
rect 225746 244608 225802 244617
rect 225746 244543 225802 244552
rect 182322 244336 182378 244345
rect 182322 244271 182378 244280
rect 182336 243490 182364 244271
rect 225760 243626 225788 244543
rect 226298 244200 226354 244209
rect 226298 244135 226354 244144
rect 226206 243928 226262 243937
rect 226206 243863 226262 243872
rect 225748 243620 225800 243626
rect 225748 243562 225800 243568
rect 226220 243558 226248 243863
rect 226208 243552 226260 243558
rect 226208 243494 226260 243500
rect 226312 243490 226340 244135
rect 226482 243520 226538 243529
rect 182324 243484 182376 243490
rect 182324 243426 182376 243432
rect 226300 243484 226352 243490
rect 226538 243478 226616 243506
rect 226482 243455 226538 243464
rect 226300 243426 226352 243432
rect 182322 243112 182378 243121
rect 182322 243047 182378 243056
rect 226298 243112 226354 243121
rect 226298 243047 226354 243056
rect 182336 242266 182364 243047
rect 226022 242704 226078 242713
rect 226022 242639 226078 242648
rect 226036 242266 226064 242639
rect 182324 242260 182376 242266
rect 182324 242202 182376 242208
rect 226024 242260 226076 242266
rect 226024 242202 226076 242208
rect 226312 242198 226340 243047
rect 226390 242296 226446 242305
rect 226390 242231 226446 242240
rect 226300 242192 226352 242198
rect 226300 242134 226352 242140
rect 226404 242130 226432 242231
rect 226392 242124 226444 242130
rect 226392 242066 226444 242072
rect 182232 242056 182284 242062
rect 182232 241998 182284 242004
rect 226022 242024 226078 242033
rect 226022 241959 226078 241968
rect 203864 239818 203892 241860
rect 226036 240702 226064 241959
rect 226024 240696 226076 240702
rect 226024 240638 226076 240644
rect 203116 239812 203168 239818
rect 203116 239754 203168 239760
rect 203852 239812 203904 239818
rect 203852 239754 203904 239760
rect 182140 239268 182192 239274
rect 182140 239210 182192 239216
rect 180392 237432 180444 237438
rect 180392 237374 180444 237380
rect 180300 236956 180352 236962
rect 180300 236898 180352 236904
rect 178920 236548 178972 236554
rect 178920 236490 178972 236496
rect 203128 233737 203156 239754
rect 226588 239274 226616 243478
rect 227968 243354 227996 245194
rect 228048 244980 228100 244986
rect 228048 244922 228100 244928
rect 228060 243422 228088 244922
rect 228140 244912 228192 244918
rect 228140 244854 228192 244860
rect 228048 243416 228100 243422
rect 228048 243358 228100 243364
rect 227956 243348 228008 243354
rect 227956 243290 228008 243296
rect 228152 242062 228180 244854
rect 233476 244844 233528 244850
rect 233476 244786 233528 244792
rect 233488 244209 233516 244786
rect 233672 244753 233700 246350
rect 233658 244744 233714 244753
rect 233658 244679 233714 244688
rect 233474 244200 233530 244209
rect 233474 244135 233530 244144
rect 233660 243620 233712 243626
rect 233660 243562 233712 243568
rect 233476 243416 233528 243422
rect 233474 243384 233476 243393
rect 233528 243384 233530 243393
rect 233474 243319 233530 243328
rect 233568 243348 233620 243354
rect 233568 243290 233620 243296
rect 233580 242849 233608 243290
rect 233566 242840 233622 242849
rect 233566 242775 233622 242784
rect 228692 242260 228744 242266
rect 228692 242202 228744 242208
rect 228600 242124 228652 242130
rect 228600 242066 228652 242072
rect 228140 242056 228192 242062
rect 228140 241998 228192 242004
rect 226576 239268 226628 239274
rect 226576 239210 226628 239216
rect 228612 237846 228640 242066
rect 228704 237914 228732 242202
rect 233568 242124 233620 242130
rect 233568 242066 233620 242072
rect 233476 242056 233528 242062
rect 233474 242024 233476 242033
rect 233528 242024 233530 242033
rect 233474 241959 233530 241968
rect 233476 239268 233528 239274
rect 233476 239210 233528 239216
rect 233488 239177 233516 239210
rect 233474 239168 233530 239177
rect 233474 239103 233530 239112
rect 233580 238769 233608 242066
rect 233672 241489 233700 243562
rect 233844 243552 233896 243558
rect 233844 243494 233896 243500
rect 233752 243484 233804 243490
rect 233752 243426 233804 243432
rect 233658 241480 233714 241489
rect 233658 241415 233714 241424
rect 233764 240673 233792 243426
rect 233750 240664 233806 240673
rect 233750 240599 233806 240608
rect 233856 240129 233884 243494
rect 264662 242296 264718 242305
rect 264662 242231 264718 242240
rect 234120 240696 234172 240702
rect 234120 240638 234172 240644
rect 233842 240120 233898 240129
rect 233842 240055 233898 240064
rect 233566 238760 233622 238769
rect 233566 238695 233622 238704
rect 228692 237908 228744 237914
rect 228692 237850 228744 237856
rect 233476 237908 233528 237914
rect 233476 237850 233528 237856
rect 228600 237840 228652 237846
rect 233488 237817 233516 237850
rect 233568 237840 233620 237846
rect 228600 237782 228652 237788
rect 233474 237808 233530 237817
rect 233568 237782 233620 237788
rect 233474 237743 233530 237752
rect 233580 237409 233608 237782
rect 233566 237400 233622 237409
rect 233566 237335 233622 237344
rect 234132 236457 234160 240638
rect 234118 236448 234174 236457
rect 234118 236383 234174 236392
rect 236892 235862 237228 235890
rect 237628 235862 237780 235890
rect 237996 235862 238332 235890
rect 238548 235862 238884 235890
rect 239192 235862 239436 235890
rect 239652 235862 239988 235890
rect 240388 235862 240540 235890
rect 240756 235862 241092 235890
rect 241584 235862 241644 235890
rect 242196 235862 242532 235890
rect 242748 235862 243084 235890
rect 243300 235862 243636 235890
rect 243852 235862 244188 235890
rect 203114 233728 203170 233737
rect 203114 233663 203170 233672
rect 231820 233216 231872 233222
rect 231820 233158 231872 233164
rect 231728 233080 231780 233086
rect 231728 233022 231780 233028
rect 231636 232672 231688 232678
rect 231636 232614 231688 232620
rect 231544 232604 231596 232610
rect 231544 232546 231596 232552
rect 231452 232536 231504 232542
rect 231452 232478 231504 232484
rect 231360 232468 231412 232474
rect 231360 232410 231412 232416
rect 220504 229680 220556 229686
rect 220504 229622 220556 229628
rect 220516 227716 220544 229622
rect 175332 225328 175384 225334
rect 175332 225270 175384 225276
rect 170180 224784 170232 224790
rect 170180 224726 170232 224732
rect 154198 222670 154488 222698
rect 154566 222670 154764 222698
rect 231082 221896 231138 221905
rect 231082 221831 231138 221840
rect 148742 221624 148798 221633
rect 148742 221559 148798 221568
rect 148756 221390 148784 221559
rect 231096 221390 231124 221831
rect 148744 221384 148796 221390
rect 148744 221326 148796 221332
rect 165120 221384 165172 221390
rect 165120 221326 165172 221332
rect 231084 221384 231136 221390
rect 231084 221326 231136 221332
rect 145614 219312 145670 219321
rect 145614 219247 145670 219256
rect 145628 218670 145656 219247
rect 145616 218664 145668 218670
rect 145616 218606 145668 218612
rect 145614 217000 145670 217009
rect 145614 216935 145670 216944
rect 145628 215882 145656 216935
rect 145616 215876 145668 215882
rect 145616 215818 145668 215824
rect 165132 215814 165160 221326
rect 230990 219040 231046 219049
rect 230990 218975 231046 218984
rect 231004 218874 231032 218975
rect 230992 218868 231044 218874
rect 230992 218810 231044 218816
rect 165120 215808 165172 215814
rect 175516 215808 175568 215814
rect 165120 215750 165172 215756
rect 175514 215776 175516 215785
rect 175568 215776 175570 215785
rect 175514 215711 175570 215720
rect 145614 214416 145670 214425
rect 145614 214351 145670 214360
rect 145628 213162 145656 214351
rect 145616 213156 145668 213162
rect 145616 213098 145668 213104
rect 145614 212240 145670 212249
rect 145614 212175 145670 212184
rect 145628 211734 145656 212175
rect 145616 211728 145668 211734
rect 145616 211670 145668 211676
rect 145614 209928 145670 209937
rect 145614 209863 145670 209872
rect 145628 209014 145656 209863
rect 145616 209008 145668 209014
rect 145616 208950 145668 208956
rect 145798 207480 145854 207489
rect 145798 207415 145854 207424
rect 138162 205168 138218 205177
rect 138162 205103 138218 205112
rect 145614 205168 145670 205177
rect 145614 205103 145670 205112
rect 145628 204866 145656 205103
rect 145616 204860 145668 204866
rect 145616 204802 145668 204808
rect 138162 203536 138218 203545
rect 138162 203471 138218 203480
rect 138072 172696 138124 172702
rect 138072 172638 138124 172644
rect 138176 172634 138204 203471
rect 145522 202856 145578 202865
rect 145522 202791 145578 202800
rect 145536 202078 145564 202791
rect 143040 202072 143092 202078
rect 143040 202014 143092 202020
rect 145524 202072 145576 202078
rect 145524 202014 145576 202020
rect 140280 197924 140332 197930
rect 140280 197866 140332 197872
rect 140292 188206 140320 197866
rect 140372 195204 140424 195210
rect 140372 195146 140424 195152
rect 140280 188200 140332 188206
rect 140280 188142 140332 188148
rect 140384 186846 140412 195146
rect 143052 191130 143080 202014
rect 144418 200544 144474 200553
rect 144418 200479 144474 200488
rect 143132 192416 143184 192422
rect 143132 192358 143184 192364
rect 143040 191124 143092 191130
rect 143040 191066 143092 191072
rect 140372 186840 140424 186846
rect 140372 186782 140424 186788
rect 143144 184262 143172 192358
rect 144432 189430 144460 200479
rect 145614 198096 145670 198105
rect 145614 198031 145670 198040
rect 145628 197930 145656 198031
rect 145616 197924 145668 197930
rect 145616 197866 145668 197872
rect 145614 195784 145670 195793
rect 145614 195719 145670 195728
rect 145628 195210 145656 195719
rect 145616 195204 145668 195210
rect 145616 195146 145668 195152
rect 145812 195142 145840 207415
rect 231372 205177 231400 232410
rect 231464 208305 231492 232478
rect 231556 211433 231584 232546
rect 231648 214561 231676 232614
rect 231740 220817 231768 233022
rect 231726 220808 231782 220817
rect 231726 220743 231782 220752
rect 231728 218732 231780 218738
rect 231728 218674 231780 218680
rect 231634 214552 231690 214561
rect 231634 214487 231690 214496
rect 231636 211728 231688 211734
rect 231636 211670 231688 211676
rect 231542 211424 231598 211433
rect 231542 211359 231598 211368
rect 231544 209008 231596 209014
rect 231544 208950 231596 208956
rect 231450 208296 231506 208305
rect 231450 208231 231506 208240
rect 231358 205168 231414 205177
rect 231358 205103 231414 205112
rect 231452 204860 231504 204866
rect 231452 204802 231504 204808
rect 231358 203536 231414 203545
rect 231358 203471 231414 203480
rect 231268 202072 231320 202078
rect 231268 202014 231320 202020
rect 145800 195136 145852 195142
rect 145800 195078 145852 195084
rect 145798 193472 145854 193481
rect 145798 193407 145854 193416
rect 145812 192422 145840 193407
rect 167878 192792 167934 192801
rect 167878 192727 167934 192736
rect 167892 192422 167920 192727
rect 145800 192416 145852 192422
rect 145800 192358 145852 192364
rect 167880 192416 167932 192422
rect 167880 192358 167932 192364
rect 175516 192416 175568 192422
rect 175516 192358 175568 192364
rect 175528 190897 175556 192358
rect 231280 191169 231308 202014
rect 231266 191160 231322 191169
rect 231266 191095 231322 191104
rect 145154 190888 145210 190897
rect 145154 190823 145210 190832
rect 175514 190888 175570 190897
rect 175514 190823 175570 190832
rect 145168 189702 145196 190823
rect 145156 189696 145208 189702
rect 145156 189638 145208 189644
rect 230808 189696 230860 189702
rect 230808 189638 230860 189644
rect 144420 189424 144472 189430
rect 144420 189366 144472 189372
rect 145614 188712 145670 188721
rect 145614 188647 145670 188656
rect 145628 188274 145656 188647
rect 145616 188268 145668 188274
rect 145616 188210 145668 188216
rect 144786 186400 144842 186409
rect 144786 186335 144842 186344
rect 143132 184256 143184 184262
rect 143132 184198 143184 184204
rect 144800 180046 144828 186335
rect 145798 183408 145854 183417
rect 145798 183343 145854 183352
rect 145156 181196 145208 181202
rect 145156 181138 145208 181144
rect 144880 180720 144932 180726
rect 144880 180662 144932 180668
rect 144788 180040 144840 180046
rect 144788 179982 144840 179988
rect 143684 179972 143736 179978
rect 143684 179914 143736 179920
rect 140280 175620 140332 175626
rect 140280 175562 140332 175568
rect 138164 172628 138216 172634
rect 138164 172570 138216 172576
rect 137980 172424 138032 172430
rect 137980 172366 138032 172372
rect 137612 172356 137664 172362
rect 137612 172298 137664 172304
rect 139636 170180 139688 170186
rect 139636 170122 139688 170128
rect 139648 169545 139676 170122
rect 139634 169536 139690 169545
rect 139634 169471 139690 169480
rect 139636 168888 139688 168894
rect 139634 168856 139636 168865
rect 139688 168856 139690 168865
rect 139634 168791 139690 168800
rect 139726 167088 139782 167097
rect 139726 167023 139782 167032
rect 139634 166544 139690 166553
rect 139634 166479 139690 166488
rect 135036 166304 135088 166310
rect 135036 166246 135088 166252
rect 134944 159300 134996 159306
rect 134944 159242 134996 159248
rect 134852 155152 134904 155158
rect 134852 155094 134904 155100
rect 134864 144074 134892 155094
rect 134956 148222 134984 159242
rect 135048 155090 135076 166246
rect 139648 166242 139676 166479
rect 139740 166310 139768 167023
rect 139728 166304 139780 166310
rect 139728 166246 139780 166252
rect 139636 166236 139688 166242
rect 139636 166178 139688 166184
rect 139082 165728 139138 165737
rect 139082 165663 139138 165672
rect 138990 165048 139046 165057
rect 138990 164983 139046 164992
rect 135312 162156 135364 162162
rect 135312 162098 135364 162104
rect 136232 162156 136284 162162
rect 136232 162098 136284 162104
rect 135220 158008 135272 158014
rect 135220 157950 135272 157956
rect 135128 155152 135180 155158
rect 135128 155094 135180 155100
rect 135036 155084 135088 155090
rect 135036 155026 135088 155032
rect 134944 148216 134996 148222
rect 134944 148158 134996 148164
rect 135140 148154 135168 155094
rect 135232 150534 135260 157950
rect 135324 155090 135352 162098
rect 136140 157940 136192 157946
rect 136140 157882 136192 157888
rect 135312 155084 135364 155090
rect 135312 155026 135364 155032
rect 135220 150528 135272 150534
rect 135220 150470 135272 150476
rect 135128 148148 135180 148154
rect 135128 148090 135180 148096
rect 136152 146794 136180 157882
rect 136244 152302 136272 162098
rect 136324 162088 136376 162094
rect 136324 162030 136376 162036
rect 136232 152296 136284 152302
rect 136232 152238 136284 152244
rect 136336 152166 136364 162030
rect 136416 160864 136468 160870
rect 136416 160806 136468 160812
rect 136428 152234 136456 160806
rect 136508 160660 136560 160666
rect 136508 160602 136560 160608
rect 136520 152370 136548 160602
rect 137520 157124 137572 157130
rect 137520 157066 137572 157072
rect 136508 152364 136560 152370
rect 136508 152306 136560 152312
rect 136416 152228 136468 152234
rect 136416 152170 136468 152176
rect 136324 152160 136376 152166
rect 136324 152102 136376 152108
rect 136140 146788 136192 146794
rect 136140 146730 136192 146736
rect 137532 145434 137560 157066
rect 138808 156988 138860 156994
rect 138808 156930 138860 156936
rect 138820 149378 138848 156930
rect 138900 156648 138952 156654
rect 138900 156590 138952 156596
rect 138808 149372 138860 149378
rect 138808 149314 138860 149320
rect 137520 145428 137572 145434
rect 137520 145370 137572 145376
rect 138912 144113 138940 156590
rect 139004 154886 139032 164983
rect 138992 154880 139044 154886
rect 138992 154822 139044 154828
rect 139096 154818 139124 165663
rect 139728 162360 139780 162366
rect 139728 162302 139780 162308
rect 139358 159744 139414 159753
rect 139358 159679 139414 159688
rect 139268 159436 139320 159442
rect 139268 159378 139320 159384
rect 139174 158112 139230 158121
rect 139174 158047 139230 158056
rect 139084 154812 139136 154818
rect 139084 154754 139136 154760
rect 139188 149446 139216 158047
rect 139280 150097 139308 159378
rect 139372 150874 139400 159679
rect 139450 159472 139506 159481
rect 139450 159407 139506 159416
rect 139360 150868 139412 150874
rect 139360 150810 139412 150816
rect 139464 150738 139492 159407
rect 139542 156752 139598 156761
rect 139740 156722 139768 162302
rect 139912 162224 139964 162230
rect 139912 162166 139964 162172
rect 139818 161104 139874 161113
rect 139818 161039 139874 161048
rect 139832 160870 139860 161039
rect 139820 160864 139872 160870
rect 139820 160806 139872 160812
rect 139542 156687 139598 156696
rect 139728 156716 139780 156722
rect 139452 150732 139504 150738
rect 139452 150674 139504 150680
rect 139266 150088 139322 150097
rect 139266 150023 139322 150032
rect 139556 149582 139584 156687
rect 139728 156658 139780 156664
rect 139818 155800 139874 155809
rect 139818 155735 139874 155744
rect 139726 155256 139782 155265
rect 139726 155191 139782 155200
rect 139740 155158 139768 155191
rect 139728 155152 139780 155158
rect 139728 155094 139780 155100
rect 139636 155084 139688 155090
rect 139636 155026 139688 155032
rect 139648 154857 139676 155026
rect 139728 155016 139780 155022
rect 139728 154958 139780 154964
rect 139634 154848 139690 154857
rect 139634 154783 139690 154792
rect 139740 154177 139768 154958
rect 139726 154168 139782 154177
rect 139726 154103 139782 154112
rect 139636 150936 139688 150942
rect 139636 150878 139688 150884
rect 139648 150777 139676 150878
rect 139634 150768 139690 150777
rect 139634 150703 139690 150712
rect 139544 149576 139596 149582
rect 139544 149518 139596 149524
rect 139832 149514 139860 155735
rect 139924 152817 139952 162166
rect 140004 160932 140056 160938
rect 140004 160874 140056 160880
rect 139910 152808 139966 152817
rect 139910 152743 139966 152752
rect 140016 152137 140044 160874
rect 140096 160728 140148 160734
rect 140096 160670 140148 160676
rect 140108 156874 140136 160670
rect 140186 157024 140242 157033
rect 140186 156959 140188 156968
rect 140240 156959 140242 156968
rect 140188 156930 140240 156936
rect 140108 156846 140228 156874
rect 140096 156716 140148 156722
rect 140096 156658 140148 156664
rect 140108 153497 140136 156658
rect 140094 153488 140150 153497
rect 140094 153423 140150 153432
rect 140002 152128 140058 152137
rect 140002 152063 140058 152072
rect 140200 151457 140228 156846
rect 140186 151448 140242 151457
rect 140186 151383 140242 151392
rect 139820 149508 139872 149514
rect 139820 149450 139872 149456
rect 139176 149440 139228 149446
rect 139176 149382 139228 149388
rect 139636 148896 139688 148902
rect 139636 148838 139688 148844
rect 138898 144104 138954 144113
rect 134760 144068 134812 144074
rect 134760 144010 134812 144016
rect 134852 144068 134904 144074
rect 138898 144039 138954 144048
rect 134852 144010 134904 144016
rect 139648 142209 139676 148838
rect 139728 148216 139780 148222
rect 139726 148184 139728 148193
rect 139780 148184 139782 148193
rect 139726 148119 139782 148128
rect 139726 146824 139782 146833
rect 139726 146759 139728 146768
rect 139780 146759 139782 146768
rect 139728 146730 139780 146736
rect 139910 145464 139966 145473
rect 139910 145399 139912 145408
rect 139964 145399 139966 145408
rect 139912 145370 139964 145376
rect 139728 144068 139780 144074
rect 139728 144010 139780 144016
rect 139740 142753 139768 144010
rect 139726 142744 139782 142753
rect 139726 142679 139782 142688
rect 139634 142200 139690 142209
rect 139634 142135 139690 142144
rect 132000 139920 132052 139926
rect 132000 139862 132052 139868
rect 140292 139858 140320 175562
rect 143696 169930 143724 179914
rect 144604 173036 144656 173042
rect 144604 172978 144656 172984
rect 143868 172968 143920 172974
rect 143868 172910 143920 172916
rect 143604 169902 143724 169930
rect 143604 169658 143632 169902
rect 143880 169794 143908 172910
rect 144616 169794 144644 172978
rect 144892 169794 144920 180662
rect 144972 180652 145024 180658
rect 144972 180594 145024 180600
rect 144984 173042 145012 180594
rect 145168 179994 145196 181138
rect 145076 179966 145196 179994
rect 144972 173036 145024 173042
rect 144972 172978 145024 172984
rect 145076 172974 145104 179966
rect 145812 179910 145840 183343
rect 230820 183281 230848 189638
rect 231268 188268 231320 188274
rect 231268 188210 231320 188216
rect 230806 183272 230862 183281
rect 230806 183207 230862 183216
rect 147732 181060 147784 181066
rect 147732 181002 147784 181008
rect 147640 180856 147692 180862
rect 147640 180798 147692 180804
rect 146444 180788 146496 180794
rect 146444 180730 146496 180736
rect 146352 180380 146404 180386
rect 146352 180322 146404 180328
rect 145800 179904 145852 179910
rect 145800 179846 145852 179852
rect 146364 173042 146392 180322
rect 145708 173036 145760 173042
rect 145708 172978 145760 172984
rect 146352 173036 146404 173042
rect 146352 172978 146404 172984
rect 145064 172968 145116 172974
rect 145064 172910 145116 172916
rect 145720 169794 145748 172978
rect 146456 169930 146484 180730
rect 146536 171948 146588 171954
rect 146536 171890 146588 171896
rect 143756 169766 143908 169794
rect 144308 169766 144644 169794
rect 144860 169766 144920 169794
rect 145412 169766 145748 169794
rect 146364 169902 146484 169930
rect 146364 169658 146392 169902
rect 146548 169794 146576 171890
rect 147652 169930 147680 180798
rect 147744 171954 147772 181002
rect 147824 180992 147876 180998
rect 147824 180934 147876 180940
rect 147732 171948 147784 171954
rect 147732 171890 147784 171896
rect 147376 169902 147680 169930
rect 147376 169794 147404 169902
rect 147836 169794 147864 180934
rect 149124 180182 149152 182836
rect 149204 181264 149256 181270
rect 149204 181206 149256 181212
rect 149112 180176 149164 180182
rect 149112 180118 149164 180124
rect 149216 173042 149244 181206
rect 149492 180930 149520 182836
rect 149480 180924 149532 180930
rect 149480 180866 149532 180872
rect 149860 180114 149888 182836
rect 150320 180522 150348 182836
rect 150688 181338 150716 182836
rect 150676 181332 150728 181338
rect 150676 181274 150728 181280
rect 150308 180516 150360 180522
rect 150308 180458 150360 180464
rect 149848 180108 149900 180114
rect 149848 180050 149900 180056
rect 151056 180046 151084 182836
rect 151424 182822 151530 182850
rect 151044 180040 151096 180046
rect 151044 179982 151096 179988
rect 151424 173110 151452 182822
rect 151688 181332 151740 181338
rect 151688 181274 151740 181280
rect 151412 173104 151464 173110
rect 151412 173046 151464 173052
rect 148468 173036 148520 173042
rect 148468 172978 148520 172984
rect 149204 173036 149256 173042
rect 149204 172978 149256 172984
rect 151320 173036 151372 173042
rect 151320 172978 151372 172984
rect 148480 169794 148508 172978
rect 150124 172900 150176 172906
rect 150124 172842 150176 172848
rect 149020 172220 149072 172226
rect 149020 172162 149072 172168
rect 149032 169794 149060 172162
rect 149572 171744 149624 171750
rect 149572 171686 149624 171692
rect 149584 169794 149612 171686
rect 150136 169794 150164 172842
rect 150584 172832 150636 172838
rect 150584 172774 150636 172780
rect 150596 169794 150624 172774
rect 151332 169794 151360 172978
rect 151700 172770 151728 181274
rect 151780 180448 151832 180454
rect 151780 180390 151832 180396
rect 151792 173042 151820 180390
rect 151780 173036 151832 173042
rect 151780 172978 151832 172984
rect 151688 172764 151740 172770
rect 151688 172706 151740 172712
rect 151884 172294 151912 182836
rect 152252 181134 152280 182836
rect 152726 182822 153016 182850
rect 152988 181218 153016 182822
rect 153080 181338 153108 182836
rect 153068 181332 153120 181338
rect 153068 181274 153120 181280
rect 152988 181190 153292 181218
rect 152240 181128 152292 181134
rect 152240 181070 152292 181076
rect 153264 180930 153292 181190
rect 153160 180924 153212 180930
rect 153160 180866 153212 180872
rect 153252 180924 153304 180930
rect 153252 180866 153304 180872
rect 152976 180516 153028 180522
rect 152976 180458 153028 180464
rect 152056 180312 152108 180318
rect 152056 180254 152108 180260
rect 152068 179858 152096 180254
rect 152884 180176 152936 180182
rect 152884 180118 152936 180124
rect 152792 180108 152844 180114
rect 152792 180050 152844 180056
rect 151976 179830 152096 179858
rect 151872 172288 151924 172294
rect 151872 172230 151924 172236
rect 151976 169794 152004 179830
rect 152804 175642 152832 180050
rect 152620 175614 152832 175642
rect 152424 172900 152476 172906
rect 152424 172842 152476 172848
rect 152436 169794 152464 172842
rect 152620 171818 152648 175614
rect 152896 175506 152924 180118
rect 152700 175484 152752 175490
rect 152700 175426 152752 175432
rect 152804 175478 152924 175506
rect 152988 175490 153016 180458
rect 152976 175484 153028 175490
rect 152712 171886 152740 175426
rect 152804 171954 152832 175478
rect 152976 175426 153028 175432
rect 153172 175370 153200 180866
rect 153448 180590 153476 182836
rect 153436 180584 153488 180590
rect 153436 180526 153488 180532
rect 153908 180386 153936 182836
rect 153896 180380 153948 180386
rect 153896 180322 153948 180328
rect 153252 180040 153304 180046
rect 153252 179982 153304 179988
rect 152896 175342 153200 175370
rect 152896 172090 152924 175342
rect 153264 175234 153292 179982
rect 153344 179972 153396 179978
rect 153344 179914 153396 179920
rect 152988 175206 153292 175234
rect 152988 172906 153016 175206
rect 153356 175098 153384 179914
rect 153080 175070 153384 175098
rect 152976 172900 153028 172906
rect 152976 172842 153028 172848
rect 152884 172084 152936 172090
rect 152884 172026 152936 172032
rect 152792 171948 152844 171954
rect 152792 171890 152844 171896
rect 152700 171880 152752 171886
rect 152700 171822 152752 171828
rect 152608 171812 152660 171818
rect 152608 171754 152660 171760
rect 153080 169794 153108 175070
rect 154276 172809 154304 182836
rect 154644 172945 154672 182836
rect 155118 182822 155408 182850
rect 155380 180402 155408 182822
rect 155472 180522 155500 182836
rect 155460 180516 155512 180522
rect 155460 180458 155512 180464
rect 155380 180374 155776 180402
rect 154630 172936 154686 172945
rect 154630 172871 154686 172880
rect 154262 172800 154318 172809
rect 153344 172764 153396 172770
rect 154262 172735 154318 172744
rect 153344 172706 153396 172712
rect 153356 169794 153384 172706
rect 154816 172696 154868 172702
rect 154816 172638 154868 172644
rect 154172 172628 154224 172634
rect 154172 172570 154224 172576
rect 154080 172220 154132 172226
rect 154080 172162 154132 172168
rect 154092 169794 154120 172162
rect 146516 169766 146576 169794
rect 147068 169766 147404 169794
rect 147620 169766 147864 169794
rect 148172 169766 148508 169794
rect 148724 169766 149060 169794
rect 149276 169766 149612 169794
rect 149828 169766 150164 169794
rect 150472 169766 150624 169794
rect 151024 169766 151360 169794
rect 151576 169766 152004 169794
rect 152128 169766 152464 169794
rect 152680 169766 153108 169794
rect 153232 169766 153384 169794
rect 153784 169766 154120 169794
rect 154184 169794 154212 172570
rect 154828 169930 154856 172638
rect 155644 172560 155696 172566
rect 155644 172502 155696 172508
rect 155092 172424 155144 172430
rect 155092 172366 155144 172372
rect 154828 169902 154902 169930
rect 154184 169766 154336 169794
rect 154874 169780 154902 169902
rect 155104 169794 155132 172366
rect 155656 169794 155684 172502
rect 155748 172430 155776 180374
rect 155840 172566 155868 182836
rect 156300 181338 156328 182836
rect 156682 182822 157064 182850
rect 156288 181332 156340 181338
rect 156288 181274 156340 181280
rect 156104 180516 156156 180522
rect 156104 180458 156156 180464
rect 156116 172634 156144 180458
rect 156840 180176 156892 180182
rect 156840 180118 156892 180124
rect 157036 180130 157064 182822
rect 157128 180250 157156 182836
rect 157220 182822 157510 182850
rect 157220 181202 157248 182822
rect 157484 181332 157536 181338
rect 157484 181274 157536 181280
rect 157208 181196 157260 181202
rect 157208 181138 157260 181144
rect 157116 180244 157168 180250
rect 157116 180186 157168 180192
rect 156852 172906 156880 180118
rect 157036 180102 157432 180130
rect 157024 180040 157076 180046
rect 157024 179982 157076 179988
rect 156840 172900 156892 172906
rect 156840 172842 156892 172848
rect 157036 172770 157064 179982
rect 157024 172764 157076 172770
rect 157024 172706 157076 172712
rect 156104 172628 156156 172634
rect 156104 172570 156156 172576
rect 155828 172560 155880 172566
rect 155828 172502 155880 172508
rect 156196 172492 156248 172498
rect 156196 172434 156248 172440
rect 155736 172424 155788 172430
rect 155736 172366 155788 172372
rect 156208 169794 156236 172434
rect 157404 172362 157432 180102
rect 157496 172498 157524 181274
rect 157864 180658 157892 182836
rect 158324 180726 158352 182836
rect 158404 181332 158456 181338
rect 158404 181274 158456 181280
rect 158312 180720 158364 180726
rect 158312 180662 158364 180668
rect 157852 180652 157904 180658
rect 157852 180594 157904 180600
rect 158220 180652 158272 180658
rect 158220 180594 158272 180600
rect 157574 172664 157630 172673
rect 157574 172599 157630 172608
rect 157484 172492 157536 172498
rect 157484 172434 157536 172440
rect 156840 172356 156892 172362
rect 156840 172298 156892 172304
rect 157392 172356 157444 172362
rect 157392 172298 157444 172304
rect 156852 169794 156880 172298
rect 157588 169794 157616 172599
rect 157942 172528 157998 172537
rect 157942 172463 157998 172472
rect 157956 169794 157984 172463
rect 158232 172226 158260 180594
rect 158416 180538 158444 181274
rect 158324 180510 158444 180538
rect 158324 172537 158352 180510
rect 158692 180318 158720 182836
rect 159060 180794 159088 182836
rect 159520 181066 159548 182836
rect 159508 181060 159560 181066
rect 159508 181002 159560 181008
rect 159888 180862 159916 182836
rect 160256 180998 160284 182836
rect 160716 181270 160744 182836
rect 160704 181264 160756 181270
rect 160704 181206 160756 181212
rect 160244 180992 160296 180998
rect 160244 180934 160296 180940
rect 159876 180856 159928 180862
rect 159876 180798 159928 180804
rect 159048 180788 159100 180794
rect 159048 180730 159100 180736
rect 158680 180312 158732 180318
rect 158680 180254 158732 180260
rect 158310 172528 158366 172537
rect 158310 172463 158366 172472
rect 158220 172220 158272 172226
rect 158220 172162 158272 172168
rect 160704 172152 160756 172158
rect 160704 172094 160756 172100
rect 159048 172084 159100 172090
rect 159048 172026 159100 172032
rect 158496 171948 158548 171954
rect 158496 171890 158548 171896
rect 158508 169794 158536 171890
rect 159060 169794 159088 172026
rect 160336 171880 160388 171886
rect 160336 171822 160388 171828
rect 159600 171812 159652 171818
rect 159600 171754 159652 171760
rect 159612 169794 159640 171754
rect 160348 169794 160376 171822
rect 160716 169794 160744 172094
rect 161084 172022 161112 182836
rect 161256 172900 161308 172906
rect 161256 172842 161308 172848
rect 161072 172016 161124 172022
rect 161072 171958 161124 171964
rect 161268 169794 161296 172842
rect 161452 171750 161480 182836
rect 161808 173036 161860 173042
rect 161808 172978 161860 172984
rect 161440 171744 161492 171750
rect 161440 171686 161492 171692
rect 161820 169794 161848 172978
rect 161912 172906 161940 182836
rect 161900 172900 161952 172906
rect 161900 172842 161952 172848
rect 162280 172838 162308 182836
rect 162452 180516 162504 180522
rect 162452 180458 162504 180464
rect 162360 180244 162412 180250
rect 162360 180186 162412 180192
rect 162372 172974 162400 180186
rect 162464 173042 162492 180458
rect 162648 180454 162676 182836
rect 163108 180794 163136 182836
rect 163096 180788 163148 180794
rect 163096 180730 163148 180736
rect 162636 180448 162688 180454
rect 162636 180390 162688 180396
rect 163476 180114 163504 182836
rect 163568 182822 163858 182850
rect 163464 180108 163516 180114
rect 163464 180050 163516 180056
rect 163568 179978 163596 182822
rect 163832 180584 163884 180590
rect 163832 180526 163884 180532
rect 163740 180380 163792 180386
rect 163740 180322 163792 180328
rect 163556 179972 163608 179978
rect 163556 179914 163608 179920
rect 162452 173036 162504 173042
rect 162452 172978 162504 172984
rect 163188 173036 163240 173042
rect 163188 172978 163240 172984
rect 162360 172968 162412 172974
rect 162360 172910 162412 172916
rect 162268 172832 162320 172838
rect 162268 172774 162320 172780
rect 162544 172288 162596 172294
rect 162544 172230 162596 172236
rect 162556 169794 162584 172230
rect 163200 169930 163228 172978
rect 163752 172974 163780 180322
rect 163844 173042 163872 180526
rect 164304 180046 164332 182836
rect 164672 180658 164700 182836
rect 231280 181785 231308 188210
rect 231266 181776 231322 181785
rect 231266 181711 231322 181720
rect 164660 180652 164712 180658
rect 164660 180594 164712 180600
rect 164292 180040 164344 180046
rect 164292 179982 164344 179988
rect 179576 175830 179604 177940
rect 179564 175824 179616 175830
rect 179564 175766 179616 175772
rect 173400 175688 173452 175694
rect 173400 175630 173452 175636
rect 170640 175144 170692 175150
rect 170640 175086 170692 175092
rect 163832 173036 163884 173042
rect 163832 172978 163884 172984
rect 164660 173036 164712 173042
rect 164660 172978 164712 172984
rect 163464 172968 163516 172974
rect 163464 172910 163516 172916
rect 163740 172968 163792 172974
rect 163740 172910 163792 172916
rect 163200 169902 163274 169930
rect 155104 169766 155440 169794
rect 155656 169766 155992 169794
rect 156208 169766 156544 169794
rect 156852 169766 157188 169794
rect 157588 169766 157740 169794
rect 157956 169766 158292 169794
rect 158508 169766 158844 169794
rect 159060 169766 159396 169794
rect 159612 169766 159948 169794
rect 160348 169766 160500 169794
rect 160716 169766 161052 169794
rect 161268 169766 161604 169794
rect 161820 169766 162156 169794
rect 162556 169766 162708 169794
rect 163246 169780 163274 169902
rect 163476 169794 163504 172910
rect 164474 172528 164530 172537
rect 164474 172463 164530 172472
rect 164488 169794 164516 172463
rect 163476 169766 163812 169794
rect 164456 169766 164516 169794
rect 164672 169794 164700 172978
rect 165212 172968 165264 172974
rect 165212 172910 165264 172916
rect 166314 172936 166370 172945
rect 165224 169794 165252 172910
rect 166314 172871 166370 172880
rect 165854 172800 165910 172809
rect 165854 172735 165910 172744
rect 165868 169794 165896 172735
rect 166328 169794 166356 172871
rect 167420 172628 167472 172634
rect 167420 172570 167472 172576
rect 167236 172424 167288 172430
rect 167236 172366 167288 172372
rect 167248 169794 167276 172366
rect 164672 169766 165008 169794
rect 165224 169766 165560 169794
rect 165868 169766 166112 169794
rect 166328 169766 166664 169794
rect 167216 169766 167276 169794
rect 167432 169794 167460 172570
rect 167972 172560 168024 172566
rect 167972 172502 168024 172508
rect 167984 169794 168012 172502
rect 168616 172492 168668 172498
rect 168616 172434 168668 172440
rect 168628 169794 168656 172434
rect 170178 172392 170234 172401
rect 169076 172356 169128 172362
rect 170178 172327 170234 172336
rect 169076 172298 169128 172304
rect 169088 169794 169116 172298
rect 169994 172256 170050 172265
rect 169994 172191 170050 172200
rect 170008 169794 170036 172191
rect 167432 169766 167768 169794
rect 167984 169766 168320 169794
rect 168628 169766 168872 169794
rect 169088 169766 169424 169794
rect 169976 169766 170036 169794
rect 170192 169794 170220 172327
rect 170192 169766 170528 169794
rect 143204 169630 143632 169658
rect 145964 169630 146392 169658
rect 140830 167768 140886 167777
rect 140830 167703 140886 167712
rect 140370 164368 140426 164377
rect 140370 164303 140426 164312
rect 140384 163454 140412 164303
rect 140554 163824 140610 163833
rect 140554 163759 140610 163768
rect 140568 163590 140596 163759
rect 140556 163584 140608 163590
rect 140556 163526 140608 163532
rect 140648 163516 140700 163522
rect 140648 163458 140700 163464
rect 140372 163448 140424 163454
rect 140660 163425 140688 163458
rect 140372 163390 140424 163396
rect 140646 163416 140702 163425
rect 140646 163351 140702 163360
rect 140462 162600 140518 162609
rect 140462 162535 140518 162544
rect 140476 162162 140504 162535
rect 140554 162192 140610 162201
rect 140464 162156 140516 162162
rect 140554 162127 140610 162136
rect 140464 162098 140516 162104
rect 140568 162094 140596 162127
rect 140556 162088 140608 162094
rect 140556 162030 140608 162036
rect 140462 160832 140518 160841
rect 140462 160767 140518 160776
rect 140476 160666 140504 160767
rect 140464 160660 140516 160666
rect 140464 160602 140516 160608
rect 140740 159368 140792 159374
rect 140740 159310 140792 159316
rect 140370 158384 140426 158393
rect 140370 158319 140426 158328
rect 140384 158014 140412 158319
rect 140648 158144 140700 158150
rect 140648 158086 140700 158092
rect 140556 158076 140608 158082
rect 140556 158018 140608 158024
rect 140372 158008 140424 158014
rect 140372 157950 140424 157956
rect 140464 156784 140516 156790
rect 140464 156726 140516 156732
rect 140372 156580 140424 156586
rect 140372 156522 140424 156528
rect 140384 143433 140412 156522
rect 140476 144793 140504 156726
rect 140568 146153 140596 158018
rect 140660 147513 140688 158086
rect 140752 148873 140780 159310
rect 140844 157198 140872 167703
rect 140924 159504 140976 159510
rect 140924 159446 140976 159452
rect 140832 157192 140884 157198
rect 140832 157134 140884 157140
rect 140936 149417 140964 159446
rect 140922 149408 140978 149417
rect 140922 149343 140978 149352
rect 140738 148864 140794 148873
rect 140738 148799 140794 148808
rect 140646 147504 140702 147513
rect 140646 147439 140702 147448
rect 140554 146144 140610 146153
rect 140554 146079 140610 146088
rect 140462 144784 140518 144793
rect 140462 144719 140518 144728
rect 140370 143424 140426 143433
rect 140370 143359 140426 143368
rect 142776 141886 143112 141914
rect 143572 141886 143632 141914
rect 144124 141886 144184 141914
rect 144676 141886 144736 141914
rect 145136 141886 145196 141914
rect 145688 141886 145748 141914
rect 146240 141886 146300 141914
rect 146792 141886 146852 141914
rect 147252 141886 147312 141914
rect 147804 141886 147864 141914
rect 148356 141886 148416 141914
rect 148908 141886 148968 141914
rect 149368 141886 149428 141914
rect 149920 141886 149980 141914
rect 150472 141886 150532 141914
rect 151024 141886 151084 141914
rect 151484 141886 151544 141914
rect 152036 141886 152096 141914
rect 152588 141886 152648 141914
rect 153048 141886 153108 141914
rect 153600 141886 153660 141914
rect 154152 141886 154212 141914
rect 154704 141886 154764 141914
rect 155164 141886 155224 141914
rect 155716 141886 155776 141914
rect 156268 141886 156328 141914
rect 156820 141886 156880 141914
rect 157280 141886 157340 141914
rect 140280 139852 140332 139858
rect 140280 139794 140332 139800
rect 75788 139444 75840 139450
rect 75788 139386 75840 139392
rect 137980 139376 138032 139382
rect 137980 139318 138032 139324
rect 69808 139240 69860 139246
rect 69808 139182 69860 139188
rect 75144 139240 75196 139246
rect 75144 139182 75196 139188
rect 137888 139240 137940 139246
rect 137888 139182 137940 139188
rect 69164 138900 69216 138906
rect 69164 138842 69216 138848
rect 137796 138832 137848 138838
rect 137796 138774 137848 138780
rect 68428 138764 68480 138770
rect 68428 138706 68480 138712
rect 137704 138764 137756 138770
rect 137704 138706 137756 138712
rect 137612 138696 137664 138702
rect 137612 138638 137664 138644
rect 137520 138628 137572 138634
rect 137520 138570 137572 138576
rect 126480 135840 126532 135846
rect 126480 135782 126532 135788
rect 126492 133740 126520 135782
rect 136876 132984 136928 132990
rect 136874 132952 136876 132961
rect 136928 132952 136930 132961
rect 136874 132887 136930 132896
rect 68336 131624 68388 131630
rect 68336 131566 68388 131572
rect 67232 131420 67284 131426
rect 67232 131362 67284 131368
rect 67968 131012 68020 131018
rect 67968 130954 68020 130960
rect 67508 130740 67560 130746
rect 67508 130682 67560 130688
rect 67140 130536 67192 130542
rect 67140 130478 67192 130484
rect 67060 128694 67166 128722
rect 67520 128708 67548 130682
rect 67980 128708 68008 130954
rect 68348 128708 68376 131566
rect 69072 131148 69124 131154
rect 69072 131090 69124 131096
rect 68704 130604 68756 130610
rect 68704 130546 68756 130552
rect 68716 128708 68744 130546
rect 69084 128708 69112 131090
rect 70268 130944 70320 130950
rect 70268 130886 70320 130892
rect 69532 130808 69584 130814
rect 69532 130750 69584 130756
rect 69544 128708 69572 130750
rect 69900 130672 69952 130678
rect 69900 130614 69952 130620
rect 69912 128708 69940 130614
rect 70280 128708 70308 130886
rect 70636 130400 70688 130406
rect 70636 130342 70688 130348
rect 70648 128708 70676 130342
rect 136876 130264 136928 130270
rect 136876 130206 136928 130212
rect 136888 130105 136916 130206
rect 136874 130096 136930 130105
rect 136874 130031 136930 130040
rect 136874 127920 136930 127929
rect 136874 127855 136930 127864
rect 136888 127550 136916 127855
rect 136876 127544 136928 127550
rect 136876 127486 136928 127492
rect 47818 123296 47874 123305
rect 47818 123231 47874 123240
rect 47832 122246 47860 123231
rect 47820 122240 47872 122246
rect 51316 122240 51368 122246
rect 47820 122182 47872 122188
rect 51314 122208 51316 122217
rect 51368 122208 51370 122217
rect 47084 109524 47136 109530
rect 47084 109466 47136 109472
rect 38250 109424 38306 109433
rect 38250 109359 38306 109368
rect 47832 108345 47860 122182
rect 51314 122143 51370 122152
rect 137334 115272 137390 115281
rect 137334 115207 137336 115216
rect 137388 115207 137390 115216
rect 137336 115178 137388 115184
rect 137428 112380 137480 112386
rect 137428 112322 137480 112328
rect 51316 109524 51368 109530
rect 51316 109466 51368 109472
rect 51328 108889 51356 109466
rect 74038 109016 74094 109025
rect 74038 108951 74094 108960
rect 51314 108880 51370 108889
rect 51314 108815 51370 108824
rect 47082 108336 47138 108345
rect 47082 108271 47138 108280
rect 47818 108336 47874 108345
rect 47818 108271 47874 108280
rect 38250 100720 38306 100729
rect 38250 100655 38306 100664
rect 38264 78522 38292 100655
rect 45796 94428 45848 94434
rect 45796 94370 45848 94376
rect 45808 93006 45836 94370
rect 38804 93000 38856 93006
rect 38802 92968 38804 92977
rect 45796 93000 45848 93006
rect 38856 92968 38858 92977
rect 45796 92942 45848 92948
rect 38802 92903 38858 92912
rect 38252 78516 38304 78522
rect 38252 78458 38304 78464
rect 47096 61969 47124 108271
rect 74052 97154 74080 108951
rect 137336 108232 137388 108238
rect 137336 108174 137388 108180
rect 74040 97148 74092 97154
rect 74040 97090 74092 97096
rect 81676 97148 81728 97154
rect 81676 97090 81728 97096
rect 81688 96921 81716 97090
rect 137348 97057 137376 108174
rect 137440 100865 137468 112322
rect 137532 111745 137560 138570
rect 137624 114873 137652 138638
rect 137716 117865 137744 138706
rect 137808 120585 137836 138774
rect 137900 127385 137928 139182
rect 137886 127376 137942 127385
rect 137886 127311 137942 127320
rect 137888 124824 137940 124830
rect 137888 124766 137940 124772
rect 137794 120576 137850 120585
rect 137794 120511 137850 120520
rect 137796 117888 137848 117894
rect 137702 117856 137758 117865
rect 137796 117830 137848 117836
rect 137702 117791 137758 117800
rect 137704 115168 137756 115174
rect 137704 115110 137756 115116
rect 137610 114864 137666 114873
rect 137610 114799 137666 114808
rect 137518 111736 137574 111745
rect 137518 111671 137574 111680
rect 137518 109696 137574 109705
rect 137518 109631 137574 109640
rect 137426 100856 137482 100865
rect 137426 100791 137482 100800
rect 137334 97048 137390 97057
rect 137334 96983 137390 96992
rect 81674 96912 81730 96921
rect 81674 96847 81730 96856
rect 51314 95552 51370 95561
rect 51314 95487 51370 95496
rect 51328 94434 51356 95487
rect 51316 94428 51368 94434
rect 51316 94370 51368 94376
rect 55100 87498 55128 88860
rect 55088 87492 55140 87498
rect 55088 87434 55140 87440
rect 53984 87288 54036 87294
rect 53984 87230 54036 87236
rect 52604 87084 52656 87090
rect 52604 87026 52656 87032
rect 51224 87016 51276 87022
rect 51224 86958 51276 86964
rect 49844 86880 49896 86886
rect 49844 86822 49896 86828
rect 49200 78516 49252 78522
rect 49200 78458 49252 78464
rect 49212 75804 49240 78458
rect 49856 75804 49884 86822
rect 51132 86812 51184 86818
rect 51132 86754 51184 86760
rect 50488 79196 50540 79202
rect 50488 79138 50540 79144
rect 50500 75804 50528 79138
rect 51144 75804 51172 86754
rect 51236 79202 51264 86958
rect 52512 86948 52564 86954
rect 52512 86890 52564 86896
rect 52524 79202 52552 86890
rect 51224 79196 51276 79202
rect 51224 79138 51276 79144
rect 51776 79196 51828 79202
rect 51776 79138 51828 79144
rect 52512 79196 52564 79202
rect 52512 79138 52564 79144
rect 51788 75804 51816 79138
rect 52616 75818 52644 87026
rect 53156 78516 53208 78522
rect 53156 78458 53208 78464
rect 52538 75790 52644 75818
rect 53168 75804 53196 78458
rect 53996 75818 54024 87230
rect 55468 86274 55496 88860
rect 55836 86342 55864 88860
rect 56100 87492 56152 87498
rect 56100 87434 56152 87440
rect 55824 86336 55876 86342
rect 55824 86278 55876 86284
rect 55456 86268 55508 86274
rect 55456 86210 55508 86216
rect 54444 79060 54496 79066
rect 54444 79002 54496 79008
rect 53826 75790 54024 75818
rect 54456 75804 54484 79002
rect 55180 78584 55232 78590
rect 55180 78526 55232 78532
rect 55192 75804 55220 78526
rect 55824 78176 55876 78182
rect 55824 78118 55876 78124
rect 55836 75804 55864 78118
rect 56112 77978 56140 87434
rect 56296 86206 56324 88860
rect 56284 86200 56336 86206
rect 56284 86142 56336 86148
rect 56664 86138 56692 88860
rect 57032 86546 57060 88860
rect 57492 86750 57520 88860
rect 57480 86744 57532 86750
rect 57480 86686 57532 86692
rect 57020 86540 57072 86546
rect 57020 86482 57072 86488
rect 57860 86410 57888 88860
rect 58228 87362 58256 88860
rect 58688 87498 58716 88860
rect 58676 87492 58728 87498
rect 58676 87434 58728 87440
rect 58216 87356 58268 87362
rect 58216 87298 58268 87304
rect 59056 86818 59084 88860
rect 59044 86812 59096 86818
rect 59044 86754 59096 86760
rect 59424 86478 59452 88860
rect 59884 87430 59912 88860
rect 59872 87424 59924 87430
rect 59872 87366 59924 87372
rect 60252 87294 60280 88860
rect 60634 88846 60832 88874
rect 60240 87288 60292 87294
rect 60240 87230 60292 87236
rect 59412 86472 59464 86478
rect 59412 86414 59464 86420
rect 57848 86404 57900 86410
rect 57848 86346 57900 86352
rect 60516 86336 60568 86342
rect 60516 86278 60568 86284
rect 60332 86268 60384 86274
rect 60332 86210 60384 86216
rect 56652 86132 56704 86138
rect 56652 86074 56704 86080
rect 60240 86132 60292 86138
rect 60240 86074 60292 86080
rect 56468 79196 56520 79202
rect 56468 79138 56520 79144
rect 56100 77972 56152 77978
rect 56100 77914 56152 77920
rect 56480 75804 56508 79138
rect 59136 78924 59188 78930
rect 59136 78866 59188 78872
rect 58492 78244 58544 78250
rect 58492 78186 58544 78192
rect 57848 78108 57900 78114
rect 57848 78050 57900 78056
rect 57112 77904 57164 77910
rect 57112 77846 57164 77852
rect 57124 75804 57152 77846
rect 57860 75804 57888 78050
rect 58504 75804 58532 78186
rect 59148 75804 59176 78866
rect 60252 78232 60280 86074
rect 60344 78590 60372 86210
rect 60424 86200 60476 86206
rect 60424 86142 60476 86148
rect 60332 78584 60384 78590
rect 60332 78526 60384 78532
rect 60436 78454 60464 86142
rect 60528 78998 60556 86278
rect 60516 78992 60568 78998
rect 60516 78934 60568 78940
rect 60804 78833 60832 88846
rect 60884 86608 60936 86614
rect 60884 86550 60936 86556
rect 60790 78824 60846 78833
rect 60790 78759 60846 78768
rect 60424 78448 60476 78454
rect 60424 78390 60476 78396
rect 60424 78244 60476 78250
rect 60252 78204 60424 78232
rect 60424 78186 60476 78192
rect 59780 78040 59832 78046
rect 59780 77982 59832 77988
rect 59792 75804 59820 77982
rect 60896 75818 60924 86550
rect 61080 86342 61108 88860
rect 61462 88846 61568 88874
rect 61830 88846 62120 88874
rect 61344 86676 61396 86682
rect 61344 86618 61396 86624
rect 61068 86336 61120 86342
rect 61068 86278 61120 86284
rect 61356 75818 61384 86618
rect 61540 78697 61568 88846
rect 61804 86744 61856 86750
rect 61804 86686 61856 86692
rect 61712 86540 61764 86546
rect 61712 86482 61764 86488
rect 61620 86404 61672 86410
rect 61620 86346 61672 86352
rect 61632 78726 61660 86346
rect 61724 78862 61752 86482
rect 61712 78856 61764 78862
rect 61712 78798 61764 78804
rect 61816 78794 61844 86686
rect 61988 86540 62040 86546
rect 61988 86482 62040 86488
rect 61896 86404 61948 86410
rect 61896 86346 61948 86352
rect 61908 79066 61936 86346
rect 62000 86342 62028 86482
rect 61988 86336 62040 86342
rect 61988 86278 62040 86284
rect 61988 86200 62040 86206
rect 61988 86142 62040 86148
rect 61896 79060 61948 79066
rect 61896 79002 61948 79008
rect 61804 78788 61856 78794
rect 61804 78730 61856 78736
rect 61620 78720 61672 78726
rect 61526 78688 61582 78697
rect 61620 78662 61672 78668
rect 62000 78658 62028 86142
rect 61526 78623 61582 78632
rect 61988 78652 62040 78658
rect 61988 78594 62040 78600
rect 62092 78561 62120 88846
rect 62184 88846 62290 88874
rect 62078 78552 62134 78561
rect 62078 78487 62134 78496
rect 62184 78425 62212 88846
rect 62264 86336 62316 86342
rect 62264 86278 62316 86284
rect 62170 78416 62226 78425
rect 62170 78351 62226 78360
rect 62276 75818 62304 86278
rect 62644 86138 62672 88860
rect 63104 86886 63132 88860
rect 63472 87022 63500 88860
rect 63840 87158 63868 88860
rect 63828 87152 63880 87158
rect 63828 87094 63880 87100
rect 63460 87016 63512 87022
rect 63460 86958 63512 86964
rect 64300 86954 64328 88860
rect 64668 87090 64696 88860
rect 64656 87084 64708 87090
rect 64656 87026 64708 87032
rect 64288 86948 64340 86954
rect 64288 86890 64340 86896
rect 63092 86880 63144 86886
rect 63092 86822 63144 86828
rect 63644 86880 63696 86886
rect 63644 86822 63696 86828
rect 62632 86132 62684 86138
rect 62632 86074 62684 86080
rect 63552 86132 63604 86138
rect 63552 86074 63604 86080
rect 62448 79196 62500 79202
rect 62448 79138 62500 79144
rect 60542 75790 60924 75818
rect 61186 75790 61384 75818
rect 61830 75790 62304 75818
rect 62460 75804 62488 79138
rect 63564 78522 63592 86074
rect 63656 79202 63684 86822
rect 64380 86268 64432 86274
rect 64380 86210 64432 86216
rect 63644 79196 63696 79202
rect 63644 79138 63696 79144
rect 63828 78584 63880 78590
rect 63828 78526 63880 78532
rect 63552 78516 63604 78522
rect 63552 78458 63604 78464
rect 63184 77972 63236 77978
rect 63184 77914 63236 77920
rect 63196 75804 63224 77914
rect 63840 75804 63868 78526
rect 64392 77910 64420 86210
rect 65036 86206 65064 88860
rect 65496 87498 65524 88860
rect 65484 87492 65536 87498
rect 65484 87434 65536 87440
rect 65864 86410 65892 88860
rect 65956 88846 66246 88874
rect 65852 86404 65904 86410
rect 65852 86346 65904 86352
rect 65956 86290 65984 88846
rect 65220 86262 65984 86290
rect 65024 86200 65076 86206
rect 65024 86142 65076 86148
rect 64472 78992 64524 78998
rect 64472 78934 64524 78940
rect 64380 77904 64432 77910
rect 64380 77846 64432 77852
rect 64484 75804 64512 78934
rect 65116 78448 65168 78454
rect 65116 78390 65168 78396
rect 65128 75804 65156 78390
rect 65220 78250 65248 86262
rect 65760 86200 65812 86206
rect 65760 86142 65812 86148
rect 65772 79066 65800 86142
rect 66692 86138 66720 88860
rect 66772 86812 66824 86818
rect 66772 86754 66824 86760
rect 66784 86138 66812 86754
rect 67060 86206 67088 88860
rect 67140 87356 67192 87362
rect 67140 87298 67192 87304
rect 67048 86200 67100 86206
rect 67048 86142 67100 86148
rect 65852 86132 65904 86138
rect 65852 86074 65904 86080
rect 66680 86132 66732 86138
rect 66680 86074 66732 86080
rect 66772 86132 66824 86138
rect 66772 86074 66824 86080
rect 65760 79060 65812 79066
rect 65760 79002 65812 79008
rect 65208 78244 65260 78250
rect 65208 78186 65260 78192
rect 65864 78182 65892 86074
rect 67152 78930 67180 87298
rect 67232 87220 67284 87226
rect 67232 87162 67284 87168
rect 67140 78924 67192 78930
rect 67140 78866 67192 78872
rect 66496 78856 66548 78862
rect 66496 78798 66548 78804
rect 65852 78176 65904 78182
rect 65852 78118 65904 78124
rect 65760 78108 65812 78114
rect 65760 78050 65812 78056
rect 65772 75804 65800 78050
rect 66508 75804 66536 78798
rect 67140 78788 67192 78794
rect 67140 78730 67192 78736
rect 67152 75804 67180 78730
rect 67244 78250 67272 87162
rect 67324 86472 67376 86478
rect 67324 86414 67376 86420
rect 67232 78244 67284 78250
rect 67232 78186 67284 78192
rect 67336 78114 67364 86414
rect 67428 86274 67456 88860
rect 67416 86268 67468 86274
rect 67416 86210 67468 86216
rect 67416 86132 67468 86138
rect 67416 86074 67468 86080
rect 67508 86132 67560 86138
rect 67508 86074 67560 86080
rect 67428 78386 67456 86074
rect 67416 78380 67468 78386
rect 67416 78322 67468 78328
rect 67324 78108 67376 78114
rect 67324 78050 67376 78056
rect 67520 78046 67548 86074
rect 67888 83894 67916 88860
rect 67980 88846 68270 88874
rect 68348 88846 68638 88874
rect 67876 83888 67928 83894
rect 67876 83830 67928 83836
rect 67784 78720 67836 78726
rect 67784 78662 67836 78668
rect 67508 78040 67560 78046
rect 67508 77982 67560 77988
rect 67796 75804 67824 78662
rect 67980 78454 68008 88846
rect 68348 83978 68376 88846
rect 69084 86138 69112 88860
rect 69452 86614 69480 88860
rect 69820 86682 69848 88860
rect 69808 86676 69860 86682
rect 69808 86618 69860 86624
rect 69440 86608 69492 86614
rect 69440 86550 69492 86556
rect 69900 86540 69952 86546
rect 69900 86482 69952 86488
rect 69072 86132 69124 86138
rect 69072 86074 69124 86080
rect 68072 83950 68376 83978
rect 68072 78862 68100 83950
rect 68244 83888 68296 83894
rect 68244 83830 68296 83836
rect 68060 78856 68112 78862
rect 68060 78798 68112 78804
rect 68256 78658 68284 83830
rect 68428 78924 68480 78930
rect 68428 78866 68480 78872
rect 68244 78652 68296 78658
rect 68244 78594 68296 78600
rect 67968 78448 68020 78454
rect 67968 78390 68020 78396
rect 68440 75804 68468 78866
rect 69912 78862 69940 86482
rect 70280 86342 70308 88860
rect 70648 86886 70676 88860
rect 70728 87424 70780 87430
rect 70728 87366 70780 87372
rect 70636 86880 70688 86886
rect 70636 86822 70688 86828
rect 70268 86336 70320 86342
rect 70268 86278 70320 86284
rect 69900 78856 69952 78862
rect 69900 78798 69952 78804
rect 69808 78380 69860 78386
rect 69808 78322 69860 78328
rect 69164 78244 69216 78250
rect 69164 78186 69216 78192
rect 69176 75804 69204 78186
rect 69820 75804 69848 78322
rect 70452 78108 70504 78114
rect 70452 78050 70504 78056
rect 70464 75804 70492 78050
rect 70740 75818 70768 87366
rect 70820 87288 70872 87294
rect 70820 87230 70872 87236
rect 70832 75920 70860 87230
rect 136874 85624 136930 85633
rect 136874 85559 136930 85568
rect 136888 85254 136916 85559
rect 136876 85248 136928 85254
rect 136876 85190 136928 85196
rect 136876 84704 136928 84710
rect 136874 84672 136876 84681
rect 136928 84672 136930 84681
rect 136874 84607 136930 84616
rect 85170 84128 85226 84137
rect 85092 84086 85170 84114
rect 85092 81990 85120 84086
rect 85226 84086 85566 84114
rect 85170 84063 85226 84072
rect 92256 84024 92308 84030
rect 92256 83966 92308 83972
rect 92268 83964 92296 83966
rect 89600 83962 89628 83964
rect 90888 83962 90916 83964
rect 116556 83962 116584 83964
rect 120604 83962 120632 83964
rect 124652 83962 124680 83964
rect 127320 83962 127348 83964
rect 89588 83956 89640 83962
rect 89588 83898 89640 83904
rect 90876 83956 90928 83962
rect 90876 83898 90928 83904
rect 116544 83956 116596 83962
rect 116544 83898 116596 83904
rect 120592 83956 120644 83962
rect 120592 83898 120644 83904
rect 124640 83956 124692 83962
rect 124640 83898 124692 83904
rect 127308 83956 127360 83962
rect 127308 83898 127360 83904
rect 132748 83894 132776 83964
rect 134852 83956 134904 83962
rect 134852 83898 134904 83904
rect 86828 83888 86880 83894
rect 86828 83830 86880 83836
rect 88208 83888 88260 83894
rect 88208 83830 88260 83836
rect 93636 83888 93688 83894
rect 93636 83830 93688 83836
rect 94924 83888 94976 83894
rect 94924 83830 94976 83836
rect 96304 83888 96356 83894
rect 96304 83830 96356 83836
rect 97684 83888 97736 83894
rect 97684 83830 97736 83836
rect 98972 83888 99024 83894
rect 98972 83830 99024 83836
rect 100352 83888 100404 83894
rect 100352 83830 100404 83836
rect 101732 83888 101784 83894
rect 101732 83830 101784 83836
rect 103020 83888 103072 83894
rect 103020 83830 103072 83836
rect 104400 83888 104452 83894
rect 104400 83830 104452 83836
rect 105780 83888 105832 83894
rect 105780 83830 105832 83836
rect 107068 83888 107120 83894
rect 107068 83830 107120 83836
rect 108448 83888 108500 83894
rect 108448 83830 108500 83836
rect 109828 83888 109880 83894
rect 109828 83830 109880 83836
rect 111116 83888 111168 83894
rect 111116 83830 111168 83836
rect 112496 83888 112548 83894
rect 112496 83830 112548 83836
rect 113876 83888 113928 83894
rect 113876 83830 113928 83836
rect 115164 83888 115216 83894
rect 115164 83830 115216 83836
rect 117924 83888 117976 83894
rect 117924 83830 117976 83836
rect 119212 83888 119264 83894
rect 119212 83830 119264 83836
rect 121972 83888 122024 83894
rect 121972 83830 122024 83836
rect 123260 83888 123312 83894
rect 123260 83830 123312 83836
rect 126020 83888 126072 83894
rect 126020 83830 126072 83836
rect 128688 83888 128740 83894
rect 128688 83830 128740 83836
rect 132736 83888 132788 83894
rect 132736 83830 132788 83836
rect 86840 83828 86868 83830
rect 88220 83828 88248 83830
rect 93648 83828 93676 83830
rect 94936 83828 94964 83830
rect 96316 83828 96344 83830
rect 97696 83828 97724 83830
rect 98984 83828 99012 83830
rect 100364 83828 100392 83830
rect 101744 83828 101772 83830
rect 103032 83828 103060 83830
rect 104412 83828 104440 83830
rect 105792 83828 105820 83830
rect 107080 83828 107108 83830
rect 108460 83828 108488 83830
rect 109840 83828 109868 83830
rect 111128 83828 111156 83830
rect 112508 83828 112536 83830
rect 113888 83828 113916 83830
rect 115176 83828 115204 83830
rect 117936 83828 117964 83830
rect 119224 83828 119252 83830
rect 121984 83828 122012 83830
rect 123272 83828 123300 83830
rect 126032 83828 126060 83830
rect 128700 83828 128728 83830
rect 91980 83820 92032 83826
rect 91980 83762 92032 83768
rect 96120 83820 96172 83826
rect 96120 83762 96172 83768
rect 99524 83820 99576 83826
rect 99524 83762 99576 83768
rect 100904 83820 100956 83826
rect 100904 83762 100956 83768
rect 102284 83820 102336 83826
rect 102284 83762 102336 83768
rect 103664 83820 103716 83826
rect 103664 83762 103716 83768
rect 105044 83820 105096 83826
rect 105044 83762 105096 83768
rect 106424 83820 106476 83826
rect 106424 83762 106476 83768
rect 107804 83820 107856 83826
rect 107804 83762 107856 83768
rect 112956 83820 113008 83826
rect 112956 83762 113008 83768
rect 125560 83820 125612 83826
rect 125560 83762 125612 83768
rect 133380 83820 133432 83826
rect 134142 83814 134800 83842
rect 133380 83762 133432 83768
rect 85080 81984 85132 81990
rect 85080 81926 85132 81932
rect 79560 81780 79612 81786
rect 79560 81722 79612 81728
rect 73120 78856 73172 78862
rect 72474 78824 72530 78833
rect 73120 78798 73172 78804
rect 72474 78759 72530 78768
rect 70832 75892 71412 75920
rect 70740 75790 71122 75818
rect 71384 75682 71412 75892
rect 72488 75804 72516 78759
rect 73132 75804 73160 78798
rect 73762 78688 73818 78697
rect 73762 78623 73818 78632
rect 73776 75804 73804 78623
rect 74498 78552 74554 78561
rect 74498 78487 74554 78496
rect 75788 78516 75840 78522
rect 74512 75804 74540 78487
rect 75788 78458 75840 78464
rect 75142 78416 75198 78425
rect 75142 78351 75198 78360
rect 75156 75804 75184 78351
rect 75800 75804 75828 78458
rect 71384 75654 71858 75682
rect 76458 75382 76564 75410
rect 47082 61960 47138 61969
rect 47082 61895 47138 61904
rect 62920 46086 62948 47924
rect 62908 46080 62960 46086
rect 62908 46022 62960 46028
rect 63644 46080 63696 46086
rect 63644 46022 63696 46028
rect 63656 37110 63684 46022
rect 63644 37104 63696 37110
rect 63644 37046 63696 37052
rect 76536 20926 76564 75382
rect 79572 71625 79600 81722
rect 79744 81712 79796 81718
rect 79744 81654 79796 81660
rect 79652 81576 79704 81582
rect 79652 81518 79704 81524
rect 79664 73257 79692 81518
rect 79650 73248 79706 73257
rect 79650 73183 79706 73192
rect 79756 72169 79784 81654
rect 79836 81644 79888 81650
rect 79836 81586 79888 81592
rect 79848 72713 79876 81586
rect 79928 81508 79980 81514
rect 79928 81450 79980 81456
rect 79940 73937 79968 81450
rect 80020 81440 80072 81446
rect 80020 81382 80072 81388
rect 80032 74481 80060 81382
rect 80112 81372 80164 81378
rect 80112 81314 80164 81320
rect 80124 75025 80152 81314
rect 80204 81304 80256 81310
rect 80204 81246 80256 81252
rect 80216 75569 80244 81246
rect 80202 75560 80258 75569
rect 80202 75495 80258 75504
rect 80110 75016 80166 75025
rect 80110 74951 80166 74960
rect 80018 74472 80074 74481
rect 80018 74407 80074 74416
rect 79926 73928 79982 73937
rect 79926 73863 79982 73872
rect 79834 72704 79890 72713
rect 79834 72639 79890 72648
rect 79742 72160 79798 72169
rect 79742 72095 79798 72104
rect 79558 71616 79614 71625
rect 79558 71551 79614 71560
rect 80202 71072 80258 71081
rect 80202 71007 80258 71016
rect 80216 70974 80244 71007
rect 80204 70968 80256 70974
rect 80204 70910 80256 70916
rect 84436 70968 84488 70974
rect 84436 70910 84488 70916
rect 84448 70294 84476 70910
rect 84436 70288 84488 70294
rect 84436 70230 84488 70236
rect 79466 69984 79522 69993
rect 79466 69919 79522 69928
rect 79480 69682 79508 69919
rect 80202 69848 80258 69857
rect 80202 69783 80258 69792
rect 79468 69676 79520 69682
rect 79468 69618 79520 69624
rect 80216 69614 80244 69783
rect 80204 69608 80256 69614
rect 80204 69550 80256 69556
rect 80202 69032 80258 69041
rect 80202 68967 80258 68976
rect 80216 68866 80244 68967
rect 80204 68860 80256 68866
rect 80204 68802 80256 68808
rect 80110 68488 80166 68497
rect 80110 68423 80166 68432
rect 80124 68322 80152 68423
rect 80112 68316 80164 68322
rect 80112 68258 80164 68264
rect 80204 68248 80256 68254
rect 80202 68216 80204 68225
rect 80256 68216 80258 68225
rect 80202 68151 80258 68160
rect 80204 67568 80256 67574
rect 80202 67536 80204 67545
rect 80256 67536 80258 67545
rect 80112 67500 80164 67506
rect 80202 67471 80258 67480
rect 80112 67442 80164 67448
rect 80124 67001 80152 67442
rect 80110 66992 80166 67001
rect 80110 66927 80166 66936
rect 80110 66448 80166 66457
rect 80110 66383 80166 66392
rect 80124 66078 80152 66383
rect 80204 66140 80256 66146
rect 80204 66082 80256 66088
rect 80112 66072 80164 66078
rect 80112 66014 80164 66020
rect 80216 65913 80244 66082
rect 80202 65904 80258 65913
rect 80202 65839 80258 65848
rect 80204 65392 80256 65398
rect 80202 65360 80204 65369
rect 80256 65360 80258 65369
rect 80202 65295 80258 65304
rect 80112 64780 80164 64786
rect 80112 64722 80164 64728
rect 80124 64145 80152 64722
rect 80204 64712 80256 64718
rect 80202 64680 80204 64689
rect 80256 64680 80258 64689
rect 80202 64615 80258 64624
rect 80110 64136 80166 64145
rect 80110 64071 80166 64080
rect 80204 64032 80256 64038
rect 80204 63974 80256 63980
rect 80216 63601 80244 63974
rect 80202 63592 80258 63601
rect 80202 63527 80258 63536
rect 80204 63352 80256 63358
rect 80204 63294 80256 63300
rect 80216 63057 80244 63294
rect 80202 63048 80258 63057
rect 80202 62983 80258 62992
rect 80204 62604 80256 62610
rect 80204 62546 80256 62552
rect 80112 62536 80164 62542
rect 80216 62513 80244 62546
rect 80112 62478 80164 62484
rect 80202 62504 80258 62513
rect 80124 61833 80152 62478
rect 80202 62439 80258 62448
rect 80110 61824 80166 61833
rect 80110 61759 80166 61768
rect 80204 61244 80256 61250
rect 80204 61186 80256 61192
rect 80112 61176 80164 61182
rect 80112 61118 80164 61124
rect 79098 60872 79154 60881
rect 79098 60807 79154 60816
rect 79112 60366 79140 60807
rect 79100 60360 79152 60366
rect 79100 60302 79152 60308
rect 80124 60201 80152 61118
rect 80216 60745 80244 61186
rect 80202 60736 80258 60745
rect 80202 60671 80258 60680
rect 80110 60192 80166 60201
rect 80110 60127 80166 60136
rect 80112 59884 80164 59890
rect 80112 59826 80164 59832
rect 80124 58977 80152 59826
rect 80204 59816 80256 59822
rect 80204 59758 80256 59764
rect 80216 59657 80244 59758
rect 80202 59648 80258 59657
rect 80202 59583 80258 59592
rect 80110 58968 80166 58977
rect 80110 58903 80166 58912
rect 80020 58592 80072 58598
rect 80020 58534 80072 58540
rect 80032 55577 80060 58534
rect 80112 58524 80164 58530
rect 80112 58466 80164 58472
rect 80124 57889 80152 58466
rect 80204 58456 80256 58462
rect 80202 58424 80204 58433
rect 80256 58424 80258 58433
rect 80202 58359 80258 58368
rect 80110 57880 80166 57889
rect 80110 57815 80166 57824
rect 80204 57368 80256 57374
rect 80202 57336 80204 57345
rect 80256 57336 80258 57345
rect 80202 57271 80258 57280
rect 80112 57096 80164 57102
rect 80112 57038 80164 57044
rect 80124 56121 80152 57038
rect 80204 57028 80256 57034
rect 80204 56970 80256 56976
rect 80216 56801 80244 56970
rect 80202 56792 80258 56801
rect 80202 56727 80258 56736
rect 80110 56112 80166 56121
rect 80110 56047 80166 56056
rect 80112 55736 80164 55742
rect 80112 55678 80164 55684
rect 80018 55568 80074 55577
rect 80018 55503 80074 55512
rect 79744 54580 79796 54586
rect 79744 54522 79796 54528
rect 79468 54512 79520 54518
rect 79468 54454 79520 54460
rect 79480 50409 79508 54454
rect 79756 51089 79784 54522
rect 80124 54489 80152 55678
rect 80204 55464 80256 55470
rect 80204 55406 80256 55412
rect 80216 55033 80244 55406
rect 80202 55024 80258 55033
rect 80202 54959 80258 54968
rect 80110 54480 80166 54489
rect 80110 54415 80166 54424
rect 80204 54240 80256 54246
rect 80204 54182 80256 54188
rect 80216 53945 80244 54182
rect 80202 53936 80258 53945
rect 80202 53871 80258 53880
rect 80204 53356 80256 53362
rect 80204 53298 80256 53304
rect 80216 53265 80244 53298
rect 80202 53256 80258 53265
rect 80202 53191 80258 53200
rect 80020 53016 80072 53022
rect 80020 52958 80072 52964
rect 79742 51080 79798 51089
rect 79742 51015 79798 51024
rect 79466 50400 79522 50409
rect 79466 50335 79522 50344
rect 80032 48777 80060 52958
rect 80112 52948 80164 52954
rect 80112 52890 80164 52896
rect 80124 52177 80152 52890
rect 80204 52880 80256 52886
rect 80204 52822 80256 52828
rect 80216 52721 80244 52822
rect 80202 52712 80258 52721
rect 80202 52647 80258 52656
rect 80110 52168 80166 52177
rect 80110 52103 80166 52112
rect 80202 51624 80258 51633
rect 80202 51559 80204 51568
rect 80256 51559 80258 51568
rect 80204 51530 80256 51536
rect 80110 49448 80166 49457
rect 80110 49383 80166 49392
rect 80124 48942 80152 49383
rect 80202 49312 80258 49321
rect 80202 49247 80204 49256
rect 80256 49247 80258 49256
rect 80204 49218 80256 49224
rect 80112 48936 80164 48942
rect 80112 48878 80164 48884
rect 80018 48768 80074 48777
rect 80018 48703 80074 48712
rect 79558 47544 79614 47553
rect 79558 47479 79614 47488
rect 79572 37246 79600 47479
rect 79560 37240 79612 37246
rect 79560 37182 79612 37188
rect 85092 25414 85120 81926
rect 89220 81848 89272 81854
rect 89220 81790 89272 81796
rect 89232 72402 89260 81790
rect 89772 77700 89824 77706
rect 89772 77642 89824 77648
rect 89784 72946 89812 77642
rect 89772 72940 89824 72946
rect 89772 72882 89824 72888
rect 91992 72674 92020 83762
rect 96132 72946 96160 83762
rect 96396 83752 96448 83758
rect 96396 83694 96448 83700
rect 97776 83752 97828 83758
rect 97776 83694 97828 83700
rect 96408 73558 96436 83694
rect 96396 73552 96448 73558
rect 96396 73494 96448 73500
rect 97788 73490 97816 83694
rect 97776 73484 97828 73490
rect 97776 73426 97828 73432
rect 99536 73354 99564 83762
rect 99616 81916 99668 81922
rect 99616 81858 99668 81864
rect 99628 81242 99656 81858
rect 99616 81236 99668 81242
rect 99616 81178 99668 81184
rect 100260 81236 100312 81242
rect 100260 81178 100312 81184
rect 100272 73694 100300 81178
rect 100260 73688 100312 73694
rect 100260 73630 100312 73636
rect 100916 73422 100944 83762
rect 101732 81168 101784 81174
rect 101732 81110 101784 81116
rect 101640 80760 101692 80766
rect 101640 80702 101692 80708
rect 100996 73688 101048 73694
rect 100996 73630 101048 73636
rect 100904 73416 100956 73422
rect 100904 73358 100956 73364
rect 99524 73348 99576 73354
rect 99524 73290 99576 73296
rect 95752 72940 95804 72946
rect 95752 72882 95804 72888
rect 96120 72940 96172 72946
rect 96120 72882 96172 72888
rect 98236 72940 98288 72946
rect 98236 72882 98288 72888
rect 91980 72668 92032 72674
rect 91980 72610 92032 72616
rect 93268 72668 93320 72674
rect 93268 72610 93320 72616
rect 89220 72396 89272 72402
rect 89220 72338 89272 72344
rect 90784 72396 90836 72402
rect 90784 72338 90836 72344
rect 87196 70288 87248 70294
rect 87196 70230 87248 70236
rect 87208 69721 87236 70230
rect 90796 69834 90824 72338
rect 93280 69834 93308 72610
rect 95764 69834 95792 72882
rect 98248 69834 98276 72882
rect 101008 69834 101036 73630
rect 101652 72742 101680 80702
rect 101640 72736 101692 72742
rect 101640 72678 101692 72684
rect 101744 72674 101772 81110
rect 102296 73286 102324 83762
rect 102284 73280 102336 73286
rect 102284 73222 102336 73228
rect 103676 73218 103704 83762
rect 103664 73212 103716 73218
rect 103664 73154 103716 73160
rect 105056 73150 105084 83762
rect 105044 73144 105096 73150
rect 105044 73086 105096 73092
rect 106436 73082 106464 83762
rect 106424 73076 106476 73082
rect 106424 73018 106476 73024
rect 107816 73014 107844 83762
rect 111208 80148 111260 80154
rect 111208 80090 111260 80096
rect 111220 75054 111248 80090
rect 112968 78425 112996 83762
rect 113968 83752 114020 83758
rect 113968 83694 114020 83700
rect 116636 83752 116688 83758
rect 116636 83694 116688 83700
rect 119304 83752 119356 83758
rect 119304 83694 119356 83700
rect 112954 78416 113010 78425
rect 112954 78351 113010 78360
rect 111208 75048 111260 75054
rect 111208 74990 111260 74996
rect 113980 74986 114008 83694
rect 113968 74980 114020 74986
rect 113968 74922 114020 74928
rect 116648 74918 116676 83694
rect 119316 76346 119344 83694
rect 125572 81281 125600 83762
rect 133392 83729 133420 83762
rect 133378 83720 133434 83729
rect 133378 83655 133434 83664
rect 133392 81922 133420 83655
rect 133380 81916 133432 81922
rect 133380 81858 133432 81864
rect 125558 81272 125614 81281
rect 125558 81207 125614 81216
rect 124732 80148 124784 80154
rect 124732 80090 124784 80096
rect 124744 76414 124772 80090
rect 124732 76408 124784 76414
rect 124732 76350 124784 76356
rect 119304 76340 119356 76346
rect 119304 76282 119356 76288
rect 116636 74912 116688 74918
rect 116636 74854 116688 74860
rect 108264 73552 108316 73558
rect 108264 73494 108316 73500
rect 107804 73008 107856 73014
rect 107804 72950 107856 72956
rect 105780 72736 105832 72742
rect 105780 72678 105832 72684
rect 101732 72668 101784 72674
rect 101732 72610 101784 72616
rect 103204 72668 103256 72674
rect 103204 72610 103256 72616
rect 103216 69834 103244 72610
rect 105792 69834 105820 72678
rect 108276 69834 108304 73494
rect 110748 73484 110800 73490
rect 110748 73426 110800 73432
rect 110760 69834 110788 73426
rect 115716 73416 115768 73422
rect 115716 73358 115768 73364
rect 113416 73348 113468 73354
rect 113416 73290 113468 73296
rect 113428 69834 113456 73290
rect 115728 69834 115756 73358
rect 118292 73280 118344 73286
rect 118292 73222 118344 73228
rect 118304 69834 118332 73222
rect 120776 73212 120828 73218
rect 120776 73154 120828 73160
rect 120788 69834 120816 73154
rect 123260 73144 123312 73150
rect 123260 73086 123312 73092
rect 123272 69834 123300 73086
rect 125836 73076 125888 73082
rect 125836 73018 125888 73024
rect 125848 69834 125876 73018
rect 128596 73008 128648 73014
rect 128596 72950 128648 72956
rect 128608 69834 128636 72950
rect 131356 70900 131408 70906
rect 131356 70842 131408 70848
rect 90796 69806 91132 69834
rect 93280 69806 93616 69834
rect 95764 69806 96100 69834
rect 98248 69806 98584 69834
rect 101008 69806 101068 69834
rect 103216 69806 103552 69834
rect 105792 69806 106128 69834
rect 108276 69806 108612 69834
rect 110760 69806 111096 69834
rect 113428 69806 113580 69834
rect 115728 69806 116064 69834
rect 118304 69806 118640 69834
rect 120788 69806 121124 69834
rect 123272 69806 123608 69834
rect 125848 69806 126092 69834
rect 128576 69806 128636 69834
rect 131368 69721 131396 70842
rect 87194 69712 87250 69721
rect 87194 69647 87250 69656
rect 131354 69712 131410 69721
rect 131354 69647 131410 69656
rect 87196 69540 87248 69546
rect 87196 69482 87248 69488
rect 131540 69540 131592 69546
rect 131540 69482 131592 69488
rect 87208 69313 87236 69482
rect 87288 69472 87340 69478
rect 87288 69414 87340 69420
rect 131356 69472 131408 69478
rect 131356 69414 131408 69420
rect 87194 69304 87250 69313
rect 87194 69239 87250 69248
rect 87300 68905 87328 69414
rect 131368 69313 131396 69414
rect 131448 69404 131500 69410
rect 131448 69346 131500 69352
rect 131354 69304 131410 69313
rect 131354 69239 131410 69248
rect 131460 68905 131488 69346
rect 87286 68896 87342 68905
rect 87196 68860 87248 68866
rect 87286 68831 87342 68840
rect 131446 68896 131502 68905
rect 131446 68831 131502 68840
rect 87196 68802 87248 68808
rect 87208 68497 87236 68802
rect 131552 68497 131580 69482
rect 87194 68488 87250 68497
rect 87194 68423 87250 68432
rect 131538 68488 131594 68497
rect 131538 68423 131594 68432
rect 87196 68180 87248 68186
rect 87196 68122 87248 68128
rect 132000 68180 132052 68186
rect 132000 68122 132052 68128
rect 87208 68089 87236 68122
rect 87288 68112 87340 68118
rect 87194 68080 87250 68089
rect 132012 68089 132040 68122
rect 132552 68112 132604 68118
rect 87288 68054 87340 68060
rect 131998 68080 132054 68089
rect 87194 68015 87250 68024
rect 87300 67681 87328 68054
rect 131816 68044 131868 68050
rect 132552 68054 132604 68060
rect 131998 68015 132054 68024
rect 131816 67986 131868 67992
rect 131356 67976 131408 67982
rect 131356 67918 131408 67924
rect 87286 67672 87342 67681
rect 87286 67607 87342 67616
rect 87196 67568 87248 67574
rect 87196 67510 87248 67516
rect 87208 67273 87236 67510
rect 87288 67500 87340 67506
rect 87288 67442 87340 67448
rect 87194 67264 87250 67273
rect 87194 67199 87250 67208
rect 87300 66865 87328 67442
rect 131368 66865 131396 67918
rect 131828 67273 131856 67986
rect 132564 67681 132592 68054
rect 132550 67672 132606 67681
rect 132550 67607 132606 67616
rect 131814 67264 131870 67273
rect 131814 67199 131870 67208
rect 133012 66956 133064 66962
rect 133012 66898 133064 66904
rect 87286 66856 87342 66865
rect 87286 66791 87342 66800
rect 131354 66856 131410 66865
rect 131354 66791 131410 66800
rect 132184 66684 132236 66690
rect 132184 66626 132236 66632
rect 131356 66616 131408 66622
rect 131356 66558 131408 66564
rect 131368 66457 131396 66558
rect 131354 66448 131410 66457
rect 131354 66383 131410 66392
rect 131356 66208 131408 66214
rect 87286 66176 87342 66185
rect 87196 66140 87248 66146
rect 131356 66150 131408 66156
rect 87286 66111 87342 66120
rect 87196 66082 87248 66088
rect 87208 66049 87236 66082
rect 87300 66078 87328 66111
rect 87288 66072 87340 66078
rect 87194 66040 87250 66049
rect 87288 66014 87340 66020
rect 87194 65975 87250 65984
rect 131368 65641 131396 66150
rect 132196 66049 132224 66626
rect 133024 66214 133052 66898
rect 133012 66208 133064 66214
rect 133012 66150 133064 66156
rect 132182 66040 132238 66049
rect 132182 65975 132238 65984
rect 87194 65632 87250 65641
rect 87194 65567 87250 65576
rect 131354 65632 131410 65641
rect 131354 65567 131410 65576
rect 87208 65398 87236 65567
rect 87196 65392 87248 65398
rect 87196 65334 87248 65340
rect 131816 65392 131868 65398
rect 131816 65334 131868 65340
rect 131448 65324 131500 65330
rect 131448 65266 131500 65272
rect 131356 65256 131408 65262
rect 131354 65224 131356 65233
rect 131408 65224 131410 65233
rect 131354 65159 131410 65168
rect 87286 64952 87342 64961
rect 87286 64887 87342 64896
rect 87194 64816 87250 64825
rect 87194 64751 87196 64760
rect 87248 64751 87250 64760
rect 87196 64722 87248 64728
rect 87300 64718 87328 64887
rect 131460 64825 131488 65266
rect 131446 64816 131502 64825
rect 131446 64751 131502 64760
rect 87288 64712 87340 64718
rect 87288 64654 87340 64660
rect 131828 64417 131856 65334
rect 87654 64408 87710 64417
rect 87654 64343 87710 64352
rect 131814 64408 131870 64417
rect 131814 64343 131870 64352
rect 87668 64038 87696 64343
rect 87656 64032 87708 64038
rect 87656 63974 87708 63980
rect 131356 64032 131408 64038
rect 131356 63974 131408 63980
rect 131814 64000 131870 64009
rect 87194 63728 87250 63737
rect 87194 63663 87250 63672
rect 87208 63358 87236 63663
rect 131368 63601 131396 63974
rect 131814 63935 131816 63944
rect 131868 63935 131870 63944
rect 131816 63906 131868 63912
rect 131354 63592 131410 63601
rect 131354 63527 131410 63536
rect 132000 63420 132052 63426
rect 132000 63362 132052 63368
rect 87196 63352 87248 63358
rect 131356 63352 131408 63358
rect 87196 63294 87248 63300
rect 87286 63320 87342 63329
rect 131356 63294 131408 63300
rect 87286 63255 87342 63264
rect 87194 62912 87250 62921
rect 87194 62847 87250 62856
rect 87010 62776 87066 62785
rect 87010 62711 87066 62720
rect 86918 60600 86974 60609
rect 86918 60535 86974 60544
rect 86826 60056 86882 60065
rect 86826 59991 86882 60000
rect 86840 57374 86868 59991
rect 86932 58462 86960 60535
rect 87024 60366 87052 62711
rect 87208 62542 87236 62847
rect 87300 62610 87328 63255
rect 131368 63193 131396 63294
rect 131354 63184 131410 63193
rect 131354 63119 131410 63128
rect 132012 62785 132040 63362
rect 131998 62776 132054 62785
rect 131998 62711 132054 62720
rect 87288 62604 87340 62610
rect 87288 62546 87340 62552
rect 87196 62536 87248 62542
rect 87196 62478 87248 62484
rect 87286 62368 87342 62377
rect 87286 62303 87342 62312
rect 131446 62368 131502 62377
rect 131446 62303 131502 62312
rect 87194 61824 87250 61833
rect 87194 61759 87250 61768
rect 87102 61416 87158 61425
rect 87102 61351 87158 61360
rect 87012 60360 87064 60366
rect 87012 60302 87064 60308
rect 87010 60192 87066 60201
rect 87010 60127 87066 60136
rect 87024 58530 87052 60127
rect 87116 59822 87144 61351
rect 87208 61182 87236 61759
rect 87300 61250 87328 62303
rect 131354 62096 131410 62105
rect 131354 62031 131410 62040
rect 131368 61930 131396 62031
rect 131460 61998 131488 62303
rect 131448 61992 131500 61998
rect 131448 61934 131500 61940
rect 131356 61924 131408 61930
rect 131356 61866 131408 61872
rect 131354 61688 131410 61697
rect 131354 61623 131410 61632
rect 131368 61318 131396 61623
rect 131356 61312 131408 61318
rect 131356 61254 131408 61260
rect 87288 61244 87340 61250
rect 87288 61186 87340 61192
rect 87196 61176 87248 61182
rect 87196 61118 87248 61124
rect 87194 61008 87250 61017
rect 87194 60943 87250 60952
rect 131446 61008 131502 61017
rect 131446 60943 131502 60952
rect 87208 59890 87236 60943
rect 131354 60872 131410 60881
rect 131354 60807 131410 60816
rect 131368 60638 131396 60807
rect 131356 60632 131408 60638
rect 131356 60574 131408 60580
rect 131460 60570 131488 60943
rect 131448 60564 131500 60570
rect 131448 60506 131500 60512
rect 131354 60192 131410 60201
rect 131354 60127 131410 60136
rect 131368 59958 131396 60127
rect 131814 60056 131870 60065
rect 131814 59991 131816 60000
rect 131868 59991 131870 60000
rect 131816 59962 131868 59968
rect 131356 59952 131408 59958
rect 131356 59894 131408 59900
rect 87196 59884 87248 59890
rect 87196 59826 87248 59832
rect 87104 59816 87156 59822
rect 87104 59758 87156 59764
rect 87378 59376 87434 59385
rect 87378 59311 87434 59320
rect 131538 59376 131594 59385
rect 131538 59311 131594 59320
rect 87286 58968 87342 58977
rect 87286 58903 87342 58912
rect 87194 58832 87250 58841
rect 87194 58767 87250 58776
rect 87208 58598 87236 58767
rect 87196 58592 87248 58598
rect 87196 58534 87248 58540
rect 87012 58524 87064 58530
rect 87012 58466 87064 58472
rect 86920 58456 86972 58462
rect 86920 58398 86972 58404
rect 87010 58152 87066 58161
rect 87010 58087 87066 58096
rect 86828 57368 86880 57374
rect 86734 57336 86790 57345
rect 86828 57310 86880 57316
rect 86734 57271 86790 57280
rect 86550 57200 86606 57209
rect 86550 57135 86606 57144
rect 85908 54444 85960 54450
rect 85908 54386 85960 54392
rect 85920 48942 85948 54386
rect 86564 53362 86592 57135
rect 86748 54246 86776 57271
rect 87024 55470 87052 58087
rect 87102 57744 87158 57753
rect 87102 57679 87158 57688
rect 87116 55742 87144 57679
rect 87300 57102 87328 58903
rect 87288 57096 87340 57102
rect 87288 57038 87340 57044
rect 87392 57034 87420 59311
rect 131446 58968 131502 58977
rect 131446 58903 131502 58912
rect 131354 58832 131410 58841
rect 131354 58767 131410 58776
rect 131368 58598 131396 58767
rect 131460 58666 131488 58903
rect 131552 58734 131580 59311
rect 131540 58728 131592 58734
rect 131540 58670 131592 58676
rect 131448 58660 131500 58666
rect 131448 58602 131500 58608
rect 131356 58592 131408 58598
rect 131356 58534 131408 58540
rect 131538 58152 131594 58161
rect 131538 58087 131594 58096
rect 131446 57608 131502 57617
rect 131446 57543 131502 57552
rect 131356 57368 131408 57374
rect 131356 57310 131408 57316
rect 131368 57209 131396 57310
rect 131460 57238 131488 57543
rect 131552 57306 131580 58087
rect 131630 57744 131686 57753
rect 131630 57679 131686 57688
rect 131540 57300 131592 57306
rect 131540 57242 131592 57248
rect 131448 57232 131500 57238
rect 131354 57200 131410 57209
rect 131448 57174 131500 57180
rect 131644 57170 131672 57679
rect 131354 57135 131410 57144
rect 131632 57164 131684 57170
rect 131632 57106 131684 57112
rect 87380 57028 87432 57034
rect 87380 56970 87432 56976
rect 88206 56520 88262 56529
rect 88206 56455 88262 56464
rect 131446 56520 131502 56529
rect 131446 56455 131502 56464
rect 87930 55976 87986 55985
rect 87930 55911 87986 55920
rect 87104 55736 87156 55742
rect 87104 55678 87156 55684
rect 87012 55464 87064 55470
rect 87012 55406 87064 55412
rect 87286 55296 87342 55305
rect 87286 55231 87342 55240
rect 87194 54888 87250 54897
rect 87194 54823 87250 54832
rect 87208 54518 87236 54823
rect 87300 54586 87328 55231
rect 87288 54580 87340 54586
rect 87288 54522 87340 54528
rect 87196 54512 87248 54518
rect 87196 54454 87248 54460
rect 87286 54480 87342 54489
rect 87286 54415 87288 54424
rect 87340 54415 87342 54424
rect 87288 54386 87340 54392
rect 87102 54344 87158 54353
rect 87102 54279 87158 54288
rect 86736 54240 86788 54246
rect 86736 54182 86788 54188
rect 86552 53356 86604 53362
rect 86552 53298 86604 53304
rect 87116 49282 87144 54279
rect 87194 53392 87250 53401
rect 87194 53327 87250 53336
rect 87208 53022 87236 53327
rect 87196 53016 87248 53022
rect 87196 52958 87248 52964
rect 87944 51594 87972 55911
rect 88220 52886 88248 56455
rect 88390 56112 88446 56121
rect 88390 56047 88446 56056
rect 88404 52954 88432 56047
rect 131354 55976 131410 55985
rect 131460 55946 131488 56455
rect 131538 56112 131594 56121
rect 131538 56047 131594 56056
rect 131354 55911 131410 55920
rect 131448 55940 131500 55946
rect 131368 55878 131396 55911
rect 131448 55882 131500 55888
rect 131356 55872 131408 55878
rect 131356 55814 131408 55820
rect 131552 55810 131580 56047
rect 131540 55804 131592 55810
rect 131540 55746 131592 55752
rect 131538 55296 131594 55305
rect 131538 55231 131594 55240
rect 131446 54888 131502 54897
rect 131446 54823 131502 54832
rect 131354 54752 131410 54761
rect 131354 54687 131410 54696
rect 131368 54586 131396 54687
rect 131356 54580 131408 54586
rect 131356 54522 131408 54528
rect 131460 54518 131488 54823
rect 131448 54512 131500 54518
rect 131448 54454 131500 54460
rect 131552 54450 131580 55231
rect 131540 54444 131592 54450
rect 131540 54386 131592 54392
rect 131446 54344 131502 54353
rect 131446 54279 131502 54288
rect 94568 53894 94904 53922
rect 104596 53894 104840 53922
rect 114868 53894 115204 53922
rect 124896 53894 125232 53922
rect 88392 52948 88444 52954
rect 88392 52890 88444 52896
rect 88208 52880 88260 52886
rect 88208 52822 88260 52828
rect 87932 51588 87984 51594
rect 87932 51530 87984 51536
rect 94568 50710 94596 53894
rect 104596 53809 104624 53894
rect 104582 53800 104638 53809
rect 104582 53735 104638 53744
rect 115176 50914 115204 53894
rect 125204 50982 125232 53894
rect 131354 53528 131410 53537
rect 131354 53463 131410 53472
rect 131368 53022 131396 53463
rect 131460 53090 131488 54279
rect 131448 53084 131500 53090
rect 131448 53026 131500 53032
rect 131356 53016 131408 53022
rect 131356 52958 131408 52964
rect 125192 50976 125244 50982
rect 125192 50918 125244 50924
rect 127032 50976 127084 50982
rect 127032 50918 127084 50924
rect 115164 50908 115216 50914
rect 115164 50850 115216 50856
rect 94004 50704 94056 50710
rect 94004 50646 94056 50652
rect 94556 50704 94608 50710
rect 94556 50646 94608 50652
rect 87104 49276 87156 49282
rect 87104 49218 87156 49224
rect 85908 48936 85960 48942
rect 85908 48878 85960 48884
rect 94016 37790 94044 50646
rect 99524 47508 99576 47514
rect 99524 47450 99576 47456
rect 99536 37790 99564 47450
rect 93084 37784 93136 37790
rect 93084 37726 93136 37732
rect 94004 37784 94056 37790
rect 94004 37726 94056 37732
rect 98788 37784 98840 37790
rect 98788 37726 98840 37732
rect 99524 37784 99576 37790
rect 99524 37726 99576 37732
rect 93096 34746 93124 37726
rect 98800 34746 98828 37726
rect 103848 37240 103900 37246
rect 103848 37182 103900 37188
rect 92788 34718 93124 34746
rect 98492 34718 98828 34746
rect 103860 34746 103888 37182
rect 120960 37172 121012 37178
rect 120960 37114 121012 37120
rect 109552 37104 109604 37110
rect 109552 37046 109604 37052
rect 115808 37104 115860 37110
rect 115808 37046 115860 37052
rect 109564 34746 109592 37046
rect 115820 34746 115848 37046
rect 103860 34718 104196 34746
rect 109564 34718 109900 34746
rect 115604 34718 115848 34746
rect 120972 34746 121000 37114
rect 127044 34746 127072 50918
rect 128596 50908 128648 50914
rect 128596 50850 128648 50856
rect 120972 34718 121308 34746
rect 127012 34718 127072 34746
rect 128608 28082 128636 50850
rect 128608 28066 128912 28082
rect 128608 28060 128924 28066
rect 128608 28054 128872 28060
rect 128872 28002 128924 28008
rect 129516 28060 129568 28066
rect 129516 28002 129568 28008
rect 129528 27561 129556 28002
rect 129514 27552 129570 27561
rect 129514 27487 129570 27496
rect 88482 26872 88538 26881
rect 88482 26807 88538 26816
rect 85080 25408 85132 25414
rect 85080 25350 85132 25356
rect 76524 20920 76576 20926
rect 76524 20862 76576 20868
rect 38160 12488 38212 12494
rect 38160 12430 38212 12436
rect 28224 12420 28276 12426
rect 28224 12362 28276 12368
rect 28236 9304 28264 12362
rect 88496 12358 88524 26807
rect 109564 18942 109900 18970
rect 109564 17118 109592 18942
rect 109552 17112 109604 17118
rect 109552 17054 109604 17060
rect 133392 12426 133420 81858
rect 134772 80562 134800 83814
rect 134760 80556 134812 80562
rect 134760 80498 134812 80504
rect 134772 50982 134800 80498
rect 134864 78561 134892 83898
rect 137532 79134 137560 109631
rect 137716 102225 137744 115110
rect 137808 103993 137836 117830
rect 137900 108209 137928 124766
rect 137992 124257 138020 139318
rect 138992 139308 139044 139314
rect 138992 139250 139044 139256
rect 138898 130912 138954 130921
rect 138898 130847 138954 130856
rect 138162 125064 138218 125073
rect 138162 124999 138218 125008
rect 138176 124898 138204 124999
rect 138164 124892 138216 124898
rect 138164 124834 138216 124840
rect 137978 124248 138034 124257
rect 137978 124183 138034 124192
rect 138164 122104 138216 122110
rect 138162 122072 138164 122081
rect 138216 122072 138218 122081
rect 137980 122036 138032 122042
rect 138162 122007 138218 122016
rect 137980 121978 138032 121984
rect 137886 108200 137942 108209
rect 137886 108135 137942 108144
rect 137992 106713 138020 121978
rect 138072 119316 138124 119322
rect 138072 119258 138124 119264
rect 137978 106704 138034 106713
rect 137978 106639 138034 106648
rect 138084 105353 138112 119258
rect 138162 118400 138218 118409
rect 138162 118335 138218 118344
rect 138176 117962 138204 118335
rect 138164 117956 138216 117962
rect 138164 117898 138216 117904
rect 138162 112688 138218 112697
rect 138162 112623 138218 112632
rect 138176 112590 138204 112623
rect 138164 112584 138216 112590
rect 138164 112526 138216 112532
rect 138164 111020 138216 111026
rect 138164 110962 138216 110968
rect 138070 105344 138126 105353
rect 138070 105279 138126 105288
rect 137794 103984 137850 103993
rect 137794 103919 137850 103928
rect 137702 102216 137758 102225
rect 137702 102151 137758 102160
rect 138176 99233 138204 110962
rect 138162 99224 138218 99233
rect 138162 99159 138218 99168
rect 138164 95788 138216 95794
rect 138164 95730 138216 95736
rect 138176 95697 138204 95730
rect 138162 95688 138218 95697
rect 138162 95623 138218 95632
rect 138162 93920 138218 93929
rect 138162 93855 138164 93864
rect 138216 93855 138218 93864
rect 138164 93826 138216 93832
rect 137796 92728 137848 92734
rect 137794 92696 137796 92705
rect 137848 92696 137850 92705
rect 137794 92631 137850 92640
rect 137612 91640 137664 91646
rect 137612 91582 137664 91588
rect 137624 91481 137652 91582
rect 137610 91472 137666 91481
rect 137610 91407 137666 91416
rect 138164 89192 138216 89198
rect 138162 89160 138164 89169
rect 138216 89160 138218 89169
rect 138162 89095 138218 89104
rect 137612 88852 137664 88858
rect 137612 88794 137664 88800
rect 137624 88217 137652 88794
rect 137610 88208 137666 88217
rect 137610 88143 137666 88152
rect 137520 79128 137572 79134
rect 137520 79070 137572 79076
rect 134850 78552 134906 78561
rect 138912 78522 138940 130847
rect 139004 130270 139032 139250
rect 142776 138634 142804 141886
rect 143604 138702 143632 141886
rect 144156 138770 144184 141886
rect 144708 138838 144736 141886
rect 145168 139382 145196 141886
rect 145156 139376 145208 139382
rect 145156 139318 145208 139324
rect 145720 139246 145748 141886
rect 146272 139314 146300 141886
rect 146260 139308 146312 139314
rect 146260 139250 146312 139256
rect 145708 139240 145760 139246
rect 145708 139182 145760 139188
rect 144696 138832 144748 138838
rect 144696 138774 144748 138780
rect 144144 138764 144196 138770
rect 144144 138706 144196 138712
rect 143592 138696 143644 138702
rect 143592 138638 143644 138644
rect 142764 138628 142816 138634
rect 142764 138570 142816 138576
rect 146824 132990 146852 141886
rect 147284 138702 147312 141886
rect 147836 138770 147864 141886
rect 147824 138764 147876 138770
rect 147824 138706 147876 138712
rect 147272 138696 147324 138702
rect 147272 138638 147324 138644
rect 148388 138634 148416 141886
rect 148376 138628 148428 138634
rect 148376 138570 148428 138576
rect 146812 132984 146864 132990
rect 146812 132926 146864 132932
rect 148940 131698 148968 141886
rect 149400 139790 149428 141886
rect 149388 139784 149440 139790
rect 149388 139726 149440 139732
rect 149112 139512 149164 139518
rect 149112 139454 149164 139460
rect 149020 138628 149072 138634
rect 149020 138570 149072 138576
rect 148928 131692 148980 131698
rect 148928 131634 148980 131640
rect 149032 131018 149060 138570
rect 149020 131012 149072 131018
rect 149020 130954 149072 130960
rect 138992 130264 139044 130270
rect 138992 130206 139044 130212
rect 149124 128708 149152 139454
rect 149952 139110 149980 141886
rect 150504 139722 150532 141886
rect 150492 139716 150544 139722
rect 150492 139658 150544 139664
rect 149940 139104 149992 139110
rect 149940 139046 149992 139052
rect 151056 138906 151084 141886
rect 151044 138900 151096 138906
rect 151044 138842 151096 138848
rect 151516 138838 151544 141886
rect 151504 138832 151556 138838
rect 151504 138774 151556 138780
rect 152068 138634 152096 141886
rect 152620 139194 152648 141886
rect 152620 139166 153016 139194
rect 152700 139036 152752 139042
rect 152700 138978 152752 138984
rect 152056 138628 152108 138634
rect 152056 138570 152108 138576
rect 149204 131692 149256 131698
rect 149204 131634 149256 131640
rect 149216 131154 149244 131634
rect 150216 131624 150268 131630
rect 150216 131566 150268 131572
rect 149848 131556 149900 131562
rect 149848 131498 149900 131504
rect 149480 131216 149532 131222
rect 149480 131158 149532 131164
rect 149204 131148 149256 131154
rect 149204 131090 149256 131096
rect 149492 128708 149520 131158
rect 149860 128708 149888 131498
rect 150228 128708 150256 131566
rect 152712 131426 152740 138978
rect 152884 138560 152936 138566
rect 152884 138502 152936 138508
rect 151044 131420 151096 131426
rect 151044 131362 151096 131368
rect 152700 131420 152752 131426
rect 152700 131362 152752 131368
rect 150584 130604 150636 130610
rect 150584 130546 150636 130552
rect 150596 128708 150624 130546
rect 151056 128708 151084 131362
rect 152608 131216 152660 131222
rect 152608 131158 152660 131164
rect 151412 130876 151464 130882
rect 151412 130818 151464 130824
rect 151424 128708 151452 130818
rect 151780 130808 151832 130814
rect 151780 130750 151832 130756
rect 151792 128708 151820 130750
rect 152148 130332 152200 130338
rect 152148 130274 152200 130280
rect 152160 128708 152188 130274
rect 152620 128708 152648 131158
rect 152896 128722 152924 138502
rect 152988 131426 153016 139166
rect 152976 131420 153028 131426
rect 152976 131362 153028 131368
rect 153080 130746 153108 141886
rect 153252 139444 153304 139450
rect 153252 139386 153304 139392
rect 153160 138628 153212 138634
rect 153160 138570 153212 138576
rect 153172 131494 153200 138570
rect 153160 131488 153212 131494
rect 153160 131430 153212 131436
rect 153068 130740 153120 130746
rect 153068 130682 153120 130688
rect 153264 128722 153292 139386
rect 153632 138974 153660 141886
rect 154184 139246 154212 141886
rect 154172 139240 154224 139246
rect 154172 139182 154224 139188
rect 154736 139110 154764 141886
rect 155000 139580 155052 139586
rect 155000 139522 155052 139528
rect 154724 139104 154776 139110
rect 154724 139046 154776 139052
rect 153620 138968 153672 138974
rect 153620 138910 153672 138916
rect 154724 138968 154776 138974
rect 154724 138910 154776 138916
rect 154264 138764 154316 138770
rect 154264 138706 154316 138712
rect 154080 138696 154132 138702
rect 154080 138638 154132 138644
rect 153712 131080 153764 131086
rect 153712 131022 153764 131028
rect 152896 128694 153002 128722
rect 153264 128694 153370 128722
rect 153724 128708 153752 131022
rect 154092 130474 154120 138638
rect 154276 130610 154304 138706
rect 154736 131358 154764 138910
rect 155012 135386 155040 139522
rect 155196 139382 155224 141886
rect 155276 139716 155328 139722
rect 155276 139658 155328 139664
rect 155184 139376 155236 139382
rect 155184 139318 155236 139324
rect 155012 135358 155224 135386
rect 154724 131352 154776 131358
rect 154724 131294 154776 131300
rect 154264 130604 154316 130610
rect 154264 130546 154316 130552
rect 154172 130536 154224 130542
rect 154172 130478 154224 130484
rect 154080 130468 154132 130474
rect 154080 130410 154132 130416
rect 154184 128708 154212 130478
rect 154540 130400 154592 130406
rect 154540 130342 154592 130348
rect 154552 128708 154580 130342
rect 154908 130332 154960 130338
rect 154908 130274 154960 130280
rect 154920 128708 154948 130274
rect 155196 130082 155224 135358
rect 155288 130338 155316 139658
rect 155748 139466 155776 141886
rect 155748 139438 156144 139466
rect 155920 139376 155972 139382
rect 155920 139318 155972 139324
rect 155552 139240 155604 139246
rect 155552 139182 155604 139188
rect 155828 139240 155880 139246
rect 155828 139182 155880 139188
rect 155368 139172 155420 139178
rect 155368 139114 155420 139120
rect 155380 131630 155408 139114
rect 155460 139104 155512 139110
rect 155460 139046 155512 139052
rect 155472 131630 155500 139046
rect 155368 131624 155420 131630
rect 155368 131566 155420 131572
rect 155460 131624 155512 131630
rect 155460 131566 155512 131572
rect 155564 130814 155592 139182
rect 155736 139104 155788 139110
rect 155736 139046 155788 139052
rect 155644 138764 155696 138770
rect 155644 138706 155696 138712
rect 155656 131562 155684 138706
rect 155644 131556 155696 131562
rect 155644 131498 155696 131504
rect 155552 130808 155604 130814
rect 155552 130750 155604 130756
rect 155748 130678 155776 139046
rect 155736 130672 155788 130678
rect 155736 130614 155788 130620
rect 155276 130332 155328 130338
rect 155276 130274 155328 130280
rect 155736 130332 155788 130338
rect 155736 130274 155788 130280
rect 155196 130054 155316 130082
rect 155288 128708 155316 130054
rect 155748 128708 155776 130274
rect 155840 128722 155868 139182
rect 155932 130746 155960 139318
rect 156012 139036 156064 139042
rect 156012 138978 156064 138984
rect 155920 130740 155972 130746
rect 155920 130682 155972 130688
rect 156024 130338 156052 138978
rect 156116 130678 156144 139438
rect 156300 138702 156328 141886
rect 156748 139036 156800 139042
rect 156748 138978 156800 138984
rect 156288 138696 156340 138702
rect 156288 138638 156340 138644
rect 156760 135386 156788 138978
rect 156852 138634 156880 141886
rect 156932 138968 156984 138974
rect 156932 138910 156984 138916
rect 156840 138628 156892 138634
rect 156840 138570 156892 138576
rect 156760 135358 156880 135386
rect 156472 131216 156524 131222
rect 156472 131158 156524 131164
rect 156104 130672 156156 130678
rect 156104 130614 156156 130620
rect 156012 130332 156064 130338
rect 156012 130274 156064 130280
rect 155840 128694 156130 128722
rect 156484 128708 156512 131158
rect 156564 130468 156616 130474
rect 156564 130410 156616 130416
rect 156576 128722 156604 130410
rect 156852 130406 156880 135358
rect 156944 130542 156972 138910
rect 157312 138786 157340 141886
rect 157818 141642 157846 141900
rect 158370 141778 158398 141900
rect 158936 141886 158996 141914
rect 159396 141886 159456 141914
rect 159948 141886 160008 141914
rect 160500 141886 160560 141914
rect 161052 141886 161112 141914
rect 161512 141886 161572 141914
rect 162064 141886 162124 141914
rect 162616 141886 162676 141914
rect 163076 141886 163136 141914
rect 163628 141886 163688 141914
rect 164180 141886 164240 141914
rect 164732 141886 164792 141914
rect 165192 141886 165252 141914
rect 165744 141886 165804 141914
rect 166296 141886 166356 141914
rect 166848 141886 166908 141914
rect 167308 141886 167368 141914
rect 167860 141886 167920 141914
rect 168412 141886 168472 141914
rect 168964 141886 169024 141914
rect 169424 141886 169484 141914
rect 169976 141886 170036 141914
rect 170528 141886 170588 141914
rect 157588 141614 157846 141642
rect 157956 141750 158398 141778
rect 157588 139518 157616 141614
rect 157956 141506 157984 141750
rect 157680 141478 157984 141506
rect 157576 139512 157628 139518
rect 157576 139454 157628 139460
rect 157576 138900 157628 138906
rect 157576 138842 157628 138848
rect 157312 138758 157432 138786
rect 157300 138628 157352 138634
rect 157300 138570 157352 138576
rect 157312 131630 157340 138570
rect 157300 131624 157352 131630
rect 157300 131566 157352 131572
rect 157404 131562 157432 138758
rect 157588 138702 157616 138842
rect 157484 138696 157536 138702
rect 157484 138638 157536 138644
rect 157576 138696 157628 138702
rect 157576 138638 157628 138644
rect 157392 131556 157444 131562
rect 157392 131498 157444 131504
rect 157496 131426 157524 138638
rect 157484 131420 157536 131426
rect 157484 131362 157536 131368
rect 157680 131290 157708 141478
rect 157852 139784 157904 139790
rect 157852 139726 157904 139732
rect 157864 131306 157892 139726
rect 158864 139308 158916 139314
rect 158864 139250 158916 139256
rect 158404 138900 158456 138906
rect 158404 138842 158456 138848
rect 158220 138832 158272 138838
rect 158220 138774 158272 138780
rect 158312 138832 158364 138838
rect 158312 138774 158364 138780
rect 157668 131284 157720 131290
rect 157864 131278 158168 131306
rect 157668 131226 157720 131232
rect 158036 131148 158088 131154
rect 158036 131090 158088 131096
rect 157668 131012 157720 131018
rect 157668 130954 157720 130960
rect 157300 130604 157352 130610
rect 157300 130546 157352 130552
rect 156932 130536 156984 130542
rect 156932 130478 156984 130484
rect 156840 130400 156892 130406
rect 156840 130342 156892 130348
rect 156576 128694 156866 128722
rect 157312 128708 157340 130546
rect 157680 128708 157708 130954
rect 158048 128708 158076 131090
rect 158140 128858 158168 131278
rect 158232 130406 158260 138774
rect 158324 130950 158352 138774
rect 158312 130944 158364 130950
rect 158312 130886 158364 130892
rect 158416 130882 158444 138842
rect 158496 138696 158548 138702
rect 158496 138638 158548 138644
rect 158404 130876 158456 130882
rect 158404 130818 158456 130824
rect 158220 130400 158272 130406
rect 158220 130342 158272 130348
rect 158508 130338 158536 138638
rect 158496 130332 158548 130338
rect 158496 130274 158548 130280
rect 158140 128830 158260 128858
rect 158232 128722 158260 128830
rect 158232 128694 158430 128722
rect 158876 128708 158904 139250
rect 158968 138770 158996 141886
rect 159232 139648 159284 139654
rect 159232 139590 159284 139596
rect 158956 138764 159008 138770
rect 158956 138706 159008 138712
rect 159244 128708 159272 139590
rect 159428 139178 159456 141886
rect 159416 139172 159468 139178
rect 159416 139114 159468 139120
rect 159980 139110 160008 141886
rect 160532 139518 160560 141886
rect 160520 139512 160572 139518
rect 160520 139454 160572 139460
rect 159968 139104 160020 139110
rect 159968 139046 160020 139052
rect 161084 138906 161112 141886
rect 161072 138900 161124 138906
rect 161072 138842 161124 138848
rect 161544 138838 161572 141886
rect 161532 138832 161584 138838
rect 161532 138774 161584 138780
rect 161072 138764 161124 138770
rect 161072 138706 161124 138712
rect 160980 138696 161032 138702
rect 160980 138638 161032 138644
rect 159600 135840 159652 135846
rect 159600 135782 159652 135788
rect 159612 131154 159640 135782
rect 160428 131488 160480 131494
rect 160428 131430 160480 131436
rect 159600 131148 159652 131154
rect 159600 131090 159652 131096
rect 159968 130400 160020 130406
rect 159968 130342 160020 130348
rect 159600 130332 159652 130338
rect 159600 130274 159652 130280
rect 159612 128708 159640 130274
rect 159980 128708 160008 130342
rect 160440 128708 160468 131430
rect 160992 131290 161020 138638
rect 160980 131284 161032 131290
rect 160980 131226 161032 131232
rect 161084 131018 161112 138706
rect 162096 138634 162124 141886
rect 162648 138702 162676 141886
rect 163108 139314 163136 141886
rect 163660 139382 163688 141886
rect 163648 139376 163700 139382
rect 163648 139318 163700 139324
rect 163096 139308 163148 139314
rect 163096 139250 163148 139256
rect 164212 138838 164240 141886
rect 164764 138974 164792 141886
rect 165224 139042 165252 141886
rect 165776 139722 165804 141886
rect 165764 139716 165816 139722
rect 165764 139658 165816 139664
rect 166328 139586 166356 141886
rect 166316 139580 166368 139586
rect 166316 139522 166368 139528
rect 166880 139450 166908 141886
rect 166868 139444 166920 139450
rect 166868 139386 166920 139392
rect 167340 139246 167368 141886
rect 167328 139240 167380 139246
rect 167328 139182 167380 139188
rect 165212 139036 165264 139042
rect 165212 138978 165264 138984
rect 164752 138968 164804 138974
rect 164752 138910 164804 138916
rect 164200 138832 164252 138838
rect 164200 138774 164252 138780
rect 167892 138770 167920 141886
rect 168444 141694 168472 141886
rect 168432 141688 168484 141694
rect 168432 141630 168484 141636
rect 168996 139926 169024 141886
rect 168984 139920 169036 139926
rect 168984 139862 169036 139868
rect 169456 139858 169484 141886
rect 170008 141762 170036 141886
rect 169996 141756 170048 141762
rect 169996 141698 170048 141704
rect 170560 139897 170588 141886
rect 170652 141762 170680 175086
rect 171376 174464 171428 174470
rect 171376 174406 171428 174412
rect 170732 170248 170784 170254
rect 170732 170190 170784 170196
rect 170744 169273 170772 170190
rect 171388 169545 171416 174406
rect 171374 169536 171430 169545
rect 171374 169471 171430 169480
rect 170730 169264 170786 169273
rect 170730 169199 170786 169208
rect 170732 166236 170784 166242
rect 170732 166178 170784 166184
rect 170640 141756 170692 141762
rect 170640 141698 170692 141704
rect 170744 141694 170772 166178
rect 171388 144754 171416 169471
rect 173306 168448 173362 168457
rect 173306 168383 173362 168392
rect 173320 167738 173348 168383
rect 173308 167732 173360 167738
rect 173308 167674 173360 167680
rect 173306 167360 173362 167369
rect 173306 167295 173362 167304
rect 173122 166816 173178 166825
rect 173122 166751 173178 166760
rect 173136 166650 173164 166751
rect 173124 166644 173176 166650
rect 173124 166586 173176 166592
rect 173122 166272 173178 166281
rect 173122 166207 173178 166216
rect 173030 164504 173086 164513
rect 173030 164439 173086 164448
rect 172938 162872 172994 162881
rect 172938 162807 172940 162816
rect 172992 162807 172994 162816
rect 172940 162778 172992 162784
rect 172938 162328 172994 162337
rect 172938 162263 172940 162272
rect 172992 162263 172994 162272
rect 172940 162234 172992 162240
rect 172754 160560 172810 160569
rect 172754 160495 172810 160504
rect 172768 159646 172796 160495
rect 173044 160394 173072 164439
rect 173136 160802 173164 166207
rect 173214 163960 173270 163969
rect 173214 163895 173270 163904
rect 173124 160796 173176 160802
rect 173124 160738 173176 160744
rect 173032 160388 173084 160394
rect 173032 160330 173084 160336
rect 173228 160274 173256 163895
rect 172860 160246 173256 160274
rect 172756 159640 172808 159646
rect 172756 159582 172808 159588
rect 172860 153526 172888 160246
rect 173320 160138 173348 167295
rect 173044 160110 173348 160138
rect 172938 157840 172994 157849
rect 172938 157775 172994 157784
rect 172952 157130 172980 157775
rect 172940 157124 172992 157130
rect 172940 157066 172992 157072
rect 172940 155084 172992 155090
rect 172940 155026 172992 155032
rect 172952 153905 172980 155026
rect 173044 154954 173072 160110
rect 173306 160016 173362 160025
rect 173306 159951 173308 159960
rect 173360 159951 173362 159960
rect 173308 159922 173360 159928
rect 173216 159572 173268 159578
rect 173216 159514 173268 159520
rect 173122 158928 173178 158937
rect 173122 158863 173178 158872
rect 173136 157946 173164 158863
rect 173228 158098 173256 159514
rect 173306 158384 173362 158393
rect 173306 158319 173362 158328
rect 173320 158218 173348 158319
rect 173308 158212 173360 158218
rect 173308 158154 173360 158160
rect 173228 158070 173348 158098
rect 173124 157940 173176 157946
rect 173124 157882 173176 157888
rect 173124 157668 173176 157674
rect 173124 157610 173176 157616
rect 173136 156761 173164 157610
rect 173216 157600 173268 157606
rect 173216 157542 173268 157548
rect 173228 157305 173256 157542
rect 173214 157296 173270 157305
rect 173214 157231 173270 157240
rect 173216 157192 173268 157198
rect 173216 157134 173268 157140
rect 173122 156752 173178 156761
rect 173122 156687 173178 156696
rect 173032 154948 173084 154954
rect 173032 154890 173084 154896
rect 173124 154472 173176 154478
rect 173122 154440 173124 154449
rect 173176 154440 173178 154449
rect 173122 154375 173178 154384
rect 172938 153896 172994 153905
rect 172938 153831 172994 153840
rect 173228 153662 173256 157134
rect 173216 153656 173268 153662
rect 173216 153598 173268 153604
rect 173320 153594 173348 158070
rect 173308 153588 173360 153594
rect 173308 153530 173360 153536
rect 172848 153520 172900 153526
rect 172848 153462 172900 153468
rect 173308 153452 173360 153458
rect 173308 153394 173360 153400
rect 173320 152817 173348 153394
rect 173306 152808 173362 152817
rect 173306 152743 173362 152752
rect 173308 151888 173360 151894
rect 173308 151830 173360 151836
rect 173320 151729 173348 151830
rect 173306 151720 173362 151729
rect 173306 151655 173362 151664
rect 172940 150868 172992 150874
rect 172940 150810 172992 150816
rect 172952 149961 172980 150810
rect 172938 149952 172994 149961
rect 172938 149887 172994 149896
rect 173308 149508 173360 149514
rect 173308 149450 173360 149456
rect 172756 147876 172808 147882
rect 172756 147818 172808 147824
rect 172768 147241 172796 147818
rect 172754 147232 172810 147241
rect 172754 147167 172810 147176
rect 172756 146380 172808 146386
rect 172756 146322 172808 146328
rect 172768 146017 172796 146322
rect 172754 146008 172810 146017
rect 172754 145943 172810 145952
rect 170824 144748 170876 144754
rect 170824 144690 170876 144696
rect 171376 144748 171428 144754
rect 171376 144690 171428 144696
rect 170732 141688 170784 141694
rect 170732 141630 170784 141636
rect 170546 139888 170602 139897
rect 169444 139852 169496 139858
rect 170546 139823 170602 139832
rect 169444 139794 169496 139800
rect 163740 138764 163792 138770
rect 163740 138706 163792 138712
rect 167880 138764 167932 138770
rect 167880 138706 167932 138712
rect 162636 138696 162688 138702
rect 162636 138638 162688 138644
rect 161164 138628 161216 138634
rect 161164 138570 161216 138576
rect 162084 138628 162136 138634
rect 162084 138570 162136 138576
rect 161072 131012 161124 131018
rect 161072 130954 161124 130960
rect 160796 130808 160848 130814
rect 160796 130750 160848 130756
rect 160808 128708 160836 130750
rect 161176 130678 161204 138570
rect 163556 131420 163608 131426
rect 163556 131362 163608 131368
rect 161532 131352 161584 131358
rect 161532 131294 161584 131300
rect 161164 130672 161216 130678
rect 161164 130614 161216 130620
rect 161164 130468 161216 130474
rect 161164 130410 161216 130416
rect 161176 128708 161204 130410
rect 161544 128708 161572 131294
rect 162360 131080 162412 131086
rect 162360 131022 162412 131028
rect 161992 130536 162044 130542
rect 161992 130478 162044 130484
rect 162004 128708 162032 130478
rect 162372 128708 162400 131022
rect 162728 130672 162780 130678
rect 162728 130614 162780 130620
rect 162740 128708 162768 130614
rect 163096 130604 163148 130610
rect 163096 130546 163148 130552
rect 163108 128708 163136 130546
rect 163568 128708 163596 131362
rect 163752 131222 163780 138706
rect 170836 138634 170864 144690
rect 173320 142753 173348 149450
rect 173306 142744 173362 142753
rect 173306 142679 173362 142688
rect 173412 142209 173440 175630
rect 173860 175620 173912 175626
rect 173860 175562 173912 175568
rect 173676 175552 173728 175558
rect 173676 175494 173728 175500
rect 173492 175484 173544 175490
rect 173492 175426 173544 175432
rect 173504 143841 173532 175426
rect 173584 175348 173636 175354
rect 173584 175290 173636 175296
rect 173596 144929 173624 175290
rect 173688 145722 173716 175494
rect 173768 175416 173820 175422
rect 173768 175358 173820 175364
rect 173780 146946 173808 175358
rect 173872 149514 173900 175562
rect 176160 175280 176212 175286
rect 176160 175222 176212 175228
rect 174780 175212 174832 175218
rect 174780 175154 174832 175160
rect 174042 167904 174098 167913
rect 174042 167839 174044 167848
rect 174096 167839 174098 167848
rect 174044 167810 174096 167816
rect 174042 165728 174098 165737
rect 174042 165663 174098 165672
rect 173950 165048 174006 165057
rect 173950 164983 174006 164992
rect 173964 163266 173992 164983
rect 174056 164814 174084 165663
rect 174044 164808 174096 164814
rect 174044 164750 174096 164756
rect 174044 163448 174096 163454
rect 174042 163416 174044 163425
rect 174096 163416 174098 163425
rect 174042 163351 174098 163360
rect 173964 163238 174084 163266
rect 173950 161784 174006 161793
rect 173950 161719 174006 161728
rect 173964 160938 173992 161719
rect 174056 161362 174084 163238
rect 174056 161334 174176 161362
rect 174042 161240 174098 161249
rect 174042 161175 174098 161184
rect 173952 160932 174004 160938
rect 173952 160874 174004 160880
rect 174056 160870 174084 161175
rect 174044 160864 174096 160870
rect 174044 160806 174096 160812
rect 173952 160796 174004 160802
rect 173952 160738 174004 160744
rect 173964 156466 173992 160738
rect 174148 160682 174176 161334
rect 174056 160654 174176 160682
rect 174056 159578 174084 160654
rect 174044 159572 174096 159578
rect 174044 159514 174096 159520
rect 174042 159472 174098 159481
rect 174042 159407 174044 159416
rect 174096 159407 174098 159416
rect 174044 159378 174096 159384
rect 173964 156438 174176 156466
rect 174044 156376 174096 156382
rect 174044 156318 174096 156324
rect 173952 156240 174004 156246
rect 174056 156217 174084 156318
rect 173952 156182 174004 156188
rect 174042 156208 174098 156217
rect 173964 155537 173992 156182
rect 174042 156143 174098 156152
rect 174148 156058 174176 156438
rect 174056 156030 174176 156058
rect 173950 155528 174006 155537
rect 173950 155463 174006 155472
rect 173952 155016 174004 155022
rect 173950 154984 173952 154993
rect 174004 154984 174006 154993
rect 173950 154919 174006 154928
rect 174056 154886 174084 156030
rect 174044 154880 174096 154886
rect 174044 154822 174096 154828
rect 174044 153384 174096 153390
rect 174042 153352 174044 153361
rect 174096 153352 174098 153361
rect 174042 153287 174098 153296
rect 174044 152296 174096 152302
rect 174042 152264 174044 152273
rect 174096 152264 174098 152273
rect 174042 152199 174098 152208
rect 173952 151480 174004 151486
rect 173952 151422 174004 151428
rect 173964 151049 173992 151422
rect 173950 151040 174006 151049
rect 173950 150975 174006 150984
rect 174044 150800 174096 150806
rect 174044 150742 174096 150748
rect 174056 150505 174084 150742
rect 174042 150496 174098 150505
rect 174042 150431 174098 150440
rect 173860 149508 173912 149514
rect 173860 149450 173912 149456
rect 174044 149440 174096 149446
rect 174042 149408 174044 149417
rect 174096 149408 174098 149417
rect 173860 149372 173912 149378
rect 174042 149343 174098 149352
rect 173860 149314 173912 149320
rect 173872 148329 173900 149314
rect 174044 148896 174096 148902
rect 174042 148864 174044 148873
rect 174096 148864 174098 148873
rect 174042 148799 174098 148808
rect 173858 148320 173914 148329
rect 173858 148255 173914 148264
rect 174044 147808 174096 147814
rect 174042 147776 174044 147785
rect 174096 147776 174098 147785
rect 174042 147711 174098 147720
rect 173780 146918 173992 146946
rect 173688 145694 173900 145722
rect 173674 145464 173730 145473
rect 173674 145399 173676 145408
rect 173728 145399 173730 145408
rect 173676 145370 173728 145376
rect 173582 144920 173638 144929
rect 173582 144855 173638 144864
rect 173490 143832 173546 143841
rect 173490 143767 173546 143776
rect 173872 143297 173900 145694
rect 173964 144385 173992 146918
rect 174044 146720 174096 146726
rect 174044 146662 174096 146668
rect 174056 146561 174084 146662
rect 174042 146552 174098 146561
rect 174042 146487 174098 146496
rect 174792 146386 174820 175154
rect 174872 160796 174924 160802
rect 174872 160738 174924 160744
rect 174884 154478 174912 160738
rect 175424 160660 175476 160666
rect 175424 160602 175476 160608
rect 175436 155090 175464 160602
rect 176068 159504 176120 159510
rect 176068 159446 176120 159452
rect 175424 155084 175476 155090
rect 175424 155026 175476 155032
rect 174872 154472 174924 154478
rect 174872 154414 174924 154420
rect 176080 153458 176108 159446
rect 176068 153452 176120 153458
rect 176068 153394 176120 153400
rect 174780 146380 174832 146386
rect 174780 146322 174832 146328
rect 176172 145434 176200 175222
rect 177540 167868 177592 167874
rect 177540 167810 177592 167816
rect 176896 159368 176948 159374
rect 176896 159310 176948 159316
rect 176344 158212 176396 158218
rect 176344 158154 176396 158160
rect 176252 157940 176304 157946
rect 176252 157882 176304 157888
rect 176264 149582 176292 157882
rect 176252 149576 176304 149582
rect 176252 149518 176304 149524
rect 176356 149514 176384 158154
rect 176908 152302 176936 159310
rect 176988 159300 177040 159306
rect 176988 159242 177040 159248
rect 176896 152296 176948 152302
rect 176896 152238 176948 152244
rect 177000 151894 177028 159242
rect 177552 156450 177580 167810
rect 180300 167732 180352 167738
rect 180300 167674 180352 167680
rect 178920 166644 178972 166650
rect 178920 166586 178972 166592
rect 177908 163584 177960 163590
rect 177908 163526 177960 163532
rect 177920 157606 177948 163526
rect 178276 157940 178328 157946
rect 178276 157882 178328 157888
rect 177908 157600 177960 157606
rect 177908 157542 177960 157548
rect 177632 157124 177684 157130
rect 177632 157066 177684 157072
rect 177540 156444 177592 156450
rect 177540 156386 177592 156392
rect 176988 151888 177040 151894
rect 176988 151830 177040 151836
rect 176344 149508 176396 149514
rect 176344 149450 176396 149456
rect 177644 148086 177672 157066
rect 178288 151486 178316 157882
rect 178932 155090 178960 166586
rect 179104 162836 179156 162842
rect 179104 162778 179156 162784
rect 179012 162292 179064 162298
rect 179012 162234 179064 162240
rect 178920 155084 178972 155090
rect 178920 155026 178972 155032
rect 179024 152302 179052 162234
rect 179116 152370 179144 162778
rect 179656 162088 179708 162094
rect 179656 162030 179708 162036
rect 179668 155022 179696 162030
rect 180116 160728 180168 160734
rect 180116 160670 180168 160676
rect 179656 155016 179708 155022
rect 179656 154958 179708 154964
rect 180128 153390 180156 160670
rect 180208 156512 180260 156518
rect 180208 156454 180260 156460
rect 180116 153384 180168 153390
rect 180116 153326 180168 153332
rect 179104 152364 179156 152370
rect 179104 152306 179156 152312
rect 179012 152296 179064 152302
rect 179012 152238 179064 152244
rect 178276 151480 178328 151486
rect 178276 151422 178328 151428
rect 180220 149378 180248 156454
rect 180312 155673 180340 167674
rect 180864 166854 180892 177940
rect 182244 166922 182272 177940
rect 183624 174470 183652 177940
rect 183612 174464 183664 174470
rect 183612 174406 183664 174412
rect 184912 174146 184940 177940
rect 186292 174810 186320 177940
rect 186280 174804 186332 174810
rect 186280 174746 186332 174752
rect 187672 174674 187700 177940
rect 188960 175830 188988 177940
rect 188948 175824 189000 175830
rect 188948 175766 189000 175772
rect 190340 175150 190368 177940
rect 190328 175144 190380 175150
rect 190328 175086 190380 175092
rect 191340 174804 191392 174810
rect 191340 174746 191392 174752
rect 187660 174668 187712 174674
rect 187660 174610 187712 174616
rect 189316 174464 189368 174470
rect 189316 174406 189368 174412
rect 184912 174118 185032 174146
rect 185004 166990 185032 174118
rect 184992 166984 185044 166990
rect 184992 166926 185044 166932
rect 182232 166916 182284 166922
rect 182232 166858 182284 166864
rect 187292 166916 187344 166922
rect 187292 166858 187344 166864
rect 180852 166848 180904 166854
rect 180852 166790 180904 166796
rect 184992 166848 185044 166854
rect 184992 166790 185044 166796
rect 181588 164808 181640 164814
rect 181588 164750 181640 164756
rect 180942 163280 180998 163289
rect 180942 163215 180998 163224
rect 180484 159980 180536 159986
rect 180484 159922 180536 159928
rect 180392 159436 180444 159442
rect 180392 159378 180444 159384
rect 180298 155664 180354 155673
rect 180298 155599 180354 155608
rect 180208 149372 180260 149378
rect 180208 149314 180260 149320
rect 180404 149145 180432 159378
rect 180496 149553 180524 159922
rect 180668 159640 180720 159646
rect 180668 159582 180720 159588
rect 180574 156752 180630 156761
rect 180574 156687 180630 156696
rect 180482 149544 180538 149553
rect 180482 149479 180538 149488
rect 180390 149136 180446 149145
rect 180390 149071 180446 149080
rect 177632 148080 177684 148086
rect 177632 148022 177684 148028
rect 180588 147814 180616 156687
rect 180680 149961 180708 159582
rect 180758 157976 180814 157985
rect 180758 157911 180814 157920
rect 180666 149952 180722 149961
rect 180666 149887 180722 149896
rect 180772 149446 180800 157911
rect 180956 157674 180984 163215
rect 181126 162872 181182 162881
rect 181126 162807 181182 162816
rect 181036 161000 181088 161006
rect 181036 160942 181088 160948
rect 181048 160870 181076 160942
rect 181036 160864 181088 160870
rect 181036 160806 181088 160812
rect 181034 159608 181090 159617
rect 181034 159543 181090 159552
rect 181048 159306 181076 159543
rect 181036 159300 181088 159306
rect 181036 159242 181088 159248
rect 180944 157668 180996 157674
rect 180944 157610 180996 157616
rect 180942 157568 180998 157577
rect 180942 157503 180998 157512
rect 180850 156344 180906 156353
rect 180850 156279 180906 156288
rect 180760 149440 180812 149446
rect 180760 149382 180812 149388
rect 180864 147882 180892 156279
rect 180956 148902 180984 157503
rect 181036 156444 181088 156450
rect 181036 156386 181088 156392
rect 181048 155265 181076 156386
rect 181140 156382 181168 162807
rect 181218 162464 181274 162473
rect 181218 162399 181274 162408
rect 181128 156376 181180 156382
rect 181128 156318 181180 156324
rect 181232 156246 181260 162399
rect 181402 161240 181458 161249
rect 181402 161175 181458 161184
rect 181416 160666 181444 161175
rect 181600 160682 181628 164750
rect 185004 163796 185032 166790
rect 187304 163796 187332 166858
rect 189328 163810 189356 174406
rect 191352 166582 191380 174746
rect 191720 174146 191748 177940
rect 192720 174668 192772 174674
rect 192720 174610 192772 174616
rect 191720 174118 192024 174146
rect 191996 167330 192024 174118
rect 191984 167324 192036 167330
rect 191984 167266 192036 167272
rect 191984 166984 192036 166990
rect 191984 166926 192036 166932
rect 191340 166576 191392 166582
rect 191340 166518 191392 166524
rect 189328 163782 189710 163810
rect 191996 163796 192024 166926
rect 192732 166718 192760 174610
rect 193008 174146 193036 177940
rect 194388 174146 194416 177940
rect 195768 174146 195796 177940
rect 197056 174470 197084 177940
rect 198240 175824 198292 175830
rect 198240 175766 198292 175772
rect 197044 174464 197096 174470
rect 197044 174406 197096 174412
rect 197504 174464 197556 174470
rect 197504 174406 197556 174412
rect 193008 174118 193404 174146
rect 194388 174118 194784 174146
rect 195768 174118 196164 174146
rect 193376 167194 193404 174118
rect 194756 167262 194784 174118
rect 194744 167256 194796 167262
rect 194744 167198 194796 167204
rect 193364 167188 193416 167194
rect 193364 167130 193416 167136
rect 196136 167126 196164 174118
rect 196124 167120 196176 167126
rect 196124 167062 196176 167068
rect 197516 167058 197544 174406
rect 197504 167052 197556 167058
rect 197504 166994 197556 167000
rect 198252 166854 198280 175766
rect 198436 174470 198464 177940
rect 199620 175144 199672 175150
rect 199620 175086 199672 175092
rect 198424 174464 198476 174470
rect 198424 174406 198476 174412
rect 198884 174464 198936 174470
rect 198884 174406 198936 174412
rect 198896 166990 198924 174406
rect 198884 166984 198936 166990
rect 198884 166926 198936 166932
rect 198240 166848 198292 166854
rect 198240 166790 198292 166796
rect 199068 166848 199120 166854
rect 199068 166790 199120 166796
rect 192720 166712 192772 166718
rect 192720 166654 192772 166660
rect 196676 166712 196728 166718
rect 196676 166654 196728 166660
rect 194376 166576 194428 166582
rect 194376 166518 194428 166524
rect 194388 163796 194416 166518
rect 196688 163796 196716 166654
rect 199080 163796 199108 166790
rect 199632 166718 199660 175086
rect 199816 174470 199844 177940
rect 201104 174470 201132 177940
rect 202484 175150 202512 177940
rect 203864 175694 203892 177940
rect 203852 175688 203904 175694
rect 203852 175630 203904 175636
rect 202472 175144 202524 175150
rect 202472 175086 202524 175092
rect 205152 174470 205180 177940
rect 206532 175626 206560 177940
rect 206520 175620 206572 175626
rect 206520 175562 206572 175568
rect 199804 174464 199856 174470
rect 199804 174406 199856 174412
rect 200264 174464 200316 174470
rect 200264 174406 200316 174412
rect 201092 174464 201144 174470
rect 201092 174406 201144 174412
rect 201644 174464 201696 174470
rect 201644 174406 201696 174412
rect 205140 174464 205192 174470
rect 205140 174406 205192 174412
rect 205784 174464 205836 174470
rect 205784 174406 205836 174412
rect 200276 166922 200304 174406
rect 200264 166916 200316 166922
rect 200264 166858 200316 166864
rect 201656 166854 201684 174406
rect 205796 168894 205824 174406
rect 207912 172265 207940 177940
rect 209200 175558 209228 177940
rect 209188 175552 209240 175558
rect 209188 175494 209240 175500
rect 210580 174470 210608 177940
rect 211960 175694 211988 177940
rect 211948 175688 212000 175694
rect 211948 175630 212000 175636
rect 213248 175558 213276 177940
rect 213236 175552 213288 175558
rect 213236 175494 213288 175500
rect 214628 175422 214656 177940
rect 216008 175422 216036 177940
rect 214616 175416 214668 175422
rect 214616 175358 214668 175364
rect 215996 175416 216048 175422
rect 215996 175358 216048 175364
rect 217296 175354 217324 177940
rect 217284 175348 217336 175354
rect 217284 175290 217336 175296
rect 210568 174464 210620 174470
rect 210568 174406 210620 174412
rect 211304 174464 211356 174470
rect 211304 174406 211356 174412
rect 207898 172256 207954 172265
rect 207898 172191 207954 172200
rect 211316 170254 211344 174406
rect 218676 172401 218704 177940
rect 220056 175286 220084 177940
rect 221344 175286 221372 177940
rect 220044 175280 220096 175286
rect 220044 175222 220096 175228
rect 221332 175280 221384 175286
rect 221332 175222 221384 175228
rect 222724 175218 222752 177940
rect 226772 175762 226800 177940
rect 226760 175756 226812 175762
rect 226760 175698 226812 175704
rect 228152 175626 228180 177940
rect 228692 175824 228744 175830
rect 228692 175766 228744 175772
rect 228704 175626 228732 175766
rect 228140 175620 228192 175626
rect 228140 175562 228192 175568
rect 228692 175620 228744 175626
rect 228692 175562 228744 175568
rect 224460 175416 224512 175422
rect 224460 175358 224512 175364
rect 222712 175212 222764 175218
rect 222712 175154 222764 175160
rect 218662 172392 218718 172401
rect 218662 172327 218718 172336
rect 211304 170248 211356 170254
rect 211304 170190 211356 170196
rect 205784 168888 205836 168894
rect 205784 168830 205836 168836
rect 203760 167324 203812 167330
rect 203760 167266 203812 167272
rect 201644 166848 201696 166854
rect 201644 166790 201696 166796
rect 199620 166712 199672 166718
rect 199620 166654 199672 166660
rect 201460 166712 201512 166718
rect 201460 166654 201512 166660
rect 201472 163796 201500 166654
rect 203772 163796 203800 167266
rect 208452 167256 208504 167262
rect 208452 167198 208504 167204
rect 206152 167188 206204 167194
rect 206152 167130 206204 167136
rect 206164 163796 206192 167130
rect 208464 163796 208492 167198
rect 210844 167120 210896 167126
rect 210844 167062 210896 167068
rect 210856 163796 210884 167062
rect 213236 167052 213288 167058
rect 213236 166994 213288 167000
rect 213248 163796 213276 166994
rect 215536 166984 215588 166990
rect 215536 166926 215588 166932
rect 215548 163796 215576 166926
rect 217928 166916 217980 166922
rect 217928 166858 217980 166864
rect 217940 163796 217968 166858
rect 220228 166848 220280 166854
rect 220228 166790 220280 166796
rect 220240 163796 220268 166790
rect 222620 166236 222672 166242
rect 222620 166178 222672 166184
rect 222632 163796 222660 166178
rect 181770 163688 181826 163697
rect 181770 163623 181826 163632
rect 181784 163590 181812 163623
rect 181772 163584 181824 163590
rect 181772 163526 181824 163532
rect 181772 163448 181824 163454
rect 181772 163390 181824 163396
rect 181404 160660 181456 160666
rect 181600 160654 181720 160682
rect 181404 160602 181456 160608
rect 181402 160424 181458 160433
rect 181402 160359 181458 160368
rect 181310 160016 181366 160025
rect 181310 159951 181366 159960
rect 181324 159374 181352 159951
rect 181416 159510 181444 160359
rect 181404 159504 181456 159510
rect 181404 159446 181456 159452
rect 181312 159368 181364 159374
rect 181312 159310 181364 159316
rect 181494 159200 181550 159209
rect 181494 159135 181550 159144
rect 181508 157946 181536 159135
rect 181496 157940 181548 157946
rect 181496 157882 181548 157888
rect 181220 156240 181272 156246
rect 181220 156182 181272 156188
rect 181034 155256 181090 155265
rect 181034 155191 181090 155200
rect 181220 155084 181272 155090
rect 181220 155026 181272 155032
rect 181036 155016 181088 155022
rect 181036 154958 181088 154964
rect 181048 154857 181076 154958
rect 181128 154880 181180 154886
rect 181034 154848 181090 154857
rect 181128 154822 181180 154828
rect 181034 154783 181090 154792
rect 181140 154041 181168 154822
rect 181232 154449 181260 155026
rect 181218 154440 181274 154449
rect 181218 154375 181274 154384
rect 181126 154032 181182 154041
rect 181126 153967 181182 153976
rect 181220 153656 181272 153662
rect 181692 153633 181720 160654
rect 181220 153598 181272 153604
rect 181678 153624 181734 153633
rect 181036 153588 181088 153594
rect 181036 153530 181088 153536
rect 181048 153225 181076 153530
rect 181128 153452 181180 153458
rect 181128 153394 181180 153400
rect 181034 153216 181090 153225
rect 181034 153151 181090 153160
rect 181140 152409 181168 153394
rect 181232 152817 181260 153598
rect 181678 153559 181734 153568
rect 181218 152808 181274 152817
rect 181218 152743 181274 152752
rect 181126 152400 181182 152409
rect 181036 152364 181088 152370
rect 181126 152335 181182 152344
rect 181036 152306 181088 152312
rect 181048 151593 181076 152306
rect 181128 152296 181180 152302
rect 181128 152238 181180 152244
rect 181034 151584 181090 151593
rect 181034 151519 181090 151528
rect 181140 151185 181168 152238
rect 181784 152001 181812 163390
rect 182324 162088 182376 162094
rect 182322 162056 182324 162065
rect 182376 162056 182378 162065
rect 182322 161991 182378 162000
rect 182322 161648 182378 161657
rect 182322 161583 182378 161592
rect 181864 161000 181916 161006
rect 181864 160942 181916 160948
rect 181770 151992 181826 152001
rect 181770 151927 181826 151936
rect 181126 151176 181182 151185
rect 181126 151111 181182 151120
rect 181876 150369 181904 160942
rect 181956 160932 182008 160938
rect 181956 160874 182008 160880
rect 181968 156330 181996 160874
rect 182138 160832 182194 160841
rect 182336 160802 182364 161583
rect 182138 160767 182194 160776
rect 182324 160796 182376 160802
rect 182152 160734 182180 160767
rect 182324 160738 182376 160744
rect 182140 160728 182192 160734
rect 182140 160670 182192 160676
rect 182138 158792 182194 158801
rect 182138 158727 182194 158736
rect 182046 157160 182102 157169
rect 182046 157095 182102 157104
rect 182060 156518 182088 157095
rect 182048 156512 182100 156518
rect 182048 156454 182100 156460
rect 181968 156302 182088 156330
rect 181954 156072 182010 156081
rect 181954 156007 182010 156016
rect 181862 150360 181918 150369
rect 181862 150295 181918 150304
rect 181772 149508 181824 149514
rect 181772 149450 181824 149456
rect 180944 148896 180996 148902
rect 180944 148838 180996 148844
rect 181784 148329 181812 149450
rect 181770 148320 181826 148329
rect 181770 148255 181826 148264
rect 180852 147876 180904 147882
rect 180852 147818 180904 147824
rect 180576 147808 180628 147814
rect 180576 147750 180628 147756
rect 181968 146726 181996 156007
rect 182060 150777 182088 156302
rect 182152 150806 182180 158727
rect 182322 158384 182378 158393
rect 182322 158319 182378 158328
rect 182336 150874 182364 158319
rect 182324 150868 182376 150874
rect 182324 150810 182376 150816
rect 182140 150800 182192 150806
rect 182046 150768 182102 150777
rect 182140 150742 182192 150748
rect 182046 150703 182102 150712
rect 182324 149576 182376 149582
rect 182324 149518 182376 149524
rect 182336 148737 182364 149518
rect 182322 148728 182378 148737
rect 182322 148663 182378 148672
rect 182324 148080 182376 148086
rect 182322 148048 182324 148057
rect 182376 148048 182378 148057
rect 182322 147983 182378 147992
rect 181956 146720 182008 146726
rect 181956 146662 182008 146668
rect 203864 145434 203892 147884
rect 176160 145428 176212 145434
rect 176160 145370 176212 145376
rect 203852 145428 203904 145434
rect 203852 145370 203904 145376
rect 173950 144376 174006 144385
rect 173950 144311 174006 144320
rect 173858 143288 173914 143297
rect 173858 143223 173914 143232
rect 173398 142200 173454 142209
rect 173398 142135 173454 142144
rect 224472 139926 224500 175358
rect 228704 168214 228732 175562
rect 231372 173042 231400 203471
rect 231464 192665 231492 204802
rect 231556 195793 231584 208950
rect 231648 197425 231676 211670
rect 231740 202049 231768 218674
rect 231832 217689 231860 233158
rect 236892 232474 236920 235862
rect 237628 232542 237656 235862
rect 237996 232610 238024 235862
rect 238548 232678 238576 235862
rect 239192 233222 239220 235862
rect 239180 233216 239232 233222
rect 239180 233158 239232 233164
rect 239652 233086 239680 235862
rect 239640 233080 239692 233086
rect 239640 233022 239692 233028
rect 238536 232672 238588 232678
rect 238536 232614 238588 232620
rect 237984 232604 238036 232610
rect 237984 232546 238036 232552
rect 237616 232536 237668 232542
rect 237616 232478 237668 232484
rect 236880 232468 236932 232474
rect 236880 232410 236932 232416
rect 232004 228252 232056 228258
rect 232004 228194 232056 228200
rect 232016 227073 232044 228194
rect 232002 227064 232058 227073
rect 232002 226999 232058 227008
rect 231910 225568 231966 225577
rect 231910 225503 231912 225512
rect 231964 225503 231966 225512
rect 234120 225532 234172 225538
rect 231912 225474 231964 225480
rect 234120 225474 234172 225480
rect 232004 224104 232056 224110
rect 232004 224046 232056 224052
rect 232016 223945 232044 224046
rect 232002 223936 232058 223945
rect 232002 223871 232058 223880
rect 232740 218868 232792 218874
rect 232740 218810 232792 218816
rect 231818 217680 231874 217689
rect 231818 217615 231874 217624
rect 232002 216048 232058 216057
rect 232002 215983 232004 215992
rect 232056 215983 232058 215992
rect 232004 215954 232056 215960
rect 231820 215876 231872 215882
rect 231820 215818 231872 215824
rect 231726 202040 231782 202049
rect 231726 201975 231782 201984
rect 231832 200553 231860 215818
rect 231912 213156 231964 213162
rect 231912 213098 231964 213104
rect 231818 200544 231874 200553
rect 231818 200479 231874 200488
rect 231728 199352 231780 199358
rect 231728 199294 231780 199300
rect 231634 197416 231690 197425
rect 231634 197351 231690 197360
rect 231542 195784 231598 195793
rect 231542 195719 231598 195728
rect 231450 192656 231506 192665
rect 231450 192591 231506 192600
rect 231740 189537 231768 199294
rect 231924 198921 231952 213098
rect 232002 212376 232058 212385
rect 232002 212311 232004 212320
rect 232056 212311 232058 212320
rect 232004 212282 232056 212288
rect 232002 209520 232058 209529
rect 232002 209455 232058 209464
rect 232016 209286 232044 209455
rect 232004 209280 232056 209286
rect 232004 209222 232056 209228
rect 232002 206528 232058 206537
rect 232002 206463 232004 206472
rect 232056 206463 232058 206472
rect 232004 206434 232056 206440
rect 232004 206220 232056 206226
rect 232004 206162 232056 206168
rect 231910 198912 231966 198921
rect 231910 198847 231966 198856
rect 231820 197924 231872 197930
rect 231820 197866 231872 197872
rect 231726 189528 231782 189537
rect 231726 189463 231782 189472
rect 231832 188041 231860 197866
rect 232016 194297 232044 206162
rect 232002 194288 232058 194297
rect 232002 194223 232058 194232
rect 231818 188032 231874 188041
rect 231818 187967 231874 187976
rect 231820 186840 231872 186846
rect 231820 186782 231872 186788
rect 231832 186409 231860 186782
rect 231818 186400 231874 186409
rect 231818 186335 231874 186344
rect 231820 185480 231872 185486
rect 231820 185422 231872 185428
rect 231832 184913 231860 185422
rect 231818 184904 231874 184913
rect 231818 184839 231874 184848
rect 231636 180924 231688 180930
rect 231636 180866 231688 180872
rect 231648 180153 231676 180866
rect 231634 180144 231690 180153
rect 231634 180079 231690 180088
rect 231636 179904 231688 179910
rect 231636 179846 231688 179852
rect 231648 178657 231676 179846
rect 231634 178648 231690 178657
rect 231634 178583 231690 178592
rect 231360 173036 231412 173042
rect 231360 172978 231412 172984
rect 232752 172022 232780 218810
rect 232832 175484 232884 175490
rect 232832 175426 232884 175432
rect 232740 172016 232792 172022
rect 232740 171958 232792 171964
rect 228692 168208 228744 168214
rect 228692 168150 228744 168156
rect 228876 168208 228928 168214
rect 228876 168150 228928 168156
rect 225932 164740 225984 164746
rect 225932 164682 225984 164688
rect 225944 163697 225972 164682
rect 225930 163688 225986 163697
rect 225930 163623 225986 163632
rect 228888 163425 228916 168150
rect 231820 166576 231872 166582
rect 231820 166518 231872 166524
rect 230900 166236 230952 166242
rect 230900 166178 230952 166184
rect 228690 163416 228746 163425
rect 226392 163380 226444 163386
rect 226392 163322 226444 163328
rect 228612 163374 228690 163402
rect 226404 163289 226432 163322
rect 226484 163312 226536 163318
rect 226390 163280 226446 163289
rect 225564 163244 225616 163250
rect 228612 163300 228640 163374
rect 228690 163351 228746 163360
rect 228874 163416 228930 163425
rect 228874 163351 228930 163360
rect 230912 163318 230940 166178
rect 231832 163386 231860 166518
rect 231820 163380 231872 163386
rect 231820 163322 231872 163328
rect 230900 163312 230952 163318
rect 228612 163272 228732 163300
rect 226484 163254 226536 163260
rect 226390 163215 226446 163224
rect 225564 163186 225616 163192
rect 225576 162473 225604 163186
rect 225932 163040 225984 163046
rect 225932 162982 225984 162988
rect 225562 162464 225618 162473
rect 225562 162399 225618 162408
rect 225944 162065 225972 162982
rect 226496 162881 226524 163254
rect 226482 162872 226538 162881
rect 226482 162807 226538 162816
rect 225930 162056 225986 162065
rect 225930 161991 225986 162000
rect 226484 161680 226536 161686
rect 226482 161648 226484 161657
rect 226536 161648 226538 161657
rect 226482 161583 226538 161592
rect 226484 161544 226536 161550
rect 226484 161486 226536 161492
rect 226496 161249 226524 161486
rect 226482 161240 226538 161249
rect 225932 161204 225984 161210
rect 226482 161175 226538 161184
rect 225932 161146 225984 161152
rect 225944 160841 225972 161146
rect 225930 160832 225986 160841
rect 225930 160767 225986 160776
rect 226484 160592 226536 160598
rect 226482 160560 226484 160569
rect 226536 160560 226538 160569
rect 225932 160524 225984 160530
rect 226482 160495 226538 160504
rect 225932 160466 225984 160472
rect 225564 160320 225616 160326
rect 225564 160262 225616 160268
rect 225576 160161 225604 160262
rect 225562 160152 225618 160161
rect 225562 160087 225618 160096
rect 225944 159753 225972 160466
rect 226484 159776 226536 159782
rect 225930 159744 225986 159753
rect 226484 159718 226536 159724
rect 225930 159679 225986 159688
rect 226496 159345 226524 159718
rect 226482 159336 226538 159345
rect 226482 159271 226538 159280
rect 226484 158960 226536 158966
rect 226482 158928 226484 158937
rect 226536 158928 226538 158937
rect 226482 158863 226538 158872
rect 225564 158688 225616 158694
rect 225564 158630 225616 158636
rect 225576 158529 225604 158630
rect 225562 158520 225618 158529
rect 225562 158455 225618 158464
rect 226392 158280 226444 158286
rect 226392 158222 226444 158228
rect 226404 158121 226432 158222
rect 226390 158112 226446 158121
rect 226390 158047 226446 158056
rect 226300 157736 226352 157742
rect 226298 157704 226300 157713
rect 226352 157704 226354 157713
rect 226298 157639 226354 157648
rect 226484 157464 226536 157470
rect 226482 157432 226484 157441
rect 226536 157432 226538 157441
rect 226482 157367 226538 157376
rect 226482 157024 226538 157033
rect 226482 156959 226484 156968
rect 226536 156959 226538 156968
rect 226484 156930 226536 156936
rect 225378 156616 225434 156625
rect 225378 156551 225380 156560
rect 225432 156551 225434 156560
rect 225380 156522 225432 156528
rect 226482 156208 226538 156217
rect 226482 156143 226538 156152
rect 226496 156042 226524 156143
rect 226484 156036 226536 156042
rect 226484 155978 226536 155984
rect 226482 155800 226538 155809
rect 226482 155735 226538 155744
rect 226496 155634 226524 155735
rect 226484 155628 226536 155634
rect 226484 155570 226536 155576
rect 225562 155392 225618 155401
rect 225562 155327 225564 155336
rect 225616 155327 225618 155336
rect 225564 155298 225616 155304
rect 225746 154984 225802 154993
rect 225746 154919 225802 154928
rect 225760 154546 225788 154919
rect 226114 154576 226170 154585
rect 225748 154540 225800 154546
rect 226114 154511 226170 154520
rect 225748 154482 225800 154488
rect 225838 154304 225894 154313
rect 225838 154239 225894 154248
rect 225852 154138 225880 154239
rect 225840 154132 225892 154138
rect 225840 154074 225892 154080
rect 226128 153866 226156 154511
rect 226482 153896 226538 153905
rect 226116 153860 226168 153866
rect 226482 153831 226538 153840
rect 226116 153802 226168 153808
rect 226496 153798 226524 153831
rect 226484 153792 226536 153798
rect 228704 153769 228732 163272
rect 230900 163254 230952 163260
rect 229336 162088 229388 162094
rect 229336 162030 229388 162036
rect 229348 160598 229376 162030
rect 229336 160592 229388 160598
rect 229336 160534 229388 160540
rect 228414 153760 228470 153769
rect 226484 153734 226536 153740
rect 228336 153718 228414 153746
rect 226114 153488 226170 153497
rect 226114 153423 226116 153432
rect 226168 153423 226170 153432
rect 226116 153394 226168 153400
rect 225746 153080 225802 153089
rect 225746 153015 225802 153024
rect 225378 152672 225434 152681
rect 225378 152607 225380 152616
rect 225432 152607 225434 152616
rect 225380 152578 225432 152584
rect 225760 152438 225788 153015
rect 225748 152432 225800 152438
rect 225748 152374 225800 152380
rect 225930 152264 225986 152273
rect 225930 152199 225986 152208
rect 225944 151758 225972 152199
rect 226114 151856 226170 151865
rect 226114 151791 226170 151800
rect 225932 151752 225984 151758
rect 225932 151694 225984 151700
rect 225378 151448 225434 151457
rect 225378 151383 225380 151392
rect 225432 151383 225434 151392
rect 225380 151354 225432 151360
rect 226128 151010 226156 151791
rect 227956 151752 228008 151758
rect 227956 151694 228008 151700
rect 226482 151176 226538 151185
rect 226482 151111 226484 151120
rect 226536 151111 226538 151120
rect 226484 151082 226536 151088
rect 226116 151004 226168 151010
rect 226116 150946 226168 150952
rect 225562 150768 225618 150777
rect 225562 150703 225618 150712
rect 225576 150126 225604 150703
rect 225746 150360 225802 150369
rect 225746 150295 225802 150304
rect 225564 150120 225616 150126
rect 225564 150062 225616 150068
rect 225760 149650 225788 150295
rect 226482 149952 226538 149961
rect 226538 149910 226616 149938
rect 226482 149887 226538 149896
rect 225748 149644 225800 149650
rect 225748 149586 225800 149592
rect 225562 149544 225618 149553
rect 225562 149479 225618 149488
rect 225378 149136 225434 149145
rect 225378 149071 225380 149080
rect 225432 149071 225434 149080
rect 225380 149042 225432 149048
rect 225576 148358 225604 149479
rect 226482 148728 226538 148737
rect 226482 148663 226484 148672
rect 226536 148663 226538 148672
rect 226484 148634 226536 148640
rect 225564 148352 225616 148358
rect 225564 148294 225616 148300
rect 226482 148320 226538 148329
rect 226482 148255 226484 148264
rect 226536 148255 226538 148264
rect 226484 148226 226536 148232
rect 225562 148048 225618 148057
rect 225562 147983 225618 147992
rect 225576 147406 225604 147983
rect 225564 147400 225616 147406
rect 225564 147342 225616 147348
rect 226588 145366 226616 149910
rect 227968 149582 227996 151694
rect 228048 151140 228100 151146
rect 228048 151082 228100 151088
rect 227956 149576 228008 149582
rect 227956 149518 228008 149524
rect 228060 148154 228088 151082
rect 228048 148148 228100 148154
rect 228048 148090 228100 148096
rect 228336 145978 228364 153718
rect 228414 153695 228470 153704
rect 228690 153760 228746 153769
rect 228690 153695 228746 153704
rect 229244 151412 229296 151418
rect 229244 151354 229296 151360
rect 229152 151004 229204 151010
rect 229152 150946 229204 150952
rect 229164 149514 229192 150946
rect 229152 149508 229204 149514
rect 229152 149450 229204 149456
rect 229256 148222 229284 151354
rect 230624 150120 230676 150126
rect 230624 150062 230676 150068
rect 230348 149644 230400 149650
rect 230348 149586 230400 149592
rect 229244 148216 229296 148222
rect 229244 148158 229296 148164
rect 230360 146386 230388 149586
rect 230636 146726 230664 150062
rect 232004 147400 232056 147406
rect 232004 147342 232056 147348
rect 230624 146720 230676 146726
rect 230624 146662 230676 146668
rect 230348 146380 230400 146386
rect 230348 146322 230400 146328
rect 228324 145972 228376 145978
rect 228324 145914 228376 145920
rect 226576 145360 226628 145366
rect 226576 145302 226628 145308
rect 228324 145292 228376 145298
rect 228324 145234 228376 145240
rect 224460 139920 224512 139926
rect 224460 139862 224512 139868
rect 167880 138628 167932 138634
rect 167880 138570 167932 138576
rect 170824 138628 170876 138634
rect 170824 138570 170876 138576
rect 163924 131624 163976 131630
rect 163924 131566 163976 131572
rect 163740 131216 163792 131222
rect 163740 131158 163792 131164
rect 163936 128708 163964 131566
rect 164292 131556 164344 131562
rect 164292 131498 164344 131504
rect 164304 128708 164332 131498
rect 164660 131148 164712 131154
rect 164660 131090 164712 131096
rect 164672 128708 164700 131090
rect 145340 127544 145392 127550
rect 145340 127486 145392 127492
rect 148742 127512 148798 127521
rect 144420 124892 144472 124898
rect 144420 124834 144472 124840
rect 143040 122104 143092 122110
rect 143040 122046 143092 122052
rect 141660 117956 141712 117962
rect 141660 117898 141712 117904
rect 140280 115236 140332 115242
rect 140280 115178 140332 115184
rect 138992 112584 139044 112590
rect 138992 112526 139044 112532
rect 139004 79202 139032 112526
rect 138992 79196 139044 79202
rect 138992 79138 139044 79144
rect 140292 78998 140320 115178
rect 140372 105512 140424 105518
rect 140372 105454 140424 105460
rect 140384 95794 140412 105454
rect 140464 101364 140516 101370
rect 140464 101306 140516 101312
rect 140372 95788 140424 95794
rect 140372 95730 140424 95736
rect 140476 92734 140504 101306
rect 140556 98576 140608 98582
rect 140556 98518 140608 98524
rect 140464 92728 140516 92734
rect 140464 92670 140516 92676
rect 140568 91646 140596 98518
rect 140556 91640 140608 91646
rect 140556 91582 140608 91588
rect 141672 79066 141700 117898
rect 142764 79128 142816 79134
rect 142764 79070 142816 79076
rect 141660 79060 141712 79066
rect 141660 79002 141712 79008
rect 140280 78992 140332 78998
rect 140280 78934 140332 78940
rect 134850 78487 134906 78496
rect 138900 78516 138952 78522
rect 138900 78458 138952 78464
rect 139636 76340 139688 76346
rect 139636 76282 139688 76288
rect 139648 75569 139676 76282
rect 142776 75818 142804 79070
rect 143052 79066 143080 122046
rect 143132 103132 143184 103138
rect 143132 103074 143184 103080
rect 143144 93890 143172 103074
rect 143776 94428 143828 94434
rect 143776 94370 143828 94376
rect 143132 93884 143184 93890
rect 143132 93826 143184 93832
rect 143684 91708 143736 91714
rect 143684 91650 143736 91656
rect 143500 88920 143552 88926
rect 143500 88862 143552 88868
rect 143512 84710 143540 88862
rect 143696 85254 143724 91650
rect 143788 88858 143816 94370
rect 143776 88852 143828 88858
rect 143776 88794 143828 88800
rect 143684 85248 143736 85254
rect 143684 85190 143736 85196
rect 143500 84704 143552 84710
rect 143500 84646 143552 84652
rect 143224 79196 143276 79202
rect 143224 79138 143276 79144
rect 143040 79060 143092 79066
rect 143040 79002 143092 79008
rect 143236 75818 143264 79138
rect 144328 79128 144380 79134
rect 144328 79070 144380 79076
rect 143776 78992 143828 78998
rect 143776 78934 143828 78940
rect 143788 75818 143816 78934
rect 144340 75818 144368 79070
rect 144432 78386 144460 124834
rect 144602 97048 144658 97057
rect 144602 96983 144658 96992
rect 144616 89198 144644 96983
rect 145246 92424 145302 92433
rect 145246 92359 145302 92368
rect 145260 91714 145288 92359
rect 145248 91708 145300 91714
rect 145248 91650 145300 91656
rect 145246 89432 145302 89441
rect 145246 89367 145302 89376
rect 144604 89192 144656 89198
rect 144604 89134 144656 89140
rect 145260 88926 145288 89367
rect 145248 88920 145300 88926
rect 145248 88862 145300 88868
rect 145352 79406 145380 127486
rect 148742 127447 148798 127456
rect 148756 126666 148784 127447
rect 148744 126660 148796 126666
rect 148744 126602 148796 126608
rect 165120 126660 165172 126666
rect 165120 126602 165172 126608
rect 145614 125336 145670 125345
rect 145614 125271 145670 125280
rect 145628 124830 145656 125271
rect 145616 124824 145668 124830
rect 145616 124766 145668 124772
rect 145614 123024 145670 123033
rect 145614 122959 145670 122968
rect 145628 122042 145656 122959
rect 145616 122036 145668 122042
rect 145616 121978 145668 121984
rect 165132 121974 165160 126602
rect 165120 121968 165172 121974
rect 165120 121910 165172 121916
rect 145614 120576 145670 120585
rect 145614 120511 145670 120520
rect 145628 119322 145656 120511
rect 145616 119316 145668 119322
rect 145616 119258 145668 119264
rect 167892 118817 167920 138570
rect 228336 137154 228364 145234
rect 232016 142714 232044 147342
rect 232004 142708 232056 142714
rect 232004 142650 232056 142656
rect 232844 139897 232872 175426
rect 234132 171954 234160 225474
rect 240388 224110 240416 235862
rect 240756 228258 240784 235862
rect 241584 232474 241612 235862
rect 242504 233018 242532 235862
rect 242492 233012 242544 233018
rect 242492 232954 242544 232960
rect 243056 232542 243084 235862
rect 243608 232950 243636 235862
rect 243596 232944 243648 232950
rect 243596 232886 243648 232892
rect 244160 232882 244188 235862
rect 244436 235862 244496 235890
rect 245048 235862 245384 235890
rect 245600 235862 245844 235890
rect 246152 235862 246488 235890
rect 246704 235862 247040 235890
rect 244148 232876 244200 232882
rect 244148 232818 244200 232824
rect 244436 232678 244464 235862
rect 245356 233222 245384 235862
rect 245344 233216 245396 233222
rect 245344 233158 245396 233164
rect 245816 233086 245844 235862
rect 245804 233080 245856 233086
rect 245804 233022 245856 233028
rect 244424 232672 244476 232678
rect 244424 232614 244476 232620
rect 245804 232604 245856 232610
rect 245804 232546 245856 232552
rect 243044 232536 243096 232542
rect 243044 232478 243096 232484
rect 241572 232468 241624 232474
rect 241572 232410 241624 232416
rect 245436 232468 245488 232474
rect 245436 232410 245488 232416
rect 240744 228252 240796 228258
rect 240744 228194 240796 228200
rect 244424 225464 244476 225470
rect 244424 225406 244476 225412
rect 244056 225396 244108 225402
rect 244056 225338 244108 225344
rect 243320 224988 243372 224994
rect 243320 224930 243372 224936
rect 240376 224104 240428 224110
rect 240376 224046 240428 224052
rect 243332 222834 243360 224930
rect 243688 224920 243740 224926
rect 243688 224862 243740 224868
rect 243700 222834 243728 224862
rect 244068 222834 244096 225338
rect 244436 222834 244464 225406
rect 245448 225266 245476 232410
rect 245436 225260 245488 225266
rect 245436 225202 245488 225208
rect 245620 225056 245672 225062
rect 245620 224998 245672 225004
rect 244884 224648 244936 224654
rect 244884 224590 244936 224596
rect 244896 222834 244924 224590
rect 245252 224580 245304 224586
rect 245252 224522 245304 224528
rect 245264 222834 245292 224522
rect 245632 222834 245660 224998
rect 245816 222834 245844 232546
rect 246460 232474 246488 235862
rect 247012 233290 247040 235862
rect 247196 235862 247256 235890
rect 247808 235862 248144 235890
rect 248360 235862 248512 235890
rect 248912 235862 249248 235890
rect 249464 235862 249800 235890
rect 247000 233284 247052 233290
rect 247000 233226 247052 233232
rect 247196 232864 247224 235862
rect 247736 233624 247788 233630
rect 247736 233566 247788 233572
rect 247644 233012 247696 233018
rect 247644 232954 247696 232960
rect 247552 232876 247604 232882
rect 247196 232836 247316 232864
rect 246724 232808 246776 232814
rect 246724 232750 246776 232756
rect 246448 232468 246500 232474
rect 246448 232410 246500 232416
rect 246448 224444 246500 224450
rect 246448 224386 246500 224392
rect 246460 222834 246488 224386
rect 246736 222834 246764 232750
rect 247184 232740 247236 232746
rect 247184 232682 247236 232688
rect 247000 232536 247052 232542
rect 247000 232478 247052 232484
rect 247012 225198 247040 232478
rect 247000 225192 247052 225198
rect 247000 225134 247052 225140
rect 247196 222834 247224 232682
rect 247288 224790 247316 232836
rect 247552 232818 247604 232824
rect 247368 232672 247420 232678
rect 247368 232614 247420 232620
rect 247276 224784 247328 224790
rect 247276 224726 247328 224732
rect 247380 224110 247408 232614
rect 247564 224858 247592 232818
rect 247656 225130 247684 232954
rect 247644 225124 247696 225130
rect 247644 225066 247696 225072
rect 247552 224852 247604 224858
rect 247552 224794 247604 224800
rect 247552 224716 247604 224722
rect 247552 224658 247604 224664
rect 247368 224104 247420 224110
rect 247368 224046 247420 224052
rect 247564 222834 247592 224658
rect 247748 222834 247776 233566
rect 248012 232808 248064 232814
rect 248012 232750 248064 232756
rect 248024 225402 248052 232750
rect 248116 232678 248144 235862
rect 248484 233306 248512 235862
rect 249116 233760 249168 233766
rect 249116 233702 249168 233708
rect 248656 233556 248708 233562
rect 248656 233498 248708 233504
rect 248392 233278 248512 233306
rect 248288 232944 248340 232950
rect 248288 232886 248340 232892
rect 248104 232672 248156 232678
rect 248104 232614 248156 232620
rect 248196 232536 248248 232542
rect 248196 232478 248248 232484
rect 248012 225396 248064 225402
rect 248012 225338 248064 225344
rect 248208 222834 248236 232478
rect 248300 225402 248328 232886
rect 248288 225396 248340 225402
rect 248288 225338 248340 225344
rect 248392 224246 248420 233278
rect 248472 233148 248524 233154
rect 248472 233090 248524 233096
rect 248484 225282 248512 233090
rect 248564 232808 248616 232814
rect 248564 232750 248616 232756
rect 248576 225470 248604 232750
rect 248564 225464 248616 225470
rect 248564 225406 248616 225412
rect 248484 225254 248604 225282
rect 248380 224240 248432 224246
rect 248380 224182 248432 224188
rect 248576 222834 248604 225254
rect 248668 224586 248696 233498
rect 248932 233488 248984 233494
rect 248932 233430 248984 233436
rect 248656 224580 248708 224586
rect 248656 224522 248708 224528
rect 248944 222834 248972 233430
rect 249024 233420 249076 233426
rect 249024 233362 249076 233368
rect 249036 224654 249064 233362
rect 249128 224722 249156 233702
rect 249220 224722 249248 235862
rect 249300 233692 249352 233698
rect 249300 233634 249352 233640
rect 249116 224716 249168 224722
rect 249116 224658 249168 224664
rect 249208 224716 249260 224722
rect 249208 224658 249260 224664
rect 249024 224648 249076 224654
rect 249024 224590 249076 224596
rect 249312 222834 249340 233634
rect 249576 233284 249628 233290
rect 249576 233226 249628 233232
rect 249392 233216 249444 233222
rect 249392 233158 249444 233164
rect 249484 233216 249536 233222
rect 249484 233158 249536 233164
rect 249404 224518 249432 233158
rect 249496 225062 249524 233158
rect 249484 225056 249536 225062
rect 249484 224998 249536 225004
rect 249392 224512 249444 224518
rect 249392 224454 249444 224460
rect 249588 224314 249616 233226
rect 249668 233080 249720 233086
rect 249668 233022 249720 233028
rect 249680 224586 249708 233022
rect 249772 224654 249800 235862
rect 249956 235862 250016 235890
rect 250568 235862 251088 235890
rect 251212 235862 251364 235890
rect 251764 235862 252100 235890
rect 252316 235862 252744 235890
rect 252868 235862 253112 235890
rect 249852 233080 249904 233086
rect 249852 233022 249904 233028
rect 249760 224648 249812 224654
rect 249760 224590 249812 224596
rect 249668 224580 249720 224586
rect 249668 224522 249720 224528
rect 249576 224308 249628 224314
rect 249576 224250 249628 224256
rect 249864 222834 249892 233022
rect 249956 232762 249984 235862
rect 250312 233216 250364 233222
rect 250312 233158 250364 233164
rect 249956 232734 250076 232762
rect 249944 232672 249996 232678
rect 249944 232614 249996 232620
rect 249956 224382 249984 232614
rect 250048 225470 250076 232734
rect 250036 225464 250088 225470
rect 250036 225406 250088 225412
rect 249944 224376 249996 224382
rect 249944 224318 249996 224324
rect 250324 222834 250352 233158
rect 250864 225260 250916 225266
rect 250864 225202 250916 225208
rect 250680 224784 250732 224790
rect 250680 224726 250732 224732
rect 250692 222834 250720 224726
rect 250876 222834 250904 225202
rect 251060 225062 251088 235862
rect 251336 225266 251364 235862
rect 252072 232678 252100 235862
rect 252060 232672 252112 232678
rect 252060 232614 252112 232620
rect 251416 232468 251468 232474
rect 251416 232410 251468 232416
rect 251324 225260 251376 225266
rect 251324 225202 251376 225208
rect 251428 225130 251456 232410
rect 252716 225402 252744 235862
rect 253084 232610 253112 235862
rect 253176 235862 253420 235890
rect 253636 235862 253972 235890
rect 254188 235862 254524 235890
rect 254740 235862 255076 235890
rect 255568 235862 255628 235890
rect 255844 235862 256180 235890
rect 256396 235862 256732 235890
rect 256948 235862 257284 235890
rect 257500 235862 257836 235890
rect 258328 235862 258480 235890
rect 258696 235862 259032 235890
rect 259248 235862 259584 235890
rect 259800 235862 260136 235890
rect 260352 235862 260688 235890
rect 261088 235862 261240 235890
rect 261456 235862 261792 235890
rect 262008 235862 262344 235890
rect 262560 235862 262896 235890
rect 263112 235862 263448 235890
rect 263848 235862 264000 235890
rect 264216 235862 264552 235890
rect 253072 232604 253124 232610
rect 253072 232546 253124 232552
rect 252060 225396 252112 225402
rect 252060 225338 252112 225344
rect 252704 225396 252756 225402
rect 252704 225338 252756 225344
rect 251692 225192 251744 225198
rect 251692 225134 251744 225140
rect 251324 225124 251376 225130
rect 251324 225066 251376 225072
rect 251416 225124 251468 225130
rect 251416 225066 251468 225072
rect 251048 225056 251100 225062
rect 251048 224998 251100 225004
rect 251336 222834 251364 225066
rect 251704 222834 251732 225134
rect 252072 222834 252100 225338
rect 253176 224994 253204 235862
rect 253164 224988 253216 224994
rect 253164 224930 253216 224936
rect 253636 224926 253664 235862
rect 254188 232882 254216 235862
rect 254176 232876 254228 232882
rect 254176 232818 254228 232824
rect 254740 232814 254768 235862
rect 255568 233426 255596 235862
rect 255844 233562 255872 235862
rect 255832 233556 255884 233562
rect 255832 233498 255884 233504
rect 255556 233420 255608 233426
rect 255556 233362 255608 233368
rect 256396 233290 256424 235862
rect 256384 233284 256436 233290
rect 256384 233226 256436 233232
rect 256948 232950 256976 235862
rect 256936 232944 256988 232950
rect 256936 232886 256988 232892
rect 254728 232808 254780 232814
rect 254728 232750 254780 232756
rect 257028 232672 257080 232678
rect 257028 232614 257080 232620
rect 256200 232468 256252 232474
rect 256200 232410 256252 232416
rect 254728 229680 254780 229686
rect 254728 229622 254780 229628
rect 254740 225470 254768 229622
rect 254728 225464 254780 225470
rect 254728 225406 254780 225412
rect 253992 225124 254044 225130
rect 253992 225066 254044 225072
rect 253624 224920 253676 224926
rect 253624 224862 253676 224868
rect 252428 224852 252480 224858
rect 252428 224794 252480 224800
rect 252440 222834 252468 224794
rect 253624 224580 253676 224586
rect 253624 224522 253676 224528
rect 253256 224512 253308 224518
rect 253256 224454 253308 224460
rect 252796 224104 252848 224110
rect 252796 224046 252848 224052
rect 252808 223106 252836 224046
rect 252808 223078 252882 223106
rect 243116 222806 243360 222834
rect 243484 222806 243728 222834
rect 243852 222806 244096 222834
rect 244220 222806 244464 222834
rect 244588 222806 244924 222834
rect 245048 222806 245292 222834
rect 245416 222806 245660 222834
rect 245784 222806 245844 222834
rect 246152 222806 246488 222834
rect 246612 222806 246764 222834
rect 246980 222806 247224 222834
rect 247348 222806 247592 222834
rect 247716 222806 247776 222834
rect 248176 222806 248236 222834
rect 248544 222806 248604 222834
rect 248912 222806 248972 222834
rect 249280 222806 249340 222834
rect 249740 222806 249892 222834
rect 250108 222806 250352 222834
rect 250476 222806 250720 222834
rect 250844 222806 250904 222834
rect 251304 222806 251364 222834
rect 251672 222806 251732 222834
rect 252040 222806 252100 222834
rect 252408 222806 252468 222834
rect 252854 222820 252882 223078
rect 253268 222834 253296 224454
rect 253636 222834 253664 224522
rect 254004 222834 254032 225066
rect 256016 224852 256068 224858
rect 256016 224794 256068 224800
rect 254452 224580 254504 224586
rect 254452 224522 254504 224528
rect 254464 222834 254492 224522
rect 255188 224376 255240 224382
rect 255188 224318 255240 224324
rect 254820 224308 254872 224314
rect 254820 224250 254872 224256
rect 254832 222834 254860 224250
rect 255200 222834 255228 224318
rect 255556 224172 255608 224178
rect 255556 224114 255608 224120
rect 255568 222834 255596 224114
rect 256028 222834 256056 224794
rect 256212 224450 256240 232410
rect 256752 224920 256804 224926
rect 256752 224862 256804 224868
rect 256384 224716 256436 224722
rect 256384 224658 256436 224664
rect 256200 224444 256252 224450
rect 256200 224386 256252 224392
rect 256396 222834 256424 224658
rect 256764 222834 256792 224862
rect 257040 223090 257068 232614
rect 257500 232474 257528 235862
rect 258328 233018 258356 235862
rect 258316 233012 258368 233018
rect 258316 232954 258368 232960
rect 258696 232746 258724 235862
rect 259248 233766 259276 235862
rect 259236 233760 259288 233766
rect 259236 233702 259288 233708
rect 259800 233698 259828 235862
rect 259788 233692 259840 233698
rect 259788 233634 259840 233640
rect 258960 233284 259012 233290
rect 258960 233226 259012 233232
rect 258684 232740 258736 232746
rect 258684 232682 258736 232688
rect 257488 232468 257540 232474
rect 257488 232410 257540 232416
rect 258684 225464 258736 225470
rect 258684 225406 258736 225412
rect 258316 225396 258368 225402
rect 258316 225338 258368 225344
rect 257580 225192 257632 225198
rect 257580 225134 257632 225140
rect 257120 224988 257172 224994
rect 257120 224930 257172 224936
rect 257028 223084 257080 223090
rect 257028 223026 257080 223032
rect 257132 222834 257160 224930
rect 257592 222834 257620 225134
rect 257902 223084 257954 223090
rect 257902 223026 257954 223032
rect 253236 222806 253296 222834
rect 253604 222806 253664 222834
rect 253972 222806 254032 222834
rect 254432 222806 254492 222834
rect 254800 222806 254860 222834
rect 255168 222806 255228 222834
rect 255536 222806 255596 222834
rect 255996 222806 256056 222834
rect 256364 222806 256424 222834
rect 256732 222806 256792 222834
rect 257100 222806 257160 222834
rect 257560 222806 257620 222834
rect 257914 222820 257942 223026
rect 258328 222834 258356 225338
rect 258696 222834 258724 225406
rect 258296 222806 258356 222834
rect 258664 222806 258724 222834
rect 239364 221384 239416 221390
rect 239364 221326 239416 221332
rect 238260 216012 238312 216018
rect 238260 215954 238312 215960
rect 236880 212340 236932 212346
rect 236880 212282 236932 212288
rect 235500 209280 235552 209286
rect 235500 209222 235552 209228
rect 234212 206492 234264 206498
rect 234212 206434 234264 206440
rect 234224 172906 234252 206434
rect 234304 195204 234356 195210
rect 234304 195146 234356 195152
rect 234316 186846 234344 195146
rect 234304 186840 234356 186846
rect 234304 186782 234356 186788
rect 235512 172974 235540 209222
rect 236892 173042 236920 212282
rect 236972 192484 237024 192490
rect 236972 192426 237024 192432
rect 236984 185486 237012 192426
rect 237616 185548 237668 185554
rect 237616 185490 237668 185496
rect 236972 185480 237024 185486
rect 236972 185422 237024 185428
rect 237628 180930 237656 185490
rect 237616 180924 237668 180930
rect 237616 180866 237668 180872
rect 236788 173036 236840 173042
rect 236788 172978 236840 172984
rect 236880 173036 236932 173042
rect 236880 172978 236932 172984
rect 235500 172968 235552 172974
rect 235500 172910 235552 172916
rect 234212 172900 234264 172906
rect 234212 172842 234264 172848
rect 234120 171948 234172 171954
rect 234120 171890 234172 171896
rect 233476 170248 233528 170254
rect 233476 170190 233528 170196
rect 233488 169545 233516 170190
rect 236800 169794 236828 172978
rect 237800 172968 237852 172974
rect 237800 172910 237852 172916
rect 237248 172900 237300 172906
rect 237248 172842 237300 172848
rect 237260 169794 237288 172842
rect 237812 169794 237840 172910
rect 238272 171750 238300 215954
rect 238352 173036 238404 173042
rect 238352 172978 238404 172984
rect 238260 171744 238312 171750
rect 238260 171686 238312 171692
rect 238364 169794 238392 172978
rect 239272 172016 239324 172022
rect 239272 171958 239324 171964
rect 238996 171744 239048 171750
rect 238996 171686 239048 171692
rect 239008 169794 239036 171686
rect 239284 169930 239312 171958
rect 239376 170050 239404 221326
rect 240926 218768 240982 218777
rect 240926 218703 240928 218712
rect 240980 218703 240982 218712
rect 240928 218674 240980 218680
rect 240466 216320 240522 216329
rect 240466 216255 240522 216264
rect 240480 215882 240508 216255
rect 240468 215876 240520 215882
rect 240468 215818 240520 215824
rect 240926 213872 240982 213881
rect 240926 213807 240982 213816
rect 240940 213162 240968 213807
rect 240928 213156 240980 213162
rect 240928 213098 240980 213104
rect 240926 211968 240982 211977
rect 240926 211903 240982 211912
rect 240940 211734 240968 211903
rect 240928 211728 240980 211734
rect 240928 211670 240980 211676
rect 240466 209248 240522 209257
rect 240466 209183 240522 209192
rect 240480 209014 240508 209183
rect 240468 209008 240520 209014
rect 240468 208950 240520 208956
rect 258972 208946 259000 233226
rect 260352 232542 260380 235862
rect 261088 233154 261116 235862
rect 261456 233494 261484 235862
rect 262008 233562 262036 235862
rect 261996 233556 262048 233562
rect 261996 233498 262048 233504
rect 261444 233488 261496 233494
rect 261444 233430 261496 233436
rect 261076 233148 261128 233154
rect 261076 233090 261128 233096
rect 262560 233086 262588 235862
rect 263112 233222 263140 235862
rect 263100 233216 263152 233222
rect 263100 233158 263152 233164
rect 262548 233080 262600 233086
rect 262548 233022 262600 233028
rect 260340 232536 260392 232542
rect 260340 232478 260392 232484
rect 263848 224790 263876 235862
rect 264216 233737 264244 235862
rect 264202 233728 264258 233737
rect 264202 233663 264258 233672
rect 263836 224784 263888 224790
rect 263836 224726 263888 224732
rect 262364 212884 262416 212890
rect 262364 212826 262416 212832
rect 262376 212793 262404 212826
rect 261166 212784 261222 212793
rect 261166 212719 261222 212728
rect 262362 212784 262418 212793
rect 262362 212719 262418 212728
rect 258960 208940 259012 208946
rect 258960 208882 259012 208888
rect 240650 206800 240706 206809
rect 240650 206735 240706 206744
rect 240664 206226 240692 206735
rect 240652 206220 240704 206226
rect 240652 206162 240704 206168
rect 240926 204896 240982 204905
rect 240926 204831 240928 204840
rect 240980 204831 240982 204840
rect 240928 204802 240980 204808
rect 240374 202448 240430 202457
rect 240374 202383 240430 202392
rect 240388 202078 240416 202383
rect 240376 202072 240428 202078
rect 240376 202014 240428 202020
rect 240466 199864 240522 199873
rect 240466 199799 240522 199808
rect 240480 199358 240508 199799
rect 240468 199352 240520 199358
rect 240468 199294 240520 199300
rect 240926 198096 240982 198105
rect 240926 198031 240982 198040
rect 240940 197930 240968 198031
rect 240928 197924 240980 197930
rect 240928 197866 240980 197872
rect 240926 195240 240982 195249
rect 240926 195175 240928 195184
rect 240980 195175 240982 195184
rect 240928 195146 240980 195152
rect 240466 192792 240522 192801
rect 240466 192727 240522 192736
rect 240480 192490 240508 192727
rect 240468 192484 240520 192490
rect 240468 192426 240520 192432
rect 240650 190344 240706 190353
rect 240650 190279 240706 190288
rect 240664 189702 240692 190279
rect 240652 189696 240704 189702
rect 240652 189638 240704 189644
rect 240742 188304 240798 188313
rect 240742 188239 240744 188248
rect 240796 188239 240798 188248
rect 240744 188210 240796 188216
rect 240926 185856 240982 185865
rect 240926 185791 240982 185800
rect 240940 185554 240968 185791
rect 240928 185548 240980 185554
rect 240928 185490 240980 185496
rect 239638 183408 239694 183417
rect 239638 183343 239694 183352
rect 239652 179910 239680 183343
rect 243116 182822 243360 182850
rect 243484 182822 243728 182850
rect 243852 182822 244188 182850
rect 244312 182822 244464 182850
rect 244680 182822 244924 182850
rect 245048 182822 245384 182850
rect 245508 182822 245752 182850
rect 245876 182822 246120 182850
rect 246244 182822 246580 182850
rect 246704 182822 246948 182850
rect 247072 182822 247224 182850
rect 247440 182822 247776 182850
rect 247900 182822 248144 182850
rect 248268 182822 248420 182850
rect 248636 182822 248972 182850
rect 249096 182822 249340 182850
rect 249464 182822 249616 182850
rect 243332 181270 243360 182822
rect 243320 181264 243372 181270
rect 243320 181206 243372 181212
rect 243044 181196 243096 181202
rect 243044 181138 243096 181144
rect 242952 180992 243004 180998
rect 242952 180934 243004 180940
rect 242860 180924 242912 180930
rect 242860 180866 242912 180872
rect 242400 180652 242452 180658
rect 242400 180594 242452 180600
rect 239640 179904 239692 179910
rect 239640 179846 239692 179852
rect 242308 173036 242360 173042
rect 242308 172978 242360 172984
rect 241572 172492 241624 172498
rect 241572 172434 241624 172440
rect 240560 171948 240612 171954
rect 240560 171890 240612 171896
rect 239364 170044 239416 170050
rect 239364 169986 239416 169992
rect 240008 170044 240060 170050
rect 240008 169986 240060 169992
rect 239284 169902 239404 169930
rect 239376 169794 239404 169902
rect 240020 169794 240048 169986
rect 240572 169794 240600 171890
rect 241584 169794 241612 172434
rect 242320 169794 242348 172978
rect 242412 172498 242440 180594
rect 242872 173042 242900 180866
rect 242860 173036 242912 173042
rect 242860 172978 242912 172984
rect 242400 172492 242452 172498
rect 242400 172434 242452 172440
rect 242964 169794 242992 180934
rect 243056 173178 243084 181138
rect 243700 180522 243728 182822
rect 243688 180516 243740 180522
rect 243688 180458 243740 180464
rect 244160 180114 244188 182822
rect 244436 181338 244464 182822
rect 244424 181332 244476 181338
rect 244424 181274 244476 181280
rect 244896 180862 244924 182822
rect 245160 181264 245212 181270
rect 245160 181206 245212 181212
rect 244884 180856 244936 180862
rect 244884 180798 244936 180804
rect 244148 180108 244200 180114
rect 244148 180050 244200 180056
rect 243044 173172 243096 173178
rect 243044 173114 243096 173120
rect 243044 173036 243096 173042
rect 243044 172978 243096 172984
rect 236800 169766 237136 169794
rect 237260 169766 237596 169794
rect 237812 169766 238148 169794
rect 238364 169766 238700 169794
rect 239008 169766 239252 169794
rect 239376 169766 239804 169794
rect 240020 169766 240356 169794
rect 240572 169766 240908 169794
rect 241460 169766 241612 169794
rect 242012 169766 242348 169794
rect 242564 169766 242992 169794
rect 243056 169794 243084 172978
rect 245068 172628 245120 172634
rect 245068 172570 245120 172576
rect 243964 171880 244016 171886
rect 243964 171822 244016 171828
rect 243976 169794 244004 171822
rect 244424 171812 244476 171818
rect 244424 171754 244476 171760
rect 244436 169794 244464 171754
rect 245080 169794 245108 172570
rect 245172 172158 245200 181206
rect 245356 181066 245384 182822
rect 245436 181332 245488 181338
rect 245436 181274 245488 181280
rect 245344 181060 245396 181066
rect 245344 181002 245396 181008
rect 245252 180516 245304 180522
rect 245252 180458 245304 180464
rect 245264 172838 245292 180458
rect 245344 180108 245396 180114
rect 245344 180050 245396 180056
rect 245356 172974 245384 180050
rect 245344 172968 245396 172974
rect 245344 172910 245396 172916
rect 245448 172906 245476 181274
rect 245724 181270 245752 182822
rect 245712 181264 245764 181270
rect 245712 181206 245764 181212
rect 245712 181128 245764 181134
rect 245712 181070 245764 181076
rect 245436 172900 245488 172906
rect 245436 172842 245488 172848
rect 245252 172832 245304 172838
rect 245252 172774 245304 172780
rect 245160 172152 245212 172158
rect 245160 172094 245212 172100
rect 245620 171948 245672 171954
rect 245620 171890 245672 171896
rect 245632 169794 245660 171890
rect 243056 169766 243116 169794
rect 243668 169766 244004 169794
rect 244220 169766 244464 169794
rect 244772 169766 245108 169794
rect 245324 169766 245660 169794
rect 245724 169794 245752 181070
rect 245804 180584 245856 180590
rect 245804 180526 245856 180532
rect 245816 172634 245844 180526
rect 246092 180522 246120 182822
rect 246080 180516 246132 180522
rect 246080 180458 246132 180464
rect 246552 180114 246580 182822
rect 246920 180726 246948 182822
rect 247196 180794 247224 182822
rect 247184 180788 247236 180794
rect 247184 180730 247236 180736
rect 246908 180720 246960 180726
rect 246908 180662 246960 180668
rect 247184 180448 247236 180454
rect 247184 180390 247236 180396
rect 246540 180108 246592 180114
rect 246540 180050 246592 180056
rect 247196 173042 247224 180390
rect 247748 180250 247776 182822
rect 247736 180244 247788 180250
rect 247736 180186 247788 180192
rect 248116 180046 248144 182822
rect 248104 180040 248156 180046
rect 248104 179982 248156 179988
rect 248392 179978 248420 182822
rect 248944 181134 248972 182822
rect 249312 181270 249340 182822
rect 249588 181338 249616 182822
rect 249680 182822 249832 182850
rect 250292 182822 250536 182850
rect 249576 181332 249628 181338
rect 249576 181274 249628 181280
rect 249300 181264 249352 181270
rect 249300 181206 249352 181212
rect 248932 181128 248984 181134
rect 248932 181070 248984 181076
rect 249208 180516 249260 180522
rect 249208 180458 249260 180464
rect 249300 180516 249352 180522
rect 249300 180458 249352 180464
rect 248840 180176 248892 180182
rect 248840 180118 248892 180124
rect 248380 179972 248432 179978
rect 248380 179914 248432 179920
rect 248852 173042 248880 180118
rect 248932 180108 248984 180114
rect 248932 180050 248984 180056
rect 246724 173036 246776 173042
rect 246724 172978 246776 172984
rect 247184 173036 247236 173042
rect 247184 172978 247236 172984
rect 248840 173036 248892 173042
rect 248840 172978 248892 172984
rect 245804 172628 245856 172634
rect 245804 172570 245856 172576
rect 246736 169794 246764 172978
rect 248380 172764 248432 172770
rect 248380 172706 248432 172712
rect 247828 172084 247880 172090
rect 247828 172026 247880 172032
rect 247092 172016 247144 172022
rect 247092 171958 247144 171964
rect 247104 169794 247132 171958
rect 247840 169794 247868 172026
rect 248392 169794 248420 172706
rect 248564 172696 248616 172702
rect 248564 172638 248616 172644
rect 245724 169766 245876 169794
rect 246428 169766 246764 169794
rect 246980 169766 247132 169794
rect 247532 169766 247868 169794
rect 248084 169766 248420 169794
rect 248576 169794 248604 172638
rect 248944 172226 248972 180050
rect 249024 179972 249076 179978
rect 249024 179914 249076 179920
rect 248932 172220 248984 172226
rect 248932 172162 248984 172168
rect 249036 171750 249064 179914
rect 249220 172362 249248 180458
rect 249208 172356 249260 172362
rect 249208 172298 249260 172304
rect 249312 171818 249340 180458
rect 249576 180244 249628 180250
rect 249576 180186 249628 180192
rect 249392 180040 249444 180046
rect 249392 179982 249444 179988
rect 249404 172498 249432 179982
rect 249588 176306 249616 180186
rect 249576 176300 249628 176306
rect 249576 176242 249628 176248
rect 249680 176186 249708 182822
rect 250508 181406 250536 182822
rect 250600 182822 250660 182850
rect 251060 182822 251120 182850
rect 251428 182822 251488 182850
rect 251612 182822 251856 182850
rect 251980 182822 252316 182850
rect 252440 182822 252684 182850
rect 252808 182822 253052 182850
rect 253176 182822 253512 182850
rect 253728 182822 253880 182850
rect 254188 182822 254248 182850
rect 254372 182822 254708 182850
rect 254832 182822 255076 182850
rect 255200 182822 255444 182850
rect 255904 182822 255964 182850
rect 256272 182822 256332 182850
rect 250496 181400 250548 181406
rect 250496 181342 250548 181348
rect 249944 181332 249996 181338
rect 249944 181274 249996 181280
rect 249760 181060 249812 181066
rect 249760 181002 249812 181008
rect 249496 176158 249708 176186
rect 249496 172537 249524 176158
rect 249576 176096 249628 176102
rect 249576 176038 249628 176044
rect 249588 172634 249616 176038
rect 249772 175234 249800 181002
rect 249852 180380 249904 180386
rect 249852 180322 249904 180328
rect 249680 175206 249800 175234
rect 249576 172628 249628 172634
rect 249576 172570 249628 172576
rect 249482 172528 249538 172537
rect 249392 172492 249444 172498
rect 249482 172463 249538 172472
rect 249392 172434 249444 172440
rect 249680 171886 249708 175206
rect 249864 175098 249892 180322
rect 249772 175070 249892 175098
rect 249668 171880 249720 171886
rect 249668 171822 249720 171828
rect 249300 171812 249352 171818
rect 249300 171754 249352 171760
rect 249024 171744 249076 171750
rect 249024 171686 249076 171692
rect 249772 169930 249800 175070
rect 249852 173036 249904 173042
rect 249852 172978 249904 172984
rect 249496 169902 249800 169930
rect 249496 169794 249524 169902
rect 249864 169794 249892 172978
rect 249956 172809 249984 181274
rect 250600 180114 250628 182822
rect 250772 181264 250824 181270
rect 250772 181206 250824 181212
rect 250864 181264 250916 181270
rect 250864 181206 250916 181212
rect 250680 181128 250732 181134
rect 250680 181070 250732 181076
rect 250588 180108 250640 180114
rect 250588 180050 250640 180056
rect 250588 173036 250640 173042
rect 250588 172978 250640 172984
rect 249942 172800 249998 172809
rect 249942 172735 249998 172744
rect 250600 169794 250628 172978
rect 250692 172430 250720 181070
rect 250784 172566 250812 181206
rect 250772 172560 250824 172566
rect 250772 172502 250824 172508
rect 250680 172424 250732 172430
rect 250680 172366 250732 172372
rect 250876 171954 250904 181206
rect 251060 180658 251088 182822
rect 251428 181202 251456 182822
rect 251416 181196 251468 181202
rect 251416 181138 251468 181144
rect 251324 181128 251376 181134
rect 251324 181070 251376 181076
rect 251140 180788 251192 180794
rect 251140 180730 251192 180736
rect 251048 180652 251100 180658
rect 251048 180594 251100 180600
rect 250956 180108 251008 180114
rect 251008 180068 251088 180096
rect 250956 180050 251008 180056
rect 251060 172673 251088 180068
rect 251046 172664 251102 172673
rect 251046 172599 251102 172608
rect 250864 171948 250916 171954
rect 250864 171890 250916 171896
rect 251152 169794 251180 180730
rect 251232 180584 251284 180590
rect 251232 180526 251284 180532
rect 248576 169766 248636 169794
rect 249188 169766 249524 169794
rect 249740 169766 249892 169794
rect 250292 169766 250628 169794
rect 250844 169766 251180 169794
rect 251244 169794 251272 180526
rect 251336 173042 251364 181070
rect 251612 180998 251640 182822
rect 251600 180992 251652 180998
rect 251600 180934 251652 180940
rect 251980 180930 252008 182822
rect 252440 181066 252468 182822
rect 252428 181060 252480 181066
rect 252428 181002 252480 181008
rect 251968 180924 252020 180930
rect 251968 180866 252020 180872
rect 252060 180924 252112 180930
rect 252060 180866 252112 180872
rect 251324 173036 251376 173042
rect 251324 172978 251376 172984
rect 252072 172022 252100 180866
rect 252808 180522 252836 182822
rect 253176 180658 253204 182822
rect 253440 181332 253492 181338
rect 253440 181274 253492 181280
rect 253624 181332 253676 181338
rect 253624 181274 253676 181280
rect 253164 180652 253216 180658
rect 253164 180594 253216 180600
rect 252796 180516 252848 180522
rect 252796 180458 252848 180464
rect 252704 180108 252756 180114
rect 252704 180050 252756 180056
rect 252716 173042 252744 180050
rect 252152 173036 252204 173042
rect 252152 172978 252204 172984
rect 252704 173036 252756 173042
rect 252704 172978 252756 172984
rect 252060 172016 252112 172022
rect 252060 171958 252112 171964
rect 252164 169794 252192 172978
rect 253164 172968 253216 172974
rect 253164 172910 253216 172916
rect 252796 172832 252848 172838
rect 252796 172774 252848 172780
rect 252244 172152 252296 172158
rect 252244 172094 252296 172100
rect 251244 169766 251304 169794
rect 251856 169766 252192 169794
rect 252256 169794 252284 172094
rect 252808 169794 252836 172774
rect 253176 169794 253204 172910
rect 253452 172906 253480 181274
rect 253532 180244 253584 180250
rect 253532 180186 253584 180192
rect 253544 172974 253572 180186
rect 253532 172968 253584 172974
rect 253532 172910 253584 172916
rect 253440 172900 253492 172906
rect 253440 172842 253492 172848
rect 253636 172090 253664 181274
rect 253728 181270 253756 182822
rect 253716 181264 253768 181270
rect 253716 181206 253768 181212
rect 254188 180862 254216 182822
rect 254176 180856 254228 180862
rect 254176 180798 254228 180804
rect 254372 180454 254400 182822
rect 254832 180930 254860 182822
rect 255200 181338 255228 182822
rect 255188 181332 255240 181338
rect 255188 181274 255240 181280
rect 254820 180924 254872 180930
rect 254820 180866 254872 180872
rect 254360 180448 254412 180454
rect 254360 180390 254412 180396
rect 253716 180312 253768 180318
rect 253716 180254 253768 180260
rect 253728 173042 253756 180254
rect 253716 173036 253768 173042
rect 253716 172978 253768 172984
rect 254268 173036 254320 173042
rect 254268 172978 254320 172984
rect 253808 172832 253860 172838
rect 253808 172774 253860 172780
rect 253624 172084 253676 172090
rect 253624 172026 253676 172032
rect 253820 169794 253848 172774
rect 254280 169794 254308 172978
rect 254820 172968 254872 172974
rect 254820 172910 254872 172916
rect 254832 169794 254860 172910
rect 255556 172900 255608 172906
rect 255556 172842 255608 172848
rect 255568 169794 255596 172842
rect 255936 172770 255964 182822
rect 255924 172764 255976 172770
rect 255924 172706 255976 172712
rect 256304 172702 256332 182822
rect 256396 182822 256640 182850
rect 257100 182822 257160 182850
rect 256396 180386 256424 182822
rect 256384 180380 256436 180386
rect 256384 180322 256436 180328
rect 257028 180176 257080 180182
rect 257028 180118 257080 180124
rect 256936 180040 256988 180046
rect 256936 179982 256988 179988
rect 256948 175082 256976 179982
rect 256936 175076 256988 175082
rect 256936 175018 256988 175024
rect 256292 172696 256344 172702
rect 256292 172638 256344 172644
rect 255924 172356 255976 172362
rect 255924 172298 255976 172304
rect 255936 169794 255964 172298
rect 256476 172220 256528 172226
rect 256476 172162 256528 172168
rect 256488 169794 256516 172162
rect 257040 169794 257068 180118
rect 257132 179978 257160 182822
rect 257224 182822 257468 182850
rect 257592 182822 257836 182850
rect 258296 182822 258356 182850
rect 257224 181134 257252 182822
rect 257212 181128 257264 181134
rect 257212 181070 257264 181076
rect 257592 180794 257620 182822
rect 257580 180788 257632 180794
rect 257580 180730 257632 180736
rect 258328 180590 258356 182822
rect 258420 182822 258664 182850
rect 258316 180584 258368 180590
rect 258316 180526 258368 180532
rect 258420 180114 258448 182822
rect 261076 180652 261128 180658
rect 261076 180594 261128 180600
rect 258408 180108 258460 180114
rect 258408 180050 258460 180056
rect 257120 179972 257172 179978
rect 257120 179914 257172 179920
rect 261088 175234 261116 180594
rect 261180 175830 261208 212719
rect 263744 196564 263796 196570
rect 263744 196506 263796 196512
rect 262362 192792 262418 192801
rect 262362 192727 262418 192736
rect 262376 192422 262404 192727
rect 262364 192416 262416 192422
rect 262364 192358 262416 192364
rect 261168 175824 261220 175830
rect 261168 175766 261220 175772
rect 261088 175206 261944 175234
rect 257580 175076 257632 175082
rect 257580 175018 257632 175024
rect 257592 169794 257620 175018
rect 261074 172800 261130 172809
rect 261074 172735 261130 172744
rect 258316 172628 258368 172634
rect 258316 172570 258368 172576
rect 258328 169794 258356 172570
rect 260340 172560 260392 172566
rect 260340 172502 260392 172508
rect 258684 172492 258736 172498
rect 258684 172434 258736 172440
rect 258696 169794 258724 172434
rect 259788 172424 259840 172430
rect 259788 172366 259840 172372
rect 259236 172356 259288 172362
rect 259236 172298 259288 172304
rect 259248 169794 259276 172298
rect 259800 169794 259828 172366
rect 260352 169794 260380 172502
rect 261088 169794 261116 172735
rect 261442 172528 261498 172537
rect 261442 172463 261498 172472
rect 261456 169794 261484 172463
rect 261916 169794 261944 175206
rect 262546 172664 262602 172673
rect 262546 172599 262602 172608
rect 262560 169794 262588 172599
rect 263756 169794 263784 196506
rect 264202 172392 264258 172401
rect 264202 172327 264258 172336
rect 263834 172256 263890 172265
rect 263834 172191 263890 172200
rect 252256 169766 252408 169794
rect 252808 169766 252960 169794
rect 253176 169766 253512 169794
rect 253820 169766 254064 169794
rect 254280 169766 254616 169794
rect 254832 169766 255168 169794
rect 255568 169766 255720 169794
rect 255936 169766 256272 169794
rect 256488 169766 256824 169794
rect 257040 169766 257376 169794
rect 257592 169766 257928 169794
rect 258328 169766 258480 169794
rect 258696 169766 259032 169794
rect 259248 169766 259584 169794
rect 259800 169766 260136 169794
rect 260352 169766 260688 169794
rect 261088 169766 261240 169794
rect 261456 169766 261792 169794
rect 261916 169766 262344 169794
rect 262560 169766 262896 169794
rect 263448 169766 263784 169794
rect 263848 169794 263876 172191
rect 264216 169794 264244 172327
rect 263848 169766 264000 169794
rect 264216 169766 264552 169794
rect 233474 169536 233530 169545
rect 233474 169471 233530 169480
rect 233476 168888 233528 168894
rect 233474 168856 233476 168865
rect 236696 168888 236748 168894
rect 233528 168856 233530 168865
rect 236696 168830 236748 168836
rect 233474 168791 233530 168800
rect 233658 168176 233714 168185
rect 233658 168111 233714 168120
rect 233474 166952 233530 166961
rect 233474 166887 233530 166896
rect 233488 166582 233516 166887
rect 233476 166576 233528 166582
rect 233476 166518 233528 166524
rect 233474 166272 233530 166281
rect 233474 166207 233476 166216
rect 233528 166207 233530 166216
rect 233476 166178 233528 166184
rect 233566 165728 233622 165737
rect 233566 165663 233622 165672
rect 233474 165048 233530 165057
rect 233474 164983 233530 164992
rect 233488 163046 233516 164983
rect 233580 163250 233608 165663
rect 233672 164746 233700 168111
rect 236708 167573 236736 168830
rect 236694 167564 236750 167573
rect 236694 167499 236750 167508
rect 233660 164740 233712 164746
rect 233660 164682 233712 164688
rect 233750 164368 233806 164377
rect 233750 164303 233806 164312
rect 233568 163244 233620 163250
rect 233568 163186 233620 163192
rect 233566 163144 233622 163153
rect 233566 163079 233622 163088
rect 233476 163040 233528 163046
rect 233476 162982 233528 162988
rect 233474 162464 233530 162473
rect 233474 162399 233530 162408
rect 233488 162094 233516 162399
rect 233476 162088 233528 162094
rect 233476 162030 233528 162036
rect 233474 161240 233530 161249
rect 233580 161210 233608 163079
rect 233658 161920 233714 161929
rect 233658 161855 233714 161864
rect 233474 161175 233530 161184
rect 233568 161204 233620 161210
rect 233488 160530 233516 161175
rect 233568 161146 233620 161152
rect 233566 160560 233622 160569
rect 233476 160524 233528 160530
rect 233566 160495 233622 160504
rect 233476 160466 233528 160472
rect 233474 160016 233530 160025
rect 233474 159951 233530 159960
rect 233488 158966 233516 159951
rect 233580 159782 233608 160495
rect 233672 160326 233700 161855
rect 233764 161686 233792 164303
rect 233842 163824 233898 163833
rect 233842 163759 233898 163768
rect 233752 161680 233804 161686
rect 233752 161622 233804 161628
rect 233856 161550 233884 163759
rect 233844 161544 233896 161550
rect 233844 161486 233896 161492
rect 233660 160320 233712 160326
rect 233660 160262 233712 160268
rect 233568 159776 233620 159782
rect 233568 159718 233620 159724
rect 233566 159336 233622 159345
rect 233566 159271 233622 159280
rect 233476 158960 233528 158966
rect 233476 158902 233528 158908
rect 233580 158694 233608 159271
rect 233568 158688 233620 158694
rect 233474 158656 233530 158665
rect 233568 158630 233620 158636
rect 233474 158591 233530 158600
rect 233488 158286 233516 158591
rect 233476 158280 233528 158286
rect 233476 158222 233528 158228
rect 233474 158112 233530 158121
rect 233474 158047 233530 158056
rect 233488 157742 233516 158047
rect 233476 157736 233528 157742
rect 233476 157678 233528 157684
rect 233476 157464 233528 157470
rect 233474 157432 233476 157441
rect 233528 157432 233530 157441
rect 233474 157367 233530 157376
rect 233476 156988 233528 156994
rect 233476 156930 233528 156936
rect 233488 156761 233516 156930
rect 233474 156752 233530 156761
rect 233474 156687 233530 156696
rect 233476 156580 233528 156586
rect 233476 156522 233528 156528
rect 233488 156217 233516 156522
rect 233474 156208 233530 156217
rect 233474 156143 233530 156152
rect 233476 156036 233528 156042
rect 233476 155978 233528 155984
rect 233488 155537 233516 155978
rect 233568 155628 233620 155634
rect 233568 155570 233620 155576
rect 233474 155528 233530 155537
rect 233474 155463 233530 155472
rect 233476 155356 233528 155362
rect 233476 155298 233528 155304
rect 233488 154177 233516 155298
rect 233580 154857 233608 155570
rect 233566 154848 233622 154857
rect 233566 154783 233622 154792
rect 233568 154540 233620 154546
rect 233568 154482 233620 154488
rect 233474 154168 233530 154177
rect 233474 154103 233530 154112
rect 233476 153860 233528 153866
rect 233476 153802 233528 153808
rect 233488 152953 233516 153802
rect 233580 153633 233608 154482
rect 233660 154132 233712 154138
rect 233660 154074 233712 154080
rect 233566 153624 233622 153633
rect 233566 153559 233622 153568
rect 233568 153452 233620 153458
rect 233568 153394 233620 153400
rect 233474 152944 233530 152953
rect 233474 152879 233530 152888
rect 233476 152432 233528 152438
rect 233476 152374 233528 152380
rect 233488 150369 233516 152374
rect 233580 151049 233608 153394
rect 233672 152273 233700 154074
rect 233752 153792 233804 153798
rect 233752 153734 233804 153740
rect 233658 152264 233714 152273
rect 233658 152199 233714 152208
rect 233764 151729 233792 153734
rect 233844 152636 233896 152642
rect 233844 152578 233896 152584
rect 233750 151720 233806 151729
rect 233750 151655 233806 151664
rect 233566 151040 233622 151049
rect 233566 150975 233622 150984
rect 233474 150360 233530 150369
rect 233474 150295 233530 150304
rect 233856 149825 233884 152578
rect 233842 149816 233898 149825
rect 233842 149751 233898 149760
rect 233476 149576 233528 149582
rect 233476 149518 233528 149524
rect 233488 149145 233516 149518
rect 233568 149508 233620 149514
rect 233568 149450 233620 149456
rect 233474 149136 233530 149145
rect 233474 149071 233530 149080
rect 233580 148465 233608 149450
rect 233752 149100 233804 149106
rect 233752 149042 233804 149048
rect 233566 148456 233622 148465
rect 233566 148391 233622 148400
rect 233660 148352 233712 148358
rect 233660 148294 233712 148300
rect 233476 148216 233528 148222
rect 233476 148158 233528 148164
rect 233488 147921 233516 148158
rect 233568 148148 233620 148154
rect 233568 148090 233620 148096
rect 233474 147912 233530 147921
rect 233474 147847 233530 147856
rect 233580 147241 233608 148090
rect 233566 147232 233622 147241
rect 233566 147167 233622 147176
rect 233476 146720 233528 146726
rect 233476 146662 233528 146668
rect 233488 146561 233516 146662
rect 233474 146552 233530 146561
rect 233474 146487 233530 146496
rect 233476 146380 233528 146386
rect 233476 146322 233528 146328
rect 233488 146017 233516 146322
rect 233474 146008 233530 146017
rect 233474 145943 233530 145952
rect 233476 145360 233528 145366
rect 233474 145328 233476 145337
rect 233528 145328 233530 145337
rect 233474 145263 233530 145272
rect 233672 144657 233700 148294
rect 233658 144648 233714 144657
rect 233658 144583 233714 144592
rect 233764 144113 233792 149042
rect 233936 148692 233988 148698
rect 233936 148634 233988 148640
rect 233844 148284 233896 148290
rect 233844 148226 233896 148232
rect 233750 144104 233806 144113
rect 233750 144039 233806 144048
rect 233856 142753 233884 148226
rect 233948 143433 233976 148634
rect 233934 143424 233990 143433
rect 233934 143359 233990 143368
rect 233842 142744 233898 142753
rect 233476 142708 233528 142714
rect 233842 142679 233898 142688
rect 233476 142650 233528 142656
rect 233488 142209 233516 142650
rect 233474 142200 233530 142209
rect 233474 142135 233530 142144
rect 236800 141886 237136 141914
rect 237260 141886 237596 141914
rect 237812 141886 238148 141914
rect 238364 141886 238700 141914
rect 239008 141886 239252 141914
rect 239468 141886 239804 141914
rect 240020 141886 240356 141914
rect 240572 141886 240816 141914
rect 241368 141886 241704 141914
rect 241920 141886 242256 141914
rect 242472 141886 242808 141914
rect 232830 139888 232886 139897
rect 232830 139823 232886 139832
rect 231820 139308 231872 139314
rect 231820 139250 231872 139256
rect 231728 139240 231780 139246
rect 231728 139182 231780 139188
rect 231360 138900 231412 138906
rect 231360 138842 231412 138848
rect 228336 137126 228548 137154
rect 220504 135840 220556 135846
rect 220504 135782 220556 135788
rect 220516 133740 220544 135782
rect 175424 131284 175476 131290
rect 175424 131226 175476 131232
rect 167234 118808 167290 118817
rect 167234 118743 167290 118752
rect 167878 118808 167934 118817
rect 167878 118743 167934 118752
rect 145614 118264 145670 118273
rect 145614 118199 145670 118208
rect 145628 117894 145656 118199
rect 145616 117888 145668 117894
rect 145616 117830 145668 117836
rect 145614 115952 145670 115961
rect 145614 115887 145670 115896
rect 145628 115174 145656 115887
rect 145616 115168 145668 115174
rect 145616 115110 145668 115116
rect 145614 113504 145670 113513
rect 145614 113439 145670 113448
rect 145628 112386 145656 113439
rect 145616 112380 145668 112386
rect 145616 112322 145668 112328
rect 145614 111192 145670 111201
rect 145614 111127 145670 111136
rect 145628 111026 145656 111127
rect 145616 111020 145668 111026
rect 145616 110962 145668 110968
rect 145614 108880 145670 108889
rect 145614 108815 145670 108824
rect 145628 108238 145656 108815
rect 145616 108232 145668 108238
rect 145616 108174 145668 108180
rect 145614 106568 145670 106577
rect 145614 106503 145670 106512
rect 145628 105518 145656 106503
rect 145616 105512 145668 105518
rect 145616 105454 145668 105460
rect 145430 103984 145486 103993
rect 145430 103919 145486 103928
rect 145444 103138 145472 103919
rect 145432 103132 145484 103138
rect 145432 103074 145484 103080
rect 145614 101808 145670 101817
rect 145614 101743 145670 101752
rect 145628 101370 145656 101743
rect 145616 101364 145668 101370
rect 145616 101306 145668 101312
rect 145614 99496 145670 99505
rect 145614 99431 145670 99440
rect 145628 98582 145656 99431
rect 145616 98576 145668 98582
rect 145616 98518 145668 98524
rect 146350 94736 146406 94745
rect 146350 94671 146406 94680
rect 146364 94434 146392 94671
rect 146352 94428 146404 94434
rect 146352 94370 146404 94376
rect 155564 88994 155854 89010
rect 155276 88988 155328 88994
rect 155276 88930 155328 88936
rect 155552 88988 155854 88994
rect 155604 88982 155854 88988
rect 155552 88930 155604 88936
rect 149124 86886 149152 88860
rect 149112 86880 149164 86886
rect 149112 86822 149164 86828
rect 149492 86138 149520 88860
rect 149860 87090 149888 88860
rect 150320 87226 150348 88860
rect 150308 87220 150360 87226
rect 150308 87162 150360 87168
rect 149848 87084 149900 87090
rect 149848 87026 149900 87032
rect 150584 86676 150636 86682
rect 150584 86618 150636 86624
rect 149480 86132 149532 86138
rect 149480 86074 149532 86080
rect 150492 86132 150544 86138
rect 150492 86074 150544 86080
rect 145340 79400 145392 79406
rect 145340 79342 145392 79348
rect 145984 79400 146036 79406
rect 145984 79342 146036 79348
rect 145248 79060 145300 79066
rect 145248 79002 145300 79008
rect 144420 78380 144472 78386
rect 144420 78322 144472 78328
rect 142776 75790 143112 75818
rect 143236 75790 143572 75818
rect 143788 75790 144124 75818
rect 144340 75790 144676 75818
rect 145260 75682 145288 79002
rect 145432 78380 145484 78386
rect 145432 78322 145484 78328
rect 145444 75818 145472 78322
rect 145996 75818 146024 79342
rect 147640 78788 147692 78794
rect 147640 78730 147692 78736
rect 146536 78516 146588 78522
rect 146536 78458 146588 78464
rect 146548 75818 146576 78458
rect 147652 75818 147680 78730
rect 150504 78522 150532 86074
rect 150492 78516 150544 78522
rect 150492 78458 150544 78464
rect 150492 78380 150544 78386
rect 150492 78322 150544 78328
rect 149756 78312 149808 78318
rect 149756 78254 149808 78260
rect 148744 78244 148796 78250
rect 148744 78186 148796 78192
rect 148192 77972 148244 77978
rect 148192 77914 148244 77920
rect 148204 75818 148232 77914
rect 148756 75818 148784 78186
rect 149204 78176 149256 78182
rect 149204 78118 149256 78124
rect 149216 75818 149244 78118
rect 149768 75818 149796 78254
rect 150400 77904 150452 77910
rect 150400 77846 150452 77852
rect 150412 75818 150440 77846
rect 150504 76090 150532 78322
rect 150596 77910 150624 86618
rect 150688 86614 150716 88860
rect 150676 86608 150728 86614
rect 150676 86550 150728 86556
rect 151056 86478 151084 88860
rect 151320 87016 151372 87022
rect 151320 86958 151372 86964
rect 151044 86472 151096 86478
rect 151044 86414 151096 86420
rect 151332 78794 151360 86958
rect 151516 86342 151544 88860
rect 151898 88846 152004 88874
rect 151504 86336 151556 86342
rect 151504 86278 151556 86284
rect 151412 78992 151464 78998
rect 151412 78934 151464 78940
rect 151320 78788 151372 78794
rect 151320 78730 151372 78736
rect 150584 77904 150636 77910
rect 150584 77846 150636 77852
rect 150504 76062 150624 76090
rect 145444 75790 145780 75818
rect 145996 75790 146332 75818
rect 146548 75790 146792 75818
rect 147344 75790 147680 75818
rect 147896 75790 148232 75818
rect 148448 75790 148784 75818
rect 149000 75790 149244 75818
rect 149552 75790 149796 75818
rect 150104 75790 150440 75818
rect 150596 75682 150624 76062
rect 151424 75818 151452 78934
rect 151976 78658 152004 88846
rect 152252 86954 152280 88860
rect 152712 87430 152740 88860
rect 152700 87424 152752 87430
rect 152700 87366 152752 87372
rect 153080 87362 153108 88860
rect 153068 87356 153120 87362
rect 153068 87298 153120 87304
rect 152700 87288 152752 87294
rect 152700 87230 152752 87236
rect 152240 86948 152292 86954
rect 152240 86890 152292 86896
rect 151964 78652 152016 78658
rect 151964 78594 152016 78600
rect 151780 78584 151832 78590
rect 151780 78526 151832 78532
rect 151792 75818 151820 78526
rect 152712 77978 152740 87230
rect 153344 86744 153396 86750
rect 153344 86686 153396 86692
rect 153160 78108 153212 78114
rect 153160 78050 153212 78056
rect 153068 78040 153120 78046
rect 153068 77982 153120 77988
rect 152700 77972 152752 77978
rect 152700 77914 152752 77920
rect 152516 77904 152568 77910
rect 152516 77846 152568 77852
rect 152528 75818 152556 77846
rect 153080 75818 153108 77982
rect 151116 75790 151452 75818
rect 151668 75790 151820 75818
rect 152220 75790 152556 75818
rect 152772 75790 153108 75818
rect 145228 75654 145288 75682
rect 150564 75654 150624 75682
rect 153172 75682 153200 78050
rect 153356 77910 153384 86686
rect 153448 86410 153476 88860
rect 153436 86404 153488 86410
rect 153436 86346 153488 86352
rect 153908 86138 153936 88860
rect 154172 87492 154224 87498
rect 154172 87434 154224 87440
rect 154080 87152 154132 87158
rect 154080 87094 154132 87100
rect 153896 86132 153948 86138
rect 153896 86074 153948 86080
rect 153988 79060 154040 79066
rect 153988 79002 154040 79008
rect 153344 77904 153396 77910
rect 153344 77846 153396 77852
rect 154000 75818 154028 79002
rect 154092 78250 154120 87094
rect 154080 78244 154132 78250
rect 154080 78186 154132 78192
rect 154184 78182 154212 87434
rect 154276 86274 154304 88860
rect 154264 86268 154316 86274
rect 154264 86210 154316 86216
rect 154644 86206 154672 88860
rect 154632 86200 154684 86206
rect 154632 86142 154684 86148
rect 155104 86138 155132 88860
rect 155184 86540 155236 86546
rect 155184 86482 155236 86488
rect 154724 86132 154776 86138
rect 154724 86074 154776 86080
rect 155092 86132 155144 86138
rect 155092 86074 155144 86080
rect 154736 78794 154764 86074
rect 154724 78788 154776 78794
rect 154724 78730 154776 78736
rect 154172 78176 154224 78182
rect 154172 78118 154224 78124
rect 155092 78176 155144 78182
rect 155092 78118 155144 78124
rect 154632 77972 154684 77978
rect 154632 77914 154684 77920
rect 154644 75818 154672 77914
rect 155104 75818 155132 78118
rect 155196 77910 155224 86482
rect 155288 78697 155316 88930
rect 155486 88846 155776 88874
rect 155644 86744 155696 86750
rect 155644 86686 155696 86692
rect 155368 86608 155420 86614
rect 155368 86550 155420 86556
rect 155380 79338 155408 86550
rect 155552 86472 155604 86478
rect 155552 86414 155604 86420
rect 155460 86336 155512 86342
rect 155460 86278 155512 86284
rect 155368 79332 155420 79338
rect 155368 79274 155420 79280
rect 155366 79232 155422 79241
rect 155366 79167 155422 79176
rect 155274 78688 155330 78697
rect 155274 78623 155330 78632
rect 155380 78318 155408 79167
rect 155368 78312 155420 78318
rect 155368 78254 155420 78260
rect 155184 77904 155236 77910
rect 155184 77846 155236 77852
rect 155472 77842 155500 86278
rect 155564 84302 155592 86414
rect 155552 84296 155604 84302
rect 155552 84238 155604 84244
rect 155656 79354 155684 86686
rect 155748 79474 155776 88846
rect 156012 86812 156064 86818
rect 156012 86754 156064 86760
rect 155920 86608 155972 86614
rect 155920 86550 155972 86556
rect 155828 86132 155880 86138
rect 155828 86074 155880 86080
rect 155736 79468 155788 79474
rect 155736 79410 155788 79416
rect 155656 79326 155776 79354
rect 155644 79264 155696 79270
rect 155644 79206 155696 79212
rect 155656 78318 155684 79206
rect 155748 78386 155776 79326
rect 155840 78386 155868 86074
rect 155736 78380 155788 78386
rect 155736 78322 155788 78328
rect 155828 78380 155880 78386
rect 155828 78322 155880 78328
rect 155644 78312 155696 78318
rect 155644 78254 155696 78260
rect 155460 77836 155512 77842
rect 155460 77778 155512 77784
rect 155932 75954 155960 86550
rect 156024 79377 156052 86754
rect 156104 86676 156156 86682
rect 156104 86618 156156 86624
rect 156010 79368 156066 79377
rect 156010 79303 156066 79312
rect 156116 78182 156144 86618
rect 156300 86138 156328 88860
rect 156668 86546 156696 88860
rect 157128 87022 157156 88860
rect 157392 87492 157444 87498
rect 157392 87434 157444 87440
rect 157404 87106 157432 87434
rect 157496 87294 157524 88860
rect 157484 87288 157536 87294
rect 157484 87230 157536 87236
rect 157484 87152 157536 87158
rect 157404 87100 157484 87106
rect 157404 87094 157536 87100
rect 157404 87078 157524 87094
rect 157116 87016 157168 87022
rect 157116 86958 157168 86964
rect 157864 86954 157892 88860
rect 158220 87356 158272 87362
rect 158220 87298 158272 87304
rect 157852 86948 157904 86954
rect 157852 86890 157904 86896
rect 157760 86880 157812 86886
rect 157760 86822 157812 86828
rect 156656 86540 156708 86546
rect 156656 86482 156708 86488
rect 157392 86472 157444 86478
rect 157392 86414 157444 86420
rect 156656 86404 156708 86410
rect 156656 86346 156708 86352
rect 156288 86132 156340 86138
rect 156288 86074 156340 86080
rect 156668 78522 156696 86346
rect 157024 86268 157076 86274
rect 157024 86210 157076 86216
rect 157116 86268 157168 86274
rect 157116 86210 157168 86216
rect 156932 86200 156984 86206
rect 156932 86142 156984 86148
rect 156944 78862 156972 86142
rect 157036 78930 157064 86210
rect 157128 78998 157156 86210
rect 157208 86200 157260 86206
rect 157208 86142 157260 86148
rect 157116 78992 157168 78998
rect 157116 78934 157168 78940
rect 157024 78924 157076 78930
rect 157024 78866 157076 78872
rect 156932 78856 156984 78862
rect 156932 78798 156984 78804
rect 157220 78590 157248 86142
rect 157300 86132 157352 86138
rect 157300 86074 157352 86080
rect 157312 78590 157340 86074
rect 157208 78584 157260 78590
rect 157208 78526 157260 78532
rect 157300 78584 157352 78590
rect 157300 78526 157352 78532
rect 156656 78516 156708 78522
rect 156656 78458 156708 78464
rect 156104 78176 156156 78182
rect 156104 78118 156156 78124
rect 157404 77910 157432 86414
rect 157484 86404 157536 86410
rect 157484 86346 157536 86352
rect 156012 77904 156064 77910
rect 156012 77846 156064 77852
rect 156840 77904 156892 77910
rect 156840 77846 156892 77852
rect 157392 77904 157444 77910
rect 157392 77846 157444 77852
rect 155840 75926 155960 75954
rect 155840 75818 155868 75926
rect 156024 75818 156052 77846
rect 156852 75818 156880 77846
rect 157496 75954 157524 86346
rect 157668 78244 157720 78250
rect 157668 78186 157720 78192
rect 157404 75926 157524 75954
rect 157404 75818 157432 75926
rect 157680 75818 157708 78186
rect 153784 75790 154028 75818
rect 154336 75790 154672 75818
rect 154888 75790 155132 75818
rect 155440 75790 155868 75818
rect 155992 75790 156052 75818
rect 156544 75790 156880 75818
rect 157096 75790 157432 75818
rect 157556 75790 157708 75818
rect 157772 75818 157800 86822
rect 158232 78998 158260 87298
rect 158324 87158 158352 88860
rect 158404 87424 158456 87430
rect 158404 87366 158456 87372
rect 158312 87152 158364 87158
rect 158312 87094 158364 87100
rect 158312 86132 158364 86138
rect 158312 86074 158364 86080
rect 158324 79134 158352 86074
rect 158416 79202 158444 87366
rect 158692 86818 158720 88860
rect 158956 87084 159008 87090
rect 158956 87026 159008 87032
rect 158864 86880 158916 86886
rect 158864 86822 158916 86828
rect 158680 86812 158732 86818
rect 158680 86754 158732 86760
rect 158404 79196 158456 79202
rect 158404 79138 158456 79144
rect 158312 79128 158364 79134
rect 158312 79070 158364 79076
rect 158220 78992 158272 78998
rect 158220 78934 158272 78940
rect 158312 78448 158364 78454
rect 158312 78390 158364 78396
rect 158324 75818 158352 78390
rect 158876 78250 158904 86822
rect 158864 78244 158916 78250
rect 158864 78186 158916 78192
rect 158968 75818 158996 87026
rect 159060 87022 159088 88860
rect 159324 87220 159376 87226
rect 159324 87162 159376 87168
rect 159048 87016 159100 87022
rect 159048 86958 159100 86964
rect 159336 75818 159364 87162
rect 159520 86750 159548 88860
rect 159600 87424 159652 87430
rect 159600 87366 159652 87372
rect 159508 86744 159560 86750
rect 159508 86686 159560 86692
rect 159612 77910 159640 87366
rect 159784 86540 159836 86546
rect 159784 86482 159836 86488
rect 159692 86132 159744 86138
rect 159692 86074 159744 86080
rect 159704 78046 159732 86074
rect 159796 79066 159824 86482
rect 159888 86274 159916 88860
rect 159876 86268 159928 86274
rect 159876 86210 159928 86216
rect 160256 86206 160284 88860
rect 160716 87498 160744 88860
rect 160704 87492 160756 87498
rect 160704 87434 160756 87440
rect 160980 87492 161032 87498
rect 160980 87434 161032 87440
rect 160244 86200 160296 86206
rect 160244 86142 160296 86148
rect 160428 84296 160480 84302
rect 160428 84238 160480 84244
rect 159784 79060 159836 79066
rect 159784 79002 159836 79008
rect 160336 78312 160388 78318
rect 160336 78254 160388 78260
rect 159692 78040 159744 78046
rect 159692 77982 159744 77988
rect 159600 77904 159652 77910
rect 159600 77846 159652 77852
rect 160348 75818 160376 78254
rect 157772 75790 158108 75818
rect 158324 75790 158660 75818
rect 158968 75790 159212 75818
rect 159336 75790 159764 75818
rect 160316 75790 160376 75818
rect 160440 75818 160468 84238
rect 160992 78266 161020 87434
rect 161084 87430 161112 88860
rect 161072 87424 161124 87430
rect 161072 87366 161124 87372
rect 161072 87288 161124 87294
rect 161072 87230 161124 87236
rect 161084 78454 161112 87230
rect 161452 86138 161480 88860
rect 161912 87294 161940 88860
rect 162280 87498 162308 88860
rect 162268 87492 162320 87498
rect 162268 87434 162320 87440
rect 161900 87288 161952 87294
rect 161900 87230 161952 87236
rect 162648 86682 162676 88860
rect 162636 86676 162688 86682
rect 162636 86618 162688 86624
rect 163108 86614 163136 88860
rect 163096 86608 163148 86614
rect 163096 86550 163148 86556
rect 163476 86342 163504 88860
rect 163844 86478 163872 88860
rect 163832 86472 163884 86478
rect 163832 86414 163884 86420
rect 164304 86410 164332 88860
rect 164672 86886 164700 88860
rect 164660 86880 164712 86886
rect 164660 86822 164712 86828
rect 164292 86404 164344 86410
rect 164292 86346 164344 86352
rect 163464 86336 163516 86342
rect 163464 86278 163516 86284
rect 161440 86132 161492 86138
rect 161440 86074 161492 86080
rect 167248 80562 167276 118743
rect 167878 98816 167934 98825
rect 167878 98751 167934 98760
rect 167892 98582 167920 98751
rect 167880 98576 167932 98582
rect 167880 98518 167932 98524
rect 174044 81780 174096 81786
rect 174044 81722 174096 81728
rect 173768 81712 173820 81718
rect 173768 81654 173820 81660
rect 173492 81644 173544 81650
rect 173492 81586 173544 81592
rect 173308 81372 173360 81378
rect 173308 81314 173360 81320
rect 167236 80556 167288 80562
rect 167236 80498 167288 80504
rect 167248 79814 167276 80498
rect 167236 79808 167288 79814
rect 167236 79750 167288 79756
rect 170180 79808 170232 79814
rect 170180 79750 170232 79756
rect 162636 79196 162688 79202
rect 162636 79138 162688 79144
rect 162084 79128 162136 79134
rect 162084 79070 162136 79076
rect 161716 78652 161768 78658
rect 161716 78594 161768 78600
rect 161072 78448 161124 78454
rect 161072 78390 161124 78396
rect 160900 78238 161020 78266
rect 160900 77978 160928 78238
rect 160888 77972 160940 77978
rect 160888 77914 160940 77920
rect 160980 77836 161032 77842
rect 160980 77778 161032 77784
rect 160992 75818 161020 77778
rect 161728 75818 161756 78594
rect 162096 75818 162124 79070
rect 162648 75818 162676 79138
rect 167972 79060 168024 79066
rect 167972 79002 168024 79008
rect 163188 78992 163240 78998
rect 163188 78934 163240 78940
rect 163200 75818 163228 78934
rect 164752 78924 164804 78930
rect 164752 78866 164804 78872
rect 164568 78788 164620 78794
rect 164568 78730 164620 78736
rect 163740 78516 163792 78522
rect 163740 78458 163792 78464
rect 163752 75818 163780 78458
rect 164580 75818 164608 78730
rect 160440 75790 160776 75818
rect 160992 75790 161328 75818
rect 161728 75790 161880 75818
rect 162096 75790 162432 75818
rect 162648 75790 162984 75818
rect 163200 75790 163536 75818
rect 163752 75790 164088 75818
rect 164548 75790 164608 75818
rect 164764 75818 164792 78866
rect 165304 78856 165356 78862
rect 165304 78798 165356 78804
rect 165316 75818 165344 78798
rect 166408 78720 166460 78726
rect 166408 78662 166460 78668
rect 167326 78688 167382 78697
rect 165856 78380 165908 78386
rect 165856 78322 165908 78328
rect 165868 75818 165896 78322
rect 166420 75818 166448 78662
rect 167326 78623 167382 78632
rect 167340 75818 167368 78623
rect 167420 78584 167472 78590
rect 167420 78526 167472 78532
rect 164764 75790 165100 75818
rect 165316 75790 165652 75818
rect 165868 75790 166204 75818
rect 166420 75790 166756 75818
rect 167308 75790 167368 75818
rect 167432 75818 167460 78526
rect 167984 75818 168012 79002
rect 170086 78552 170142 78561
rect 170086 78487 170142 78496
rect 169074 78416 169130 78425
rect 169074 78351 169130 78360
rect 168614 77872 168670 77881
rect 168614 77807 168670 77816
rect 168628 75818 168656 77807
rect 169088 75818 169116 78351
rect 169996 76408 170048 76414
rect 169996 76350 170048 76356
rect 170008 76113 170036 76350
rect 169994 76104 170050 76113
rect 169994 76039 170050 76048
rect 170100 75818 170128 78487
rect 167432 75790 167768 75818
rect 167984 75790 168320 75818
rect 168628 75790 168872 75818
rect 169088 75790 169424 75818
rect 169976 75790 170128 75818
rect 170192 75818 170220 79750
rect 170192 75790 170528 75818
rect 153172 75654 153324 75682
rect 139634 75560 139690 75569
rect 139634 75495 139690 75504
rect 170732 75048 170784 75054
rect 170732 74990 170784 74996
rect 170640 74912 170692 74918
rect 140922 74880 140978 74889
rect 170640 74854 170692 74860
rect 140922 74815 140978 74824
rect 139634 74200 139690 74209
rect 139634 74135 139690 74144
rect 139648 73762 139676 74135
rect 138072 73756 138124 73762
rect 138072 73698 138124 73704
rect 139636 73756 139688 73762
rect 139636 73698 139688 73704
rect 136508 72464 136560 72470
rect 136508 72406 136560 72412
rect 135956 70968 136008 70974
rect 135956 70910 136008 70916
rect 135968 69546 135996 70910
rect 136416 69744 136468 69750
rect 136416 69686 136468 69692
rect 135956 69540 136008 69546
rect 135956 69482 136008 69488
rect 136428 68118 136456 69686
rect 136520 69478 136548 72406
rect 136784 72396 136836 72402
rect 136784 72338 136836 72344
rect 136600 69676 136652 69682
rect 136600 69618 136652 69624
rect 136508 69472 136560 69478
rect 136508 69414 136560 69420
rect 136508 68316 136560 68322
rect 136508 68258 136560 68264
rect 136416 68112 136468 68118
rect 136416 68054 136468 68060
rect 136520 66622 136548 68258
rect 136612 68050 136640 69618
rect 136692 69608 136744 69614
rect 136692 69550 136744 69556
rect 136600 68044 136652 68050
rect 136600 67986 136652 67992
rect 136704 67982 136732 69550
rect 136796 69410 136824 72338
rect 138084 70906 138112 73698
rect 139726 73520 139782 73529
rect 139726 73455 139782 73464
rect 139634 72976 139690 72985
rect 139634 72911 139690 72920
rect 139648 72402 139676 72911
rect 139740 72470 139768 73455
rect 139728 72464 139780 72470
rect 139728 72406 139780 72412
rect 139636 72396 139688 72402
rect 139636 72338 139688 72344
rect 139634 72296 139690 72305
rect 139634 72231 139690 72240
rect 139648 70974 139676 72231
rect 139910 71616 139966 71625
rect 139910 71551 139966 71560
rect 139636 70968 139688 70974
rect 139636 70910 139688 70916
rect 139818 70936 139874 70945
rect 138072 70900 138124 70906
rect 139818 70871 139874 70880
rect 138072 70842 138124 70848
rect 139726 70256 139782 70265
rect 139726 70191 139782 70200
rect 139634 69712 139690 69721
rect 139740 69682 139768 70191
rect 139832 69750 139860 70871
rect 139820 69744 139872 69750
rect 139820 69686 139872 69692
rect 139634 69647 139690 69656
rect 139728 69676 139780 69682
rect 139648 69614 139676 69647
rect 139728 69618 139780 69624
rect 139636 69608 139688 69614
rect 139636 69550 139688 69556
rect 136784 69404 136836 69410
rect 136784 69346 136836 69352
rect 139726 69032 139782 69041
rect 139726 68967 139782 68976
rect 139634 68352 139690 68361
rect 139740 68322 139768 68967
rect 139634 68287 139690 68296
rect 139728 68316 139780 68322
rect 139648 68254 139676 68287
rect 139728 68258 139780 68264
rect 136784 68248 136836 68254
rect 136784 68190 136836 68196
rect 139636 68248 139688 68254
rect 139636 68190 139688 68196
rect 136692 67976 136744 67982
rect 136692 67918 136744 67924
rect 136692 66820 136744 66826
rect 136692 66762 136744 66768
rect 136508 66616 136560 66622
rect 136508 66558 136560 66564
rect 136704 65262 136732 66762
rect 136796 66690 136824 68190
rect 139924 68186 139952 71551
rect 139912 68180 139964 68186
rect 139912 68122 139964 68128
rect 139634 67672 139690 67681
rect 139634 67607 139690 67616
rect 139648 66962 139676 67607
rect 139726 66992 139782 67001
rect 139636 66956 139688 66962
rect 139726 66927 139782 66936
rect 139636 66898 139688 66904
rect 139740 66826 139768 66927
rect 139728 66820 139780 66826
rect 139728 66762 139780 66768
rect 136784 66684 136836 66690
rect 136784 66626 136836 66632
rect 139726 66448 139782 66457
rect 139726 66383 139782 66392
rect 139634 65768 139690 65777
rect 139634 65703 139690 65712
rect 139648 65398 139676 65703
rect 139636 65392 139688 65398
rect 139636 65334 139688 65340
rect 139740 65330 139768 66383
rect 139728 65324 139780 65330
rect 139728 65266 139780 65272
rect 136692 65256 136744 65262
rect 136692 65198 136744 65204
rect 139726 65088 139782 65097
rect 139726 65023 139782 65032
rect 139634 64408 139690 64417
rect 139634 64343 139690 64352
rect 139648 64038 139676 64343
rect 139636 64032 139688 64038
rect 139636 63974 139688 63980
rect 139740 63970 139768 65023
rect 139728 63964 139780 63970
rect 139728 63906 139780 63912
rect 139726 63728 139782 63737
rect 139726 63663 139782 63672
rect 139636 63420 139688 63426
rect 139636 63362 139688 63368
rect 139648 63193 139676 63362
rect 139740 63358 139768 63663
rect 139728 63352 139780 63358
rect 139728 63294 139780 63300
rect 139634 63184 139690 63193
rect 139634 63119 139690 63128
rect 139726 62504 139782 62513
rect 139726 62439 139782 62448
rect 139740 61998 139768 62439
rect 139728 61992 139780 61998
rect 139728 61934 139780 61940
rect 139636 61924 139688 61930
rect 139636 61866 139688 61872
rect 139648 61833 139676 61866
rect 139634 61824 139690 61833
rect 139634 61759 139690 61768
rect 139636 61244 139688 61250
rect 139636 61186 139688 61192
rect 139648 61153 139676 61186
rect 139634 61144 139690 61153
rect 139634 61079 139690 61088
rect 139728 60632 139780 60638
rect 139634 60600 139690 60609
rect 139728 60574 139780 60580
rect 139634 60535 139636 60544
rect 139688 60535 139690 60544
rect 139636 60506 139688 60512
rect 137244 60020 137296 60026
rect 137244 59962 137296 59968
rect 137256 59278 137284 59962
rect 139740 59929 139768 60574
rect 139726 59920 139782 59929
rect 139636 59884 139688 59890
rect 139726 59855 139782 59864
rect 139636 59826 139688 59832
rect 137244 59272 137296 59278
rect 139648 59249 139676 59826
rect 139728 59272 139780 59278
rect 137244 59214 137296 59220
rect 139634 59240 139690 59249
rect 139728 59214 139780 59220
rect 139634 59175 139690 59184
rect 139740 58569 139768 59214
rect 139820 58796 139872 58802
rect 139820 58738 139872 58744
rect 139726 58560 139782 58569
rect 139636 58524 139688 58530
rect 139726 58495 139782 58504
rect 139636 58466 139688 58472
rect 139648 57889 139676 58466
rect 139728 58456 139780 58462
rect 139728 58398 139780 58404
rect 139634 57880 139690 57889
rect 139634 57815 139690 57824
rect 136232 57368 136284 57374
rect 139740 57345 139768 58398
rect 136232 57310 136284 57316
rect 139726 57336 139782 57345
rect 136244 54246 136272 57310
rect 137336 57300 137388 57306
rect 139726 57271 139782 57280
rect 137336 57242 137388 57248
rect 137348 56626 137376 57242
rect 139728 57164 139780 57170
rect 139728 57106 139780 57112
rect 137336 56620 137388 56626
rect 137336 56562 137388 56568
rect 139636 56620 139688 56626
rect 139636 56562 139688 56568
rect 139648 55985 139676 56562
rect 139634 55976 139690 55985
rect 138072 55940 138124 55946
rect 139634 55911 139690 55920
rect 138072 55882 138124 55888
rect 136784 54580 136836 54586
rect 136784 54522 136836 54528
rect 136232 54240 136284 54246
rect 136232 54182 136284 54188
rect 134760 50976 134812 50982
rect 134760 50918 134812 50924
rect 136796 50234 136824 54522
rect 138084 53974 138112 55882
rect 139452 55872 139504 55878
rect 139452 55814 139504 55820
rect 138072 53968 138124 53974
rect 138072 53910 138124 53916
rect 139464 52041 139492 55814
rect 139544 55804 139596 55810
rect 139544 55746 139596 55752
rect 139556 52721 139584 55746
rect 139740 55305 139768 57106
rect 139832 56665 139860 58738
rect 139912 57368 139964 57374
rect 139912 57310 139964 57316
rect 139818 56656 139874 56665
rect 139818 56591 139874 56600
rect 139726 55296 139782 55305
rect 139726 55231 139782 55240
rect 139924 54625 139952 57310
rect 139910 54616 139966 54625
rect 139910 54551 139966 54560
rect 139912 54512 139964 54518
rect 139912 54454 139964 54460
rect 139636 54444 139688 54450
rect 139636 54386 139688 54392
rect 139542 52712 139598 52721
rect 139542 52647 139598 52656
rect 139450 52032 139506 52041
rect 139450 51967 139506 51976
rect 139648 51361 139676 54386
rect 139728 54240 139780 54246
rect 139728 54182 139780 54188
rect 139740 54081 139768 54182
rect 139726 54072 139782 54081
rect 139726 54007 139782 54016
rect 139728 53084 139780 53090
rect 139728 53026 139780 53032
rect 139634 51352 139690 51361
rect 139634 51287 139690 51296
rect 136784 50228 136836 50234
rect 136784 50170 136836 50176
rect 139636 50228 139688 50234
rect 139636 50170 139688 50176
rect 139648 50137 139676 50170
rect 139634 50128 139690 50137
rect 139634 50063 139690 50072
rect 139740 49457 139768 53026
rect 139820 53016 139872 53022
rect 139820 52958 139872 52964
rect 139726 49448 139782 49457
rect 139726 49383 139782 49392
rect 139832 48777 139860 52958
rect 139924 50817 139952 54454
rect 140004 53968 140056 53974
rect 140004 53910 140056 53916
rect 140016 53401 140044 53910
rect 140002 53392 140058 53401
rect 140002 53327 140058 53336
rect 139910 50808 139966 50817
rect 139910 50743 139966 50752
rect 139818 48768 139874 48777
rect 139818 48703 139874 48712
rect 139634 48224 139690 48233
rect 139634 48159 139690 48168
rect 139648 47514 139676 48159
rect 139636 47508 139688 47514
rect 139636 47450 139688 47456
rect 140936 37178 140964 74815
rect 170652 74753 170680 74854
rect 170638 74744 170694 74753
rect 170638 74679 170694 74688
rect 170744 74209 170772 74990
rect 170824 74980 170876 74986
rect 170824 74922 170876 74928
rect 170836 74753 170864 74922
rect 170822 74744 170878 74753
rect 170822 74679 170878 74688
rect 170730 74200 170786 74209
rect 170730 74135 170786 74144
rect 173320 73393 173348 81314
rect 173306 73384 173362 73393
rect 173306 73319 173362 73328
rect 173504 71353 173532 81586
rect 173676 81508 173728 81514
rect 173676 81450 173728 81456
rect 173584 81304 173636 81310
rect 173584 81246 173636 81252
rect 173490 71344 173546 71353
rect 173490 71279 173546 71288
rect 173596 70265 173624 81246
rect 173688 72305 173716 81450
rect 173674 72296 173730 72305
rect 173674 72231 173730 72240
rect 173780 70809 173808 81654
rect 173860 81576 173912 81582
rect 173860 81518 173912 81524
rect 173872 71761 173900 81518
rect 173952 81440 174004 81446
rect 173952 81382 174004 81388
rect 173964 72849 173992 81382
rect 173950 72840 174006 72849
rect 173950 72775 174006 72784
rect 173858 71752 173914 71761
rect 173858 71687 173914 71696
rect 173766 70800 173822 70809
rect 173766 70735 173822 70744
rect 173582 70256 173638 70265
rect 173582 70191 173638 70200
rect 174056 69721 174084 81722
rect 174042 69712 174098 69721
rect 174042 69647 174098 69656
rect 173308 69540 173360 69546
rect 173308 69482 173360 69488
rect 173320 69177 173348 69482
rect 173306 69168 173362 69177
rect 173306 69103 173362 69112
rect 172848 68860 172900 68866
rect 172848 68802 172900 68808
rect 172860 68633 172888 68802
rect 172846 68624 172902 68633
rect 172846 68559 172902 68568
rect 174044 68180 174096 68186
rect 174044 68122 174096 68128
rect 173952 68112 174004 68118
rect 174056 68089 174084 68122
rect 173952 68054 174004 68060
rect 174042 68080 174098 68089
rect 173964 67545 173992 68054
rect 174042 68015 174098 68024
rect 173950 67536 174006 67545
rect 173492 67500 173544 67506
rect 173950 67471 174006 67480
rect 173492 67442 173544 67448
rect 173504 67001 173532 67442
rect 173490 66992 173546 67001
rect 173490 66927 173546 66936
rect 173860 66752 173912 66758
rect 173860 66694 173912 66700
rect 173584 66684 173636 66690
rect 173584 66626 173636 66632
rect 173596 66049 173624 66626
rect 173582 66040 173638 66049
rect 173582 65975 173638 65984
rect 173872 65505 173900 66694
rect 174044 66616 174096 66622
rect 174042 66584 174044 66593
rect 174096 66584 174098 66593
rect 174042 66519 174098 66528
rect 173858 65496 173914 65505
rect 173858 65431 173914 65440
rect 173492 65392 173544 65398
rect 173492 65334 173544 65340
rect 173504 64961 173532 65334
rect 173768 65324 173820 65330
rect 173768 65266 173820 65272
rect 173490 64952 173546 64961
rect 173490 64887 173546 64896
rect 173780 64417 173808 65266
rect 173766 64408 173822 64417
rect 173766 64343 173822 64352
rect 173860 64032 173912 64038
rect 173860 63974 173912 63980
rect 173872 63329 173900 63974
rect 173952 63964 174004 63970
rect 173952 63906 174004 63912
rect 173858 63320 173914 63329
rect 173858 63255 173914 63264
rect 173964 62785 173992 63906
rect 174044 63896 174096 63902
rect 174042 63864 174044 63873
rect 174096 63864 174098 63873
rect 174042 63799 174098 63808
rect 173950 62776 174006 62785
rect 173950 62711 174006 62720
rect 173768 62604 173820 62610
rect 173768 62546 173820 62552
rect 173308 62536 173360 62542
rect 173308 62478 173360 62484
rect 173320 62241 173348 62478
rect 173306 62232 173362 62241
rect 173306 62167 173362 62176
rect 173780 61833 173808 62546
rect 173766 61824 173822 61833
rect 173766 61759 173822 61768
rect 173950 61280 174006 61289
rect 173676 61244 173728 61250
rect 173950 61215 174006 61224
rect 173676 61186 173728 61192
rect 173688 60201 173716 61186
rect 173964 61114 173992 61215
rect 174044 61176 174096 61182
rect 174044 61118 174096 61124
rect 173952 61108 174004 61114
rect 173952 61050 174004 61056
rect 174056 60745 174084 61118
rect 174042 60736 174098 60745
rect 174042 60671 174098 60680
rect 173674 60192 173730 60201
rect 173674 60127 173730 60136
rect 173860 59884 173912 59890
rect 173860 59826 173912 59832
rect 173676 59816 173728 59822
rect 173676 59758 173728 59764
rect 173688 59113 173716 59758
rect 173674 59104 173730 59113
rect 173674 59039 173730 59048
rect 173872 58569 173900 59826
rect 174044 59748 174096 59754
rect 174044 59690 174096 59696
rect 174056 59657 174084 59690
rect 174042 59648 174098 59657
rect 174042 59583 174098 59592
rect 173858 58560 173914 58569
rect 173768 58524 173820 58530
rect 173858 58495 173914 58504
rect 173768 58466 173820 58472
rect 173780 57481 173808 58466
rect 174044 58456 174096 58462
rect 174044 58398 174096 58404
rect 174056 58025 174084 58398
rect 174042 58016 174098 58025
rect 174042 57951 174098 57960
rect 173766 57472 173822 57481
rect 173766 57407 173822 57416
rect 172940 57096 172992 57102
rect 172940 57038 172992 57044
rect 174042 57064 174098 57073
rect 172952 55985 172980 57038
rect 174042 56999 174044 57008
rect 174096 56999 174098 57008
rect 174044 56970 174096 56976
rect 174044 56824 174096 56830
rect 174044 56766 174096 56772
rect 174056 56529 174084 56766
rect 174042 56520 174098 56529
rect 174042 56455 174098 56464
rect 172938 55976 172994 55985
rect 172938 55911 172994 55920
rect 173308 55736 173360 55742
rect 173308 55678 173360 55684
rect 173320 55441 173348 55678
rect 173768 55668 173820 55674
rect 173768 55610 173820 55616
rect 173306 55432 173362 55441
rect 173306 55367 173362 55376
rect 173780 54897 173808 55610
rect 173766 54888 173822 54897
rect 173766 54823 173822 54832
rect 175240 54512 175292 54518
rect 175240 54454 175292 54460
rect 174044 54376 174096 54382
rect 174042 54344 174044 54353
rect 174096 54344 174098 54353
rect 174042 54279 174098 54288
rect 174044 53832 174096 53838
rect 174042 53800 174044 53809
rect 174096 53800 174098 53809
rect 173492 53764 173544 53770
rect 174042 53735 174098 53744
rect 173492 53706 173544 53712
rect 173504 53265 173532 53706
rect 173490 53256 173546 53265
rect 173490 53191 173546 53200
rect 172848 52948 172900 52954
rect 172848 52890 172900 52896
rect 172860 51769 172888 52890
rect 174044 52880 174096 52886
rect 174044 52822 174096 52828
rect 173952 52744 174004 52750
rect 173950 52712 173952 52721
rect 174004 52712 174006 52721
rect 173950 52647 174006 52656
rect 174056 52313 174084 52822
rect 174042 52304 174098 52313
rect 174042 52239 174098 52248
rect 172846 51760 172902 51769
rect 172846 51695 172902 51704
rect 173952 51588 174004 51594
rect 173952 51530 174004 51536
rect 172940 51248 172992 51254
rect 172938 51216 172940 51225
rect 172992 51216 172994 51225
rect 172938 51151 172994 51160
rect 173964 50681 173992 51530
rect 173950 50672 174006 50681
rect 173950 50607 174006 50616
rect 175252 50166 175280 54454
rect 175332 54444 175384 54450
rect 175332 54386 175384 54392
rect 173308 50160 173360 50166
rect 173306 50128 173308 50137
rect 175240 50160 175292 50166
rect 173360 50128 173362 50137
rect 172756 50092 172808 50098
rect 175240 50102 175292 50108
rect 175344 50098 175372 54386
rect 173306 50063 173362 50072
rect 175332 50092 175384 50098
rect 172756 50034 172808 50040
rect 175332 50034 175384 50040
rect 172768 49593 172796 50034
rect 172754 49584 172810 49593
rect 172754 49519 172810 49528
rect 173124 49208 173176 49214
rect 173124 49150 173176 49156
rect 173136 49049 173164 49150
rect 173122 49040 173178 49049
rect 173122 48975 173178 48984
rect 173308 48664 173360 48670
rect 173308 48606 173360 48612
rect 173320 48505 173348 48606
rect 173306 48496 173362 48505
rect 173306 48431 173362 48440
rect 173398 48088 173454 48097
rect 173398 48023 173454 48032
rect 156576 47910 156912 47938
rect 156576 46057 156604 47910
rect 156562 46048 156618 46057
rect 156562 45983 156618 45992
rect 173412 37246 173440 48023
rect 173400 37240 173452 37246
rect 173400 37182 173452 37188
rect 140924 37172 140976 37178
rect 140924 37114 140976 37120
rect 138440 12488 138492 12494
rect 138440 12430 138492 12436
rect 133380 12420 133432 12426
rect 133380 12362 133432 12368
rect 88484 12352 88536 12358
rect 88484 12294 88536 12300
rect 64932 12284 64984 12290
rect 64932 12226 64984 12232
rect 64944 9304 64972 12226
rect 101730 12184 101786 12193
rect 101730 12119 101786 12128
rect 101744 9304 101772 12119
rect 138452 9304 138480 12430
rect 175436 9434 175464 131226
rect 228520 127618 228548 137126
rect 230714 127920 230770 127929
rect 230714 127855 230770 127864
rect 228508 127612 228560 127618
rect 228508 127554 228560 127560
rect 230728 127550 230756 127855
rect 230716 127544 230768 127550
rect 230716 127486 230768 127492
rect 228416 127476 228468 127482
rect 228416 127418 228468 127424
rect 228428 124762 228456 127418
rect 228416 124756 228468 124762
rect 228416 124698 228468 124704
rect 175516 121968 175568 121974
rect 175514 121936 175516 121945
rect 175568 121936 175570 121945
rect 175514 121871 175570 121880
rect 228508 120540 228560 120546
rect 228508 120482 228560 120488
rect 228520 120313 228548 120482
rect 228506 120304 228562 120313
rect 228506 120239 228562 120248
rect 228520 108238 228548 120239
rect 231266 115272 231322 115281
rect 231266 115207 231268 115216
rect 231320 115207 231322 115216
rect 231268 115178 231320 115184
rect 231372 114873 231400 138842
rect 231636 138832 231688 138838
rect 231636 138774 231688 138780
rect 231544 138764 231596 138770
rect 231544 138706 231596 138712
rect 231452 138696 231504 138702
rect 231452 138638 231504 138644
rect 231358 114864 231414 114873
rect 231358 114799 231414 114808
rect 231358 112416 231414 112425
rect 231268 112380 231320 112386
rect 231358 112351 231414 112360
rect 231268 112322 231320 112328
rect 228508 108232 228560 108238
rect 228508 108174 228560 108180
rect 228508 108096 228560 108102
rect 228508 108038 228560 108044
rect 175516 98576 175568 98582
rect 175516 98518 175568 98524
rect 175528 97057 175556 98518
rect 175514 97048 175570 97057
rect 175514 96983 175570 96992
rect 228520 95794 228548 108038
rect 231280 100865 231308 112322
rect 231266 100856 231322 100865
rect 231266 100791 231322 100800
rect 228508 95788 228560 95794
rect 228508 95730 228560 95736
rect 228508 90892 228560 90898
rect 228508 90834 228560 90840
rect 228520 84114 228548 90834
rect 228166 84100 228548 84114
rect 228152 84086 228548 84100
rect 179576 81990 179604 83828
rect 179564 81984 179616 81990
rect 179564 81926 179616 81932
rect 180864 80630 180892 83828
rect 182140 83820 182192 83826
rect 182140 83762 182192 83768
rect 182152 83729 182180 83762
rect 182138 83720 182194 83729
rect 182138 83655 182194 83664
rect 182244 80698 182272 83828
rect 183624 83706 183652 83828
rect 183624 83678 183744 83706
rect 182232 80692 182284 80698
rect 182232 80634 182284 80640
rect 180852 80624 180904 80630
rect 180852 80566 180904 80572
rect 183060 80624 183112 80630
rect 183060 80566 183112 80572
rect 183072 72402 183100 80566
rect 183716 73694 183744 83678
rect 184912 80630 184940 83828
rect 186292 81990 186320 83828
rect 186280 81984 186332 81990
rect 186280 81926 186332 81932
rect 187672 81242 187700 83828
rect 187660 81236 187712 81242
rect 187660 81178 187712 81184
rect 188960 81174 188988 83828
rect 190340 81530 190368 83828
rect 191720 81530 191748 83828
rect 190340 81502 190644 81530
rect 191720 81502 192024 81530
rect 188948 81168 189000 81174
rect 188948 81110 189000 81116
rect 185820 80692 185872 80698
rect 185820 80634 185872 80640
rect 184900 80624 184952 80630
rect 184900 80566 184952 80572
rect 183704 73688 183756 73694
rect 183704 73630 183756 73636
rect 185832 72402 185860 80634
rect 190616 73694 190644 81502
rect 191340 80624 191392 80630
rect 191340 80566 191392 80572
rect 190144 73688 190196 73694
rect 190144 73630 190196 73636
rect 190604 73688 190656 73694
rect 190604 73630 190656 73636
rect 183060 72396 183112 72402
rect 183060 72338 183112 72344
rect 184716 72396 184768 72402
rect 184716 72338 184768 72344
rect 185820 72396 185872 72402
rect 185820 72338 185872 72344
rect 187660 72396 187712 72402
rect 187660 72338 187712 72344
rect 181770 69712 181826 69721
rect 184728 69698 184756 72338
rect 187672 69834 187700 72338
rect 190156 69834 190184 73630
rect 191352 72402 191380 80566
rect 191996 73490 192024 81502
rect 193008 79354 193036 83828
rect 194100 81984 194152 81990
rect 194100 81926 194152 81932
rect 193008 79326 193404 79354
rect 191984 73484 192036 73490
rect 191984 73426 192036 73432
rect 193376 73422 193404 79326
rect 193364 73416 193416 73422
rect 193364 73358 193416 73364
rect 194112 72402 194140 81926
rect 194388 79490 194416 83828
rect 195768 81530 195796 83828
rect 197056 81786 197084 83828
rect 198436 81786 198464 83828
rect 199816 81786 199844 83828
rect 201104 81786 201132 83828
rect 197044 81780 197096 81786
rect 197044 81722 197096 81728
rect 197504 81780 197556 81786
rect 197504 81722 197556 81728
rect 198424 81780 198476 81786
rect 198424 81722 198476 81728
rect 198884 81780 198936 81786
rect 198884 81722 198936 81728
rect 199804 81780 199856 81786
rect 199804 81722 199856 81728
rect 200264 81780 200316 81786
rect 200264 81722 200316 81728
rect 201092 81780 201144 81786
rect 201092 81722 201144 81728
rect 201644 81780 201696 81786
rect 201644 81722 201696 81728
rect 195768 81502 196164 81530
rect 195572 81236 195624 81242
rect 195572 81178 195624 81184
rect 195480 81168 195532 81174
rect 195480 81110 195532 81116
rect 194388 79462 194784 79490
rect 194756 73354 194784 79462
rect 194744 73348 194796 73354
rect 194744 73290 194796 73296
rect 195492 72470 195520 81110
rect 195480 72464 195532 72470
rect 195480 72406 195532 72412
rect 195584 72402 195612 81178
rect 196136 73286 196164 81502
rect 196124 73280 196176 73286
rect 196124 73222 196176 73228
rect 197516 73218 197544 81722
rect 197504 73212 197556 73218
rect 197504 73154 197556 73160
rect 198896 73150 198924 81722
rect 198884 73144 198936 73150
rect 198884 73086 198936 73092
rect 200276 73082 200304 81722
rect 200264 73076 200316 73082
rect 200264 73018 200316 73024
rect 201656 73014 201684 81722
rect 202484 81281 202512 83828
rect 203864 81990 203892 83828
rect 203852 81984 203904 81990
rect 203852 81926 203904 81932
rect 202470 81272 202526 81281
rect 202470 81207 202526 81216
rect 205152 75054 205180 83828
rect 206532 81310 206560 83828
rect 207912 81310 207940 83828
rect 209200 81718 209228 83828
rect 209188 81712 209240 81718
rect 209188 81654 209240 81660
rect 210580 81417 210608 83828
rect 211960 81650 211988 83828
rect 211948 81644 212000 81650
rect 211948 81586 212000 81592
rect 210566 81408 210622 81417
rect 210566 81343 210622 81352
rect 206520 81304 206572 81310
rect 206520 81246 206572 81252
rect 207900 81304 207952 81310
rect 207900 81246 207952 81252
rect 205140 75048 205192 75054
rect 205140 74990 205192 74996
rect 213248 74986 213276 83828
rect 214628 81582 214656 83828
rect 214616 81576 214668 81582
rect 214616 81518 214668 81524
rect 213236 74980 213288 74986
rect 213236 74922 213288 74928
rect 216008 74918 216036 83828
rect 217296 81514 217324 83828
rect 217284 81508 217336 81514
rect 217284 81450 217336 81456
rect 218676 76414 218704 83828
rect 220056 81446 220084 83828
rect 221344 81446 221372 83828
rect 220044 81440 220096 81446
rect 220044 81382 220096 81388
rect 221332 81440 221384 81446
rect 221332 81382 221384 81388
rect 222724 81378 222752 83828
rect 226772 81922 226800 83828
rect 226760 81916 226812 81922
rect 226760 81858 226812 81864
rect 222712 81372 222764 81378
rect 222712 81314 222764 81320
rect 218664 76408 218716 76414
rect 218664 76350 218716 76356
rect 215996 74912 216048 74918
rect 215996 74854 216048 74860
rect 202656 73552 202708 73558
rect 202656 73494 202708 73500
rect 201644 73008 201696 73014
rect 201644 72950 201696 72956
rect 200172 72464 200224 72470
rect 200172 72406 200224 72412
rect 191340 72396 191392 72402
rect 191340 72338 191392 72344
rect 192628 72396 192680 72402
rect 192628 72338 192680 72344
rect 194100 72396 194152 72402
rect 194100 72338 194152 72344
rect 195112 72396 195164 72402
rect 195112 72338 195164 72344
rect 195572 72396 195624 72402
rect 195572 72338 195624 72344
rect 197504 72396 197556 72402
rect 197504 72338 197556 72344
rect 192640 69834 192668 72338
rect 195124 69834 195152 72338
rect 197516 69970 197544 72338
rect 197516 69942 197636 69970
rect 197608 69834 197636 69942
rect 200184 69834 200212 72406
rect 202668 69834 202696 73494
rect 205140 73484 205192 73490
rect 205140 73426 205192 73432
rect 205152 69834 205180 73426
rect 207624 73416 207676 73422
rect 207624 73358 207676 73364
rect 207636 69834 207664 73358
rect 210108 73348 210160 73354
rect 210108 73290 210160 73296
rect 210120 69834 210148 73290
rect 212684 73280 212736 73286
rect 212684 73222 212736 73228
rect 212696 69834 212724 73222
rect 215168 73212 215220 73218
rect 215168 73154 215220 73160
rect 215180 69834 215208 73154
rect 217652 73144 217704 73150
rect 217652 73086 217704 73092
rect 217664 69834 217692 73086
rect 220136 73076 220188 73082
rect 220136 73018 220188 73024
rect 220148 69834 220176 73018
rect 222620 73008 222672 73014
rect 222620 72950 222672 72956
rect 222632 69834 222660 72950
rect 226024 70900 226076 70906
rect 226024 70842 226076 70848
rect 187594 69806 187700 69834
rect 190078 69806 190184 69834
rect 192562 69806 192668 69834
rect 195046 69806 195152 69834
rect 197530 69806 197636 69834
rect 200106 69806 200212 69834
rect 202590 69806 202696 69834
rect 205074 69806 205180 69834
rect 207558 69806 207664 69834
rect 210042 69806 210148 69834
rect 212618 69806 212724 69834
rect 215102 69806 215208 69834
rect 217586 69806 217692 69834
rect 220070 69806 220176 69834
rect 222554 69806 222660 69834
rect 226036 69721 226064 70842
rect 226022 69712 226078 69721
rect 184728 69670 185110 69698
rect 181770 69647 181826 69656
rect 226022 69647 226078 69656
rect 181784 69546 181812 69647
rect 181772 69540 181824 69546
rect 181772 69482 181824 69488
rect 226024 69540 226076 69546
rect 226024 69482 226076 69488
rect 225748 69472 225800 69478
rect 225748 69414 225800 69420
rect 182322 69032 182378 69041
rect 182322 68967 182378 68976
rect 182336 68866 182364 68967
rect 225760 68905 225788 69414
rect 226036 69313 226064 69482
rect 226022 69304 226078 69313
rect 226022 69239 226078 69248
rect 225746 68896 225802 68905
rect 182324 68860 182376 68866
rect 225746 68831 225802 68840
rect 182324 68802 182376 68808
rect 226300 68792 226352 68798
rect 226300 68734 226352 68740
rect 181770 68624 181826 68633
rect 181770 68559 181826 68568
rect 181586 68216 181642 68225
rect 181784 68186 181812 68559
rect 226312 68497 226340 68734
rect 226298 68488 226354 68497
rect 226298 68423 226354 68432
rect 181586 68151 181642 68160
rect 181772 68180 181824 68186
rect 181600 68118 181628 68151
rect 181772 68122 181824 68128
rect 225472 68180 225524 68186
rect 225472 68122 225524 68128
rect 181588 68112 181640 68118
rect 181588 68054 181640 68060
rect 182322 67808 182378 67817
rect 182322 67743 182378 67752
rect 182336 67506 182364 67743
rect 182324 67500 182376 67506
rect 182324 67442 182376 67448
rect 182230 67400 182286 67409
rect 182230 67335 182286 67344
rect 181402 66856 181458 66865
rect 181402 66791 181458 66800
rect 181416 66758 181444 66791
rect 181404 66752 181456 66758
rect 181404 66694 181456 66700
rect 182244 66622 182272 67335
rect 225484 67273 225512 68122
rect 225564 68112 225616 68118
rect 225564 68054 225616 68060
rect 226298 68080 226354 68089
rect 225576 67681 225604 68054
rect 225840 68044 225892 68050
rect 226298 68015 226354 68024
rect 225840 67986 225892 67992
rect 225562 67672 225618 67681
rect 225562 67607 225618 67616
rect 225470 67264 225526 67273
rect 225470 67199 225526 67208
rect 182322 66992 182378 67001
rect 182322 66927 182378 66936
rect 182336 66690 182364 66927
rect 225852 66865 225880 67986
rect 226312 67982 226340 68015
rect 226300 67976 226352 67982
rect 226300 67918 226352 67924
rect 225838 66856 225894 66865
rect 225838 66791 225894 66800
rect 226300 66752 226352 66758
rect 226300 66694 226352 66700
rect 182324 66684 182376 66690
rect 182324 66626 182376 66632
rect 226024 66684 226076 66690
rect 226024 66626 226076 66632
rect 182232 66616 182284 66622
rect 182232 66558 182284 66564
rect 226036 66457 226064 66626
rect 226022 66448 226078 66457
rect 226022 66383 226078 66392
rect 182322 66176 182378 66185
rect 182322 66111 182378 66120
rect 181402 65768 181458 65777
rect 181402 65703 181458 65712
rect 181310 65632 181366 65641
rect 181310 65567 181366 65576
rect 181034 64952 181090 64961
rect 181034 64887 181090 64896
rect 181048 64038 181076 64887
rect 181126 64544 181182 64553
rect 181126 64479 181182 64488
rect 181036 64032 181088 64038
rect 181036 63974 181088 63980
rect 181140 63970 181168 64479
rect 181128 63964 181180 63970
rect 181128 63906 181180 63912
rect 181324 63902 181352 65567
rect 181416 65330 181444 65703
rect 182336 65398 182364 66111
rect 226312 66049 226340 66694
rect 226392 66072 226444 66078
rect 226298 66040 226354 66049
rect 226392 66014 226444 66020
rect 226298 65975 226354 65984
rect 226404 65641 226432 66014
rect 226390 65632 226446 65641
rect 226390 65567 226446 65576
rect 182324 65392 182376 65398
rect 182324 65334 182376 65340
rect 226300 65392 226352 65398
rect 226300 65334 226352 65340
rect 181404 65324 181456 65330
rect 181404 65266 181456 65272
rect 226312 65233 226340 65334
rect 226298 65224 226354 65233
rect 226298 65159 226354 65168
rect 226298 64816 226354 64825
rect 226298 64751 226300 64760
rect 226352 64751 226354 64760
rect 226300 64722 226352 64728
rect 226392 64712 226444 64718
rect 226392 64654 226444 64660
rect 226404 64417 226432 64654
rect 181402 64408 181458 64417
rect 181402 64343 181458 64352
rect 226390 64408 226446 64417
rect 226390 64343 226446 64352
rect 181312 63896 181364 63902
rect 181312 63838 181364 63844
rect 181416 62542 181444 64343
rect 226390 64000 226446 64009
rect 226390 63935 226446 63944
rect 182322 63728 182378 63737
rect 182322 63663 182378 63672
rect 182046 63320 182102 63329
rect 182046 63255 182102 63264
rect 181404 62536 181456 62542
rect 181404 62478 181456 62484
rect 181770 62368 181826 62377
rect 181770 62303 181826 62312
rect 181678 61008 181734 61017
rect 181678 60943 181734 60952
rect 176896 60020 176948 60026
rect 176896 59962 176948 59968
rect 176908 57034 176936 59962
rect 176988 59952 177040 59958
rect 176988 59894 177040 59900
rect 176896 57028 176948 57034
rect 176896 56970 176948 56976
rect 177000 56830 177028 59894
rect 180942 59648 180998 59657
rect 180942 59583 180998 59592
rect 180298 57744 180354 57753
rect 178000 57708 178052 57714
rect 180298 57679 180354 57688
rect 178000 57650 178052 57656
rect 177632 57572 177684 57578
rect 177632 57514 177684 57520
rect 176988 56824 177040 56830
rect 176988 56766 177040 56772
rect 177356 55804 177408 55810
rect 177356 55746 177408 55752
rect 176896 53016 176948 53022
rect 176896 52958 176948 52964
rect 176908 49214 176936 52958
rect 177368 51254 177396 55746
rect 177644 53838 177672 57514
rect 177724 57300 177776 57306
rect 177724 57242 177776 57248
rect 177632 53832 177684 53838
rect 177632 53774 177684 53780
rect 177736 53770 177764 57242
rect 178012 54382 178040 57650
rect 178000 54376 178052 54382
rect 178000 54318 178052 54324
rect 177724 53764 177776 53770
rect 177724 53706 177776 53712
rect 180312 52750 180340 57679
rect 180956 57102 180984 59583
rect 181692 58462 181720 60943
rect 181784 59754 181812 62303
rect 181862 61824 181918 61833
rect 181862 61759 181918 61768
rect 181876 59822 181904 61759
rect 181954 61416 182010 61425
rect 181954 61351 182010 61360
rect 181968 59890 181996 61351
rect 182060 61114 182088 63255
rect 182138 62912 182194 62921
rect 182138 62847 182194 62856
rect 182152 61182 182180 62847
rect 182230 62776 182286 62785
rect 182230 62711 182286 62720
rect 182244 61250 182272 62711
rect 182336 62610 182364 63663
rect 226298 63592 226354 63601
rect 226298 63527 226354 63536
rect 226312 63494 226340 63527
rect 226300 63488 226352 63494
rect 226300 63430 226352 63436
rect 226404 63426 226432 63935
rect 226392 63420 226444 63426
rect 226392 63362 226444 63368
rect 226300 63352 226352 63358
rect 226300 63294 226352 63300
rect 226312 63193 226340 63294
rect 226298 63184 226354 63193
rect 226298 63119 226354 63128
rect 226298 62776 226354 62785
rect 226298 62711 226354 62720
rect 226312 62678 226340 62711
rect 226300 62672 226352 62678
rect 226300 62614 226352 62620
rect 182324 62604 182376 62610
rect 182324 62546 182376 62552
rect 226390 62368 226446 62377
rect 226390 62303 226446 62312
rect 226206 62096 226262 62105
rect 226206 62031 226262 62040
rect 226220 61386 226248 62031
rect 226404 61930 226432 62303
rect 226392 61924 226444 61930
rect 226392 61866 226444 61872
rect 226298 61688 226354 61697
rect 226298 61623 226354 61632
rect 226208 61380 226260 61386
rect 226208 61322 226260 61328
rect 226312 61318 226340 61623
rect 226300 61312 226352 61318
rect 225746 61280 225802 61289
rect 182232 61244 182284 61250
rect 226300 61254 226352 61260
rect 225746 61215 225802 61224
rect 182232 61186 182284 61192
rect 182140 61176 182192 61182
rect 182140 61118 182192 61124
rect 182048 61108 182100 61114
rect 182048 61050 182100 61056
rect 182138 60600 182194 60609
rect 182138 60535 182194 60544
rect 181956 59884 182008 59890
rect 181956 59826 182008 59832
rect 181864 59816 181916 59822
rect 181864 59758 181916 59764
rect 181772 59748 181824 59754
rect 181772 59690 181824 59696
rect 182046 58560 182102 58569
rect 182152 58530 182180 60535
rect 182230 60192 182286 60201
rect 182230 60127 182286 60136
rect 182244 60026 182272 60127
rect 182322 60056 182378 60065
rect 182232 60020 182284 60026
rect 225760 60026 225788 61215
rect 225930 60872 225986 60881
rect 225930 60807 225986 60816
rect 182322 59991 182378 60000
rect 225748 60020 225800 60026
rect 182232 59962 182284 59968
rect 182336 59958 182364 59991
rect 225748 59962 225800 59968
rect 225944 59958 225972 60807
rect 226390 60464 226446 60473
rect 226390 60399 226446 60408
rect 226404 60162 226432 60399
rect 226392 60156 226444 60162
rect 226392 60098 226444 60104
rect 226300 60088 226352 60094
rect 226298 60056 226300 60065
rect 226352 60056 226354 60065
rect 226298 59991 226354 60000
rect 182324 59952 182376 59958
rect 182324 59894 182376 59900
rect 225932 59952 225984 59958
rect 225932 59894 225984 59900
rect 226206 59648 226262 59657
rect 226206 59583 226262 59592
rect 182230 58968 182286 58977
rect 182230 58903 182286 58912
rect 182046 58495 182102 58504
rect 182140 58524 182192 58530
rect 181680 58456 181732 58462
rect 181680 58398 181732 58404
rect 181678 57744 181734 57753
rect 181678 57679 181734 57688
rect 181692 57578 181720 57679
rect 181680 57572 181732 57578
rect 181680 57514 181732 57520
rect 181586 57336 181642 57345
rect 181586 57271 181588 57280
rect 181640 57271 181642 57280
rect 181588 57242 181640 57248
rect 180944 57096 180996 57102
rect 180944 57038 180996 57044
rect 181310 56520 181366 56529
rect 181310 56455 181366 56464
rect 181218 56112 181274 56121
rect 181218 56047 181274 56056
rect 181126 55296 181182 55305
rect 181126 55231 181182 55240
rect 180942 53120 180998 53129
rect 180942 53055 180998 53064
rect 180300 52744 180352 52750
rect 180300 52686 180352 52692
rect 177356 51248 177408 51254
rect 177356 51190 177408 51196
rect 176896 49208 176948 49214
rect 176896 49150 176948 49156
rect 180956 48670 180984 53055
rect 181140 51594 181168 55231
rect 181232 52954 181260 56047
rect 181220 52948 181272 52954
rect 181220 52890 181272 52896
rect 181324 52886 181352 56455
rect 182060 55674 182088 58495
rect 182140 58466 182192 58472
rect 182244 55742 182272 58903
rect 226220 58734 226248 59583
rect 226390 59240 226446 59249
rect 226390 59175 226446 59184
rect 226298 58832 226354 58841
rect 226298 58767 226354 58776
rect 226208 58728 226260 58734
rect 226208 58670 226260 58676
rect 226312 58598 226340 58767
rect 226404 58666 226432 59175
rect 226392 58660 226444 58666
rect 226392 58602 226444 58608
rect 226300 58592 226352 58598
rect 226300 58534 226352 58540
rect 225746 58424 225802 58433
rect 225746 58359 225802 58368
rect 182322 58152 182378 58161
rect 182322 58087 182378 58096
rect 182336 57714 182364 58087
rect 182324 57708 182376 57714
rect 182324 57650 182376 57656
rect 183702 57472 183758 57481
rect 183702 57407 183758 57416
rect 183716 57141 183744 57407
rect 225760 57374 225788 58359
rect 225930 58016 225986 58025
rect 225930 57951 225986 57960
rect 225838 57608 225894 57617
rect 225838 57543 225894 57552
rect 225748 57368 225800 57374
rect 225748 57310 225800 57316
rect 225852 57306 225880 57543
rect 225840 57300 225892 57306
rect 225840 57242 225892 57248
rect 225944 57170 225972 57951
rect 228048 57368 228100 57374
rect 228048 57310 228100 57316
rect 226484 57232 226536 57238
rect 226482 57200 226484 57209
rect 226536 57200 226538 57209
rect 225932 57164 225984 57170
rect 183702 57132 183758 57141
rect 226482 57135 226538 57144
rect 227956 57164 228008 57170
rect 225932 57106 225984 57112
rect 227956 57106 228008 57112
rect 183702 57067 183758 57076
rect 225930 56792 225986 56801
rect 225930 56727 225986 56736
rect 182322 55976 182378 55985
rect 182322 55911 182378 55920
rect 182336 55810 182364 55911
rect 225944 55810 225972 56727
rect 226298 56384 226354 56393
rect 226298 56319 226354 56328
rect 226312 56218 226340 56319
rect 226300 56212 226352 56218
rect 226300 56154 226352 56160
rect 226298 55976 226354 55985
rect 226298 55911 226300 55920
rect 226352 55911 226354 55920
rect 226300 55882 226352 55888
rect 182324 55804 182376 55810
rect 182324 55746 182376 55752
rect 225932 55804 225984 55810
rect 225932 55746 225984 55752
rect 227968 55742 227996 57106
rect 182232 55736 182284 55742
rect 182232 55678 182284 55684
rect 227956 55736 228008 55742
rect 227956 55678 228008 55684
rect 228060 55674 228088 57310
rect 182048 55668 182100 55674
rect 182048 55610 182100 55616
rect 228048 55668 228100 55674
rect 228048 55610 228100 55616
rect 225746 55568 225802 55577
rect 225746 55503 225802 55512
rect 181678 54888 181734 54897
rect 181678 54823 181734 54832
rect 181692 54518 181720 54823
rect 225760 54518 225788 55503
rect 226390 55160 226446 55169
rect 226390 55095 226446 55104
rect 226298 54752 226354 54761
rect 226298 54687 226300 54696
rect 226352 54687 226354 54696
rect 226300 54658 226352 54664
rect 181680 54512 181732 54518
rect 181586 54480 181642 54489
rect 181680 54454 181732 54460
rect 225748 54512 225800 54518
rect 225748 54454 225800 54460
rect 226404 54450 226432 55095
rect 181586 54415 181588 54424
rect 181640 54415 181642 54424
rect 226392 54444 226444 54450
rect 181588 54386 181640 54392
rect 226392 54386 226444 54392
rect 182322 54344 182378 54353
rect 182322 54279 182378 54288
rect 226298 54344 226354 54353
rect 226298 54279 226354 54288
rect 182336 53022 182364 54279
rect 226312 54246 226340 54279
rect 226300 54240 226352 54246
rect 226300 54182 226352 54188
rect 225838 54072 225894 54081
rect 225838 54007 225894 54016
rect 182324 53016 182376 53022
rect 182324 52958 182376 52964
rect 181312 52880 181364 52886
rect 181312 52822 181364 52828
rect 181128 51588 181180 51594
rect 181128 51530 181180 51536
rect 188868 50302 188896 53908
rect 198804 51594 198832 53908
rect 198792 51588 198844 51594
rect 198792 51530 198844 51536
rect 208832 50914 208860 53908
rect 208820 50908 208872 50914
rect 208820 50850 208872 50856
rect 218860 50438 218888 53908
rect 225852 53022 225880 54007
rect 225840 53016 225892 53022
rect 225840 52958 225892 52964
rect 222436 50908 222488 50914
rect 222436 50850 222488 50856
rect 218848 50432 218900 50438
rect 218848 50374 218900 50380
rect 220964 50432 221016 50438
rect 220964 50374 221016 50380
rect 187844 50296 187896 50302
rect 187844 50238 187896 50244
rect 188856 50296 188908 50302
rect 188856 50238 188908 50244
rect 180944 48664 180996 48670
rect 180944 48606 180996 48612
rect 187856 37450 187884 50238
rect 193364 47508 193416 47514
rect 193364 47450 193416 47456
rect 193376 37790 193404 47450
rect 220976 47446 221004 50374
rect 220964 47440 221016 47446
rect 220964 47382 221016 47388
rect 192444 37784 192496 37790
rect 192444 37726 192496 37732
rect 193364 37784 193416 37790
rect 193364 37726 193416 37732
rect 186740 37444 186792 37450
rect 186740 37386 186792 37392
rect 187844 37444 187896 37450
rect 187844 37386 187896 37392
rect 186752 34732 186780 37386
rect 192456 34732 192484 37726
rect 198148 37240 198200 37246
rect 198148 37182 198200 37188
rect 198160 34732 198188 37182
rect 203852 37172 203904 37178
rect 203852 37114 203904 37120
rect 209556 37172 209608 37178
rect 209556 37114 209608 37120
rect 203864 34732 203892 37114
rect 209568 34732 209596 37114
rect 220976 34732 221004 47382
rect 215534 34488 215590 34497
rect 215286 34446 215534 34474
rect 215534 34423 215590 34432
rect 222448 28082 222476 50850
rect 228152 47446 228180 84086
rect 231372 79202 231400 112351
rect 231464 111745 231492 138638
rect 231556 117593 231584 138706
rect 231648 125322 231676 138774
rect 231740 127113 231768 139182
rect 231726 127104 231782 127113
rect 231726 127039 231782 127048
rect 231648 125294 231768 125322
rect 231634 125200 231690 125209
rect 231634 125135 231690 125144
rect 231648 125034 231676 125135
rect 231636 125028 231688 125034
rect 231636 124970 231688 124976
rect 231636 122104 231688 122110
rect 231634 122072 231636 122081
rect 231688 122072 231690 122081
rect 231634 122007 231690 122016
rect 231740 120585 231768 125294
rect 231832 124257 231860 139250
rect 236800 138702 236828 141886
rect 237260 138906 237288 141886
rect 237248 138900 237300 138906
rect 237248 138842 237300 138848
rect 237812 138770 237840 141886
rect 238364 138838 238392 141886
rect 239008 139314 239036 141886
rect 238996 139308 239048 139314
rect 238996 139250 239048 139256
rect 239468 139246 239496 141886
rect 239456 139240 239508 139246
rect 239456 139182 239508 139188
rect 238352 138832 238404 138838
rect 238352 138774 238404 138780
rect 237800 138764 237852 138770
rect 237800 138706 237852 138712
rect 236788 138696 236840 138702
rect 236788 138638 236840 138644
rect 240020 138634 240048 141886
rect 232924 138628 232976 138634
rect 232924 138570 232976 138576
rect 240008 138628 240060 138634
rect 240008 138570 240060 138576
rect 231912 132984 231964 132990
rect 231910 132952 231912 132961
rect 231964 132952 231966 132961
rect 231910 132887 231966 132896
rect 232738 130912 232794 130921
rect 232738 130847 232794 130856
rect 232004 130264 232056 130270
rect 232002 130232 232004 130241
rect 232056 130232 232058 130241
rect 232002 130167 232058 130176
rect 231912 124824 231964 124830
rect 231912 124766 231964 124772
rect 231818 124248 231874 124257
rect 231818 124183 231874 124192
rect 231726 120576 231782 120585
rect 231726 120511 231782 120520
rect 231924 120426 231952 124766
rect 232004 122036 232056 122042
rect 232004 121978 232056 121984
rect 231740 120398 231952 120426
rect 231634 118808 231690 118817
rect 231634 118743 231690 118752
rect 231648 118506 231676 118743
rect 231636 118500 231688 118506
rect 231636 118442 231688 118448
rect 231636 117888 231688 117894
rect 231636 117830 231688 117836
rect 231542 117584 231598 117593
rect 231542 117519 231598 117528
rect 231544 115168 231596 115174
rect 231544 115110 231596 115116
rect 231450 111736 231506 111745
rect 231450 111671 231506 111680
rect 231556 109818 231584 115110
rect 231464 109790 231584 109818
rect 231464 109410 231492 109790
rect 231542 109696 231598 109705
rect 231542 109631 231598 109640
rect 231556 109598 231584 109631
rect 231544 109592 231596 109598
rect 231544 109534 231596 109540
rect 231464 109382 231584 109410
rect 231452 108232 231504 108238
rect 231452 108174 231504 108180
rect 231464 97057 231492 108174
rect 231556 102361 231584 109382
rect 231648 103993 231676 117830
rect 231740 108073 231768 120398
rect 232016 119882 232044 121978
rect 231832 119854 232044 119882
rect 231726 108064 231782 108073
rect 231726 107999 231782 108008
rect 231832 106713 231860 119854
rect 231912 119316 231964 119322
rect 231912 119258 231964 119264
rect 231818 106704 231874 106713
rect 231818 106639 231874 106648
rect 231728 105512 231780 105518
rect 231728 105454 231780 105460
rect 231634 103984 231690 103993
rect 231634 103919 231690 103928
rect 231542 102352 231598 102361
rect 231542 102287 231598 102296
rect 231450 97048 231506 97057
rect 231450 96983 231506 96992
rect 231740 95697 231768 105454
rect 231924 105353 231952 119258
rect 232004 111020 232056 111026
rect 232004 110962 232056 110968
rect 231910 105344 231966 105353
rect 231910 105279 231966 105288
rect 232016 99233 232044 110962
rect 232002 99224 232058 99233
rect 232002 99159 232058 99168
rect 231726 95688 231782 95697
rect 231726 95623 231782 95632
rect 231820 94224 231872 94230
rect 231818 94192 231820 94201
rect 231872 94192 231874 94201
rect 231818 94127 231874 94136
rect 231452 93000 231504 93006
rect 231450 92968 231452 92977
rect 231504 92968 231506 92977
rect 231450 92903 231506 92912
rect 231452 91640 231504 91646
rect 231452 91582 231504 91588
rect 231464 91481 231492 91582
rect 231450 91472 231506 91481
rect 231450 91407 231506 91416
rect 231636 90076 231688 90082
rect 231636 90018 231688 90024
rect 231648 89849 231676 90018
rect 231634 89840 231690 89849
rect 231634 89775 231690 89784
rect 231636 88512 231688 88518
rect 231636 88454 231688 88460
rect 231648 88353 231676 88454
rect 231634 88344 231690 88353
rect 231634 88279 231690 88288
rect 231636 86064 231688 86070
rect 231634 86032 231636 86041
rect 231688 86032 231690 86041
rect 231634 85967 231690 85976
rect 231636 84704 231688 84710
rect 231634 84672 231636 84681
rect 231688 84672 231690 84681
rect 231634 84607 231690 84616
rect 231360 79196 231412 79202
rect 231360 79138 231412 79144
rect 232752 78930 232780 130847
rect 232936 130270 232964 138570
rect 240572 132990 240600 141886
rect 240560 132984 240612 132990
rect 240560 132926 240612 132932
rect 241676 130950 241704 141886
rect 242228 139518 242256 141886
rect 242780 139722 242808 141886
rect 243010 141642 243038 141900
rect 243576 141886 243912 141914
rect 244128 141886 244464 141914
rect 244588 141886 244924 141914
rect 245140 141886 245476 141914
rect 245692 141886 245844 141914
rect 246244 141886 246580 141914
rect 246796 141886 247132 141914
rect 247348 141886 247684 141914
rect 247808 141886 248052 141914
rect 248360 141886 248512 141914
rect 248912 141886 249248 141914
rect 249464 141886 249800 141914
rect 243010 141614 243084 141642
rect 242768 139716 242820 139722
rect 242768 139658 242820 139664
rect 243056 139586 243084 141614
rect 243044 139580 243096 139586
rect 243044 139522 243096 139528
rect 242216 139512 242268 139518
rect 242216 139454 242268 139460
rect 243884 138974 243912 141886
rect 243872 138968 243924 138974
rect 243872 138910 243924 138916
rect 244436 138702 244464 141886
rect 244896 139654 244924 141886
rect 244884 139648 244936 139654
rect 244884 139590 244936 139596
rect 245344 139376 245396 139382
rect 245344 139318 245396 139324
rect 244424 138696 244476 138702
rect 244424 138638 244476 138644
rect 245356 131630 245384 139318
rect 245448 139314 245476 141886
rect 245816 139586 245844 141886
rect 245804 139580 245856 139586
rect 245804 139522 245856 139528
rect 245436 139308 245488 139314
rect 245436 139250 245488 139256
rect 245712 139240 245764 139246
rect 245712 139182 245764 139188
rect 245620 138900 245672 138906
rect 245620 138842 245672 138848
rect 244884 131624 244936 131630
rect 244884 131566 244936 131572
rect 245344 131624 245396 131630
rect 245344 131566 245396 131572
rect 243320 131556 243372 131562
rect 243320 131498 243372 131504
rect 241664 130944 241716 130950
rect 241664 130886 241716 130892
rect 232924 130264 232976 130270
rect 232924 130206 232976 130212
rect 243332 128722 243360 131498
rect 243688 130808 243740 130814
rect 243688 130750 243740 130756
rect 243700 128722 243728 130750
rect 244056 130740 244108 130746
rect 244056 130682 244108 130688
rect 244068 128722 244096 130682
rect 244332 130604 244384 130610
rect 244332 130546 244384 130552
rect 244344 128722 244372 130546
rect 244896 128722 244924 131566
rect 245252 130740 245304 130746
rect 245252 130682 245304 130688
rect 245264 128722 245292 130682
rect 245632 128722 245660 138842
rect 245724 130746 245752 139182
rect 246552 139042 246580 141886
rect 246540 139036 246592 139042
rect 246540 138978 246592 138984
rect 247104 138702 247132 141886
rect 247656 139790 247684 141886
rect 247644 139784 247696 139790
rect 247644 139726 247696 139732
rect 247920 139512 247972 139518
rect 247920 139454 247972 139460
rect 246540 138696 246592 138702
rect 246540 138638 246592 138644
rect 247092 138696 247144 138702
rect 247092 138638 247144 138644
rect 245804 138628 245856 138634
rect 245804 138570 245856 138576
rect 245712 130740 245764 130746
rect 245712 130682 245764 130688
rect 245816 128722 245844 138570
rect 246552 131154 246580 138638
rect 246540 131148 246592 131154
rect 246540 131090 246592 131096
rect 247184 130876 247236 130882
rect 247184 130818 247236 130824
rect 246816 130740 246868 130746
rect 246816 130682 246868 130688
rect 246448 130604 246500 130610
rect 246448 130546 246500 130552
rect 246460 128722 246488 130546
rect 246828 128722 246856 130682
rect 247196 128722 247224 130818
rect 247552 130468 247604 130474
rect 247552 130410 247604 130416
rect 247564 128722 247592 130410
rect 247932 130406 247960 139454
rect 248024 131630 248052 141886
rect 248380 138832 248432 138838
rect 248380 138774 248432 138780
rect 248012 131624 248064 131630
rect 248012 131566 248064 131572
rect 248012 131352 248064 131358
rect 248012 131294 248064 131300
rect 247920 130400 247972 130406
rect 247920 130342 247972 130348
rect 248024 128722 248052 131294
rect 248392 128722 248420 138774
rect 248484 131426 248512 141886
rect 249220 139586 249248 141886
rect 249668 139716 249720 139722
rect 249668 139658 249720 139664
rect 249392 139648 249444 139654
rect 249392 139590 249444 139596
rect 249116 139580 249168 139586
rect 249116 139522 249168 139528
rect 249208 139580 249260 139586
rect 249208 139522 249260 139528
rect 248932 139172 248984 139178
rect 248932 139114 248984 139120
rect 248564 131624 248616 131630
rect 248564 131566 248616 131572
rect 248472 131420 248524 131426
rect 248472 131362 248524 131368
rect 248576 128722 248604 131566
rect 248944 128722 248972 139114
rect 249024 138968 249076 138974
rect 249024 138910 249076 138916
rect 249036 131086 249064 138910
rect 249024 131080 249076 131086
rect 249024 131022 249076 131028
rect 249128 130542 249156 139522
rect 249300 139308 249352 139314
rect 249300 139250 249352 139256
rect 249208 138900 249260 138906
rect 249208 138842 249260 138848
rect 249220 130610 249248 138842
rect 249208 130604 249260 130610
rect 249208 130546 249260 130552
rect 249116 130536 249168 130542
rect 249116 130478 249168 130484
rect 249312 130338 249340 139250
rect 249404 131222 249432 139590
rect 249576 139240 249628 139246
rect 249576 139182 249628 139188
rect 249484 139036 249536 139042
rect 249484 138978 249536 138984
rect 249496 131562 249524 138978
rect 249484 131556 249536 131562
rect 249484 131498 249536 131504
rect 249392 131216 249444 131222
rect 249392 131158 249444 131164
rect 249588 130746 249616 139182
rect 249576 130740 249628 130746
rect 249576 130682 249628 130688
rect 249300 130332 249352 130338
rect 249300 130274 249352 130280
rect 249680 128994 249708 139658
rect 249772 139382 249800 141886
rect 249956 141886 250016 141914
rect 250324 141886 250568 141914
rect 251120 141886 251272 141914
rect 251580 141886 251916 141914
rect 249760 139376 249812 139382
rect 249760 139318 249812 139324
rect 249852 139104 249904 139110
rect 249852 139046 249904 139052
rect 249588 128966 249708 128994
rect 249588 128722 249616 128966
rect 249864 128722 249892 139046
rect 249956 131154 249984 141886
rect 250036 139648 250088 139654
rect 250036 139590 250088 139596
rect 250048 131766 250076 139590
rect 250128 139444 250180 139450
rect 250128 139386 250180 139392
rect 250036 131760 250088 131766
rect 250036 131702 250088 131708
rect 250140 131578 250168 139386
rect 250220 139036 250272 139042
rect 250220 138978 250272 138984
rect 250048 131550 250168 131578
rect 250048 131494 250076 131550
rect 250036 131488 250088 131494
rect 250036 131430 250088 131436
rect 249944 131148 249996 131154
rect 249944 131090 249996 131096
rect 250232 130814 250260 138978
rect 250324 131018 250352 141886
rect 250772 139852 250824 139858
rect 250772 139794 250824 139800
rect 250680 139580 250732 139586
rect 250680 139522 250732 139528
rect 250496 139308 250548 139314
rect 250496 139250 250548 139256
rect 250404 138764 250456 138770
rect 250404 138706 250456 138712
rect 250312 131012 250364 131018
rect 250312 130954 250364 130960
rect 250220 130808 250272 130814
rect 250220 130750 250272 130756
rect 250312 130740 250364 130746
rect 250312 130682 250364 130688
rect 250324 128722 250352 130682
rect 250416 128994 250444 138706
rect 250508 131630 250536 139250
rect 250496 131624 250548 131630
rect 250496 131566 250548 131572
rect 250588 130944 250640 130950
rect 250588 130886 250640 130892
rect 250416 128966 250490 128994
rect 243116 128694 243360 128722
rect 243484 128694 243728 128722
rect 243852 128694 244096 128722
rect 244220 128694 244372 128722
rect 244588 128694 244924 128722
rect 245048 128694 245292 128722
rect 245416 128694 245660 128722
rect 245784 128694 245844 128722
rect 246152 128694 246488 128722
rect 246612 128694 246856 128722
rect 246980 128694 247224 128722
rect 247348 128694 247592 128722
rect 247716 128694 248052 128722
rect 248176 128694 248420 128722
rect 248544 128694 248604 128722
rect 248912 128694 248972 128722
rect 249280 128694 249616 128722
rect 249740 128694 249892 128722
rect 250108 128694 250352 128722
rect 250462 128708 250490 128966
rect 250600 128722 250628 130886
rect 250692 130814 250720 139522
rect 250680 130808 250732 130814
rect 250680 130750 250732 130756
rect 250784 130610 250812 139794
rect 250864 139784 250916 139790
rect 250864 139726 250916 139732
rect 250772 130604 250824 130610
rect 250772 130546 250824 130552
rect 250876 130542 250904 139726
rect 251048 139512 251100 139518
rect 251048 139454 251100 139460
rect 250864 130536 250916 130542
rect 250864 130478 250916 130484
rect 251060 130406 251088 139454
rect 251244 130678 251272 141886
rect 251888 139586 251916 141886
rect 251980 141886 252132 141914
rect 252256 141886 252684 141914
rect 252900 141886 253236 141914
rect 253452 141886 253788 141914
rect 254188 141886 254340 141914
rect 254464 141886 254800 141914
rect 255016 141886 255352 141914
rect 255568 141886 255904 141914
rect 256120 141886 256456 141914
rect 256948 141886 257008 141914
rect 257224 141886 257560 141914
rect 257776 141886 258112 141914
rect 258328 141886 258572 141914
rect 258788 141886 259124 141914
rect 259340 141886 259676 141914
rect 259892 141886 260228 141914
rect 260444 141886 260780 141914
rect 261180 141886 261332 141914
rect 261456 141886 261792 141914
rect 262008 141886 262344 141914
rect 262896 141886 263232 141914
rect 251980 139654 252008 141886
rect 251968 139648 252020 139654
rect 252256 139602 252284 141886
rect 251968 139590 252020 139596
rect 251876 139580 251928 139586
rect 251876 139522 251928 139528
rect 252072 139574 252284 139602
rect 252704 139580 252756 139586
rect 251324 139512 251376 139518
rect 251324 139454 251376 139460
rect 251336 130746 251364 139454
rect 252072 131426 252100 139574
rect 252704 139522 252756 139528
rect 252152 139376 252204 139382
rect 252152 139318 252204 139324
rect 252060 131420 252112 131426
rect 252060 131362 252112 131368
rect 251324 130740 251376 130746
rect 251324 130682 251376 130688
rect 251232 130672 251284 130678
rect 251232 130614 251284 130620
rect 251784 130604 251836 130610
rect 251784 130546 251836 130552
rect 250956 130400 251008 130406
rect 250956 130342 251008 130348
rect 251048 130400 251100 130406
rect 251048 130342 251100 130348
rect 251416 130400 251468 130406
rect 251416 130342 251468 130348
rect 250968 128722 250996 130342
rect 251428 128722 251456 130342
rect 251796 128722 251824 130546
rect 252164 130406 252192 139318
rect 252716 131426 252744 139522
rect 252900 139042 252928 141886
rect 253452 139450 253480 141886
rect 254188 139858 254216 141886
rect 254176 139852 254228 139858
rect 254176 139794 254228 139800
rect 254464 139790 254492 141886
rect 254452 139784 254504 139790
rect 254452 139726 254504 139732
rect 253440 139444 253492 139450
rect 253440 139386 253492 139392
rect 255016 139178 255044 141886
rect 255568 139654 255596 141886
rect 255556 139648 255608 139654
rect 255556 139590 255608 139596
rect 255004 139172 255056 139178
rect 255004 139114 255056 139120
rect 252888 139036 252940 139042
rect 252888 138978 252940 138984
rect 256120 138906 256148 141886
rect 256948 139246 256976 141886
rect 256936 139240 256988 139246
rect 256936 139182 256988 139188
rect 256108 138900 256160 138906
rect 256108 138842 256160 138848
rect 254820 138832 254872 138838
rect 254820 138774 254872 138780
rect 253440 138696 253492 138702
rect 253440 138638 253492 138644
rect 252704 131420 252756 131426
rect 252704 131362 252756 131368
rect 252980 131216 253032 131222
rect 252980 131158 253032 131164
rect 252244 131080 252296 131086
rect 252244 131022 252296 131028
rect 252152 130400 252204 130406
rect 252152 130342 252204 130348
rect 252256 128722 252284 131022
rect 252888 130944 252940 130950
rect 252888 130886 252940 130892
rect 250600 128694 250844 128722
rect 250968 128694 251304 128722
rect 251428 128694 251672 128722
rect 251796 128694 252040 128722
rect 252256 128694 252408 128722
rect 252900 128586 252928 130886
rect 252992 128722 253020 131158
rect 253452 130338 253480 138638
rect 254268 131624 254320 131630
rect 254268 131566 254320 131572
rect 253716 130876 253768 130882
rect 253716 130818 253768 130824
rect 253348 130332 253400 130338
rect 253348 130274 253400 130280
rect 253440 130332 253492 130338
rect 253440 130274 253492 130280
rect 253360 128722 253388 130274
rect 253728 128722 253756 130818
rect 254280 128722 254308 131566
rect 254832 131358 254860 138774
rect 254912 138696 254964 138702
rect 254912 138638 254964 138644
rect 254820 131352 254872 131358
rect 254820 131294 254872 131300
rect 254924 130626 254952 138638
rect 257224 138634 257252 141886
rect 257776 138702 257804 141886
rect 258328 138838 258356 141886
rect 258788 139382 258816 141886
rect 258776 139376 258828 139382
rect 258776 139318 258828 139324
rect 259340 139314 259368 141886
rect 259892 139450 259920 141886
rect 260444 139654 260472 141886
rect 260432 139648 260484 139654
rect 260432 139590 260484 139596
rect 259880 139444 259932 139450
rect 259880 139386 259932 139392
rect 259328 139308 259380 139314
rect 259328 139250 259380 139256
rect 261180 139246 261208 141886
rect 261456 139518 261484 141886
rect 261444 139512 261496 139518
rect 261444 139454 261496 139460
rect 261168 139240 261220 139246
rect 261168 139182 261220 139188
rect 258316 138832 258368 138838
rect 258316 138774 258368 138780
rect 257764 138696 257816 138702
rect 257764 138638 257816 138644
rect 262008 138634 262036 141886
rect 263204 138634 263232 141886
rect 263296 141886 263448 141914
rect 263848 141886 264000 141914
rect 263296 139897 263324 141886
rect 263848 139926 263876 141886
rect 264538 141642 264566 141900
rect 264538 141614 264612 141642
rect 263836 139920 263888 139926
rect 263282 139888 263338 139897
rect 263836 139862 263888 139868
rect 263282 139823 263338 139832
rect 264584 138673 264612 141614
rect 264570 138664 264626 138673
rect 255004 138628 255056 138634
rect 255004 138570 255056 138576
rect 257212 138628 257264 138634
rect 257212 138570 257264 138576
rect 261996 138628 262048 138634
rect 261996 138570 262048 138576
rect 263192 138628 263244 138634
rect 263192 138570 263244 138576
rect 263744 138628 263796 138634
rect 264570 138599 264626 138608
rect 263744 138570 263796 138576
rect 255016 131562 255044 138570
rect 255464 135840 255516 135846
rect 255464 135782 255516 135788
rect 255476 131630 255504 135782
rect 255464 131624 255516 131630
rect 255464 131566 255516 131572
rect 258408 131624 258460 131630
rect 258408 131566 258460 131572
rect 255004 131556 255056 131562
rect 255004 131498 255056 131504
rect 255648 131488 255700 131494
rect 255648 131430 255700 131436
rect 255556 130740 255608 130746
rect 255556 130682 255608 130688
rect 254832 130598 254952 130626
rect 254832 130474 254860 130598
rect 254912 130536 254964 130542
rect 254912 130478 254964 130484
rect 254820 130468 254872 130474
rect 254820 130410 254872 130416
rect 254544 130332 254596 130338
rect 254544 130274 254596 130280
rect 254556 128722 254584 130274
rect 254924 128722 254952 130478
rect 255568 128722 255596 130682
rect 252992 128694 253236 128722
rect 253360 128694 253604 128722
rect 253728 128694 253972 128722
rect 254280 128694 254432 128722
rect 254556 128694 254800 128722
rect 254924 128694 255168 128722
rect 255536 128694 255596 128722
rect 255660 128722 255688 131430
rect 258316 131420 258368 131426
rect 258316 131362 258368 131368
rect 256936 131148 256988 131154
rect 256936 131090 256988 131096
rect 256108 130672 256160 130678
rect 256108 130614 256160 130620
rect 256120 128722 256148 130614
rect 256476 130400 256528 130406
rect 256476 130342 256528 130348
rect 256488 128722 256516 130342
rect 256948 128722 256976 131090
rect 257212 131012 257264 131018
rect 257212 130954 257264 130960
rect 257224 128722 257252 130954
rect 257672 130604 257724 130610
rect 257672 130546 257724 130552
rect 257684 128722 257712 130546
rect 258328 128722 258356 131362
rect 255660 128694 255996 128722
rect 256120 128694 256364 128722
rect 256488 128694 256732 128722
rect 256948 128694 257100 128722
rect 257224 128694 257560 128722
rect 257684 128694 257928 128722
rect 258296 128694 258356 128722
rect 258420 128722 258448 131566
rect 258420 128694 258664 128722
rect 252868 128558 252928 128586
rect 239640 127544 239692 127550
rect 239640 127486 239692 127492
rect 238260 125028 238312 125034
rect 238260 124970 238312 124976
rect 236880 122104 236932 122110
rect 236880 122046 236932 122052
rect 235500 118500 235552 118506
rect 235500 118442 235552 118448
rect 234120 115236 234172 115242
rect 234120 115178 234172 115184
rect 232832 109592 232884 109598
rect 232832 109534 232884 109540
rect 232740 78924 232792 78930
rect 232740 78866 232792 78872
rect 232844 78114 232872 109534
rect 234132 78522 234160 115178
rect 234212 101364 234264 101370
rect 234212 101306 234264 101312
rect 234224 93006 234252 101306
rect 234304 98576 234356 98582
rect 234304 98518 234356 98524
rect 234212 93000 234264 93006
rect 234212 92942 234264 92948
rect 234316 91646 234344 98518
rect 234304 91640 234356 91646
rect 234304 91582 234356 91588
rect 234120 78516 234172 78522
rect 234120 78458 234172 78464
rect 235512 78386 235540 118442
rect 236328 91708 236380 91714
rect 236328 91650 236380 91656
rect 236236 88920 236288 88926
rect 236236 88862 236288 88868
rect 236248 84710 236276 88862
rect 236340 86070 236368 91650
rect 236328 86064 236380 86070
rect 236328 86006 236380 86012
rect 236236 84704 236288 84710
rect 236236 84646 236288 84652
rect 236892 79066 236920 122046
rect 236972 102724 237024 102730
rect 236972 102666 237024 102672
rect 236984 94230 237012 102666
rect 237616 94428 237668 94434
rect 237616 94370 237668 94376
rect 236972 94224 237024 94230
rect 236972 94166 237024 94172
rect 237628 88518 237656 94370
rect 237616 88512 237668 88518
rect 237616 88454 237668 88460
rect 238272 79202 238300 124970
rect 238352 95856 238404 95862
rect 238352 95798 238404 95804
rect 238364 90082 238392 95798
rect 238352 90076 238404 90082
rect 238352 90018 238404 90024
rect 237616 79196 237668 79202
rect 237616 79138 237668 79144
rect 238260 79196 238312 79202
rect 238260 79138 238312 79144
rect 236880 79060 236932 79066
rect 236880 79002 236932 79008
rect 235500 78380 235552 78386
rect 235500 78322 235552 78328
rect 232832 78108 232884 78114
rect 232832 78050 232884 78056
rect 236880 78108 236932 78114
rect 236880 78050 236932 78056
rect 233476 76408 233528 76414
rect 233476 76350 233528 76356
rect 233488 75569 233516 76350
rect 236892 75818 236920 78050
rect 237628 75818 237656 79138
rect 239180 79060 239232 79066
rect 239180 79002 239232 79008
rect 237984 78516 238036 78522
rect 237984 78458 238036 78464
rect 237996 75818 238024 78458
rect 238536 78380 238588 78386
rect 238536 78322 238588 78328
rect 238548 75818 238576 78322
rect 239192 75818 239220 79002
rect 239652 78114 239680 127486
rect 240926 125200 240982 125209
rect 240926 125135 240982 125144
rect 240940 124830 240968 125135
rect 240928 124824 240980 124830
rect 240928 124766 240980 124772
rect 240926 122888 240982 122897
rect 240926 122823 240982 122832
rect 240940 122042 240968 122823
rect 240928 122036 240980 122042
rect 240928 121978 240980 121984
rect 261074 120712 261130 120721
rect 261074 120647 261130 120656
rect 240926 120440 240982 120449
rect 240926 120375 240982 120384
rect 240940 119322 240968 120375
rect 240928 119316 240980 119322
rect 240928 119258 240980 119264
rect 261088 118817 261116 120647
rect 261074 118808 261130 118817
rect 261074 118743 261130 118752
rect 240926 118128 240982 118137
rect 240926 118063 240982 118072
rect 240940 117894 240968 118063
rect 240928 117888 240980 117894
rect 240928 117830 240980 117836
rect 240926 115816 240982 115825
rect 240926 115751 240982 115760
rect 240940 115174 240968 115751
rect 240928 115168 240980 115174
rect 240928 115110 240980 115116
rect 263756 115106 263784 138570
rect 263744 115100 263796 115106
rect 263744 115042 263796 115048
rect 240742 113368 240798 113377
rect 240742 113303 240798 113312
rect 240756 112386 240784 113303
rect 240744 112380 240796 112386
rect 240744 112322 240796 112328
rect 240926 111056 240982 111065
rect 240926 110991 240928 111000
rect 240980 110991 240982 111000
rect 240928 110962 240980 110968
rect 240834 108744 240890 108753
rect 240834 108679 240890 108688
rect 240848 108238 240876 108679
rect 240836 108232 240888 108238
rect 240836 108174 240888 108180
rect 240926 106432 240982 106441
rect 240926 106367 240982 106376
rect 240940 105518 240968 106367
rect 240928 105512 240980 105518
rect 240928 105454 240980 105460
rect 240742 103984 240798 103993
rect 240742 103919 240798 103928
rect 240756 102730 240784 103919
rect 240744 102724 240796 102730
rect 240744 102666 240796 102672
rect 240374 101672 240430 101681
rect 240374 101607 240430 101616
rect 240388 101370 240416 101607
rect 240376 101364 240428 101370
rect 240376 101306 240428 101312
rect 240834 99360 240890 99369
rect 240834 99295 240890 99304
rect 240848 98582 240876 99295
rect 262362 98816 262418 98825
rect 262362 98751 262418 98760
rect 262376 98582 262404 98751
rect 240836 98576 240888 98582
rect 240836 98518 240888 98524
rect 262364 98576 262416 98582
rect 262364 98518 262416 98524
rect 240926 96912 240982 96921
rect 240926 96847 240982 96856
rect 240940 95862 240968 96847
rect 240928 95856 240980 95862
rect 240928 95798 240980 95804
rect 240926 94600 240982 94609
rect 240926 94535 240982 94544
rect 240940 94434 240968 94535
rect 240928 94428 240980 94434
rect 240928 94370 240980 94376
rect 240926 92288 240982 92297
rect 240926 92223 240982 92232
rect 240940 91714 240968 92223
rect 240928 91708 240980 91714
rect 240928 91650 240980 91656
rect 240926 89976 240982 89985
rect 240926 89911 240982 89920
rect 240940 88926 240968 89911
rect 240928 88920 240980 88926
rect 240928 88862 240980 88868
rect 243116 88846 243360 88874
rect 243484 88846 243728 88874
rect 243852 88846 244188 88874
rect 244312 88846 244464 88874
rect 244680 88846 244924 88874
rect 245048 88846 245384 88874
rect 245508 88846 245752 88874
rect 245876 88846 246120 88874
rect 246244 88846 246580 88874
rect 246704 88846 246948 88874
rect 247072 88846 247132 88874
rect 247440 88846 247776 88874
rect 247900 88846 248144 88874
rect 248268 88846 248420 88874
rect 248636 88846 248972 88874
rect 249096 88846 249340 88874
rect 249464 88846 249708 88874
rect 249832 88846 249892 88874
rect 250292 88846 250536 88874
rect 250660 88846 250996 88874
rect 251120 88846 251180 88874
rect 251488 88846 251548 88874
rect 243332 86342 243360 88846
rect 243320 86336 243372 86342
rect 243320 86278 243372 86284
rect 243700 86206 243728 88846
rect 243688 86200 243740 86206
rect 243688 86142 243740 86148
rect 244160 86138 244188 88846
rect 244436 86274 244464 88846
rect 244896 86546 244924 88846
rect 245356 86818 245384 88846
rect 245724 86886 245752 88846
rect 246092 87362 246120 88846
rect 246080 87356 246132 87362
rect 246080 87298 246132 87304
rect 246552 87294 246580 88846
rect 246540 87288 246592 87294
rect 246540 87230 246592 87236
rect 246920 87226 246948 88846
rect 246908 87220 246960 87226
rect 246908 87162 246960 87168
rect 247000 86948 247052 86954
rect 247000 86890 247052 86896
rect 245712 86880 245764 86886
rect 245712 86822 245764 86828
rect 245344 86812 245396 86818
rect 245344 86754 245396 86760
rect 245160 86744 245212 86750
rect 245160 86686 245212 86692
rect 244884 86540 244936 86546
rect 244884 86482 244936 86488
rect 244424 86268 244476 86274
rect 244424 86210 244476 86216
rect 244148 86132 244200 86138
rect 244148 86074 244200 86080
rect 245172 79202 245200 86686
rect 247012 79202 247040 86890
rect 239732 79196 239784 79202
rect 239732 79138 239784 79144
rect 241572 79196 241624 79202
rect 241572 79138 241624 79144
rect 245160 79196 245212 79202
rect 245160 79138 245212 79144
rect 246448 79196 246500 79202
rect 246448 79138 246500 79144
rect 247000 79196 247052 79202
rect 247000 79138 247052 79144
rect 239640 78108 239692 78114
rect 239640 78050 239692 78056
rect 239744 75818 239772 79138
rect 240744 78924 240796 78930
rect 240744 78866 240796 78872
rect 240376 78108 240428 78114
rect 240376 78050 240428 78056
rect 240388 75818 240416 78050
rect 240756 75818 240784 78866
rect 236892 75790 237228 75818
rect 237628 75790 237780 75818
rect 237996 75790 238332 75818
rect 238548 75790 238884 75818
rect 239192 75790 239436 75818
rect 239744 75790 239988 75818
rect 240388 75790 240540 75818
rect 240756 75790 241092 75818
rect 241584 75682 241612 79138
rect 242492 79128 242544 79134
rect 242492 79070 242544 79076
rect 242504 75818 242532 79070
rect 244424 79060 244476 79066
rect 244424 79002 244476 79008
rect 244148 78924 244200 78930
rect 244148 78866 244200 78872
rect 243044 78788 243096 78794
rect 243044 78730 243096 78736
rect 243056 75818 243084 78730
rect 243596 78652 243648 78658
rect 243596 78594 243648 78600
rect 243608 75818 243636 78594
rect 244160 75818 244188 78866
rect 242196 75790 242532 75818
rect 242748 75790 243084 75818
rect 243300 75790 243636 75818
rect 243852 75790 244188 75818
rect 244436 75818 244464 79002
rect 245344 78244 245396 78250
rect 245344 78186 245396 78192
rect 245356 75818 245384 78186
rect 245804 78176 245856 78182
rect 245804 78118 245856 78124
rect 245816 75818 245844 78118
rect 246460 75818 246488 79138
rect 246908 78992 246960 78998
rect 246908 78934 246960 78940
rect 246920 75818 246948 78934
rect 247000 78720 247052 78726
rect 247104 78697 247132 88846
rect 247748 87090 247776 88846
rect 248116 87158 248144 88846
rect 248104 87152 248156 87158
rect 248104 87094 248156 87100
rect 247736 87084 247788 87090
rect 247736 87026 247788 87032
rect 247184 87016 247236 87022
rect 247184 86958 247236 86964
rect 247196 78998 247224 86958
rect 247920 86676 247972 86682
rect 247920 86618 247972 86624
rect 247828 86608 247880 86614
rect 247828 86550 247880 86556
rect 247840 79134 247868 86550
rect 247828 79128 247880 79134
rect 247828 79070 247880 79076
rect 247184 78992 247236 78998
rect 247184 78934 247236 78940
rect 247932 78794 247960 86618
rect 248392 86426 248420 88846
rect 248944 86478 248972 88846
rect 248932 86472 248984 86478
rect 248392 86398 248604 86426
rect 248932 86414 248984 86420
rect 248380 86336 248432 86342
rect 248380 86278 248432 86284
rect 248288 86268 248340 86274
rect 248288 86210 248340 86216
rect 248012 86200 248064 86206
rect 248012 86142 248064 86148
rect 247920 78788 247972 78794
rect 247920 78730 247972 78736
rect 247000 78662 247052 78668
rect 247090 78688 247146 78697
rect 244436 75790 244496 75818
rect 245048 75790 245384 75818
rect 245600 75790 245844 75818
rect 246152 75790 246488 75818
rect 246704 75790 246948 75818
rect 247012 75682 247040 78662
rect 247090 78623 247146 78632
rect 248024 78386 248052 86142
rect 248196 86132 248248 86138
rect 248196 86074 248248 86080
rect 248104 78992 248156 78998
rect 248104 78934 248156 78940
rect 248012 78380 248064 78386
rect 248012 78322 248064 78328
rect 248116 75818 248144 78934
rect 248208 78318 248236 86074
rect 248300 78454 248328 86210
rect 248288 78448 248340 78454
rect 248288 78390 248340 78396
rect 248196 78312 248248 78318
rect 248196 78254 248248 78260
rect 248392 78114 248420 86278
rect 248576 78969 248604 86398
rect 249116 86336 249168 86342
rect 249116 86278 249168 86284
rect 248562 78960 248618 78969
rect 248562 78895 248618 78904
rect 248472 78584 248524 78590
rect 248472 78526 248524 78532
rect 248380 78108 248432 78114
rect 248380 78050 248432 78056
rect 248484 75818 248512 78526
rect 249128 78425 249156 86278
rect 249312 86206 249340 88846
rect 249484 86540 249536 86546
rect 249484 86482 249536 86488
rect 249392 86404 249444 86410
rect 249392 86346 249444 86352
rect 249300 86200 249352 86206
rect 249300 86142 249352 86148
rect 249300 86064 249352 86070
rect 249300 86006 249352 86012
rect 249208 79128 249260 79134
rect 249208 79070 249260 79076
rect 249114 78416 249170 78425
rect 249114 78351 249170 78360
rect 249220 75818 249248 79070
rect 249312 79066 249340 86006
rect 249300 79060 249352 79066
rect 249300 79002 249352 79008
rect 249404 78930 249432 86346
rect 249392 78924 249444 78930
rect 249392 78866 249444 78872
rect 249496 78590 249524 86482
rect 249576 86268 249628 86274
rect 249576 86210 249628 86216
rect 249588 78658 249616 86210
rect 249576 78652 249628 78658
rect 249576 78594 249628 78600
rect 249484 78584 249536 78590
rect 249680 78561 249708 88846
rect 249864 86342 249892 88846
rect 249944 87424 249996 87430
rect 249944 87366 249996 87372
rect 249852 86336 249904 86342
rect 249852 86278 249904 86284
rect 249852 86200 249904 86206
rect 249852 86142 249904 86148
rect 249760 79196 249812 79202
rect 249760 79138 249812 79144
rect 249484 78526 249536 78532
rect 249666 78552 249722 78561
rect 249666 78487 249722 78496
rect 249772 75818 249800 79138
rect 249864 78833 249892 86142
rect 249850 78824 249906 78833
rect 249850 78759 249906 78768
rect 247808 75790 248144 75818
rect 248360 75790 248512 75818
rect 248912 75790 249248 75818
rect 249464 75790 249800 75818
rect 249956 75818 249984 87366
rect 250508 83894 250536 88846
rect 250968 86546 250996 88846
rect 251048 87016 251100 87022
rect 251048 86958 251100 86964
rect 250956 86540 251008 86546
rect 250956 86482 251008 86488
rect 250680 86336 250732 86342
rect 250680 86278 250732 86284
rect 250496 83888 250548 83894
rect 250496 83830 250548 83836
rect 250692 78182 250720 86278
rect 250772 86132 250824 86138
rect 250772 86074 250824 86080
rect 250784 78250 250812 86074
rect 250772 78244 250824 78250
rect 250772 78186 250824 78192
rect 250680 78176 250732 78182
rect 250680 78118 250732 78124
rect 249956 75790 250016 75818
rect 251060 75682 251088 86958
rect 251152 86750 251180 88846
rect 251324 86948 251376 86954
rect 251324 86890 251376 86896
rect 251140 86744 251192 86750
rect 251140 86686 251192 86692
rect 251232 86540 251284 86546
rect 251232 86482 251284 86488
rect 251140 83888 251192 83894
rect 251140 83830 251192 83836
rect 251152 78522 251180 83830
rect 251244 78658 251272 86482
rect 251232 78652 251284 78658
rect 251232 78594 251284 78600
rect 251140 78516 251192 78522
rect 251140 78458 251192 78464
rect 251336 75818 251364 86890
rect 251520 86614 251548 88846
rect 251612 88846 251856 88874
rect 251980 88846 252316 88874
rect 252440 88846 252684 88874
rect 252808 88846 253052 88874
rect 253176 88846 253512 88874
rect 253636 88846 253880 88874
rect 254248 88846 254308 88874
rect 251612 86682 251640 88846
rect 251600 86676 251652 86682
rect 251600 86618 251652 86624
rect 251508 86608 251560 86614
rect 251508 86550 251560 86556
rect 251416 86472 251468 86478
rect 251414 86440 251416 86449
rect 251468 86440 251470 86449
rect 251414 86375 251470 86384
rect 251980 86274 252008 88846
rect 252440 86410 252468 88846
rect 252704 86676 252756 86682
rect 252704 86618 252756 86624
rect 252428 86404 252480 86410
rect 252428 86346 252480 86352
rect 251968 86268 252020 86274
rect 251968 86210 252020 86216
rect 252612 86268 252664 86274
rect 252612 86210 252664 86216
rect 252060 78108 252112 78114
rect 252060 78050 252112 78056
rect 252072 75818 252100 78050
rect 252624 75818 252652 86210
rect 252716 78114 252744 86618
rect 252808 86206 252836 88846
rect 252796 86200 252848 86206
rect 252796 86142 252848 86148
rect 253176 86138 253204 88846
rect 253636 86342 253664 88846
rect 254280 86750 254308 88846
rect 254372 88846 254708 88874
rect 254832 88846 255076 88874
rect 255200 88846 255444 88874
rect 255660 88846 255904 88874
rect 256028 88846 256272 88874
rect 256396 88846 256640 88874
rect 256948 88846 257100 88874
rect 257224 88846 257468 88874
rect 257592 88846 257836 88874
rect 258296 88846 258356 88874
rect 254372 87498 254400 88846
rect 254360 87492 254412 87498
rect 254360 87434 254412 87440
rect 254268 86744 254320 86750
rect 254268 86686 254320 86692
rect 253624 86336 253676 86342
rect 253624 86278 253676 86284
rect 253440 86200 253492 86206
rect 253440 86142 253492 86148
rect 253164 86132 253216 86138
rect 253164 86074 253216 86080
rect 253452 78998 253480 86142
rect 254832 86138 254860 88846
rect 255200 86206 255228 88846
rect 255188 86200 255240 86206
rect 255188 86142 255240 86148
rect 253532 86132 253584 86138
rect 253532 86074 253584 86080
rect 254820 86132 254872 86138
rect 254820 86074 254872 86080
rect 255556 86132 255608 86138
rect 255556 86074 255608 86080
rect 253440 78992 253492 78998
rect 253440 78934 253492 78940
rect 253544 78726 253572 86074
rect 255568 79202 255596 86074
rect 255556 79196 255608 79202
rect 255556 79138 255608 79144
rect 255660 78794 255688 88846
rect 255740 87356 255792 87362
rect 255740 87298 255792 87304
rect 255752 79066 255780 87298
rect 256028 86154 256056 88846
rect 256292 87152 256344 87158
rect 256292 87094 256344 87100
rect 256200 86880 256252 86886
rect 256200 86822 256252 86828
rect 256108 86812 256160 86818
rect 256108 86754 256160 86760
rect 255844 86126 256056 86154
rect 255844 79134 255872 86126
rect 256120 86018 256148 86754
rect 255936 85990 256148 86018
rect 255832 79128 255884 79134
rect 255832 79070 255884 79076
rect 255740 79060 255792 79066
rect 255740 79002 255792 79008
rect 255648 78788 255700 78794
rect 255648 78730 255700 78736
rect 253532 78720 253584 78726
rect 253532 78662 253584 78668
rect 254728 78584 254780 78590
rect 254728 78526 254780 78532
rect 254176 78448 254228 78454
rect 254176 78390 254228 78396
rect 253072 78380 253124 78386
rect 253072 78322 253124 78328
rect 252796 78176 252848 78182
rect 252796 78118 252848 78124
rect 252704 78108 252756 78114
rect 252704 78050 252756 78056
rect 251212 75790 251364 75818
rect 251764 75790 252100 75818
rect 252316 75790 252652 75818
rect 252808 75818 252836 78118
rect 253084 75818 253112 78322
rect 253624 78312 253676 78318
rect 253624 78254 253676 78260
rect 253636 75818 253664 78254
rect 254188 75818 254216 78390
rect 254740 75818 254768 78526
rect 255936 75818 255964 85990
rect 256212 85934 256240 86822
rect 256016 85928 256068 85934
rect 256016 85870 256068 85876
rect 256200 85928 256252 85934
rect 256200 85870 256252 85876
rect 252808 75790 252868 75818
rect 253084 75790 253420 75818
rect 253636 75790 253972 75818
rect 254188 75790 254524 75818
rect 254740 75790 255076 75818
rect 255628 75790 255964 75818
rect 256028 75818 256056 85870
rect 256304 85746 256332 87094
rect 256396 86138 256424 88846
rect 256948 87430 256976 88846
rect 256936 87424 256988 87430
rect 256936 87366 256988 87372
rect 256936 87288 256988 87294
rect 256936 87230 256988 87236
rect 256476 87084 256528 87090
rect 256476 87026 256528 87032
rect 256384 86132 256436 86138
rect 256384 86074 256436 86080
rect 256488 86018 256516 87026
rect 256566 86440 256622 86449
rect 256566 86375 256622 86384
rect 256212 85718 256332 85746
rect 256396 85990 256516 86018
rect 256212 78998 256240 85718
rect 256292 85656 256344 85662
rect 256292 85598 256344 85604
rect 256304 79134 256332 85598
rect 256396 79202 256424 85990
rect 256580 85662 256608 86375
rect 256568 85656 256620 85662
rect 256568 85598 256620 85604
rect 256384 79196 256436 79202
rect 256384 79138 256436 79144
rect 256292 79128 256344 79134
rect 256292 79070 256344 79076
rect 256568 79128 256620 79134
rect 256568 79070 256620 79076
rect 256384 79060 256436 79066
rect 256384 79002 256436 79008
rect 256200 78992 256252 78998
rect 256200 78934 256252 78940
rect 256396 75818 256424 79002
rect 256580 78998 256608 79070
rect 256568 78992 256620 78998
rect 256568 78934 256620 78940
rect 256948 75818 256976 87230
rect 257028 87220 257080 87226
rect 257028 87162 257080 87168
rect 257040 79406 257068 87162
rect 257224 87022 257252 88846
rect 257212 87016 257264 87022
rect 257212 86958 257264 86964
rect 257592 86954 257620 88846
rect 257580 86948 257632 86954
rect 257580 86890 257632 86896
rect 258328 86682 258356 88846
rect 258420 88846 258664 88874
rect 258316 86676 258368 86682
rect 258316 86618 258368 86624
rect 258420 86274 258448 88846
rect 258408 86268 258460 86274
rect 258408 86210 258460 86216
rect 257028 79400 257080 79406
rect 257028 79342 257080 79348
rect 257488 79400 257540 79406
rect 257488 79342 257540 79348
rect 257500 75818 257528 79342
rect 258684 79196 258736 79202
rect 258684 79138 258736 79144
rect 264296 79196 264348 79202
rect 264296 79138 264348 79144
rect 258314 78688 258370 78697
rect 258314 78623 258370 78632
rect 258328 75818 258356 78623
rect 258696 75818 258724 79138
rect 259236 79128 259288 79134
rect 259236 79070 259288 79076
rect 259248 75818 259276 79070
rect 260340 79060 260392 79066
rect 260340 79002 260392 79008
rect 259786 78960 259842 78969
rect 259786 78895 259842 78904
rect 259800 75818 259828 78895
rect 260352 75818 260380 79002
rect 261074 78824 261130 78833
rect 261074 78759 261130 78768
rect 261088 75818 261116 78759
rect 263100 78652 263152 78658
rect 263100 78594 263152 78600
rect 261442 78552 261498 78561
rect 261442 78487 261498 78496
rect 262548 78516 262600 78522
rect 261456 75818 261484 78487
rect 262548 78458 262600 78464
rect 261994 78416 262050 78425
rect 261994 78351 262050 78360
rect 262008 75818 262036 78351
rect 262560 75818 262588 78458
rect 263112 75818 263140 78594
rect 264308 75818 264336 79138
rect 264480 78516 264532 78522
rect 264480 78458 264532 78464
rect 256028 75790 256180 75818
rect 256396 75790 256732 75818
rect 256948 75790 257284 75818
rect 257500 75790 257836 75818
rect 258328 75790 258480 75818
rect 258696 75790 259032 75818
rect 259248 75790 259584 75818
rect 259800 75790 260136 75818
rect 260352 75790 260688 75818
rect 261088 75790 261240 75818
rect 261456 75790 261792 75818
rect 262008 75790 262344 75818
rect 262560 75790 262896 75818
rect 263112 75790 263448 75818
rect 264000 75790 264336 75818
rect 241584 75654 241644 75682
rect 247012 75654 247256 75682
rect 250568 75654 251088 75682
rect 264492 75682 264520 78458
rect 264492 75654 264552 75682
rect 233474 75560 233530 75569
rect 233474 75495 233530 75504
rect 233660 75048 233712 75054
rect 233474 75016 233530 75025
rect 233660 74990 233712 74996
rect 233474 74951 233530 74960
rect 233568 74980 233620 74986
rect 233488 74918 233516 74951
rect 233568 74922 233620 74928
rect 233476 74912 233528 74918
rect 233476 74854 233528 74860
rect 233580 74345 233608 74922
rect 233566 74336 233622 74345
rect 233566 74271 233622 74280
rect 233672 73801 233700 74990
rect 233658 73792 233714 73801
rect 233658 73727 233714 73736
rect 234118 72704 234174 72713
rect 234118 72639 234174 72648
rect 233474 72568 233530 72577
rect 233474 72503 233530 72512
rect 233488 72402 233516 72503
rect 230624 72396 230676 72402
rect 230624 72338 230676 72344
rect 233476 72396 233528 72402
rect 233476 72338 233528 72344
rect 230636 70906 230664 72338
rect 233566 71480 233622 71489
rect 233566 71415 233622 71424
rect 233474 71072 233530 71081
rect 233474 71007 233530 71016
rect 230624 70900 230676 70906
rect 230624 70842 230676 70848
rect 229888 69744 229940 69750
rect 229888 69686 229940 69692
rect 229900 68798 229928 69686
rect 233488 69478 233516 71007
rect 233580 69546 233608 71415
rect 233658 70256 233714 70265
rect 233658 70191 233714 70200
rect 233672 69750 233700 70191
rect 233660 69744 233712 69750
rect 233660 69686 233712 69692
rect 233750 69576 233806 69585
rect 233568 69540 233620 69546
rect 233750 69511 233806 69520
rect 233568 69482 233620 69488
rect 233476 69472 233528 69478
rect 233476 69414 233528 69420
rect 233658 69032 233714 69041
rect 233658 68967 233714 68976
rect 229888 68792 229940 68798
rect 229888 68734 229940 68740
rect 233566 68352 233622 68361
rect 233566 68287 233622 68296
rect 233474 68216 233530 68225
rect 233580 68186 233608 68287
rect 233474 68151 233530 68160
rect 233568 68180 233620 68186
rect 233488 68050 233516 68151
rect 233568 68122 233620 68128
rect 233672 68118 233700 68967
rect 233660 68112 233712 68118
rect 233660 68054 233712 68060
rect 233476 68044 233528 68050
rect 233476 67986 233528 67992
rect 233764 67982 233792 69511
rect 233752 67976 233804 67982
rect 233752 67918 233804 67924
rect 233566 67128 233622 67137
rect 233566 67063 233622 67072
rect 233474 66992 233530 67001
rect 233474 66927 233530 66936
rect 233488 66758 233516 66927
rect 233476 66752 233528 66758
rect 233476 66694 233528 66700
rect 233580 66690 233608 67063
rect 233568 66684 233620 66690
rect 233568 66626 233620 66632
rect 233474 66176 233530 66185
rect 233474 66111 233530 66120
rect 233488 66078 233516 66111
rect 233476 66072 233528 66078
rect 233476 66014 233528 66020
rect 233474 65496 233530 65505
rect 233474 65431 233530 65440
rect 233488 65398 233516 65431
rect 233476 65392 233528 65398
rect 233476 65334 233528 65340
rect 233566 64816 233622 64825
rect 233566 64751 233568 64760
rect 233620 64751 233622 64760
rect 233568 64722 233620 64728
rect 233476 64712 233528 64718
rect 233476 64654 233528 64660
rect 233488 64553 233516 64654
rect 233474 64544 233530 64553
rect 233474 64479 233530 64488
rect 233660 63488 233712 63494
rect 233474 63456 233530 63465
rect 233660 63430 233712 63436
rect 233474 63391 233476 63400
rect 233528 63391 233530 63400
rect 233476 63362 233528 63368
rect 233568 63352 233620 63358
rect 233672 63329 233700 63430
rect 233568 63294 233620 63300
rect 233658 63320 233714 63329
rect 233580 62785 233608 63294
rect 233658 63255 233714 63264
rect 233566 62776 233622 62785
rect 233566 62711 233622 62720
rect 233476 62672 233528 62678
rect 233476 62614 233528 62620
rect 233488 62241 233516 62614
rect 233474 62232 233530 62241
rect 233474 62167 233530 62176
rect 233476 61924 233528 61930
rect 233476 61866 233528 61872
rect 233488 61561 233516 61866
rect 233474 61552 233530 61561
rect 233474 61487 233530 61496
rect 233476 61380 233528 61386
rect 233476 61322 233528 61328
rect 233488 61017 233516 61322
rect 233568 61312 233620 61318
rect 233568 61254 233620 61260
rect 233474 61008 233530 61017
rect 233474 60943 233530 60952
rect 233580 60337 233608 61254
rect 233566 60328 233622 60337
rect 233566 60263 233622 60272
rect 233752 60156 233804 60162
rect 233752 60098 233804 60104
rect 233476 60020 233528 60026
rect 233476 59962 233528 59968
rect 233488 59793 233516 59962
rect 233568 59952 233620 59958
rect 233568 59894 233620 59900
rect 233474 59784 233530 59793
rect 233474 59719 233530 59728
rect 233580 59113 233608 59894
rect 233566 59104 233622 59113
rect 233566 59039 233622 59048
rect 233476 58728 233528 58734
rect 233476 58670 233528 58676
rect 233488 57345 233516 58670
rect 233568 58660 233620 58666
rect 233568 58602 233620 58608
rect 233474 57336 233530 57345
rect 228600 57300 228652 57306
rect 233474 57271 233530 57280
rect 228600 57242 228652 57248
rect 228612 54382 228640 57242
rect 228692 57232 228744 57238
rect 228692 57174 228744 57180
rect 228600 54376 228652 54382
rect 228600 54318 228652 54324
rect 228704 54314 228732 57174
rect 233580 56665 233608 58602
rect 233660 58592 233712 58598
rect 233764 58569 233792 60098
rect 233844 60088 233896 60094
rect 233844 60030 233896 60036
rect 233660 58534 233712 58540
rect 233750 58560 233806 58569
rect 233566 56656 233622 56665
rect 233566 56591 233622 56600
rect 229428 56212 229480 56218
rect 229428 56154 229480 56160
rect 229336 55940 229388 55946
rect 229336 55882 229388 55888
rect 228692 54308 228744 54314
rect 228692 54250 228744 54256
rect 229348 52818 229376 55882
rect 229440 52886 229468 56154
rect 233672 56121 233700 58534
rect 233750 58495 233806 58504
rect 233856 57889 233884 60030
rect 233842 57880 233898 57889
rect 233842 57815 233898 57824
rect 233658 56112 233714 56121
rect 233658 56047 233714 56056
rect 229612 55804 229664 55810
rect 229612 55746 229664 55752
rect 229520 54716 229572 54722
rect 229520 54658 229572 54664
rect 229428 52880 229480 52886
rect 229428 52822 229480 52828
rect 229336 52812 229388 52818
rect 229336 52754 229388 52760
rect 229532 50166 229560 54658
rect 229624 52954 229652 55746
rect 233568 55736 233620 55742
rect 233568 55678 233620 55684
rect 233476 55668 233528 55674
rect 233476 55610 233528 55616
rect 233488 55441 233516 55610
rect 233474 55432 233530 55441
rect 233474 55367 233530 55376
rect 233580 54897 233608 55678
rect 233566 54888 233622 54897
rect 233566 54823 233622 54832
rect 230900 54512 230952 54518
rect 230900 54454 230952 54460
rect 230716 54444 230768 54450
rect 230716 54386 230768 54392
rect 229612 52948 229664 52954
rect 229612 52890 229664 52896
rect 230728 51458 230756 54386
rect 230912 51594 230940 54454
rect 233476 54376 233528 54382
rect 233476 54318 233528 54324
rect 231728 54240 231780 54246
rect 233488 54217 233516 54318
rect 233568 54308 233620 54314
rect 233568 54250 233620 54256
rect 231728 54182 231780 54188
rect 233474 54208 233530 54217
rect 230900 51588 230952 51594
rect 230900 51530 230952 51536
rect 230716 51452 230768 51458
rect 230716 51394 230768 51400
rect 231740 50234 231768 54182
rect 233474 54143 233530 54152
rect 233580 53673 233608 54250
rect 233566 53664 233622 53673
rect 233566 53599 233622 53608
rect 233568 53016 233620 53022
rect 233474 52984 233530 52993
rect 233568 52958 233620 52964
rect 233474 52919 233476 52928
rect 233528 52919 233530 52928
rect 233476 52890 233528 52896
rect 233476 52812 233528 52818
rect 233476 52754 233528 52760
rect 233488 51769 233516 52754
rect 233474 51760 233530 51769
rect 233474 51695 233530 51704
rect 233476 51588 233528 51594
rect 233476 51530 233528 51536
rect 233488 51225 233516 51530
rect 233474 51216 233530 51225
rect 233474 51151 233530 51160
rect 231728 50228 231780 50234
rect 231728 50170 231780 50176
rect 233476 50228 233528 50234
rect 233476 50170 233528 50176
rect 229520 50160 229572 50166
rect 229520 50102 229572 50108
rect 233488 49321 233516 50170
rect 233474 49312 233530 49321
rect 233474 49247 233530 49256
rect 233580 48777 233608 52958
rect 233660 52880 233712 52886
rect 233660 52822 233712 52828
rect 233672 52449 233700 52822
rect 233658 52440 233714 52449
rect 233658 52375 233714 52384
rect 234132 51526 234160 72639
rect 234120 51520 234172 51526
rect 234120 51462 234172 51468
rect 233660 51452 233712 51458
rect 233660 51394 233712 51400
rect 233672 50545 233700 51394
rect 233658 50536 233714 50545
rect 233658 50471 233714 50480
rect 233660 50160 233712 50166
rect 233660 50102 233712 50108
rect 233672 50001 233700 50102
rect 233658 49992 233714 50001
rect 233658 49927 233714 49936
rect 233566 48768 233622 48777
rect 233566 48703 233622 48712
rect 241216 47910 241552 47938
rect 250508 47910 250844 47938
rect 260136 47910 260472 47938
rect 233474 47680 233530 47689
rect 233474 47615 233530 47624
rect 233488 47514 233516 47615
rect 241216 47553 241244 47910
rect 241202 47544 241258 47553
rect 233476 47508 233528 47514
rect 241202 47479 241258 47488
rect 233476 47450 233528 47456
rect 228140 47440 228192 47446
rect 228140 47382 228192 47388
rect 250508 45921 250536 47910
rect 260444 47446 260472 47910
rect 260432 47440 260484 47446
rect 260432 47382 260484 47388
rect 250494 45912 250550 45921
rect 250494 45847 250550 45856
rect 260444 45406 260472 47382
rect 260432 45400 260484 45406
rect 260432 45342 260484 45348
rect 222448 28066 222844 28082
rect 222448 28060 222856 28066
rect 222448 28054 222804 28060
rect 222804 28002 222856 28008
rect 223540 28060 223592 28066
rect 223540 28002 223592 28008
rect 223552 27561 223580 28002
rect 223538 27552 223594 27561
rect 223538 27487 223594 27496
rect 203864 17118 203892 18956
rect 203852 17112 203904 17118
rect 203852 17054 203904 17060
rect 248748 12352 248800 12358
rect 211946 12320 212002 12329
rect 248748 12294 248800 12300
rect 211946 12255 212002 12264
rect 175240 9428 175292 9434
rect 175240 9370 175292 9376
rect 175424 9428 175476 9434
rect 175424 9370 175476 9376
rect 175252 9304 175280 9370
rect 211960 9304 211988 12255
rect 248760 9304 248788 12294
rect 264676 12290 264704 242231
rect 264768 242062 264796 294630
rect 265860 294620 265912 294626
rect 265860 294562 265912 294568
rect 265872 266882 265900 294562
rect 265860 266876 265912 266882
rect 265860 266818 265912 266824
rect 264756 242056 264808 242062
rect 264756 241998 264808 242004
rect 267252 224790 267280 299390
rect 285468 299318 285496 302344
rect 292540 299380 292592 299386
rect 292540 299322 292592 299328
rect 285456 299312 285508 299318
rect 285456 299254 285508 299260
rect 281868 225328 281920 225334
rect 281868 225270 281920 225276
rect 267240 224784 267292 224790
rect 267240 224726 267292 224732
rect 281880 222820 281908 225270
rect 289872 224784 289924 224790
rect 289872 224726 289924 224732
rect 289884 222820 289912 224726
rect 276162 217680 276218 217689
rect 276162 217615 276218 217624
rect 265214 216592 265270 216601
rect 265214 216527 265270 216536
rect 265228 212890 265256 216527
rect 265216 212884 265268 212890
rect 265216 212826 265268 212832
rect 274876 208940 274928 208946
rect 274876 208882 274928 208888
rect 274888 208441 274916 208882
rect 274874 208432 274930 208441
rect 274874 208367 274930 208376
rect 274874 197688 274930 197697
rect 274874 197623 274930 197632
rect 274888 196570 274916 197623
rect 274876 196564 274928 196570
rect 274876 196506 274928 196512
rect 275520 192416 275572 192422
rect 275520 192358 275572 192364
rect 275532 188177 275560 192358
rect 275518 188168 275574 188177
rect 275518 188103 275574 188112
rect 264848 175280 264900 175286
rect 264848 175222 264900 175228
rect 264756 175144 264808 175150
rect 264756 175086 264808 175092
rect 264768 149417 264796 175086
rect 264860 163289 264888 175222
rect 265860 167596 265912 167602
rect 265860 167538 265912 167544
rect 264846 163280 264902 163289
rect 264846 163215 264902 163224
rect 264754 149408 264810 149417
rect 264754 149343 264810 149352
rect 265124 102724 265176 102730
rect 265124 102666 265176 102672
rect 264848 81440 264900 81446
rect 264848 81382 264900 81388
rect 264756 81304 264808 81310
rect 264756 81246 264808 81252
rect 264768 55441 264796 81246
rect 264860 69449 264888 81382
rect 265136 79202 265164 102666
rect 265124 79196 265176 79202
rect 265124 79138 265176 79144
rect 264846 69440 264902 69449
rect 264846 69375 264902 69384
rect 264754 55432 264810 55441
rect 264754 55367 264810 55376
rect 265872 17118 265900 167538
rect 276070 123704 276126 123713
rect 276070 123639 276126 123648
rect 274876 115100 274928 115106
rect 274876 115042 274928 115048
rect 274888 114465 274916 115042
rect 274874 114456 274930 114465
rect 274874 114391 274930 114400
rect 274874 103712 274930 103721
rect 274874 103647 274930 103656
rect 274888 102730 274916 103647
rect 274876 102724 274928 102730
rect 274876 102666 274928 102672
rect 272760 98576 272812 98582
rect 272760 98518 272812 98524
rect 272772 94366 272800 98518
rect 272760 94360 272812 94366
rect 274876 94360 274928 94366
rect 272760 94302 272812 94308
rect 274874 94328 274876 94337
rect 274928 94328 274930 94337
rect 274874 94263 274930 94272
rect 276084 46086 276112 123639
rect 276176 70906 276204 217615
rect 285928 181241 285956 182836
rect 285914 181232 285970 181241
rect 285914 181167 285970 181176
rect 281868 131284 281920 131290
rect 281868 131226 281920 131232
rect 281880 128708 281908 131226
rect 289870 130368 289926 130377
rect 289870 130303 289926 130312
rect 289884 128708 289912 130303
rect 292552 112402 292580 299322
rect 292632 294552 292684 294558
rect 292632 294494 292684 294500
rect 292644 217258 292672 294494
rect 300358 290576 300414 290585
rect 300358 290511 300414 290520
rect 300084 266876 300136 266882
rect 300084 266818 300136 266824
rect 300096 266105 300124 266818
rect 300082 266096 300138 266105
rect 300082 266031 300138 266040
rect 300176 242056 300228 242062
rect 300176 241998 300228 242004
rect 300188 241625 300216 241998
rect 300174 241616 300230 241625
rect 300174 241551 300230 241560
rect 292644 217230 292856 217258
rect 292828 217174 292856 217230
rect 292816 217168 292868 217174
rect 300176 217168 300228 217174
rect 292816 217110 292868 217116
rect 300174 217136 300176 217145
rect 300228 217136 300230 217145
rect 300174 217071 300230 217080
rect 296218 202856 296274 202865
rect 296218 202791 296274 202800
rect 293550 188984 293606 188993
rect 292816 188948 292868 188954
rect 293550 188919 293552 188928
rect 292816 188890 292868 188896
rect 293604 188919 293606 188928
rect 293552 188890 293604 188896
rect 292828 188834 292856 188890
rect 292644 188806 292856 188834
rect 292644 168894 292672 188806
rect 292632 168888 292684 168894
rect 292632 168830 292684 168836
rect 296232 144074 296260 202791
rect 300174 168176 300230 168185
rect 300174 168111 300230 168120
rect 300188 167602 300216 168111
rect 300176 167596 300228 167602
rect 300176 167538 300228 167544
rect 296220 144068 296272 144074
rect 296220 144010 296272 144016
rect 300176 144068 300228 144074
rect 300176 144010 300228 144016
rect 300188 143569 300216 144010
rect 300174 143560 300230 143569
rect 300174 143495 300230 143504
rect 300174 119080 300230 119089
rect 300174 119015 300230 119024
rect 300188 117894 300216 119015
rect 292816 117888 292868 117894
rect 292644 117836 292816 117842
rect 292644 117830 292868 117836
rect 300176 117888 300228 117894
rect 300176 117830 300228 117836
rect 292644 117814 292856 117830
rect 292644 112538 292672 117814
rect 292644 112522 292856 112538
rect 292644 112516 292868 112522
rect 292644 112510 292816 112516
rect 292816 112458 292868 112464
rect 292552 112374 292856 112402
rect 292828 111978 292856 112374
rect 292816 111972 292868 111978
rect 292816 111914 292868 111920
rect 293552 111972 293604 111978
rect 293552 111914 293604 111920
rect 292816 110272 292868 110278
rect 292816 110214 292868 110220
rect 292828 109138 292856 110214
rect 293564 109569 293592 111914
rect 293550 109560 293606 109569
rect 293550 109495 293606 109504
rect 292644 109110 292856 109138
rect 285928 87401 285956 88860
rect 292540 88172 292592 88178
rect 292540 88114 292592 88120
rect 285914 87392 285970 87401
rect 285914 87327 285970 87336
rect 276164 70900 276216 70906
rect 276164 70842 276216 70848
rect 276072 46080 276124 46086
rect 276072 46022 276124 46028
rect 284536 45400 284588 45406
rect 284536 45342 284588 45348
rect 265860 17112 265912 17118
rect 265860 17054 265912 17060
rect 264664 12284 264716 12290
rect 264664 12226 264716 12232
rect 284548 9434 284576 45342
rect 292552 37110 292580 88114
rect 292644 37178 292672 109110
rect 295574 95552 295630 95561
rect 295574 95487 295630 95496
rect 292816 94428 292868 94434
rect 292816 94370 292868 94376
rect 292828 94314 292856 94370
rect 292736 94286 292856 94314
rect 292736 88178 292764 94286
rect 292724 88172 292776 88178
rect 292724 88114 292776 88120
rect 295588 78522 295616 95487
rect 299714 94600 299770 94609
rect 299714 94535 299770 94544
rect 299728 94434 299756 94535
rect 299716 94428 299768 94434
rect 299716 94370 299768 94376
rect 300372 84302 300400 290511
rect 300450 202312 300506 202321
rect 300450 202247 300506 202256
rect 300464 192665 300492 202247
rect 300450 192656 300506 192665
rect 300450 192591 300506 192600
rect 300360 84296 300412 84302
rect 300360 84238 300412 84244
rect 295576 78516 295628 78522
rect 295576 78458 295628 78464
rect 300176 70900 300228 70906
rect 300176 70842 300228 70848
rect 300188 70129 300216 70842
rect 300174 70120 300230 70129
rect 300174 70055 300230 70064
rect 300176 46080 300228 46086
rect 300176 46022 300228 46028
rect 300188 45649 300216 46022
rect 300174 45640 300230 45649
rect 300174 45575 300230 45584
rect 292632 37172 292684 37178
rect 292632 37114 292684 37120
rect 292540 37104 292592 37110
rect 292540 37046 292592 37052
rect 299806 21160 299862 21169
rect 299806 21095 299862 21104
rect 299820 20926 299848 21095
rect 299808 20920 299860 20926
rect 299808 20862 299860 20868
rect 284536 9428 284588 9434
rect 284536 9370 284588 9376
rect 285456 9428 285508 9434
rect 285456 9370 285508 9376
rect 285468 9304 285496 9370
rect 28222 8824 28278 9304
rect 64930 8824 64986 9304
rect 101730 8824 101786 9304
rect 138438 8824 138494 9304
rect 175238 8824 175294 9304
rect 211946 8824 212002 9304
rect 248746 8824 248802 9304
rect 285454 8824 285510 9304
<< via2 >>
rect 13318 287800 13374 287856
rect 13226 286440 13282 286496
rect 12950 221160 13006 221216
rect 13686 253800 13742 253856
rect 13502 188520 13558 188576
rect 13410 123104 13466 123160
rect 13318 57824 13374 57880
rect 13594 155744 13650 155800
rect 13318 25184 13374 25240
rect 24174 224152 24230 224208
rect 13686 131536 13742 131592
rect 23898 130312 23954 130368
rect 13778 90464 13834 90520
rect 88482 284808 88538 284864
rect 62906 265496 62962 265552
rect 78914 263728 78970 263784
rect 79558 263320 79614 263376
rect 80110 262096 80166 262152
rect 80202 261436 80258 261472
rect 80202 261416 80204 261436
rect 80204 261416 80256 261436
rect 80256 261416 80258 261436
rect 80110 260736 80166 260792
rect 80202 260092 80204 260112
rect 80204 260092 80256 260112
rect 80256 260092 80258 260112
rect 80202 260056 80258 260092
rect 79834 259376 79890 259432
rect 80202 258716 80258 258752
rect 80202 258696 80204 258716
rect 80204 258696 80256 258716
rect 80256 258696 80258 258716
rect 80018 258016 80074 258072
rect 80202 257336 80258 257392
rect 80110 256792 80166 256848
rect 80202 256112 80258 256168
rect 80110 255432 80166 255488
rect 80202 254752 80258 254808
rect 87194 258288 87250 258344
rect 131354 280728 131410 280784
rect 182322 284808 182378 284864
rect 139634 263456 139690 263512
rect 131354 257608 131410 257664
rect 87286 257472 87342 257528
rect 129514 257472 129570 257528
rect 143038 263184 143094 263240
rect 173398 262776 173454 262832
rect 139634 262676 139636 262696
rect 139636 262676 139688 262696
rect 139688 262676 139690 262696
rect 139634 262640 139690 262676
rect 173674 262096 173730 262152
rect 140278 261416 140334 261472
rect 173582 261452 173584 261472
rect 173584 261452 173636 261472
rect 173636 261452 173638 261472
rect 173582 261416 173638 261452
rect 140094 259512 140150 259568
rect 139910 258832 139966 258888
rect 139818 258152 139874 258208
rect 139634 257608 139690 257664
rect 87286 256792 87342 256848
rect 131354 256792 131410 256848
rect 87562 256656 87618 256712
rect 131446 256656 131502 256712
rect 87194 256248 87250 256304
rect 131538 256248 131594 256304
rect 87194 255432 87250 255488
rect 131354 255704 131410 255760
rect 87378 255568 87434 255624
rect 131446 255296 131502 255352
rect 131538 255160 131594 255216
rect 87286 255024 87342 255080
rect 131630 254752 131686 254808
rect 80110 254072 80166 254128
rect 87194 254344 87250 254400
rect 87286 254208 87342 254264
rect 131354 254072 131410 254128
rect 87378 253800 87434 253856
rect 131538 253800 131594 253856
rect 131446 253664 131502 253720
rect 80202 253392 80258 253448
rect 87194 253392 87250 253448
rect 87194 253020 87196 253040
rect 87196 253020 87248 253040
rect 87248 253020 87250 253040
rect 87194 252984 87250 253020
rect 131354 252984 131410 253040
rect 80202 252712 80258 252768
rect 131446 252848 131502 252904
rect 87286 252576 87342 252632
rect 131538 252440 131594 252496
rect 87194 252168 87250 252224
rect 80202 252032 80258 252088
rect 131354 251896 131410 251952
rect 87194 251488 87250 251544
rect 131354 251488 131410 251544
rect 80202 251352 80258 251408
rect 87194 251100 87250 251136
rect 87194 251080 87196 251100
rect 87196 251080 87248 251100
rect 87248 251080 87250 251100
rect 131354 251100 131410 251136
rect 131354 251080 131356 251100
rect 131356 251080 131408 251100
rect 131408 251080 131410 251100
rect 87286 250980 87288 251000
rect 87288 250980 87340 251000
rect 87340 250980 87342 251000
rect 87286 250944 87342 250980
rect 80110 250672 80166 250728
rect 131446 250672 131502 250728
rect 87194 250264 87250 250320
rect 131354 250284 131410 250320
rect 131354 250264 131356 250284
rect 131356 250264 131408 250284
rect 131408 250264 131410 250284
rect 80110 250128 80166 250184
rect 47082 249856 47138 249912
rect 87286 249992 87342 250048
rect 131354 249992 131410 250048
rect 87378 249584 87434 249640
rect 131814 249620 131816 249640
rect 131816 249620 131868 249640
rect 131868 249620 131870 249640
rect 80202 249448 80258 249504
rect 87194 249176 87250 249232
rect 131814 249584 131870 249620
rect 131354 249176 131410 249232
rect 80202 248804 80204 248824
rect 80204 248804 80256 248824
rect 80256 248804 80258 248824
rect 80202 248768 80258 248804
rect 88298 248768 88354 248824
rect 131354 248768 131410 248824
rect 79282 248496 79338 248552
rect 88022 247952 88078 248008
rect 80202 247444 80204 247464
rect 80204 247444 80256 247464
rect 80256 247444 80258 247464
rect 80202 247408 80258 247444
rect 79282 247136 79338 247192
rect 79282 245776 79338 245832
rect 79098 241288 79154 241344
rect 80202 246048 80258 246104
rect 87194 247580 87196 247600
rect 87196 247580 87248 247600
rect 87248 247580 87250 247600
rect 87194 247544 87250 247580
rect 88390 248360 88446 248416
rect 131446 248360 131502 248416
rect 132550 247952 132606 248008
rect 131814 247716 131816 247736
rect 131816 247716 131868 247736
rect 131868 247716 131870 247736
rect 131814 247680 131870 247716
rect 131446 247272 131502 247328
rect 87010 247136 87066 247192
rect 86918 245912 86974 245968
rect 86826 245504 86882 245560
rect 80202 244708 80258 244744
rect 80202 244688 80204 244708
rect 80204 244688 80256 244708
rect 80256 244688 80258 244708
rect 80110 244416 80166 244472
rect 80018 243328 80074 243384
rect 80202 243056 80258 243112
rect 87102 246728 87158 246784
rect 131354 246456 131410 246512
rect 87194 246356 87196 246376
rect 87196 246356 87248 246376
rect 87248 246356 87250 246376
rect 87194 246320 87250 246356
rect 132182 246864 132238 246920
rect 131998 246048 132054 246104
rect 131446 245776 131502 245832
rect 131354 245368 131410 245424
rect 87654 245096 87710 245152
rect 87562 244688 87618 244744
rect 87286 244280 87342 244336
rect 87194 243872 87250 243928
rect 87470 243464 87526 243520
rect 87194 243056 87250 243112
rect 86550 242648 86606 242704
rect 80202 242376 80258 242432
rect 86458 242240 86514 242296
rect 80202 241696 80258 241752
rect 80110 240608 80166 240664
rect 79926 239928 79982 239984
rect 80202 238976 80258 239032
rect 79282 238568 79338 238624
rect 80202 237616 80258 237672
rect 80202 236936 80258 236992
rect 80202 236120 80258 236176
rect 60698 232992 60754 233048
rect 61158 224288 61214 224344
rect 62906 224288 62962 224344
rect 87378 241968 87434 242024
rect 131814 244996 131816 245016
rect 131816 244996 131868 245016
rect 131868 244996 131870 245016
rect 131814 244960 131870 244996
rect 131630 244552 131686 244608
rect 131538 244144 131594 244200
rect 131354 243872 131410 243928
rect 131446 243464 131502 243520
rect 131538 243056 131594 243112
rect 131446 242648 131502 242704
rect 131354 242260 131410 242296
rect 131354 242240 131356 242260
rect 131356 242240 131408 242260
rect 131408 242240 131410 242260
rect 131354 241968 131410 242024
rect 73670 232992 73726 233048
rect 51958 216128 52014 216184
rect 38250 211232 38306 211288
rect 38158 203344 38214 203400
rect 139726 256248 139782 256304
rect 139634 255568 139690 255624
rect 140002 256928 140058 256984
rect 139910 254888 139966 254944
rect 139818 254344 139874 254400
rect 139634 253664 139690 253720
rect 140370 260872 140426 260928
rect 172846 260736 172902 260792
rect 140554 260192 140610 260248
rect 173582 260076 173638 260112
rect 173582 260056 173584 260076
rect 173584 260056 173636 260076
rect 173636 260056 173638 260076
rect 173398 259396 173454 259432
rect 173398 259376 173400 259396
rect 173400 259376 173452 259396
rect 173452 259376 173454 259396
rect 173582 258716 173638 258752
rect 173582 258696 173584 258716
rect 173584 258696 173636 258716
rect 173636 258696 173638 258716
rect 173306 258036 173362 258072
rect 173306 258016 173308 258036
rect 173308 258016 173360 258036
rect 173360 258016 173362 258036
rect 173582 257356 173638 257392
rect 173582 257336 173584 257356
rect 173584 257336 173636 257356
rect 173636 257336 173638 257356
rect 173122 256792 173178 256848
rect 173306 256132 173362 256168
rect 173306 256112 173308 256132
rect 173308 256112 173360 256132
rect 173360 256112 173362 256132
rect 173214 255432 173270 255488
rect 173490 254752 173546 254808
rect 181770 258288 181826 258344
rect 225194 280728 225250 280784
rect 233474 263864 233530 263920
rect 234302 262640 234358 262696
rect 234118 261960 234174 262016
rect 233474 260600 233530 260656
rect 225286 257608 225342 257664
rect 181954 257472 182010 257528
rect 223538 257472 223594 257528
rect 182322 257064 182378 257120
rect 182230 256656 182286 256712
rect 226206 256792 226262 256848
rect 225378 256384 225434 256440
rect 182046 256248 182102 256304
rect 226298 255976 226354 256032
rect 181862 255432 181918 255488
rect 182322 255568 182378 255624
rect 182230 255024 182286 255080
rect 226298 255724 226354 255760
rect 226298 255704 226300 255724
rect 226300 255704 226352 255724
rect 226352 255704 226354 255724
rect 225562 254888 225618 254944
rect 226390 255296 226446 255352
rect 225930 254480 225986 254536
rect 173214 254072 173270 254128
rect 182230 254344 182286 254400
rect 182046 253800 182102 253856
rect 182322 253936 182378 253992
rect 226298 254108 226300 254128
rect 226300 254108 226352 254128
rect 226352 254108 226354 254128
rect 226298 254072 226354 254108
rect 233842 259920 233898 259976
rect 233566 258560 233622 258616
rect 233474 257880 233530 257936
rect 233474 257236 233476 257256
rect 233476 257236 233528 257256
rect 233528 257236 233530 257256
rect 233474 257200 233530 257236
rect 233474 256520 233530 256576
rect 234670 261280 234726 261336
rect 234762 259240 234818 259296
rect 233934 255840 233990 255896
rect 233750 255160 233806 255216
rect 233566 254480 233622 254536
rect 226298 253800 226354 253856
rect 233474 253800 233530 253856
rect 173490 253392 173546 253448
rect 182138 253392 182194 253448
rect 225930 253392 225986 253448
rect 140554 252984 140610 253040
rect 182322 253020 182324 253040
rect 182324 253020 182376 253040
rect 182376 253020 182378 253040
rect 182322 252984 182378 253020
rect 226298 253020 226300 253040
rect 226300 253020 226352 253040
rect 226352 253020 226354 253040
rect 226298 252984 226354 253020
rect 173582 252712 173638 252768
rect 181402 252576 181458 252632
rect 140186 252304 140242 252360
rect 173490 252032 173546 252088
rect 226298 252576 226354 252632
rect 226390 252168 226446 252224
rect 182322 251896 182378 251952
rect 225654 251896 225710 251952
rect 140646 251624 140702 251680
rect 140554 251080 140610 251136
rect 181770 251488 181826 251544
rect 173490 251352 173546 251408
rect 226298 251524 226300 251544
rect 226300 251524 226352 251544
rect 226352 251524 226354 251544
rect 226298 251488 226354 251524
rect 182322 251100 182378 251136
rect 182322 251080 182324 251100
rect 182324 251080 182376 251100
rect 182376 251080 182378 251100
rect 225378 251080 225434 251136
rect 182230 250980 182232 251000
rect 182232 250980 182284 251000
rect 182284 250980 182286 251000
rect 182230 250944 182286 250980
rect 233658 253140 233714 253176
rect 233658 253120 233660 253140
rect 233660 253120 233712 253140
rect 233712 253120 233714 253140
rect 233566 252440 233622 252496
rect 233474 251760 233530 251816
rect 233566 251080 233622 251136
rect 173582 250672 173638 250728
rect 226390 250672 226446 250728
rect 140554 250400 140610 250456
rect 233474 250400 233530 250456
rect 173674 250128 173730 250184
rect 140002 249720 140058 249776
rect 140462 249620 140464 249640
rect 140464 249620 140516 249640
rect 140516 249620 140518 249640
rect 140462 249584 140518 249620
rect 173582 249448 173638 249504
rect 140370 248768 140426 248824
rect 173214 248768 173270 248824
rect 140370 248088 140426 248144
rect 173582 248088 173638 248144
rect 140370 247408 140426 247464
rect 173214 247408 173270 247464
rect 140646 247000 140702 247056
rect 173582 246728 173638 246784
rect 139358 240336 139414 240392
rect 139634 243192 139690 243248
rect 140554 246084 140556 246104
rect 140556 246084 140608 246104
rect 140608 246084 140610 246104
rect 140554 246048 140610 246084
rect 140370 245504 140426 245560
rect 173582 246084 173584 246104
rect 173584 246084 173636 246104
rect 173636 246084 173638 246104
rect 173582 246048 173638 246084
rect 173490 245368 173546 245424
rect 173582 244724 173584 244744
rect 173584 244724 173636 244744
rect 173636 244724 173638 244744
rect 173582 244688 173638 244724
rect 140646 244552 140702 244608
rect 140186 244416 140242 244472
rect 172846 244008 172902 244064
rect 139726 243056 139782 243112
rect 172846 242104 172902 242160
rect 140554 242004 140556 242024
rect 140556 242004 140608 242024
rect 140608 242004 140610 242024
rect 140554 241968 140610 242004
rect 140186 241832 140242 241888
rect 139542 240608 139598 240664
rect 141014 240492 141070 240528
rect 141014 240472 141016 240492
rect 141016 240472 141068 240492
rect 141068 240472 141070 240492
rect 173582 242784 173638 242840
rect 173582 241424 173638 241480
rect 173674 240744 173730 240800
rect 173490 240064 173546 240120
rect 140554 239268 140610 239304
rect 140554 239248 140556 239268
rect 140556 239248 140608 239268
rect 140608 239248 140610 239268
rect 140646 239148 140648 239168
rect 140648 239148 140700 239168
rect 140700 239148 140702 239168
rect 140646 239112 140702 239148
rect 173674 238704 173730 238760
rect 139450 238568 139506 238624
rect 182230 250264 182286 250320
rect 226298 250284 226354 250320
rect 226298 250264 226300 250284
rect 226300 250264 226352 250284
rect 226352 250264 226354 250284
rect 181586 249584 181642 249640
rect 182322 249992 182378 250048
rect 225930 249992 225986 250048
rect 233474 249720 233530 249776
rect 226298 249604 226354 249640
rect 233566 249620 233568 249640
rect 233568 249620 233620 249640
rect 233620 249620 233622 249640
rect 226298 249584 226300 249604
rect 226300 249584 226352 249604
rect 226352 249584 226354 249604
rect 233566 249584 233622 249620
rect 182322 249176 182378 249232
rect 225562 249176 225618 249232
rect 181126 248768 181182 248824
rect 226390 248768 226446 248824
rect 181034 248360 181090 248416
rect 180850 247952 180906 248008
rect 180758 247136 180814 247192
rect 180666 246728 180722 246784
rect 180942 247544 180998 247600
rect 180850 245912 180906 245968
rect 173950 243328 174006 243384
rect 173858 239384 173914 239440
rect 173766 238024 173822 238080
rect 140554 237344 140610 237400
rect 173582 237380 173584 237400
rect 173584 237380 173636 237400
rect 173636 237380 173638 237400
rect 173582 237344 173638 237380
rect 140278 237208 140334 237264
rect 173398 236664 173454 236720
rect 139266 236392 139322 236448
rect 173582 236120 173638 236176
rect 137518 225512 137574 225568
rect 74038 202800 74094 202856
rect 51958 202120 52014 202176
rect 38158 194640 38214 194696
rect 81674 190424 81730 190480
rect 51314 189472 51370 189528
rect 38802 186788 38804 186808
rect 38804 186788 38856 186808
rect 38856 186788 38858 186808
rect 38802 186752 38858 186788
rect 59502 172608 59558 172664
rect 60698 172472 60754 172528
rect 60882 172744 60938 172800
rect 61894 172336 61950 172392
rect 62170 172200 62226 172256
rect 134574 211776 134630 211832
rect 137150 198856 137206 198912
rect 137426 201984 137482 202040
rect 137334 200488 137390 200544
rect 137242 197360 137298 197416
rect 137058 195728 137114 195784
rect 137426 194232 137482 194288
rect 136966 192600 137022 192656
rect 137426 191124 137482 191160
rect 137426 191104 137428 191124
rect 137428 191104 137480 191124
rect 137480 191104 137482 191124
rect 137426 189472 137482 189528
rect 137058 183216 137114 183272
rect 137426 187976 137482 188032
rect 137426 186344 137482 186400
rect 137426 184576 137482 184632
rect 137334 181720 137390 181776
rect 137426 180088 137482 180144
rect 137426 178592 137482 178648
rect 71002 172608 71058 172664
rect 73026 172744 73082 172800
rect 72382 172472 72438 172528
rect 75786 172336 75842 172392
rect 75050 172200 75106 172256
rect 46990 162816 47046 162872
rect 79650 166624 79706 166680
rect 79558 165944 79614 166000
rect 80018 169480 80074 169536
rect 79926 168392 79982 168448
rect 85538 174648 85594 174704
rect 80202 168936 80258 168992
rect 80110 167712 80166 167768
rect 79834 167168 79890 167224
rect 79742 165400 79798 165456
rect 80202 164856 80258 164912
rect 87194 164312 87250 164368
rect 80202 164040 80258 164096
rect 80202 163632 80258 163688
rect 132734 174648 132790 174704
rect 127306 174512 127362 174568
rect 113874 172336 113930 172392
rect 108446 172200 108502 172256
rect 131998 163632 132054 163688
rect 80110 163088 80166 163144
rect 87286 163260 87288 163280
rect 87288 163260 87340 163280
rect 87340 163260 87342 163280
rect 87286 163224 87342 163260
rect 87194 162816 87250 162872
rect 80202 162544 80258 162600
rect 87194 162408 87250 162464
rect 87286 162000 87342 162056
rect 80018 161592 80074 161648
rect 87286 161592 87342 161648
rect 80202 161320 80258 161376
rect 87194 161184 87250 161240
rect 80110 160776 80166 160832
rect 87378 160776 87434 160832
rect 47082 148808 47138 148864
rect 46990 144048 47046 144104
rect 38158 124736 38214 124792
rect 38342 117392 38398 117448
rect 87286 160368 87342 160424
rect 80202 160232 80258 160288
rect 87194 159980 87250 160016
rect 87194 159960 87196 159980
rect 87196 159960 87248 159980
rect 87248 159960 87250 159980
rect 80110 159552 80166 159608
rect 87194 159552 87250 159608
rect 87286 159144 87342 159200
rect 80202 159008 80258 159064
rect 87378 158736 87434 158792
rect 80202 158500 80204 158520
rect 80204 158500 80256 158520
rect 80256 158500 80258 158520
rect 80202 158464 80258 158500
rect 87286 158328 87342 158384
rect 87194 157920 87250 157976
rect 79466 157784 79522 157840
rect 87286 157512 87342 157568
rect 80202 157240 80258 157296
rect 87194 157104 87250 157160
rect 80110 156696 80166 156752
rect 87102 156696 87158 156752
rect 80202 156152 80258 156208
rect 87010 155608 87066 155664
rect 80110 155472 80166 155528
rect 86918 155200 86974 155256
rect 80202 154928 80258 154984
rect 86826 154792 86882 154848
rect 80110 154384 80166 154440
rect 80018 153704 80074 153760
rect 80202 153196 80204 153216
rect 80204 153196 80256 153216
rect 80256 153196 80258 153216
rect 80202 153160 80258 153196
rect 80202 152616 80258 152672
rect 80202 151664 80258 151720
rect 80110 151392 80166 151448
rect 80110 150848 80166 150904
rect 79742 147856 79798 147912
rect 79374 147312 79430 147368
rect 79282 146768 79338 146824
rect 80202 150304 80258 150360
rect 87378 156288 87434 156344
rect 87194 156016 87250 156072
rect 131814 156152 131870 156208
rect 131538 155336 131594 155392
rect 131354 154928 131410 154984
rect 87102 154384 87158 154440
rect 87194 153976 87250 154032
rect 131446 154248 131502 154304
rect 131354 153840 131410 153896
rect 87930 153568 87986 153624
rect 87562 153160 87618 153216
rect 87746 152752 87802 152808
rect 87378 151936 87434 151992
rect 87286 151528 87342 151584
rect 87194 151120 87250 151176
rect 87378 150712 87434 150768
rect 87286 150304 87342 150360
rect 87194 149896 87250 149952
rect 80110 149624 80166 149680
rect 88114 152344 88170 152400
rect 87470 149488 87526 149544
rect 131354 152244 131356 152264
rect 131356 152244 131408 152264
rect 131408 152244 131410 152264
rect 131354 152208 131410 152244
rect 131354 151800 131410 151856
rect 131446 151392 131502 151448
rect 131538 151120 131594 151176
rect 131354 150712 131410 150768
rect 131446 150304 131502 150360
rect 131354 149896 131410 149952
rect 80202 149080 80258 149136
rect 87194 148672 87250 148728
rect 80110 148536 80166 148592
rect 80018 146224 80074 146280
rect 79926 145544 79982 145600
rect 79834 145000 79890 145056
rect 80202 144456 80258 144512
rect 87286 148264 87342 148320
rect 80018 143232 80074 143288
rect 87378 147992 87434 148048
rect 80202 143776 80258 143832
rect 80110 142688 80166 142744
rect 131446 149488 131502 149544
rect 87562 149080 87618 149136
rect 131354 149080 131410 149136
rect 131630 148672 131686 148728
rect 131538 148264 131594 148320
rect 131354 147992 131410 148048
rect 109550 143912 109606 143968
rect 80202 142144 80258 142200
rect 58766 131128 58822 131184
rect 60514 131420 60570 131456
rect 60514 131400 60516 131420
rect 60516 131400 60568 131420
rect 60568 131400 60570 131420
rect 60882 131128 60938 131184
rect 61618 131420 61674 131456
rect 61618 131400 61620 131420
rect 61620 131400 61672 131420
rect 61672 131400 61674 131420
rect 132458 163224 132514 163280
rect 132550 162816 132606 162872
rect 132642 162408 132698 162464
rect 132642 162000 132698 162056
rect 132642 161592 132698 161648
rect 132550 161184 132606 161240
rect 133378 160776 133434 160832
rect 132458 160504 132514 160560
rect 132642 160096 132698 160152
rect 132550 159688 132606 159744
rect 132642 159300 132698 159336
rect 132642 159280 132644 159300
rect 132644 159280 132696 159300
rect 132696 159280 132698 159300
rect 132550 158872 132606 158928
rect 132458 158464 132514 158520
rect 132642 158076 132698 158112
rect 132642 158056 132644 158076
rect 132644 158056 132696 158076
rect 132696 158056 132698 158076
rect 132090 154520 132146 154576
rect 132274 155744 132330 155800
rect 132182 153432 132238 153488
rect 132550 157648 132606 157704
rect 132642 157376 132698 157432
rect 132550 156968 132606 157024
rect 132642 156580 132698 156616
rect 132642 156560 132644 156580
rect 132644 156560 132696 156580
rect 132696 156560 132698 156580
rect 132550 153024 132606 153080
rect 132458 152616 132514 152672
rect 137702 227008 137758 227064
rect 137702 223880 137758 223936
rect 137702 221704 137758 221760
rect 137610 220752 137666 220808
rect 137610 218848 137666 218904
rect 137518 172472 137574 172528
rect 137794 217624 137850 217680
rect 137794 215856 137850 215912
rect 137702 172608 137758 172664
rect 137886 214496 137942 214552
rect 137886 212320 137942 212376
rect 137978 211368 138034 211424
rect 137978 209328 138034 209384
rect 138070 208240 138126 208296
rect 138070 206200 138126 206256
rect 152974 230952 153030 231008
rect 153158 230952 153214 231008
rect 156010 232992 156066 233048
rect 169994 232992 170050 233048
rect 226298 248360 226354 248416
rect 233474 248360 233530 248416
rect 233566 248260 233568 248280
rect 233568 248260 233620 248280
rect 233620 248260 233622 248280
rect 233566 248224 233622 248260
rect 226390 247952 226446 248008
rect 226298 247700 226354 247736
rect 226298 247680 226300 247700
rect 226300 247680 226352 247700
rect 226352 247680 226354 247700
rect 225654 247272 225710 247328
rect 182322 246356 182324 246376
rect 182324 246356 182376 246376
rect 182376 246356 182378 246376
rect 182322 246320 182378 246356
rect 234486 247272 234542 247328
rect 226390 246864 226446 246920
rect 234394 246864 234450 246920
rect 226298 246456 226354 246512
rect 226298 246048 226354 246104
rect 226206 245776 226262 245832
rect 180942 245504 180998 245560
rect 225562 245368 225618 245424
rect 182230 245096 182286 245152
rect 182046 244688 182102 244744
rect 181218 243872 181274 243928
rect 180390 242648 180446 242704
rect 180298 242240 180354 242296
rect 181586 241968 181642 242024
rect 182138 243464 182194 243520
rect 233474 245912 233530 245968
rect 233566 245504 233622 245560
rect 226390 244960 226446 245016
rect 225746 244552 225802 244608
rect 182322 244280 182378 244336
rect 226298 244144 226354 244200
rect 226206 243872 226262 243928
rect 226482 243464 226538 243520
rect 182322 243056 182378 243112
rect 226298 243056 226354 243112
rect 226022 242648 226078 242704
rect 226390 242240 226446 242296
rect 226022 241968 226078 242024
rect 233658 244688 233714 244744
rect 233474 244144 233530 244200
rect 233474 243364 233476 243384
rect 233476 243364 233528 243384
rect 233528 243364 233530 243384
rect 233474 243328 233530 243364
rect 233566 242784 233622 242840
rect 233474 242004 233476 242024
rect 233476 242004 233528 242024
rect 233528 242004 233530 242024
rect 233474 241968 233530 242004
rect 233474 239112 233530 239168
rect 233658 241424 233714 241480
rect 233750 240608 233806 240664
rect 264662 242240 264718 242296
rect 233842 240064 233898 240120
rect 233566 238704 233622 238760
rect 233474 237752 233530 237808
rect 233566 237344 233622 237400
rect 234118 236392 234174 236448
rect 203114 233672 203170 233728
rect 231082 221840 231138 221896
rect 148742 221568 148798 221624
rect 145614 219256 145670 219312
rect 145614 216944 145670 217000
rect 230990 218984 231046 219040
rect 175514 215756 175516 215776
rect 175516 215756 175568 215776
rect 175568 215756 175570 215776
rect 175514 215720 175570 215756
rect 145614 214360 145670 214416
rect 145614 212184 145670 212240
rect 145614 209872 145670 209928
rect 145798 207424 145854 207480
rect 138162 205112 138218 205168
rect 145614 205112 145670 205168
rect 138162 203480 138218 203536
rect 145522 202800 145578 202856
rect 144418 200488 144474 200544
rect 145614 198040 145670 198096
rect 145614 195728 145670 195784
rect 231726 220752 231782 220808
rect 231634 214496 231690 214552
rect 231542 211368 231598 211424
rect 231450 208240 231506 208296
rect 231358 205112 231414 205168
rect 231358 203480 231414 203536
rect 145798 193416 145854 193472
rect 167878 192736 167934 192792
rect 231266 191104 231322 191160
rect 145154 190832 145210 190888
rect 175514 190832 175570 190888
rect 145614 188656 145670 188712
rect 144786 186344 144842 186400
rect 145798 183352 145854 183408
rect 139634 169480 139690 169536
rect 139634 168836 139636 168856
rect 139636 168836 139688 168856
rect 139688 168836 139690 168856
rect 139634 168800 139690 168836
rect 139726 167032 139782 167088
rect 139634 166488 139690 166544
rect 139082 165672 139138 165728
rect 138990 164992 139046 165048
rect 139358 159688 139414 159744
rect 139174 158056 139230 158112
rect 139450 159416 139506 159472
rect 139542 156696 139598 156752
rect 139818 161048 139874 161104
rect 139266 150032 139322 150088
rect 139818 155744 139874 155800
rect 139726 155200 139782 155256
rect 139634 154792 139690 154848
rect 139726 154112 139782 154168
rect 139634 150712 139690 150768
rect 139910 152752 139966 152808
rect 140186 156988 140242 157024
rect 140186 156968 140188 156988
rect 140188 156968 140240 156988
rect 140240 156968 140242 156988
rect 140094 153432 140150 153488
rect 140002 152072 140058 152128
rect 140186 151392 140242 151448
rect 138898 144048 138954 144104
rect 139726 148164 139728 148184
rect 139728 148164 139780 148184
rect 139780 148164 139782 148184
rect 139726 148128 139782 148164
rect 139726 146788 139782 146824
rect 139726 146768 139728 146788
rect 139728 146768 139780 146788
rect 139780 146768 139782 146788
rect 139910 145428 139966 145464
rect 139910 145408 139912 145428
rect 139912 145408 139964 145428
rect 139964 145408 139966 145428
rect 139726 142688 139782 142744
rect 139634 142144 139690 142200
rect 230806 183216 230862 183272
rect 154630 172880 154686 172936
rect 154262 172744 154318 172800
rect 157574 172608 157630 172664
rect 157942 172472 157998 172528
rect 158310 172472 158366 172528
rect 231266 181720 231322 181776
rect 164474 172472 164530 172528
rect 166314 172880 166370 172936
rect 165854 172744 165910 172800
rect 170178 172336 170234 172392
rect 169994 172200 170050 172256
rect 140830 167712 140886 167768
rect 140370 164312 140426 164368
rect 140554 163768 140610 163824
rect 140646 163360 140702 163416
rect 140462 162544 140518 162600
rect 140554 162136 140610 162192
rect 140462 160776 140518 160832
rect 140370 158328 140426 158384
rect 140922 149352 140978 149408
rect 140738 148808 140794 148864
rect 140646 147448 140702 147504
rect 140554 146088 140610 146144
rect 140462 144728 140518 144784
rect 140370 143368 140426 143424
rect 136874 132932 136876 132952
rect 136876 132932 136928 132952
rect 136928 132932 136930 132952
rect 136874 132896 136930 132932
rect 136874 130040 136930 130096
rect 136874 127864 136930 127920
rect 47818 123240 47874 123296
rect 51314 122188 51316 122208
rect 51316 122188 51368 122208
rect 51368 122188 51370 122208
rect 38250 109368 38306 109424
rect 51314 122152 51370 122188
rect 137334 115236 137390 115272
rect 137334 115216 137336 115236
rect 137336 115216 137388 115236
rect 137388 115216 137390 115236
rect 74038 108960 74094 109016
rect 51314 108824 51370 108880
rect 47082 108280 47138 108336
rect 47818 108280 47874 108336
rect 38250 100664 38306 100720
rect 38802 92948 38804 92968
rect 38804 92948 38856 92968
rect 38856 92948 38858 92968
rect 38802 92912 38858 92948
rect 137886 127320 137942 127376
rect 137794 120520 137850 120576
rect 137702 117800 137758 117856
rect 137610 114808 137666 114864
rect 137518 111680 137574 111736
rect 137518 109640 137574 109696
rect 137426 100800 137482 100856
rect 137334 96992 137390 97048
rect 81674 96856 81730 96912
rect 51314 95496 51370 95552
rect 60790 78768 60846 78824
rect 61526 78632 61582 78688
rect 62078 78496 62134 78552
rect 62170 78360 62226 78416
rect 136874 85568 136930 85624
rect 136874 84652 136876 84672
rect 136876 84652 136928 84672
rect 136928 84652 136930 84672
rect 136874 84616 136930 84652
rect 85170 84072 85226 84128
rect 72474 78768 72530 78824
rect 73762 78632 73818 78688
rect 74498 78496 74554 78552
rect 75142 78360 75198 78416
rect 47082 61904 47138 61960
rect 79650 73192 79706 73248
rect 80202 75504 80258 75560
rect 80110 74960 80166 75016
rect 80018 74416 80074 74472
rect 79926 73872 79982 73928
rect 79834 72648 79890 72704
rect 79742 72104 79798 72160
rect 79558 71560 79614 71616
rect 80202 71016 80258 71072
rect 79466 69928 79522 69984
rect 80202 69792 80258 69848
rect 80202 68976 80258 69032
rect 80110 68432 80166 68488
rect 80202 68196 80204 68216
rect 80204 68196 80256 68216
rect 80256 68196 80258 68216
rect 80202 68160 80258 68196
rect 80202 67516 80204 67536
rect 80204 67516 80256 67536
rect 80256 67516 80258 67536
rect 80202 67480 80258 67516
rect 80110 66936 80166 66992
rect 80110 66392 80166 66448
rect 80202 65848 80258 65904
rect 80202 65340 80204 65360
rect 80204 65340 80256 65360
rect 80256 65340 80258 65360
rect 80202 65304 80258 65340
rect 80202 64660 80204 64680
rect 80204 64660 80256 64680
rect 80256 64660 80258 64680
rect 80202 64624 80258 64660
rect 80110 64080 80166 64136
rect 80202 63536 80258 63592
rect 80202 62992 80258 63048
rect 80202 62448 80258 62504
rect 80110 61768 80166 61824
rect 79098 60816 79154 60872
rect 80202 60680 80258 60736
rect 80110 60136 80166 60192
rect 80202 59592 80258 59648
rect 80110 58912 80166 58968
rect 80202 58404 80204 58424
rect 80204 58404 80256 58424
rect 80256 58404 80258 58424
rect 80202 58368 80258 58404
rect 80110 57824 80166 57880
rect 80202 57316 80204 57336
rect 80204 57316 80256 57336
rect 80256 57316 80258 57336
rect 80202 57280 80258 57316
rect 80202 56736 80258 56792
rect 80110 56056 80166 56112
rect 80018 55512 80074 55568
rect 80202 54968 80258 55024
rect 80110 54424 80166 54480
rect 80202 53880 80258 53936
rect 80202 53200 80258 53256
rect 79742 51024 79798 51080
rect 79466 50344 79522 50400
rect 80202 52656 80258 52712
rect 80110 52112 80166 52168
rect 80202 51588 80258 51624
rect 80202 51568 80204 51588
rect 80204 51568 80256 51588
rect 80256 51568 80258 51588
rect 80110 49392 80166 49448
rect 80202 49276 80258 49312
rect 80202 49256 80204 49276
rect 80204 49256 80256 49276
rect 80256 49256 80258 49276
rect 80018 48712 80074 48768
rect 79558 47488 79614 47544
rect 112954 78360 113010 78416
rect 133378 83664 133434 83720
rect 125558 81216 125614 81272
rect 87194 69656 87250 69712
rect 131354 69656 131410 69712
rect 87194 69248 87250 69304
rect 131354 69248 131410 69304
rect 87286 68840 87342 68896
rect 131446 68840 131502 68896
rect 87194 68432 87250 68488
rect 131538 68432 131594 68488
rect 87194 68024 87250 68080
rect 131998 68024 132054 68080
rect 87286 67616 87342 67672
rect 87194 67208 87250 67264
rect 132550 67616 132606 67672
rect 131814 67208 131870 67264
rect 87286 66800 87342 66856
rect 131354 66800 131410 66856
rect 131354 66392 131410 66448
rect 87286 66120 87342 66176
rect 87194 65984 87250 66040
rect 132182 65984 132238 66040
rect 87194 65576 87250 65632
rect 131354 65576 131410 65632
rect 131354 65204 131356 65224
rect 131356 65204 131408 65224
rect 131408 65204 131410 65224
rect 131354 65168 131410 65204
rect 87286 64896 87342 64952
rect 87194 64780 87250 64816
rect 87194 64760 87196 64780
rect 87196 64760 87248 64780
rect 87248 64760 87250 64780
rect 131446 64760 131502 64816
rect 87654 64352 87710 64408
rect 131814 64352 131870 64408
rect 87194 63672 87250 63728
rect 131814 63964 131870 64000
rect 131814 63944 131816 63964
rect 131816 63944 131868 63964
rect 131868 63944 131870 63964
rect 131354 63536 131410 63592
rect 87286 63264 87342 63320
rect 87194 62856 87250 62912
rect 87010 62720 87066 62776
rect 86918 60544 86974 60600
rect 86826 60000 86882 60056
rect 131354 63128 131410 63184
rect 131998 62720 132054 62776
rect 87286 62312 87342 62368
rect 131446 62312 131502 62368
rect 87194 61768 87250 61824
rect 87102 61360 87158 61416
rect 87010 60136 87066 60192
rect 131354 62040 131410 62096
rect 131354 61632 131410 61688
rect 87194 60952 87250 61008
rect 131446 60952 131502 61008
rect 131354 60816 131410 60872
rect 131354 60136 131410 60192
rect 131814 60020 131870 60056
rect 131814 60000 131816 60020
rect 131816 60000 131868 60020
rect 131868 60000 131870 60020
rect 87378 59320 87434 59376
rect 131538 59320 131594 59376
rect 87286 58912 87342 58968
rect 87194 58776 87250 58832
rect 87010 58096 87066 58152
rect 86734 57280 86790 57336
rect 86550 57144 86606 57200
rect 87102 57688 87158 57744
rect 131446 58912 131502 58968
rect 131354 58776 131410 58832
rect 131538 58096 131594 58152
rect 131446 57552 131502 57608
rect 131630 57688 131686 57744
rect 131354 57144 131410 57200
rect 88206 56464 88262 56520
rect 131446 56464 131502 56520
rect 87930 55920 87986 55976
rect 87286 55240 87342 55296
rect 87194 54832 87250 54888
rect 87286 54444 87342 54480
rect 87286 54424 87288 54444
rect 87288 54424 87340 54444
rect 87340 54424 87342 54444
rect 87102 54288 87158 54344
rect 87194 53336 87250 53392
rect 88390 56056 88446 56112
rect 131354 55920 131410 55976
rect 131538 56056 131594 56112
rect 131538 55240 131594 55296
rect 131446 54832 131502 54888
rect 131354 54696 131410 54752
rect 131446 54288 131502 54344
rect 104582 53744 104638 53800
rect 131354 53472 131410 53528
rect 129514 27496 129570 27552
rect 88482 26816 88538 26872
rect 138898 130856 138954 130912
rect 138162 125008 138218 125064
rect 137978 124192 138034 124248
rect 138162 122052 138164 122072
rect 138164 122052 138216 122072
rect 138216 122052 138218 122072
rect 138162 122016 138218 122052
rect 137886 108144 137942 108200
rect 137978 106648 138034 106704
rect 138162 118344 138218 118400
rect 138162 112632 138218 112688
rect 138070 105288 138126 105344
rect 137794 103928 137850 103984
rect 137702 102160 137758 102216
rect 138162 99168 138218 99224
rect 138162 95632 138218 95688
rect 138162 93884 138218 93920
rect 138162 93864 138164 93884
rect 138164 93864 138216 93884
rect 138216 93864 138218 93884
rect 137794 92676 137796 92696
rect 137796 92676 137848 92696
rect 137848 92676 137850 92696
rect 137794 92640 137850 92676
rect 137610 91416 137666 91472
rect 138162 89140 138164 89160
rect 138164 89140 138216 89160
rect 138216 89140 138218 89160
rect 138162 89104 138218 89140
rect 137610 88152 137666 88208
rect 134850 78496 134906 78552
rect 171374 169480 171430 169536
rect 170730 169208 170786 169264
rect 173306 168392 173362 168448
rect 173306 167304 173362 167360
rect 173122 166760 173178 166816
rect 173122 166216 173178 166272
rect 173030 164448 173086 164504
rect 172938 162836 172994 162872
rect 172938 162816 172940 162836
rect 172940 162816 172992 162836
rect 172992 162816 172994 162836
rect 172938 162292 172994 162328
rect 172938 162272 172940 162292
rect 172940 162272 172992 162292
rect 172992 162272 172994 162292
rect 172754 160504 172810 160560
rect 173214 163904 173270 163960
rect 172938 157784 172994 157840
rect 173306 159980 173362 160016
rect 173306 159960 173308 159980
rect 173308 159960 173360 159980
rect 173360 159960 173362 159980
rect 173122 158872 173178 158928
rect 173306 158328 173362 158384
rect 173214 157240 173270 157296
rect 173122 156696 173178 156752
rect 173122 154420 173124 154440
rect 173124 154420 173176 154440
rect 173176 154420 173178 154440
rect 173122 154384 173178 154420
rect 172938 153840 172994 153896
rect 173306 152752 173362 152808
rect 173306 151664 173362 151720
rect 172938 149896 172994 149952
rect 172754 147176 172810 147232
rect 172754 145952 172810 146008
rect 170546 139832 170602 139888
rect 173306 142688 173362 142744
rect 174042 167868 174098 167904
rect 174042 167848 174044 167868
rect 174044 167848 174096 167868
rect 174096 167848 174098 167868
rect 174042 165672 174098 165728
rect 173950 164992 174006 165048
rect 174042 163396 174044 163416
rect 174044 163396 174096 163416
rect 174096 163396 174098 163416
rect 174042 163360 174098 163396
rect 173950 161728 174006 161784
rect 174042 161184 174098 161240
rect 174042 159436 174098 159472
rect 174042 159416 174044 159436
rect 174044 159416 174096 159436
rect 174096 159416 174098 159436
rect 174042 156152 174098 156208
rect 173950 155472 174006 155528
rect 173950 154964 173952 154984
rect 173952 154964 174004 154984
rect 174004 154964 174006 154984
rect 173950 154928 174006 154964
rect 174042 153332 174044 153352
rect 174044 153332 174096 153352
rect 174096 153332 174098 153352
rect 174042 153296 174098 153332
rect 174042 152244 174044 152264
rect 174044 152244 174096 152264
rect 174096 152244 174098 152264
rect 174042 152208 174098 152244
rect 173950 150984 174006 151040
rect 174042 150440 174098 150496
rect 174042 149388 174044 149408
rect 174044 149388 174096 149408
rect 174096 149388 174098 149408
rect 174042 149352 174098 149388
rect 174042 148844 174044 148864
rect 174044 148844 174096 148864
rect 174096 148844 174098 148864
rect 174042 148808 174098 148844
rect 173858 148264 173914 148320
rect 174042 147756 174044 147776
rect 174044 147756 174096 147776
rect 174096 147756 174098 147776
rect 174042 147720 174098 147756
rect 173674 145428 173730 145464
rect 173674 145408 173676 145428
rect 173676 145408 173728 145428
rect 173728 145408 173730 145428
rect 173582 144864 173638 144920
rect 173490 143776 173546 143832
rect 174042 146496 174098 146552
rect 180942 163224 180998 163280
rect 180298 155608 180354 155664
rect 180574 156696 180630 156752
rect 180482 149488 180538 149544
rect 180390 149080 180446 149136
rect 180758 157920 180814 157976
rect 180666 149896 180722 149952
rect 181126 162816 181182 162872
rect 181034 159552 181090 159608
rect 180942 157512 180998 157568
rect 180850 156288 180906 156344
rect 181218 162408 181274 162464
rect 181402 161184 181458 161240
rect 207898 172200 207954 172256
rect 218662 172336 218718 172392
rect 181770 163632 181826 163688
rect 181402 160368 181458 160424
rect 181310 159960 181366 160016
rect 181494 159144 181550 159200
rect 181034 155200 181090 155256
rect 181034 154792 181090 154848
rect 181218 154384 181274 154440
rect 181126 153976 181182 154032
rect 181034 153160 181090 153216
rect 181678 153568 181734 153624
rect 181218 152752 181274 152808
rect 181126 152344 181182 152400
rect 181034 151528 181090 151584
rect 182322 162036 182324 162056
rect 182324 162036 182376 162056
rect 182376 162036 182378 162056
rect 182322 162000 182378 162036
rect 182322 161592 182378 161648
rect 181770 151936 181826 151992
rect 181126 151120 181182 151176
rect 182138 160776 182194 160832
rect 182138 158736 182194 158792
rect 182046 157104 182102 157160
rect 181954 156016 182010 156072
rect 181862 150304 181918 150360
rect 181770 148264 181826 148320
rect 182322 158328 182378 158384
rect 182046 150712 182102 150768
rect 182322 148672 182378 148728
rect 182322 148028 182324 148048
rect 182324 148028 182376 148048
rect 182376 148028 182378 148048
rect 182322 147992 182378 148028
rect 173950 144320 174006 144376
rect 173858 143232 173914 143288
rect 173398 142144 173454 142200
rect 232002 227008 232058 227064
rect 231910 225532 231966 225568
rect 231910 225512 231912 225532
rect 231912 225512 231964 225532
rect 231964 225512 231966 225532
rect 232002 223880 232058 223936
rect 231818 217624 231874 217680
rect 232002 216012 232058 216048
rect 232002 215992 232004 216012
rect 232004 215992 232056 216012
rect 232056 215992 232058 216012
rect 231726 201984 231782 202040
rect 231818 200488 231874 200544
rect 231634 197360 231690 197416
rect 231542 195728 231598 195784
rect 231450 192600 231506 192656
rect 232002 212340 232058 212376
rect 232002 212320 232004 212340
rect 232004 212320 232056 212340
rect 232056 212320 232058 212340
rect 232002 209464 232058 209520
rect 232002 206492 232058 206528
rect 232002 206472 232004 206492
rect 232004 206472 232056 206492
rect 232056 206472 232058 206492
rect 231910 198856 231966 198912
rect 231726 189472 231782 189528
rect 232002 194232 232058 194288
rect 231818 187976 231874 188032
rect 231818 186344 231874 186400
rect 231818 184848 231874 184904
rect 231634 180088 231690 180144
rect 231634 178592 231690 178648
rect 225930 163632 225986 163688
rect 226390 163224 226446 163280
rect 228690 163360 228746 163416
rect 228874 163360 228930 163416
rect 225562 162408 225618 162464
rect 226482 162816 226538 162872
rect 225930 162000 225986 162056
rect 226482 161628 226484 161648
rect 226484 161628 226536 161648
rect 226536 161628 226538 161648
rect 226482 161592 226538 161628
rect 226482 161184 226538 161240
rect 225930 160776 225986 160832
rect 226482 160540 226484 160560
rect 226484 160540 226536 160560
rect 226536 160540 226538 160560
rect 226482 160504 226538 160540
rect 225562 160096 225618 160152
rect 225930 159688 225986 159744
rect 226482 159280 226538 159336
rect 226482 158908 226484 158928
rect 226484 158908 226536 158928
rect 226536 158908 226538 158928
rect 226482 158872 226538 158908
rect 225562 158464 225618 158520
rect 226390 158056 226446 158112
rect 226298 157684 226300 157704
rect 226300 157684 226352 157704
rect 226352 157684 226354 157704
rect 226298 157648 226354 157684
rect 226482 157412 226484 157432
rect 226484 157412 226536 157432
rect 226536 157412 226538 157432
rect 226482 157376 226538 157412
rect 226482 156988 226538 157024
rect 226482 156968 226484 156988
rect 226484 156968 226536 156988
rect 226536 156968 226538 156988
rect 225378 156580 225434 156616
rect 225378 156560 225380 156580
rect 225380 156560 225432 156580
rect 225432 156560 225434 156580
rect 226482 156152 226538 156208
rect 226482 155744 226538 155800
rect 225562 155356 225618 155392
rect 225562 155336 225564 155356
rect 225564 155336 225616 155356
rect 225616 155336 225618 155356
rect 225746 154928 225802 154984
rect 226114 154520 226170 154576
rect 225838 154248 225894 154304
rect 226482 153840 226538 153896
rect 226114 153452 226170 153488
rect 226114 153432 226116 153452
rect 226116 153432 226168 153452
rect 226168 153432 226170 153452
rect 225746 153024 225802 153080
rect 225378 152636 225434 152672
rect 225378 152616 225380 152636
rect 225380 152616 225432 152636
rect 225432 152616 225434 152636
rect 225930 152208 225986 152264
rect 226114 151800 226170 151856
rect 225378 151412 225434 151448
rect 225378 151392 225380 151412
rect 225380 151392 225432 151412
rect 225432 151392 225434 151412
rect 226482 151140 226538 151176
rect 226482 151120 226484 151140
rect 226484 151120 226536 151140
rect 226536 151120 226538 151140
rect 225562 150712 225618 150768
rect 225746 150304 225802 150360
rect 226482 149896 226538 149952
rect 225562 149488 225618 149544
rect 225378 149100 225434 149136
rect 225378 149080 225380 149100
rect 225380 149080 225432 149100
rect 225432 149080 225434 149100
rect 226482 148692 226538 148728
rect 226482 148672 226484 148692
rect 226484 148672 226536 148692
rect 226536 148672 226538 148692
rect 226482 148284 226538 148320
rect 226482 148264 226484 148284
rect 226484 148264 226536 148284
rect 226536 148264 226538 148284
rect 225562 147992 225618 148048
rect 228414 153704 228470 153760
rect 228690 153704 228746 153760
rect 144602 96992 144658 97048
rect 145246 92368 145302 92424
rect 145246 89376 145302 89432
rect 148742 127456 148798 127512
rect 145614 125280 145670 125336
rect 145614 122968 145670 123024
rect 145614 120520 145670 120576
rect 240926 218732 240982 218768
rect 240926 218712 240928 218732
rect 240928 218712 240980 218732
rect 240980 218712 240982 218732
rect 240466 216264 240522 216320
rect 240926 213816 240982 213872
rect 240926 211912 240982 211968
rect 240466 209192 240522 209248
rect 264202 233672 264258 233728
rect 261166 212728 261222 212784
rect 262362 212728 262418 212784
rect 240650 206744 240706 206800
rect 240926 204860 240982 204896
rect 240926 204840 240928 204860
rect 240928 204840 240980 204860
rect 240980 204840 240982 204860
rect 240374 202392 240430 202448
rect 240466 199808 240522 199864
rect 240926 198040 240982 198096
rect 240926 195204 240982 195240
rect 240926 195184 240928 195204
rect 240928 195184 240980 195204
rect 240980 195184 240982 195204
rect 240466 192736 240522 192792
rect 240650 190288 240706 190344
rect 240742 188268 240798 188304
rect 240742 188248 240744 188268
rect 240744 188248 240796 188268
rect 240796 188248 240798 188268
rect 240926 185800 240982 185856
rect 239638 183352 239694 183408
rect 249482 172472 249538 172528
rect 249942 172744 249998 172800
rect 251046 172608 251102 172664
rect 262362 192736 262418 192792
rect 261074 172744 261130 172800
rect 261442 172472 261498 172528
rect 262546 172608 262602 172664
rect 264202 172336 264258 172392
rect 263834 172200 263890 172256
rect 233474 169480 233530 169536
rect 233474 168836 233476 168856
rect 233476 168836 233528 168856
rect 233528 168836 233530 168856
rect 233474 168800 233530 168836
rect 233658 168120 233714 168176
rect 233474 166896 233530 166952
rect 233474 166236 233530 166272
rect 233474 166216 233476 166236
rect 233476 166216 233528 166236
rect 233528 166216 233530 166236
rect 233566 165672 233622 165728
rect 233474 164992 233530 165048
rect 236694 167508 236750 167564
rect 233750 164312 233806 164368
rect 233566 163088 233622 163144
rect 233474 162408 233530 162464
rect 233474 161184 233530 161240
rect 233658 161864 233714 161920
rect 233566 160504 233622 160560
rect 233474 159960 233530 160016
rect 233842 163768 233898 163824
rect 233566 159280 233622 159336
rect 233474 158600 233530 158656
rect 233474 158056 233530 158112
rect 233474 157412 233476 157432
rect 233476 157412 233528 157432
rect 233528 157412 233530 157432
rect 233474 157376 233530 157412
rect 233474 156696 233530 156752
rect 233474 156152 233530 156208
rect 233474 155472 233530 155528
rect 233566 154792 233622 154848
rect 233474 154112 233530 154168
rect 233566 153568 233622 153624
rect 233474 152888 233530 152944
rect 233658 152208 233714 152264
rect 233750 151664 233806 151720
rect 233566 150984 233622 151040
rect 233474 150304 233530 150360
rect 233842 149760 233898 149816
rect 233474 149080 233530 149136
rect 233566 148400 233622 148456
rect 233474 147856 233530 147912
rect 233566 147176 233622 147232
rect 233474 146496 233530 146552
rect 233474 145952 233530 146008
rect 233474 145308 233476 145328
rect 233476 145308 233528 145328
rect 233528 145308 233530 145328
rect 233474 145272 233530 145308
rect 233658 144592 233714 144648
rect 233750 144048 233806 144104
rect 233934 143368 233990 143424
rect 233842 142688 233898 142744
rect 233474 142144 233530 142200
rect 232830 139832 232886 139888
rect 167234 118752 167290 118808
rect 167878 118752 167934 118808
rect 145614 118208 145670 118264
rect 145614 115896 145670 115952
rect 145614 113448 145670 113504
rect 145614 111136 145670 111192
rect 145614 108824 145670 108880
rect 145614 106512 145670 106568
rect 145430 103928 145486 103984
rect 145614 101752 145670 101808
rect 145614 99440 145670 99496
rect 146350 94680 146406 94736
rect 155366 79176 155422 79232
rect 155274 78632 155330 78688
rect 156010 79312 156066 79368
rect 167878 98760 167934 98816
rect 167326 78632 167382 78688
rect 170086 78496 170142 78552
rect 169074 78360 169130 78416
rect 168614 77816 168670 77872
rect 169994 76048 170050 76104
rect 139634 75504 139690 75560
rect 140922 74824 140978 74880
rect 139634 74144 139690 74200
rect 139726 73464 139782 73520
rect 139634 72920 139690 72976
rect 139634 72240 139690 72296
rect 139910 71560 139966 71616
rect 139818 70880 139874 70936
rect 139726 70200 139782 70256
rect 139634 69656 139690 69712
rect 139726 68976 139782 69032
rect 139634 68296 139690 68352
rect 139634 67616 139690 67672
rect 139726 66936 139782 66992
rect 139726 66392 139782 66448
rect 139634 65712 139690 65768
rect 139726 65032 139782 65088
rect 139634 64352 139690 64408
rect 139726 63672 139782 63728
rect 139634 63128 139690 63184
rect 139726 62448 139782 62504
rect 139634 61768 139690 61824
rect 139634 61088 139690 61144
rect 139634 60564 139690 60600
rect 139634 60544 139636 60564
rect 139636 60544 139688 60564
rect 139688 60544 139690 60564
rect 139726 59864 139782 59920
rect 139634 59184 139690 59240
rect 139726 58504 139782 58560
rect 139634 57824 139690 57880
rect 139726 57280 139782 57336
rect 139634 55920 139690 55976
rect 139818 56600 139874 56656
rect 139726 55240 139782 55296
rect 139910 54560 139966 54616
rect 139542 52656 139598 52712
rect 139450 51976 139506 52032
rect 139726 54016 139782 54072
rect 139634 51296 139690 51352
rect 139634 50072 139690 50128
rect 139726 49392 139782 49448
rect 140002 53336 140058 53392
rect 139910 50752 139966 50808
rect 139818 48712 139874 48768
rect 139634 48168 139690 48224
rect 170638 74688 170694 74744
rect 170822 74688 170878 74744
rect 170730 74144 170786 74200
rect 173306 73328 173362 73384
rect 173490 71288 173546 71344
rect 173674 72240 173730 72296
rect 173950 72784 174006 72840
rect 173858 71696 173914 71752
rect 173766 70744 173822 70800
rect 173582 70200 173638 70256
rect 174042 69656 174098 69712
rect 173306 69112 173362 69168
rect 172846 68568 172902 68624
rect 174042 68024 174098 68080
rect 173950 67480 174006 67536
rect 173490 66936 173546 66992
rect 173582 65984 173638 66040
rect 174042 66564 174044 66584
rect 174044 66564 174096 66584
rect 174096 66564 174098 66584
rect 174042 66528 174098 66564
rect 173858 65440 173914 65496
rect 173490 64896 173546 64952
rect 173766 64352 173822 64408
rect 173858 63264 173914 63320
rect 174042 63844 174044 63864
rect 174044 63844 174096 63864
rect 174096 63844 174098 63864
rect 174042 63808 174098 63844
rect 173950 62720 174006 62776
rect 173306 62176 173362 62232
rect 173766 61768 173822 61824
rect 173950 61224 174006 61280
rect 174042 60680 174098 60736
rect 173674 60136 173730 60192
rect 173674 59048 173730 59104
rect 174042 59592 174098 59648
rect 173858 58504 173914 58560
rect 174042 57960 174098 58016
rect 173766 57416 173822 57472
rect 174042 57028 174098 57064
rect 174042 57008 174044 57028
rect 174044 57008 174096 57028
rect 174096 57008 174098 57028
rect 174042 56464 174098 56520
rect 172938 55920 172994 55976
rect 173306 55376 173362 55432
rect 173766 54832 173822 54888
rect 174042 54324 174044 54344
rect 174044 54324 174096 54344
rect 174096 54324 174098 54344
rect 174042 54288 174098 54324
rect 174042 53780 174044 53800
rect 174044 53780 174096 53800
rect 174096 53780 174098 53800
rect 174042 53744 174098 53780
rect 173490 53200 173546 53256
rect 173950 52692 173952 52712
rect 173952 52692 174004 52712
rect 174004 52692 174006 52712
rect 173950 52656 174006 52692
rect 174042 52248 174098 52304
rect 172846 51704 172902 51760
rect 172938 51196 172940 51216
rect 172940 51196 172992 51216
rect 172992 51196 172994 51216
rect 172938 51160 172994 51196
rect 173950 50616 174006 50672
rect 173306 50108 173308 50128
rect 173308 50108 173360 50128
rect 173360 50108 173362 50128
rect 173306 50072 173362 50108
rect 172754 49528 172810 49584
rect 173122 48984 173178 49040
rect 173306 48440 173362 48496
rect 173398 48032 173454 48088
rect 156562 45992 156618 46048
rect 101730 12128 101786 12184
rect 230714 127864 230770 127920
rect 175514 121916 175516 121936
rect 175516 121916 175568 121936
rect 175568 121916 175570 121936
rect 175514 121880 175570 121916
rect 228506 120248 228562 120304
rect 231266 115236 231322 115272
rect 231266 115216 231268 115236
rect 231268 115216 231320 115236
rect 231320 115216 231322 115236
rect 231358 114808 231414 114864
rect 231358 112360 231414 112416
rect 175514 96992 175570 97048
rect 231266 100800 231322 100856
rect 182138 83664 182194 83720
rect 181770 69656 181826 69712
rect 202470 81216 202526 81272
rect 210566 81352 210622 81408
rect 226022 69656 226078 69712
rect 182322 68976 182378 69032
rect 226022 69248 226078 69304
rect 225746 68840 225802 68896
rect 181770 68568 181826 68624
rect 181586 68160 181642 68216
rect 226298 68432 226354 68488
rect 182322 67752 182378 67808
rect 182230 67344 182286 67400
rect 181402 66800 181458 66856
rect 226298 68024 226354 68080
rect 225562 67616 225618 67672
rect 225470 67208 225526 67264
rect 182322 66936 182378 66992
rect 225838 66800 225894 66856
rect 226022 66392 226078 66448
rect 182322 66120 182378 66176
rect 181402 65712 181458 65768
rect 181310 65576 181366 65632
rect 181034 64896 181090 64952
rect 181126 64488 181182 64544
rect 226298 65984 226354 66040
rect 226390 65576 226446 65632
rect 226298 65168 226354 65224
rect 226298 64780 226354 64816
rect 226298 64760 226300 64780
rect 226300 64760 226352 64780
rect 226352 64760 226354 64780
rect 181402 64352 181458 64408
rect 226390 64352 226446 64408
rect 226390 63944 226446 64000
rect 182322 63672 182378 63728
rect 182046 63264 182102 63320
rect 181770 62312 181826 62368
rect 181678 60952 181734 61008
rect 180942 59592 180998 59648
rect 180298 57688 180354 57744
rect 181862 61768 181918 61824
rect 181954 61360 182010 61416
rect 182138 62856 182194 62912
rect 182230 62720 182286 62776
rect 226298 63536 226354 63592
rect 226298 63128 226354 63184
rect 226298 62720 226354 62776
rect 226390 62312 226446 62368
rect 226206 62040 226262 62096
rect 226298 61632 226354 61688
rect 225746 61224 225802 61280
rect 182138 60544 182194 60600
rect 182046 58504 182102 58560
rect 182230 60136 182286 60192
rect 182322 60000 182378 60056
rect 225930 60816 225986 60872
rect 226390 60408 226446 60464
rect 226298 60036 226300 60056
rect 226300 60036 226352 60056
rect 226352 60036 226354 60056
rect 226298 60000 226354 60036
rect 226206 59592 226262 59648
rect 182230 58912 182286 58968
rect 181678 57688 181734 57744
rect 181586 57300 181642 57336
rect 181586 57280 181588 57300
rect 181588 57280 181640 57300
rect 181640 57280 181642 57300
rect 181310 56464 181366 56520
rect 181218 56056 181274 56112
rect 181126 55240 181182 55296
rect 180942 53064 180998 53120
rect 226390 59184 226446 59240
rect 226298 58776 226354 58832
rect 225746 58368 225802 58424
rect 182322 58096 182378 58152
rect 183702 57416 183758 57472
rect 225930 57960 225986 58016
rect 225838 57552 225894 57608
rect 226482 57180 226484 57200
rect 226484 57180 226536 57200
rect 226536 57180 226538 57200
rect 183702 57076 183758 57132
rect 226482 57144 226538 57180
rect 225930 56736 225986 56792
rect 182322 55920 182378 55976
rect 226298 56328 226354 56384
rect 226298 55940 226354 55976
rect 226298 55920 226300 55940
rect 226300 55920 226352 55940
rect 226352 55920 226354 55940
rect 225746 55512 225802 55568
rect 181678 54832 181734 54888
rect 226390 55104 226446 55160
rect 226298 54716 226354 54752
rect 226298 54696 226300 54716
rect 226300 54696 226352 54716
rect 226352 54696 226354 54716
rect 181586 54444 181642 54480
rect 181586 54424 181588 54444
rect 181588 54424 181640 54444
rect 181640 54424 181642 54444
rect 182322 54288 182378 54344
rect 226298 54288 226354 54344
rect 225838 54016 225894 54072
rect 215534 34432 215590 34488
rect 231726 127048 231782 127104
rect 231634 125144 231690 125200
rect 231634 122052 231636 122072
rect 231636 122052 231688 122072
rect 231688 122052 231690 122072
rect 231634 122016 231690 122052
rect 231910 132932 231912 132952
rect 231912 132932 231964 132952
rect 231964 132932 231966 132952
rect 231910 132896 231966 132932
rect 232738 130856 232794 130912
rect 232002 130212 232004 130232
rect 232004 130212 232056 130232
rect 232056 130212 232058 130232
rect 232002 130176 232058 130212
rect 231818 124192 231874 124248
rect 231726 120520 231782 120576
rect 231634 118752 231690 118808
rect 231542 117528 231598 117584
rect 231450 111680 231506 111736
rect 231542 109640 231598 109696
rect 231726 108008 231782 108064
rect 231818 106648 231874 106704
rect 231634 103928 231690 103984
rect 231542 102296 231598 102352
rect 231450 96992 231506 97048
rect 231910 105288 231966 105344
rect 232002 99168 232058 99224
rect 231726 95632 231782 95688
rect 231818 94172 231820 94192
rect 231820 94172 231872 94192
rect 231872 94172 231874 94192
rect 231818 94136 231874 94172
rect 231450 92948 231452 92968
rect 231452 92948 231504 92968
rect 231504 92948 231506 92968
rect 231450 92912 231506 92948
rect 231450 91416 231506 91472
rect 231634 89784 231690 89840
rect 231634 88288 231690 88344
rect 231634 86012 231636 86032
rect 231636 86012 231688 86032
rect 231688 86012 231690 86032
rect 231634 85976 231690 86012
rect 231634 84652 231636 84672
rect 231636 84652 231688 84672
rect 231688 84652 231690 84672
rect 231634 84616 231690 84652
rect 263282 139832 263338 139888
rect 264570 138608 264626 138664
rect 240926 125144 240982 125200
rect 240926 122832 240982 122888
rect 261074 120656 261130 120712
rect 240926 120384 240982 120440
rect 261074 118752 261130 118808
rect 240926 118072 240982 118128
rect 240926 115760 240982 115816
rect 240742 113312 240798 113368
rect 240926 111020 240982 111056
rect 240926 111000 240928 111020
rect 240928 111000 240980 111020
rect 240980 111000 240982 111020
rect 240834 108688 240890 108744
rect 240926 106376 240982 106432
rect 240742 103928 240798 103984
rect 240374 101616 240430 101672
rect 240834 99304 240890 99360
rect 262362 98760 262418 98816
rect 240926 96856 240982 96912
rect 240926 94544 240982 94600
rect 240926 92232 240982 92288
rect 240926 89920 240982 89976
rect 247090 78632 247146 78688
rect 248562 78904 248618 78960
rect 249114 78360 249170 78416
rect 249666 78496 249722 78552
rect 249850 78768 249906 78824
rect 251414 86420 251416 86440
rect 251416 86420 251468 86440
rect 251468 86420 251470 86440
rect 251414 86384 251470 86420
rect 256566 86384 256622 86440
rect 258314 78632 258370 78688
rect 259786 78904 259842 78960
rect 261074 78768 261130 78824
rect 261442 78496 261498 78552
rect 261994 78360 262050 78416
rect 233474 75504 233530 75560
rect 233474 74960 233530 75016
rect 233566 74280 233622 74336
rect 233658 73736 233714 73792
rect 234118 72648 234174 72704
rect 233474 72512 233530 72568
rect 233566 71424 233622 71480
rect 233474 71016 233530 71072
rect 233658 70200 233714 70256
rect 233750 69520 233806 69576
rect 233658 68976 233714 69032
rect 233566 68296 233622 68352
rect 233474 68160 233530 68216
rect 233566 67072 233622 67128
rect 233474 66936 233530 66992
rect 233474 66120 233530 66176
rect 233474 65440 233530 65496
rect 233566 64780 233622 64816
rect 233566 64760 233568 64780
rect 233568 64760 233620 64780
rect 233620 64760 233622 64780
rect 233474 64488 233530 64544
rect 233474 63420 233530 63456
rect 233474 63400 233476 63420
rect 233476 63400 233528 63420
rect 233528 63400 233530 63420
rect 233658 63264 233714 63320
rect 233566 62720 233622 62776
rect 233474 62176 233530 62232
rect 233474 61496 233530 61552
rect 233474 60952 233530 61008
rect 233566 60272 233622 60328
rect 233474 59728 233530 59784
rect 233566 59048 233622 59104
rect 233474 57280 233530 57336
rect 233566 56600 233622 56656
rect 233750 58504 233806 58560
rect 233842 57824 233898 57880
rect 233658 56056 233714 56112
rect 233474 55376 233530 55432
rect 233566 54832 233622 54888
rect 233474 54152 233530 54208
rect 233566 53608 233622 53664
rect 233474 52948 233530 52984
rect 233474 52928 233476 52948
rect 233476 52928 233528 52948
rect 233528 52928 233530 52948
rect 233474 51704 233530 51760
rect 233474 51160 233530 51216
rect 233474 49256 233530 49312
rect 233658 52384 233714 52440
rect 233658 50480 233714 50536
rect 233658 49936 233714 49992
rect 233566 48712 233622 48768
rect 233474 47624 233530 47680
rect 241202 47488 241258 47544
rect 250494 45856 250550 45912
rect 223538 27496 223594 27552
rect 211946 12264 212002 12320
rect 276162 217624 276218 217680
rect 265214 216536 265270 216592
rect 274874 208376 274930 208432
rect 274874 197632 274930 197688
rect 275518 188112 275574 188168
rect 264846 163224 264902 163280
rect 264754 149352 264810 149408
rect 264846 69384 264902 69440
rect 264754 55376 264810 55432
rect 276070 123648 276126 123704
rect 274874 114400 274930 114456
rect 274874 103656 274930 103712
rect 274874 94308 274876 94328
rect 274876 94308 274928 94328
rect 274928 94308 274930 94328
rect 274874 94272 274930 94308
rect 285914 181176 285970 181232
rect 289870 130312 289926 130368
rect 300358 290520 300414 290576
rect 300082 266040 300138 266096
rect 300174 241560 300230 241616
rect 300174 217116 300176 217136
rect 300176 217116 300228 217136
rect 300228 217116 300230 217136
rect 300174 217080 300230 217116
rect 296218 202800 296274 202856
rect 293550 188948 293606 188984
rect 293550 188928 293552 188948
rect 293552 188928 293604 188948
rect 293604 188928 293606 188948
rect 300174 168120 300230 168176
rect 300174 143504 300230 143560
rect 300174 119024 300230 119080
rect 293550 109504 293606 109560
rect 285914 87336 285970 87392
rect 295574 95496 295630 95552
rect 299714 94544 299770 94600
rect 300450 202256 300506 202312
rect 300450 192600 300506 192656
rect 300174 70064 300230 70120
rect 300174 45584 300230 45640
rect 299806 21104 299862 21160
<< metal3 >>
rect 300353 290578 300419 290581
rect 303416 290578 303896 290608
rect 300353 290576 303896 290578
rect 300353 290520 300358 290576
rect 300414 290520 303896 290576
rect 300353 290518 303896 290520
rect 300353 290515 300419 290518
rect 303416 290488 303896 290518
rect 129742 288266 129802 288848
rect 223582 288268 223642 288848
rect 131390 288266 131396 288268
rect 129742 288206 131396 288266
rect 131390 288204 131396 288206
rect 131460 288204 131466 288268
rect 223574 288204 223580 288268
rect 223644 288204 223650 288268
rect 13313 287858 13379 287861
rect 90174 287858 90180 287860
rect 13313 287856 90180 287858
rect 13313 287800 13318 287856
rect 13374 287800 90180 287856
rect 13313 287798 90180 287800
rect 13313 287795 13379 287798
rect 90174 287796 90180 287798
rect 90244 287796 90250 287860
rect 129550 287796 129556 287860
rect 129620 287858 129626 287860
rect 184198 287858 184204 287860
rect 129620 287798 184204 287858
rect 129620 287796 129626 287798
rect 184198 287796 184204 287798
rect 184268 287796 184274 287860
rect 9896 286498 10376 286528
rect 13221 286498 13287 286501
rect 9896 286496 13287 286498
rect 9896 286440 13226 286496
rect 13282 286440 13287 286496
rect 9896 286438 13287 286440
rect 9896 286408 10376 286438
rect 13221 286435 13287 286438
rect 88477 284866 88543 284869
rect 89998 284866 90058 284904
rect 88477 284864 90058 284866
rect 88477 284808 88482 284864
rect 88538 284808 90058 284864
rect 88477 284806 90058 284808
rect 182317 284866 182383 284869
rect 184022 284866 184082 284904
rect 182317 284864 184082 284866
rect 182317 284808 182322 284864
rect 182378 284808 184082 284864
rect 182317 284806 184082 284808
rect 88477 284803 88543 284806
rect 182317 284803 182383 284806
rect 129742 280786 129802 280824
rect 131349 280786 131415 280789
rect 129742 280784 131415 280786
rect 129742 280728 131354 280784
rect 131410 280728 131415 280784
rect 129742 280726 131415 280728
rect 223766 280786 223826 280824
rect 225189 280786 225255 280789
rect 223766 280784 225255 280786
rect 223766 280728 225194 280784
rect 225250 280728 225255 280784
rect 223766 280726 225255 280728
rect 131349 280723 131415 280726
rect 225189 280723 225255 280726
rect 300077 266098 300143 266101
rect 303416 266098 303896 266128
rect 300077 266096 303896 266098
rect 300077 266040 300082 266096
rect 300138 266040 303896 266096
rect 300077 266038 303896 266040
rect 300077 266035 300143 266038
rect 303416 266008 303896 266038
rect 52454 265492 52460 265556
rect 52524 265554 52530 265556
rect 62901 265554 62967 265557
rect 52524 265552 62967 265554
rect 52524 265496 62906 265552
rect 62962 265496 62967 265552
rect 52524 265494 62967 265496
rect 52524 265492 52530 265494
rect 62901 265491 62967 265494
rect 233469 263922 233535 263925
rect 233469 263920 237074 263922
rect 233469 263864 233474 263920
rect 233530 263864 237074 263920
rect 233469 263862 237074 263864
rect 233469 263859 233535 263862
rect 52270 263724 52276 263788
rect 52340 263786 52346 263788
rect 78909 263786 78975 263789
rect 52340 263784 78975 263786
rect 52340 263728 78914 263784
rect 78970 263728 78975 263784
rect 52340 263726 78975 263728
rect 52340 263724 52346 263726
rect 76750 263552 76810 263726
rect 78909 263723 78975 263726
rect 142246 263724 142252 263788
rect 142316 263786 142322 263788
rect 142316 263726 170466 263786
rect 142316 263724 142322 263726
rect 139629 263514 139695 263517
rect 139629 263512 143020 263514
rect 139629 263456 139634 263512
rect 139690 263456 143020 263512
rect 170406 263484 170466 263726
rect 139629 263454 143020 263456
rect 139629 263451 139695 263454
rect 237014 263416 237074 263862
rect 79553 263378 79619 263381
rect 76750 263376 79619 263378
rect 76750 263320 79558 263376
rect 79614 263320 79619 263376
rect 76750 263318 79619 263320
rect 76750 262872 76810 263318
rect 79553 263315 79619 263318
rect 143033 263242 143099 263245
rect 142990 263240 143099 263242
rect 142990 263184 143038 263240
rect 143094 263184 143099 263240
rect 142990 263179 143099 263184
rect 142990 262872 143050 263179
rect 173393 262834 173459 262837
rect 170804 262832 173459 262834
rect 170804 262776 173398 262832
rect 173454 262776 173459 262832
rect 170804 262774 173459 262776
rect 173393 262771 173459 262774
rect 139629 262698 139695 262701
rect 234297 262698 234363 262701
rect 139629 262696 143050 262698
rect 139629 262640 139634 262696
rect 139690 262640 143050 262696
rect 139629 262638 143050 262640
rect 139629 262635 139695 262638
rect 142990 262192 143050 262638
rect 234297 262696 237044 262698
rect 234297 262640 234302 262696
rect 234358 262640 237044 262696
rect 234297 262638 237044 262640
rect 234297 262635 234363 262638
rect 80105 262154 80171 262157
rect 173669 262154 173735 262157
rect 76780 262152 80171 262154
rect 76780 262096 80110 262152
rect 80166 262096 80171 262152
rect 76780 262094 80171 262096
rect 170804 262152 173735 262154
rect 170804 262096 173674 262152
rect 173730 262096 173735 262152
rect 170804 262094 173735 262096
rect 80105 262091 80171 262094
rect 173669 262091 173735 262094
rect 234113 262018 234179 262021
rect 234113 262016 237044 262018
rect 234113 261960 234118 262016
rect 234174 261960 237044 262016
rect 234113 261958 237044 261960
rect 234113 261955 234179 261958
rect 80197 261474 80263 261477
rect 76780 261472 80263 261474
rect 76780 261416 80202 261472
rect 80258 261416 80263 261472
rect 76780 261414 80263 261416
rect 80197 261411 80263 261414
rect 140273 261474 140339 261477
rect 173577 261474 173643 261477
rect 140273 261472 143020 261474
rect 140273 261416 140278 261472
rect 140334 261416 143020 261472
rect 140273 261414 143020 261416
rect 170804 261472 173643 261474
rect 170804 261416 173582 261472
rect 173638 261416 173643 261472
rect 170804 261414 173643 261416
rect 140273 261411 140339 261414
rect 173577 261411 173643 261414
rect 234665 261338 234731 261341
rect 234665 261336 237044 261338
rect 234665 261280 234670 261336
rect 234726 261280 237044 261336
rect 234665 261278 237044 261280
rect 234665 261275 234731 261278
rect 140365 260930 140431 260933
rect 140365 260928 143020 260930
rect 140365 260872 140370 260928
rect 140426 260872 143020 260928
rect 140365 260870 143020 260872
rect 140365 260867 140431 260870
rect 80105 260794 80171 260797
rect 172841 260794 172907 260797
rect 76780 260792 80171 260794
rect 76780 260736 80110 260792
rect 80166 260736 80171 260792
rect 76780 260734 80171 260736
rect 170804 260792 172907 260794
rect 170804 260736 172846 260792
rect 172902 260736 172907 260792
rect 170804 260734 172907 260736
rect 80105 260731 80171 260734
rect 172841 260731 172907 260734
rect 233469 260658 233535 260661
rect 233469 260656 237044 260658
rect 233469 260600 233474 260656
rect 233530 260600 237044 260656
rect 233469 260598 237044 260600
rect 233469 260595 233535 260598
rect 140549 260250 140615 260253
rect 140549 260248 143020 260250
rect 140549 260192 140554 260248
rect 140610 260192 143020 260248
rect 140549 260190 143020 260192
rect 140549 260187 140615 260190
rect 80197 260114 80263 260117
rect 173577 260114 173643 260117
rect 76780 260112 80263 260114
rect 76780 260056 80202 260112
rect 80258 260056 80263 260112
rect 76780 260054 80263 260056
rect 170804 260112 173643 260114
rect 170804 260056 173582 260112
rect 173638 260056 173643 260112
rect 170804 260054 173643 260056
rect 80197 260051 80263 260054
rect 173577 260051 173643 260054
rect 233837 259978 233903 259981
rect 233837 259976 237044 259978
rect 233837 259920 233842 259976
rect 233898 259920 237044 259976
rect 233837 259918 237044 259920
rect 233837 259915 233903 259918
rect 140089 259570 140155 259573
rect 140089 259568 143020 259570
rect 140089 259512 140094 259568
rect 140150 259512 143020 259568
rect 140089 259510 143020 259512
rect 140089 259507 140155 259510
rect 79829 259434 79895 259437
rect 173393 259434 173459 259437
rect 76780 259432 79895 259434
rect 76780 259376 79834 259432
rect 79890 259376 79895 259432
rect 76780 259374 79895 259376
rect 170804 259432 173459 259434
rect 170804 259376 173398 259432
rect 173454 259376 173459 259432
rect 170804 259374 173459 259376
rect 79829 259371 79895 259374
rect 173393 259371 173459 259374
rect 234757 259298 234823 259301
rect 234757 259296 237044 259298
rect 234757 259240 234762 259296
rect 234818 259240 237044 259296
rect 234757 259238 237044 259240
rect 234757 259235 234823 259238
rect 139905 258890 139971 258893
rect 139905 258888 143020 258890
rect 139905 258832 139910 258888
rect 139966 258832 143020 258888
rect 139905 258830 143020 258832
rect 139905 258827 139971 258830
rect 80197 258754 80263 258757
rect 173577 258754 173643 258757
rect 76780 258752 80263 258754
rect 76780 258696 80202 258752
rect 80258 258696 80263 258752
rect 76780 258694 80263 258696
rect 170804 258752 173643 258754
rect 170804 258696 173582 258752
rect 173638 258696 173643 258752
rect 170804 258694 173643 258696
rect 80197 258691 80263 258694
rect 173577 258691 173643 258694
rect 233561 258618 233627 258621
rect 233561 258616 237044 258618
rect 233561 258560 233566 258616
rect 233622 258560 237044 258616
rect 233561 258558 237044 258560
rect 233561 258555 233627 258558
rect 87189 258346 87255 258349
rect 181765 258346 181831 258349
rect 87189 258344 90058 258346
rect 87189 258288 87194 258344
rect 87250 258288 90058 258344
rect 87189 258286 90058 258288
rect 87189 258283 87255 258286
rect 80013 258074 80079 258077
rect 76780 258072 80079 258074
rect 76780 258016 80018 258072
rect 80074 258016 80079 258072
rect 76780 258014 80079 258016
rect 80013 258011 80079 258014
rect 89998 257704 90058 258286
rect 181765 258344 184082 258346
rect 181765 258288 181770 258344
rect 181826 258288 184082 258344
rect 181765 258286 184082 258288
rect 181765 258283 181831 258286
rect 139813 258210 139879 258213
rect 139813 258208 143020 258210
rect 139813 258152 139818 258208
rect 139874 258152 143020 258208
rect 139813 258150 143020 258152
rect 139813 258147 139879 258150
rect 173301 258074 173367 258077
rect 170804 258072 173367 258074
rect 170804 258016 173306 258072
rect 173362 258016 173367 258072
rect 170804 258014 173367 258016
rect 173301 258011 173367 258014
rect 184022 257704 184082 258286
rect 233469 257938 233535 257941
rect 233469 257936 237044 257938
rect 233469 257880 233474 257936
rect 233530 257880 237044 257936
rect 233469 257878 237044 257880
rect 233469 257875 233535 257878
rect 131349 257666 131415 257669
rect 129772 257664 131415 257666
rect 129772 257608 131354 257664
rect 131410 257608 131415 257664
rect 129772 257606 131415 257608
rect 131349 257603 131415 257606
rect 139629 257666 139695 257669
rect 225281 257666 225347 257669
rect 226334 257666 226340 257668
rect 139629 257664 143020 257666
rect 139629 257608 139634 257664
rect 139690 257608 143020 257664
rect 139629 257606 143020 257608
rect 223796 257664 226340 257666
rect 223796 257608 225286 257664
rect 225342 257608 226340 257664
rect 223796 257606 226340 257608
rect 139629 257603 139695 257606
rect 225281 257603 225347 257606
rect 226334 257604 226340 257606
rect 226404 257604 226410 257668
rect 87281 257530 87347 257533
rect 129509 257530 129575 257533
rect 181949 257530 182015 257533
rect 223533 257530 223599 257533
rect 87281 257528 90058 257530
rect 87281 257472 87286 257528
rect 87342 257472 90058 257528
rect 87281 257470 90058 257472
rect 87281 257467 87347 257470
rect 80197 257394 80263 257397
rect 76780 257392 80263 257394
rect 76780 257336 80202 257392
rect 80258 257336 80263 257392
rect 76780 257334 80263 257336
rect 80197 257331 80263 257334
rect 89998 257296 90058 257470
rect 129509 257528 129618 257530
rect 129509 257472 129514 257528
rect 129570 257472 129618 257528
rect 129509 257467 129618 257472
rect 181949 257528 184082 257530
rect 181949 257472 181954 257528
rect 182010 257472 184082 257528
rect 181949 257470 184082 257472
rect 181949 257467 182015 257470
rect 129558 257296 129618 257467
rect 173577 257394 173643 257397
rect 170804 257392 173643 257394
rect 170804 257336 173582 257392
rect 173638 257336 173643 257392
rect 170804 257334 173643 257336
rect 173577 257331 173643 257334
rect 184022 257296 184082 257470
rect 223533 257528 223642 257530
rect 223533 257472 223538 257528
rect 223594 257472 223642 257528
rect 223533 257467 223642 257472
rect 223582 257228 223642 257467
rect 233469 257258 233535 257261
rect 233469 257256 237044 257258
rect 233469 257200 233474 257256
rect 233530 257200 237044 257256
rect 233469 257198 237044 257200
rect 233469 257195 233535 257198
rect 182317 257122 182383 257125
rect 182317 257120 184082 257122
rect 182317 257064 182322 257120
rect 182378 257064 184082 257120
rect 182317 257062 184082 257064
rect 182317 257059 182383 257062
rect 139997 256986 140063 256989
rect 139997 256984 143020 256986
rect 139997 256928 140002 256984
rect 140058 256928 143020 256984
rect 139997 256926 143020 256928
rect 139997 256923 140063 256926
rect 184022 256888 184082 257062
rect 80105 256850 80171 256853
rect 76780 256848 80171 256850
rect 76780 256792 80110 256848
rect 80166 256792 80171 256848
rect 76780 256790 80171 256792
rect 80105 256787 80171 256790
rect 87281 256850 87347 256853
rect 131349 256850 131415 256853
rect 173117 256850 173183 256853
rect 226201 256850 226267 256853
rect 265158 256850 265164 256852
rect 87281 256848 90028 256850
rect 87281 256792 87286 256848
rect 87342 256792 90028 256848
rect 87281 256790 90028 256792
rect 129772 256848 131415 256850
rect 129772 256792 131354 256848
rect 131410 256792 131415 256848
rect 129772 256790 131415 256792
rect 170804 256848 173183 256850
rect 170804 256792 173122 256848
rect 173178 256792 173183 256848
rect 170804 256790 173183 256792
rect 223796 256848 226267 256850
rect 223796 256792 226206 256848
rect 226262 256792 226267 256848
rect 223796 256790 226267 256792
rect 264828 256790 265164 256850
rect 87281 256787 87347 256790
rect 131349 256787 131415 256790
rect 173117 256787 173183 256790
rect 226201 256787 226267 256790
rect 265158 256788 265164 256790
rect 265228 256788 265234 256852
rect 87557 256714 87623 256717
rect 131441 256714 131507 256717
rect 87557 256712 90058 256714
rect 87557 256656 87562 256712
rect 87618 256656 90058 256712
rect 87557 256654 90058 256656
rect 87557 256651 87623 256654
rect 89998 256480 90058 256654
rect 129742 256712 131507 256714
rect 129742 256656 131446 256712
rect 131502 256656 131507 256712
rect 129742 256654 131507 256656
rect 129742 256480 129802 256654
rect 131441 256651 131507 256654
rect 182225 256714 182291 256717
rect 182225 256712 184082 256714
rect 182225 256656 182230 256712
rect 182286 256656 184082 256712
rect 182225 256654 184082 256656
rect 182225 256651 182291 256654
rect 184022 256480 184082 256654
rect 233469 256578 233535 256581
rect 233469 256576 237044 256578
rect 233469 256520 233474 256576
rect 233530 256520 237044 256576
rect 233469 256518 237044 256520
rect 233469 256515 233535 256518
rect 225373 256442 225439 256445
rect 223796 256440 225439 256442
rect 223796 256384 225378 256440
rect 225434 256384 225439 256440
rect 223796 256382 225439 256384
rect 225373 256379 225439 256382
rect 87189 256306 87255 256309
rect 131533 256306 131599 256309
rect 87189 256304 90058 256306
rect 87189 256248 87194 256304
rect 87250 256248 90058 256304
rect 87189 256246 90058 256248
rect 87189 256243 87255 256246
rect 80197 256170 80263 256173
rect 76780 256168 80263 256170
rect 76780 256112 80202 256168
rect 80258 256112 80263 256168
rect 76780 256110 80263 256112
rect 80197 256107 80263 256110
rect 89998 256072 90058 256246
rect 129742 256304 131599 256306
rect 129742 256248 131538 256304
rect 131594 256248 131599 256304
rect 129742 256246 131599 256248
rect 129742 256072 129802 256246
rect 131533 256243 131599 256246
rect 139721 256306 139787 256309
rect 182041 256306 182107 256309
rect 139721 256304 143020 256306
rect 139721 256248 139726 256304
rect 139782 256248 143020 256304
rect 139721 256246 143020 256248
rect 182041 256304 184082 256306
rect 182041 256248 182046 256304
rect 182102 256248 184082 256304
rect 182041 256246 184082 256248
rect 139721 256243 139787 256246
rect 182041 256243 182107 256246
rect 173301 256170 173367 256173
rect 170804 256168 173367 256170
rect 170804 256112 173306 256168
rect 173362 256112 173367 256168
rect 170804 256110 173367 256112
rect 173301 256107 173367 256110
rect 184022 256072 184082 256246
rect 226293 256034 226359 256037
rect 223796 256032 226359 256034
rect 223796 255976 226298 256032
rect 226354 255976 226359 256032
rect 223796 255974 226359 255976
rect 226293 255971 226359 255974
rect 233929 255898 233995 255901
rect 233929 255896 237044 255898
rect 233929 255840 233934 255896
rect 233990 255840 237044 255896
rect 233929 255838 237044 255840
rect 233929 255835 233995 255838
rect 131349 255762 131415 255765
rect 226293 255762 226359 255765
rect 129772 255760 131415 255762
rect 129772 255704 131354 255760
rect 131410 255704 131415 255760
rect 129772 255702 131415 255704
rect 223796 255760 226359 255762
rect 223796 255704 226298 255760
rect 226354 255704 226359 255760
rect 223796 255702 226359 255704
rect 131349 255699 131415 255702
rect 226293 255699 226359 255702
rect 87373 255626 87439 255629
rect 139629 255626 139695 255629
rect 182317 255626 182383 255629
rect 87373 255624 90028 255626
rect 87373 255568 87378 255624
rect 87434 255568 90028 255624
rect 87373 255566 90028 255568
rect 139629 255624 143020 255626
rect 139629 255568 139634 255624
rect 139690 255568 143020 255624
rect 139629 255566 143020 255568
rect 182317 255624 184052 255626
rect 182317 255568 182322 255624
rect 182378 255568 184052 255624
rect 182317 255566 184052 255568
rect 87373 255563 87439 255566
rect 139629 255563 139695 255566
rect 182317 255563 182383 255566
rect 80105 255490 80171 255493
rect 76780 255488 80171 255490
rect 76780 255432 80110 255488
rect 80166 255432 80171 255488
rect 76780 255430 80171 255432
rect 80105 255427 80171 255430
rect 87189 255490 87255 255493
rect 173209 255490 173275 255493
rect 87189 255488 90058 255490
rect 87189 255432 87194 255488
rect 87250 255432 90058 255488
rect 87189 255430 90058 255432
rect 170804 255488 173275 255490
rect 170804 255432 173214 255488
rect 173270 255432 173275 255488
rect 170804 255430 173275 255432
rect 87189 255427 87255 255430
rect 89998 255256 90058 255430
rect 173209 255427 173275 255430
rect 181857 255490 181923 255493
rect 181857 255488 184082 255490
rect 181857 255432 181862 255488
rect 181918 255432 184082 255488
rect 181857 255430 184082 255432
rect 181857 255427 181923 255430
rect 131441 255354 131507 255357
rect 129772 255352 131507 255354
rect 129772 255296 131446 255352
rect 131502 255296 131507 255352
rect 129772 255294 131507 255296
rect 131441 255291 131507 255294
rect 184022 255256 184082 255430
rect 226385 255354 226451 255357
rect 223796 255352 226451 255354
rect 223796 255296 226390 255352
rect 226446 255296 226451 255352
rect 223796 255294 226451 255296
rect 226385 255291 226451 255294
rect 131533 255218 131599 255221
rect 129742 255216 131599 255218
rect 129742 255160 131538 255216
rect 131594 255160 131599 255216
rect 129742 255158 131599 255160
rect 87281 255082 87347 255085
rect 87281 255080 90058 255082
rect 87281 255024 87286 255080
rect 87342 255024 90058 255080
rect 87281 255022 90058 255024
rect 87281 255019 87347 255022
rect 89998 254848 90058 255022
rect 129742 254984 129802 255158
rect 131533 255155 131599 255158
rect 233745 255218 233811 255221
rect 233745 255216 237044 255218
rect 233745 255160 233750 255216
rect 233806 255160 237044 255216
rect 233745 255158 237044 255160
rect 233745 255155 233811 255158
rect 182225 255082 182291 255085
rect 182225 255080 184082 255082
rect 182225 255024 182230 255080
rect 182286 255024 184082 255080
rect 182225 255022 184082 255024
rect 182225 255019 182291 255022
rect 139905 254946 139971 254949
rect 139905 254944 143020 254946
rect 139905 254888 139910 254944
rect 139966 254888 143020 254944
rect 139905 254886 143020 254888
rect 139905 254883 139971 254886
rect 184022 254848 184082 255022
rect 225557 254946 225623 254949
rect 223796 254944 225623 254946
rect 223796 254888 225562 254944
rect 225618 254888 225623 254944
rect 223796 254886 225623 254888
rect 225557 254883 225623 254886
rect 80197 254810 80263 254813
rect 131625 254810 131691 254813
rect 173485 254810 173551 254813
rect 76780 254808 80263 254810
rect 76780 254752 80202 254808
rect 80258 254752 80263 254808
rect 76780 254750 80263 254752
rect 80197 254747 80263 254750
rect 129742 254808 131691 254810
rect 129742 254752 131630 254808
rect 131686 254752 131691 254808
rect 129742 254750 131691 254752
rect 170804 254808 173551 254810
rect 170804 254752 173490 254808
rect 173546 254752 173551 254808
rect 170804 254750 173551 254752
rect 129742 254576 129802 254750
rect 131625 254747 131691 254750
rect 173485 254747 173551 254750
rect 225925 254538 225991 254541
rect 223796 254536 225991 254538
rect 223796 254480 225930 254536
rect 225986 254480 225991 254536
rect 223796 254478 225991 254480
rect 225925 254475 225991 254478
rect 233561 254538 233627 254541
rect 233561 254536 237044 254538
rect 233561 254480 233566 254536
rect 233622 254480 237044 254536
rect 233561 254478 237044 254480
rect 233561 254475 233627 254478
rect 87189 254402 87255 254405
rect 139813 254402 139879 254405
rect 182225 254402 182291 254405
rect 87189 254400 90028 254402
rect 87189 254344 87194 254400
rect 87250 254344 90028 254400
rect 87189 254342 90028 254344
rect 139813 254400 143020 254402
rect 139813 254344 139818 254400
rect 139874 254344 143020 254400
rect 139813 254342 143020 254344
rect 182225 254400 184052 254402
rect 182225 254344 182230 254400
rect 182286 254344 184052 254400
rect 182225 254342 184052 254344
rect 87189 254339 87255 254342
rect 139813 254339 139879 254342
rect 182225 254339 182291 254342
rect 87281 254266 87347 254269
rect 87281 254264 90058 254266
rect 87281 254208 87286 254264
rect 87342 254208 90058 254264
rect 87281 254206 90058 254208
rect 87281 254203 87347 254206
rect 80105 254130 80171 254133
rect 76780 254128 80171 254130
rect 76780 254072 80110 254128
rect 80166 254072 80171 254128
rect 76780 254070 80171 254072
rect 80105 254067 80171 254070
rect 89998 254032 90058 254206
rect 131349 254130 131415 254133
rect 173209 254130 173275 254133
rect 226293 254130 226359 254133
rect 129772 254128 131415 254130
rect 129772 254072 131354 254128
rect 131410 254072 131415 254128
rect 129772 254070 131415 254072
rect 170804 254128 173275 254130
rect 170804 254072 173214 254128
rect 173270 254072 173275 254128
rect 170804 254070 173275 254072
rect 223796 254128 226359 254130
rect 223796 254072 226298 254128
rect 226354 254072 226359 254128
rect 223796 254070 226359 254072
rect 131349 254067 131415 254070
rect 173209 254067 173275 254070
rect 226293 254067 226359 254070
rect 182317 253994 182383 253997
rect 182317 253992 184052 253994
rect 182317 253936 182322 253992
rect 182378 253936 184052 253992
rect 182317 253934 184052 253936
rect 182317 253931 182383 253934
rect 9896 253858 10376 253888
rect 13681 253858 13747 253861
rect 9896 253856 13747 253858
rect 9896 253800 13686 253856
rect 13742 253800 13747 253856
rect 9896 253798 13747 253800
rect 9896 253768 10376 253798
rect 13681 253795 13747 253798
rect 87373 253858 87439 253861
rect 131533 253858 131599 253861
rect 87373 253856 90058 253858
rect 87373 253800 87378 253856
rect 87434 253800 90058 253856
rect 87373 253798 90058 253800
rect 129772 253856 131599 253858
rect 129772 253800 131538 253856
rect 131594 253800 131599 253856
rect 129772 253798 131599 253800
rect 87373 253795 87439 253798
rect 89998 253624 90058 253798
rect 131533 253795 131599 253798
rect 182041 253858 182107 253861
rect 226293 253858 226359 253861
rect 182041 253856 184082 253858
rect 182041 253800 182046 253856
rect 182102 253800 184082 253856
rect 182041 253798 184082 253800
rect 223796 253856 226359 253858
rect 223796 253800 226298 253856
rect 226354 253800 226359 253856
rect 223796 253798 226359 253800
rect 182041 253795 182107 253798
rect 131441 253722 131507 253725
rect 129742 253720 131507 253722
rect 129742 253664 131446 253720
rect 131502 253664 131507 253720
rect 129742 253662 131507 253664
rect 129742 253488 129802 253662
rect 131441 253659 131507 253662
rect 139629 253722 139695 253725
rect 139629 253720 143020 253722
rect 139629 253664 139634 253720
rect 139690 253664 143020 253720
rect 139629 253662 143020 253664
rect 139629 253659 139695 253662
rect 184022 253624 184082 253798
rect 226293 253795 226359 253798
rect 233469 253858 233535 253861
rect 233469 253856 237044 253858
rect 233469 253800 233474 253856
rect 233530 253800 237044 253856
rect 233469 253798 237044 253800
rect 233469 253795 233535 253798
rect 80197 253450 80263 253453
rect 76780 253448 80263 253450
rect 76780 253392 80202 253448
rect 80258 253392 80263 253448
rect 76780 253390 80263 253392
rect 80197 253387 80263 253390
rect 87189 253450 87255 253453
rect 173485 253450 173551 253453
rect 87189 253448 90058 253450
rect 87189 253392 87194 253448
rect 87250 253392 90058 253448
rect 87189 253390 90058 253392
rect 170804 253448 173551 253450
rect 170804 253392 173490 253448
rect 173546 253392 173551 253448
rect 170804 253390 173551 253392
rect 87189 253387 87255 253390
rect 89998 253216 90058 253390
rect 173485 253387 173551 253390
rect 182133 253450 182199 253453
rect 225925 253450 225991 253453
rect 182133 253448 184082 253450
rect 182133 253392 182138 253448
rect 182194 253392 184082 253448
rect 182133 253390 184082 253392
rect 223796 253448 225991 253450
rect 223796 253392 225930 253448
rect 225986 253392 225991 253448
rect 223796 253390 225991 253392
rect 182133 253387 182199 253390
rect 184022 253216 184082 253390
rect 225925 253387 225991 253390
rect 233653 253178 233719 253181
rect 233653 253176 237044 253178
rect 233653 253120 233658 253176
rect 233714 253120 237044 253176
rect 233653 253118 237044 253120
rect 233653 253115 233719 253118
rect 87189 253042 87255 253045
rect 131349 253042 131415 253045
rect 87189 253040 90058 253042
rect 87189 252984 87194 253040
rect 87250 252984 90058 253040
rect 87189 252982 90058 252984
rect 129772 253040 131415 253042
rect 129772 252984 131354 253040
rect 131410 252984 131415 253040
rect 129772 252982 131415 252984
rect 87189 252979 87255 252982
rect 89998 252808 90058 252982
rect 131349 252979 131415 252982
rect 140549 253042 140615 253045
rect 182317 253042 182383 253045
rect 226293 253042 226359 253045
rect 140549 253040 143020 253042
rect 140549 252984 140554 253040
rect 140610 252984 143020 253040
rect 140549 252982 143020 252984
rect 182317 253040 184082 253042
rect 182317 252984 182322 253040
rect 182378 252984 184082 253040
rect 182317 252982 184082 252984
rect 223796 253040 226359 253042
rect 223796 252984 226298 253040
rect 226354 252984 226359 253040
rect 223796 252982 226359 252984
rect 140549 252979 140615 252982
rect 182317 252979 182383 252982
rect 131441 252906 131507 252909
rect 129742 252904 131507 252906
rect 129742 252848 131446 252904
rect 131502 252848 131507 252904
rect 129742 252846 131507 252848
rect 80197 252770 80263 252773
rect 76780 252768 80263 252770
rect 76780 252712 80202 252768
rect 80258 252712 80263 252768
rect 76780 252710 80263 252712
rect 80197 252707 80263 252710
rect 129742 252672 129802 252846
rect 131441 252843 131507 252846
rect 184022 252808 184082 252982
rect 226293 252979 226359 252982
rect 173577 252770 173643 252773
rect 170804 252768 173643 252770
rect 170804 252712 173582 252768
rect 173638 252712 173643 252768
rect 170804 252710 173643 252712
rect 173577 252707 173643 252710
rect 87281 252634 87347 252637
rect 181397 252634 181463 252637
rect 226293 252634 226359 252637
rect 87281 252632 90058 252634
rect 87281 252576 87286 252632
rect 87342 252576 90058 252632
rect 87281 252574 90058 252576
rect 87281 252571 87347 252574
rect 89998 252400 90058 252574
rect 181397 252632 184082 252634
rect 181397 252576 181402 252632
rect 181458 252576 184082 252632
rect 181397 252574 184082 252576
rect 223796 252632 226359 252634
rect 223796 252576 226298 252632
rect 226354 252576 226359 252632
rect 223796 252574 226359 252576
rect 181397 252571 181463 252574
rect 131533 252498 131599 252501
rect 129742 252496 131599 252498
rect 129742 252440 131538 252496
rect 131594 252440 131599 252496
rect 129742 252438 131599 252440
rect 129742 252264 129802 252438
rect 131533 252435 131599 252438
rect 184022 252400 184082 252574
rect 226293 252571 226359 252574
rect 233561 252498 233627 252501
rect 233561 252496 237044 252498
rect 233561 252440 233566 252496
rect 233622 252440 237044 252496
rect 233561 252438 237044 252440
rect 233561 252435 233627 252438
rect 140181 252362 140247 252365
rect 140181 252360 143020 252362
rect 140181 252304 140186 252360
rect 140242 252304 143020 252360
rect 140181 252302 143020 252304
rect 140181 252299 140247 252302
rect 87189 252226 87255 252229
rect 226385 252226 226451 252229
rect 87189 252224 90058 252226
rect 87189 252168 87194 252224
rect 87250 252168 90058 252224
rect 87189 252166 90058 252168
rect 223796 252224 226451 252226
rect 223796 252168 226390 252224
rect 226446 252168 226451 252224
rect 223796 252166 226451 252168
rect 87189 252163 87255 252166
rect 80197 252090 80263 252093
rect 76780 252088 80263 252090
rect 76780 252032 80202 252088
rect 80258 252032 80263 252088
rect 76780 252030 80263 252032
rect 80197 252027 80263 252030
rect 89998 251992 90058 252166
rect 226385 252163 226451 252166
rect 173485 252090 173551 252093
rect 170804 252088 173551 252090
rect 170804 252032 173490 252088
rect 173546 252032 173551 252088
rect 170804 252030 173551 252032
rect 173485 252027 173551 252030
rect 131349 251954 131415 251957
rect 129772 251952 131415 251954
rect 129772 251896 131354 251952
rect 131410 251896 131415 251952
rect 129772 251894 131415 251896
rect 131349 251891 131415 251894
rect 182317 251954 182383 251957
rect 225649 251954 225715 251957
rect 182317 251952 184052 251954
rect 182317 251896 182322 251952
rect 182378 251896 184052 251952
rect 182317 251894 184052 251896
rect 223796 251952 225715 251954
rect 223796 251896 225654 251952
rect 225710 251896 225715 251952
rect 223796 251894 225715 251896
rect 182317 251891 182383 251894
rect 225649 251891 225715 251894
rect 233469 251818 233535 251821
rect 233469 251816 237044 251818
rect 233469 251760 233474 251816
rect 233530 251760 237044 251816
rect 233469 251758 237044 251760
rect 233469 251755 233535 251758
rect 140641 251682 140707 251685
rect 140641 251680 143020 251682
rect 140641 251624 140646 251680
rect 140702 251624 143020 251680
rect 140641 251622 143020 251624
rect 140641 251619 140707 251622
rect 87189 251546 87255 251549
rect 131349 251546 131415 251549
rect 87189 251544 90028 251546
rect 87189 251488 87194 251544
rect 87250 251488 90028 251544
rect 87189 251486 90028 251488
rect 129772 251544 131415 251546
rect 129772 251488 131354 251544
rect 131410 251488 131415 251544
rect 129772 251486 131415 251488
rect 87189 251483 87255 251486
rect 131349 251483 131415 251486
rect 181765 251546 181831 251549
rect 226293 251546 226359 251549
rect 181765 251544 184052 251546
rect 181765 251488 181770 251544
rect 181826 251488 184052 251544
rect 181765 251486 184052 251488
rect 223796 251544 226359 251546
rect 223796 251488 226298 251544
rect 226354 251488 226359 251544
rect 223796 251486 226359 251488
rect 181765 251483 181831 251486
rect 226293 251483 226359 251486
rect 80197 251410 80263 251413
rect 173485 251410 173551 251413
rect 76780 251408 80263 251410
rect 76780 251352 80202 251408
rect 80258 251352 80263 251408
rect 76780 251350 80263 251352
rect 170804 251408 173551 251410
rect 170804 251352 173490 251408
rect 173546 251352 173551 251408
rect 170804 251350 173551 251352
rect 80197 251347 80263 251350
rect 173485 251347 173551 251350
rect 87189 251138 87255 251141
rect 131349 251138 131415 251141
rect 87189 251136 90028 251138
rect 87189 251080 87194 251136
rect 87250 251080 90028 251136
rect 87189 251078 90028 251080
rect 129772 251136 131415 251138
rect 129772 251080 131354 251136
rect 131410 251080 131415 251136
rect 129772 251078 131415 251080
rect 87189 251075 87255 251078
rect 131349 251075 131415 251078
rect 140549 251138 140615 251141
rect 182317 251138 182383 251141
rect 225373 251138 225439 251141
rect 140549 251136 143020 251138
rect 140549 251080 140554 251136
rect 140610 251080 143020 251136
rect 140549 251078 143020 251080
rect 182317 251136 184052 251138
rect 182317 251080 182322 251136
rect 182378 251080 184052 251136
rect 182317 251078 184052 251080
rect 223796 251136 225439 251138
rect 223796 251080 225378 251136
rect 225434 251080 225439 251136
rect 223796 251078 225439 251080
rect 140549 251075 140615 251078
rect 182317 251075 182383 251078
rect 225373 251075 225439 251078
rect 233561 251138 233627 251141
rect 233561 251136 237044 251138
rect 233561 251080 233566 251136
rect 233622 251080 237044 251136
rect 233561 251078 237044 251080
rect 233561 251075 233627 251078
rect 87281 251002 87347 251005
rect 182225 251002 182291 251005
rect 87281 251000 90058 251002
rect 87281 250944 87286 251000
rect 87342 250944 90058 251000
rect 87281 250942 90058 250944
rect 87281 250939 87347 250942
rect 89998 250768 90058 250942
rect 182225 251000 184082 251002
rect 182225 250944 182230 251000
rect 182286 250944 184082 251000
rect 182225 250942 184082 250944
rect 182225 250939 182291 250942
rect 184022 250768 184082 250942
rect 80105 250730 80171 250733
rect 131441 250730 131507 250733
rect 173577 250730 173643 250733
rect 226385 250730 226451 250733
rect 76780 250728 80171 250730
rect 76780 250672 80110 250728
rect 80166 250672 80171 250728
rect 76780 250670 80171 250672
rect 129772 250728 131507 250730
rect 129772 250672 131446 250728
rect 131502 250672 131507 250728
rect 129772 250670 131507 250672
rect 170804 250728 173643 250730
rect 170804 250672 173582 250728
rect 173638 250672 173643 250728
rect 170804 250670 173643 250672
rect 223796 250728 226451 250730
rect 223796 250672 226390 250728
rect 226446 250672 226451 250728
rect 223796 250670 226451 250672
rect 80105 250667 80171 250670
rect 131441 250667 131507 250670
rect 173577 250667 173643 250670
rect 226385 250667 226451 250670
rect 140549 250458 140615 250461
rect 233469 250458 233535 250461
rect 140549 250456 143020 250458
rect 140549 250400 140554 250456
rect 140610 250400 143020 250456
rect 140549 250398 143020 250400
rect 233469 250456 237044 250458
rect 233469 250400 233474 250456
rect 233530 250400 237044 250456
rect 233469 250398 237044 250400
rect 140549 250395 140615 250398
rect 233469 250395 233535 250398
rect 87189 250322 87255 250325
rect 131349 250322 131415 250325
rect 87189 250320 90028 250322
rect 87189 250264 87194 250320
rect 87250 250264 90028 250320
rect 87189 250262 90028 250264
rect 129772 250320 131415 250322
rect 129772 250264 131354 250320
rect 131410 250264 131415 250320
rect 129772 250262 131415 250264
rect 87189 250259 87255 250262
rect 131349 250259 131415 250262
rect 182225 250322 182291 250325
rect 226293 250322 226359 250325
rect 182225 250320 184052 250322
rect 182225 250264 182230 250320
rect 182286 250264 184052 250320
rect 182225 250262 184052 250264
rect 223796 250320 226359 250322
rect 223796 250264 226298 250320
rect 226354 250264 226359 250320
rect 223796 250262 226359 250264
rect 182225 250259 182291 250262
rect 226293 250259 226359 250262
rect 80105 250186 80171 250189
rect 173669 250186 173735 250189
rect 76780 250184 80171 250186
rect 76780 250128 80110 250184
rect 80166 250128 80171 250184
rect 76780 250126 80171 250128
rect 170804 250184 173735 250186
rect 170804 250128 173674 250184
rect 173730 250128 173735 250184
rect 170804 250126 173735 250128
rect 80105 250123 80171 250126
rect 173669 250123 173735 250126
rect 87281 250050 87347 250053
rect 131349 250050 131415 250053
rect 87281 250048 90028 250050
rect 87281 249992 87286 250048
rect 87342 249992 90028 250048
rect 87281 249990 90028 249992
rect 129772 250048 131415 250050
rect 129772 249992 131354 250048
rect 131410 249992 131415 250048
rect 129772 249990 131415 249992
rect 87281 249987 87347 249990
rect 131349 249987 131415 249990
rect 182317 250050 182383 250053
rect 225925 250050 225991 250053
rect 182317 250048 184052 250050
rect 182317 249992 182322 250048
rect 182378 249992 184052 250048
rect 182317 249990 184052 249992
rect 223796 250048 225991 250050
rect 223796 249992 225930 250048
rect 225986 249992 225991 250048
rect 223796 249990 225991 249992
rect 182317 249987 182383 249990
rect 225925 249987 225991 249990
rect 47077 249914 47143 249917
rect 47077 249912 48996 249914
rect 47077 249856 47082 249912
rect 47138 249856 48996 249912
rect 47077 249854 48996 249856
rect 47077 249851 47143 249854
rect 139997 249778 140063 249781
rect 233469 249778 233535 249781
rect 139997 249776 143020 249778
rect 139997 249720 140002 249776
rect 140058 249720 143020 249776
rect 139997 249718 143020 249720
rect 233469 249776 237044 249778
rect 233469 249720 233474 249776
rect 233530 249720 237044 249776
rect 233469 249718 237044 249720
rect 139997 249715 140063 249718
rect 233469 249715 233535 249718
rect 87373 249642 87439 249645
rect 131809 249642 131875 249645
rect 87373 249640 90028 249642
rect 87373 249584 87378 249640
rect 87434 249584 90028 249640
rect 87373 249582 90028 249584
rect 129772 249640 131875 249642
rect 129772 249584 131814 249640
rect 131870 249584 131875 249640
rect 129772 249582 131875 249584
rect 87373 249579 87439 249582
rect 131809 249579 131875 249582
rect 140457 249642 140523 249645
rect 181581 249642 181647 249645
rect 226293 249642 226359 249645
rect 140457 249640 143050 249642
rect 140457 249584 140462 249640
rect 140518 249584 143050 249640
rect 140457 249582 143050 249584
rect 140457 249579 140523 249582
rect 80197 249506 80263 249509
rect 76780 249504 80263 249506
rect 76780 249448 80202 249504
rect 80258 249448 80263 249504
rect 76780 249446 80263 249448
rect 80197 249443 80263 249446
rect 87189 249234 87255 249237
rect 131349 249234 131415 249237
rect 87189 249232 90028 249234
rect 87189 249176 87194 249232
rect 87250 249176 90028 249232
rect 87189 249174 90028 249176
rect 129772 249232 131415 249234
rect 129772 249176 131354 249232
rect 131410 249176 131415 249232
rect 129772 249174 131415 249176
rect 87189 249171 87255 249174
rect 131349 249171 131415 249174
rect 142990 249136 143050 249582
rect 181581 249640 184052 249642
rect 181581 249584 181586 249640
rect 181642 249584 184052 249640
rect 181581 249582 184052 249584
rect 223796 249640 226359 249642
rect 223796 249584 226298 249640
rect 226354 249584 226359 249640
rect 223796 249582 226359 249584
rect 181581 249579 181647 249582
rect 226293 249579 226359 249582
rect 233561 249642 233627 249645
rect 233561 249640 237074 249642
rect 233561 249584 233566 249640
rect 233622 249584 237074 249640
rect 233561 249582 237074 249584
rect 233561 249579 233627 249582
rect 173577 249506 173643 249509
rect 170804 249504 173643 249506
rect 170804 249448 173582 249504
rect 173638 249448 173643 249504
rect 170804 249446 173643 249448
rect 173577 249443 173643 249446
rect 182317 249234 182383 249237
rect 225557 249234 225623 249237
rect 182317 249232 184052 249234
rect 182317 249176 182322 249232
rect 182378 249176 184052 249232
rect 182317 249174 184052 249176
rect 223796 249232 225623 249234
rect 223796 249176 225562 249232
rect 225618 249176 225623 249232
rect 223796 249174 225623 249176
rect 182317 249171 182383 249174
rect 225557 249171 225623 249174
rect 237014 249136 237074 249582
rect 80197 248826 80263 248829
rect 76780 248824 80263 248826
rect 76780 248768 80202 248824
rect 80258 248768 80263 248824
rect 76780 248766 80263 248768
rect 80197 248763 80263 248766
rect 88293 248826 88359 248829
rect 131349 248826 131415 248829
rect 88293 248824 90028 248826
rect 88293 248768 88298 248824
rect 88354 248768 90028 248824
rect 88293 248766 90028 248768
rect 129772 248824 131415 248826
rect 129772 248768 131354 248824
rect 131410 248768 131415 248824
rect 129772 248766 131415 248768
rect 88293 248763 88359 248766
rect 131349 248763 131415 248766
rect 140365 248826 140431 248829
rect 173209 248826 173275 248829
rect 140365 248824 143050 248826
rect 140365 248768 140370 248824
rect 140426 248768 143050 248824
rect 140365 248766 143050 248768
rect 170804 248824 173275 248826
rect 170804 248768 173214 248824
rect 173270 248768 173275 248824
rect 170804 248766 173275 248768
rect 140365 248763 140431 248766
rect 142990 248592 143050 248766
rect 173209 248763 173275 248766
rect 181121 248826 181187 248829
rect 226385 248826 226451 248829
rect 181121 248824 184052 248826
rect 181121 248768 181126 248824
rect 181182 248768 184052 248824
rect 181121 248766 184052 248768
rect 223796 248824 226451 248826
rect 223796 248768 226390 248824
rect 226446 248768 226451 248824
rect 223796 248766 226451 248768
rect 181121 248763 181187 248766
rect 226385 248763 226451 248766
rect 79277 248554 79343 248557
rect 76750 248552 79343 248554
rect 76750 248496 79282 248552
rect 79338 248496 79343 248552
rect 76750 248494 79343 248496
rect 76750 248184 76810 248494
rect 79277 248491 79343 248494
rect 88385 248418 88451 248421
rect 131441 248418 131507 248421
rect 88385 248416 90028 248418
rect 88385 248360 88390 248416
rect 88446 248360 90028 248416
rect 88385 248358 90028 248360
rect 129772 248416 131507 248418
rect 129772 248360 131446 248416
rect 131502 248360 131507 248416
rect 129772 248358 131507 248360
rect 88385 248355 88451 248358
rect 131441 248355 131507 248358
rect 181029 248418 181095 248421
rect 226293 248418 226359 248421
rect 181029 248416 184052 248418
rect 181029 248360 181034 248416
rect 181090 248360 184052 248416
rect 181029 248358 184052 248360
rect 223796 248416 226359 248418
rect 223796 248360 226298 248416
rect 226354 248360 226359 248416
rect 223796 248358 226359 248360
rect 181029 248355 181095 248358
rect 226293 248355 226359 248358
rect 233469 248418 233535 248421
rect 233469 248416 237044 248418
rect 233469 248360 233474 248416
rect 233530 248360 237044 248416
rect 233469 248358 237044 248360
rect 233469 248355 233535 248358
rect 233561 248282 233627 248285
rect 233561 248280 237074 248282
rect 233561 248224 233566 248280
rect 233622 248224 237074 248280
rect 233561 248222 237074 248224
rect 233561 248219 233627 248222
rect 140365 248146 140431 248149
rect 173577 248146 173643 248149
rect 140365 248144 143050 248146
rect 140365 248088 140370 248144
rect 140426 248088 143050 248144
rect 140365 248086 143050 248088
rect 170804 248144 173643 248146
rect 170804 248088 173582 248144
rect 173638 248088 173643 248144
rect 170804 248086 173643 248088
rect 140365 248083 140431 248086
rect 88017 248010 88083 248013
rect 132545 248010 132611 248013
rect 88017 248008 90028 248010
rect 88017 247952 88022 248008
rect 88078 247952 90028 248008
rect 88017 247950 90028 247952
rect 129772 248008 132611 248010
rect 129772 247952 132550 248008
rect 132606 247952 132611 248008
rect 129772 247950 132611 247952
rect 88017 247947 88083 247950
rect 132545 247947 132611 247950
rect 142990 247912 143050 248086
rect 173577 248083 173643 248086
rect 180845 248010 180911 248013
rect 226385 248010 226451 248013
rect 180845 248008 184052 248010
rect 180845 247952 180850 248008
rect 180906 247952 184052 248008
rect 180845 247950 184052 247952
rect 223796 248008 226451 248010
rect 223796 247952 226390 248008
rect 226446 247952 226451 248008
rect 223796 247950 226451 247952
rect 180845 247947 180911 247950
rect 226385 247947 226451 247950
rect 237014 247776 237074 248222
rect 131809 247738 131875 247741
rect 226293 247738 226359 247741
rect 129772 247736 131875 247738
rect 129772 247680 131814 247736
rect 131870 247680 131875 247736
rect 129772 247678 131875 247680
rect 223796 247736 226359 247738
rect 223796 247680 226298 247736
rect 226354 247680 226359 247736
rect 223796 247678 226359 247680
rect 131809 247675 131875 247678
rect 226293 247675 226359 247678
rect 87189 247602 87255 247605
rect 180937 247602 181003 247605
rect 87189 247600 90028 247602
rect 87189 247544 87194 247600
rect 87250 247544 90028 247600
rect 87189 247542 90028 247544
rect 180937 247600 184052 247602
rect 180937 247544 180942 247600
rect 180998 247544 184052 247600
rect 180937 247542 184052 247544
rect 87189 247539 87255 247542
rect 180937 247539 181003 247542
rect 80197 247466 80263 247469
rect 76780 247464 80263 247466
rect 76780 247408 80202 247464
rect 80258 247408 80263 247464
rect 76780 247406 80263 247408
rect 80197 247403 80263 247406
rect 140365 247466 140431 247469
rect 173209 247466 173275 247469
rect 140365 247464 143050 247466
rect 140365 247408 140370 247464
rect 140426 247408 143050 247464
rect 140365 247406 143050 247408
rect 170804 247464 173275 247466
rect 170804 247408 173214 247464
rect 173270 247408 173275 247464
rect 170804 247406 173275 247408
rect 140365 247403 140431 247406
rect 131441 247330 131507 247333
rect 129772 247328 131507 247330
rect 129772 247272 131446 247328
rect 131502 247272 131507 247328
rect 129772 247270 131507 247272
rect 131441 247267 131507 247270
rect 142990 247232 143050 247406
rect 173209 247403 173275 247406
rect 225649 247330 225715 247333
rect 223796 247328 225715 247330
rect 223796 247272 225654 247328
rect 225710 247272 225715 247328
rect 223796 247270 225715 247272
rect 225649 247267 225715 247270
rect 234481 247330 234547 247333
rect 234481 247328 237074 247330
rect 234481 247272 234486 247328
rect 234542 247272 237074 247328
rect 234481 247270 237074 247272
rect 234481 247267 234547 247270
rect 79277 247194 79343 247197
rect 76750 247192 79343 247194
rect 76750 247136 79282 247192
rect 79338 247136 79343 247192
rect 76750 247134 79343 247136
rect 76750 246824 76810 247134
rect 79277 247131 79343 247134
rect 87005 247194 87071 247197
rect 180753 247194 180819 247197
rect 87005 247192 90028 247194
rect 87005 247136 87010 247192
rect 87066 247136 90028 247192
rect 87005 247134 90028 247136
rect 180753 247192 184052 247194
rect 180753 247136 180758 247192
rect 180814 247136 184052 247192
rect 180753 247134 184052 247136
rect 87005 247131 87071 247134
rect 180753 247131 180819 247134
rect 237014 247096 237074 247270
rect 140641 247058 140707 247061
rect 140641 247056 143050 247058
rect 140641 247000 140646 247056
rect 140702 247000 143050 247056
rect 140641 246998 143050 247000
rect 140641 246995 140707 246998
rect 132177 246922 132243 246925
rect 129772 246920 132243 246922
rect 129772 246864 132182 246920
rect 132238 246864 132243 246920
rect 129772 246862 132243 246864
rect 132177 246859 132243 246862
rect 87097 246786 87163 246789
rect 87097 246784 90028 246786
rect 87097 246728 87102 246784
rect 87158 246728 90028 246784
rect 87097 246726 90028 246728
rect 87097 246723 87163 246726
rect 142990 246552 143050 246998
rect 226385 246922 226451 246925
rect 223796 246920 226451 246922
rect 223796 246864 226390 246920
rect 226446 246864 226451 246920
rect 223796 246862 226451 246864
rect 226385 246859 226451 246862
rect 234389 246922 234455 246925
rect 234389 246920 237074 246922
rect 234389 246864 234394 246920
rect 234450 246864 237074 246920
rect 234389 246862 237074 246864
rect 234389 246859 234455 246862
rect 173577 246786 173643 246789
rect 170804 246784 173643 246786
rect 170804 246728 173582 246784
rect 173638 246728 173643 246784
rect 170804 246726 173643 246728
rect 173577 246723 173643 246726
rect 180661 246786 180727 246789
rect 180661 246784 184052 246786
rect 180661 246728 180666 246784
rect 180722 246728 184052 246784
rect 180661 246726 184052 246728
rect 180661 246723 180727 246726
rect 131349 246514 131415 246517
rect 226293 246514 226359 246517
rect 129772 246512 131415 246514
rect 129772 246456 131354 246512
rect 131410 246456 131415 246512
rect 129772 246454 131415 246456
rect 223796 246512 226359 246514
rect 223796 246456 226298 246512
rect 226354 246456 226359 246512
rect 223796 246454 226359 246456
rect 131349 246451 131415 246454
rect 226293 246451 226359 246454
rect 237014 246416 237074 246862
rect 87189 246378 87255 246381
rect 182317 246378 182383 246381
rect 87189 246376 90028 246378
rect 87189 246320 87194 246376
rect 87250 246320 90028 246376
rect 87189 246318 90028 246320
rect 182317 246376 184052 246378
rect 182317 246320 182322 246376
rect 182378 246320 184052 246376
rect 182317 246318 184052 246320
rect 87189 246315 87255 246318
rect 182317 246315 182383 246318
rect 80197 246106 80263 246109
rect 131993 246106 132059 246109
rect 76780 246104 80263 246106
rect 76780 246048 80202 246104
rect 80258 246048 80263 246104
rect 76780 246046 80263 246048
rect 129772 246104 132059 246106
rect 129772 246048 131998 246104
rect 132054 246048 132059 246104
rect 129772 246046 132059 246048
rect 80197 246043 80263 246046
rect 131993 246043 132059 246046
rect 140549 246106 140615 246109
rect 173577 246106 173643 246109
rect 226293 246106 226359 246109
rect 140549 246104 143050 246106
rect 140549 246048 140554 246104
rect 140610 246048 143050 246104
rect 140549 246046 143050 246048
rect 170804 246104 173643 246106
rect 170804 246048 173582 246104
rect 173638 246048 173643 246104
rect 170804 246046 173643 246048
rect 223796 246104 226359 246106
rect 223796 246048 226298 246104
rect 226354 246048 226359 246104
rect 223796 246046 226359 246048
rect 140549 246043 140615 246046
rect 86913 245970 86979 245973
rect 86913 245968 90028 245970
rect 86913 245912 86918 245968
rect 86974 245912 90028 245968
rect 86913 245910 90028 245912
rect 86913 245907 86979 245910
rect 142990 245872 143050 246046
rect 173577 246043 173643 246046
rect 226293 246043 226359 246046
rect 180845 245970 180911 245973
rect 233469 245970 233535 245973
rect 180845 245968 184052 245970
rect 180845 245912 180850 245968
rect 180906 245912 184052 245968
rect 180845 245910 184052 245912
rect 233469 245968 237074 245970
rect 233469 245912 233474 245968
rect 233530 245912 237074 245968
rect 233469 245910 237074 245912
rect 180845 245907 180911 245910
rect 233469 245907 233535 245910
rect 79277 245834 79343 245837
rect 131441 245834 131507 245837
rect 226201 245834 226267 245837
rect 76750 245832 79343 245834
rect 76750 245776 79282 245832
rect 79338 245776 79343 245832
rect 76750 245774 79343 245776
rect 129772 245832 131507 245834
rect 129772 245776 131446 245832
rect 131502 245776 131507 245832
rect 129772 245774 131507 245776
rect 223796 245832 226267 245834
rect 223796 245776 226206 245832
rect 226262 245776 226267 245832
rect 223796 245774 226267 245776
rect 76750 245464 76810 245774
rect 79277 245771 79343 245774
rect 131441 245771 131507 245774
rect 226201 245771 226267 245774
rect 237014 245736 237074 245910
rect 86821 245562 86887 245565
rect 140365 245562 140431 245565
rect 180937 245562 181003 245565
rect 233561 245562 233627 245565
rect 86821 245560 90028 245562
rect 86821 245504 86826 245560
rect 86882 245504 90028 245560
rect 86821 245502 90028 245504
rect 140365 245560 143050 245562
rect 140365 245504 140370 245560
rect 140426 245504 143050 245560
rect 140365 245502 143050 245504
rect 86821 245499 86887 245502
rect 140365 245499 140431 245502
rect 131349 245426 131415 245429
rect 129772 245424 131415 245426
rect 129772 245368 131354 245424
rect 131410 245368 131415 245424
rect 129772 245366 131415 245368
rect 131349 245363 131415 245366
rect 142990 245328 143050 245502
rect 180937 245560 184052 245562
rect 180937 245504 180942 245560
rect 180998 245504 184052 245560
rect 180937 245502 184052 245504
rect 233561 245560 237074 245562
rect 233561 245504 233566 245560
rect 233622 245504 237074 245560
rect 233561 245502 237074 245504
rect 180937 245499 181003 245502
rect 233561 245499 233627 245502
rect 173485 245426 173551 245429
rect 225557 245426 225623 245429
rect 170804 245424 173551 245426
rect 170804 245368 173490 245424
rect 173546 245368 173551 245424
rect 170804 245366 173551 245368
rect 223796 245424 225623 245426
rect 223796 245368 225562 245424
rect 225618 245368 225623 245424
rect 223796 245366 225623 245368
rect 173485 245363 173551 245366
rect 225557 245363 225623 245366
rect 87649 245154 87715 245157
rect 182225 245154 182291 245157
rect 87649 245152 90028 245154
rect 87649 245096 87654 245152
rect 87710 245096 90028 245152
rect 87649 245094 90028 245096
rect 182225 245152 184052 245154
rect 182225 245096 182230 245152
rect 182286 245096 184052 245152
rect 182225 245094 184052 245096
rect 87649 245091 87715 245094
rect 182225 245091 182291 245094
rect 237014 245056 237074 245502
rect 131809 245018 131875 245021
rect 226385 245018 226451 245021
rect 129772 245016 131875 245018
rect 129772 244960 131814 245016
rect 131870 244960 131875 245016
rect 129772 244958 131875 244960
rect 223796 245016 226451 245018
rect 223796 244960 226390 245016
rect 226446 244960 226451 245016
rect 223796 244958 226451 244960
rect 131809 244955 131875 244958
rect 226385 244955 226451 244958
rect 80197 244746 80263 244749
rect 76780 244744 80263 244746
rect 76780 244688 80202 244744
rect 80258 244688 80263 244744
rect 76780 244686 80263 244688
rect 80197 244683 80263 244686
rect 87557 244746 87623 244749
rect 173577 244746 173643 244749
rect 87557 244744 90028 244746
rect 87557 244688 87562 244744
rect 87618 244688 90028 244744
rect 87557 244686 90028 244688
rect 170804 244744 173643 244746
rect 170804 244688 173582 244744
rect 173638 244688 173643 244744
rect 170804 244686 173643 244688
rect 87557 244683 87623 244686
rect 173577 244683 173643 244686
rect 182041 244746 182107 244749
rect 233653 244746 233719 244749
rect 182041 244744 184052 244746
rect 182041 244688 182046 244744
rect 182102 244688 184052 244744
rect 182041 244686 184052 244688
rect 233653 244744 237074 244746
rect 233653 244688 233658 244744
rect 233714 244688 237074 244744
rect 233653 244686 237074 244688
rect 182041 244683 182107 244686
rect 233653 244683 233719 244686
rect 131625 244610 131691 244613
rect 129772 244608 131691 244610
rect 129772 244552 131630 244608
rect 131686 244552 131691 244608
rect 129772 244550 131691 244552
rect 131625 244547 131691 244550
rect 140641 244610 140707 244613
rect 225741 244610 225807 244613
rect 140641 244608 143020 244610
rect 140641 244552 140646 244608
rect 140702 244552 143020 244608
rect 140641 244550 143020 244552
rect 223796 244608 225807 244610
rect 223796 244552 225746 244608
rect 225802 244552 225807 244608
rect 223796 244550 225807 244552
rect 140641 244547 140707 244550
rect 225741 244547 225807 244550
rect 80105 244474 80171 244477
rect 76750 244472 80171 244474
rect 76750 244416 80110 244472
rect 80166 244416 80171 244472
rect 76750 244414 80171 244416
rect 76750 244104 76810 244414
rect 80105 244411 80171 244414
rect 140181 244474 140247 244477
rect 140181 244472 143050 244474
rect 140181 244416 140186 244472
rect 140242 244416 143050 244472
rect 140181 244414 143050 244416
rect 140181 244411 140247 244414
rect 87281 244338 87347 244341
rect 87281 244336 90028 244338
rect 87281 244280 87286 244336
rect 87342 244280 90028 244336
rect 87281 244278 90028 244280
rect 87281 244275 87347 244278
rect 131533 244202 131599 244205
rect 129772 244200 131599 244202
rect 129772 244144 131538 244200
rect 131594 244144 131599 244200
rect 129772 244142 131599 244144
rect 131533 244139 131599 244142
rect 142990 243968 143050 244414
rect 237014 244376 237074 244686
rect 182317 244338 182383 244341
rect 182317 244336 184052 244338
rect 182317 244280 182322 244336
rect 182378 244280 184052 244336
rect 182317 244278 184052 244280
rect 182317 244275 182383 244278
rect 226293 244202 226359 244205
rect 223796 244200 226359 244202
rect 223796 244144 226298 244200
rect 226354 244144 226359 244200
rect 223796 244142 226359 244144
rect 226293 244139 226359 244142
rect 233469 244202 233535 244205
rect 233469 244200 237074 244202
rect 233469 244144 233474 244200
rect 233530 244144 237074 244200
rect 233469 244142 237074 244144
rect 233469 244139 233535 244142
rect 172841 244066 172907 244069
rect 170804 244064 172907 244066
rect 170804 244008 172846 244064
rect 172902 244008 172907 244064
rect 170804 244006 172907 244008
rect 172841 244003 172907 244006
rect 87189 243930 87255 243933
rect 131349 243930 131415 243933
rect 87189 243928 90028 243930
rect 87189 243872 87194 243928
rect 87250 243872 90028 243928
rect 87189 243870 90028 243872
rect 129772 243928 131415 243930
rect 129772 243872 131354 243928
rect 131410 243872 131415 243928
rect 129772 243870 131415 243872
rect 87189 243867 87255 243870
rect 131349 243867 131415 243870
rect 181213 243930 181279 243933
rect 226201 243930 226267 243933
rect 181213 243928 184052 243930
rect 181213 243872 181218 243928
rect 181274 243872 184052 243928
rect 181213 243870 184052 243872
rect 223796 243928 226267 243930
rect 223796 243872 226206 243928
rect 226262 243872 226267 243928
rect 223796 243870 226267 243872
rect 181213 243867 181279 243870
rect 226201 243867 226267 243870
rect 237014 243696 237074 244142
rect 87465 243522 87531 243525
rect 131441 243522 131507 243525
rect 87465 243520 90028 243522
rect 87465 243464 87470 243520
rect 87526 243464 90028 243520
rect 87465 243462 90028 243464
rect 129772 243520 131507 243522
rect 129772 243464 131446 243520
rect 131502 243464 131507 243520
rect 129772 243462 131507 243464
rect 87465 243459 87531 243462
rect 131441 243459 131507 243462
rect 182133 243522 182199 243525
rect 226477 243522 226543 243525
rect 182133 243520 184052 243522
rect 182133 243464 182138 243520
rect 182194 243464 184052 243520
rect 182133 243462 184052 243464
rect 223796 243520 226543 243522
rect 223796 243464 226482 243520
rect 226538 243464 226543 243520
rect 223796 243462 226543 243464
rect 182133 243459 182199 243462
rect 226477 243459 226543 243462
rect 80013 243386 80079 243389
rect 173945 243386 174011 243389
rect 76780 243384 80079 243386
rect 76780 243328 80018 243384
rect 80074 243328 80079 243384
rect 76780 243326 80079 243328
rect 170804 243384 174011 243386
rect 170804 243328 173950 243384
rect 174006 243328 174011 243384
rect 170804 243326 174011 243328
rect 80013 243323 80079 243326
rect 173945 243323 174011 243326
rect 233469 243386 233535 243389
rect 233469 243384 237074 243386
rect 233469 243328 233474 243384
rect 233530 243328 237074 243384
rect 233469 243326 237074 243328
rect 233469 243323 233535 243326
rect 139629 243250 139695 243253
rect 139629 243248 143020 243250
rect 139629 243192 139634 243248
rect 139690 243192 143020 243248
rect 139629 243190 143020 243192
rect 139629 243187 139695 243190
rect 80197 243114 80263 243117
rect 76750 243112 80263 243114
rect 76750 243056 80202 243112
rect 80258 243056 80263 243112
rect 76750 243054 80263 243056
rect 76750 242880 76810 243054
rect 80197 243051 80263 243054
rect 87189 243114 87255 243117
rect 131533 243114 131599 243117
rect 87189 243112 90028 243114
rect 87189 243056 87194 243112
rect 87250 243056 90028 243112
rect 87189 243054 90028 243056
rect 129772 243112 131599 243114
rect 129772 243056 131538 243112
rect 131594 243056 131599 243112
rect 129772 243054 131599 243056
rect 87189 243051 87255 243054
rect 131533 243051 131599 243054
rect 139721 243114 139787 243117
rect 182317 243114 182383 243117
rect 226293 243114 226359 243117
rect 139721 243112 143050 243114
rect 139721 243056 139726 243112
rect 139782 243056 143050 243112
rect 139721 243054 143050 243056
rect 139721 243051 139787 243054
rect 86545 242706 86611 242709
rect 131441 242706 131507 242709
rect 86545 242704 90028 242706
rect 86545 242648 86550 242704
rect 86606 242648 90028 242704
rect 86545 242646 90028 242648
rect 129772 242704 131507 242706
rect 129772 242648 131446 242704
rect 131502 242648 131507 242704
rect 129772 242646 131507 242648
rect 86545 242643 86611 242646
rect 131441 242643 131507 242646
rect 142990 242608 143050 243054
rect 182317 243112 184052 243114
rect 182317 243056 182322 243112
rect 182378 243056 184052 243112
rect 182317 243054 184052 243056
rect 223796 243112 226359 243114
rect 223796 243056 226298 243112
rect 226354 243056 226359 243112
rect 223796 243054 226359 243056
rect 182317 243051 182383 243054
rect 226293 243051 226359 243054
rect 237014 243016 237074 243326
rect 173577 242842 173643 242845
rect 170804 242840 173643 242842
rect 170804 242784 173582 242840
rect 173638 242784 173643 242840
rect 170804 242782 173643 242784
rect 173577 242779 173643 242782
rect 233561 242842 233627 242845
rect 233561 242840 237074 242842
rect 233561 242784 233566 242840
rect 233622 242784 237074 242840
rect 233561 242782 237074 242784
rect 233561 242779 233627 242782
rect 180385 242706 180451 242709
rect 226017 242706 226083 242709
rect 180385 242704 184052 242706
rect 180385 242648 180390 242704
rect 180446 242648 184052 242704
rect 180385 242646 184052 242648
rect 223796 242704 226083 242706
rect 223796 242648 226022 242704
rect 226078 242648 226083 242704
rect 223796 242646 226083 242648
rect 180385 242643 180451 242646
rect 226017 242643 226083 242646
rect 80197 242434 80263 242437
rect 76750 242432 80263 242434
rect 76750 242376 80202 242432
rect 80258 242376 80263 242432
rect 76750 242374 80263 242376
rect 76750 242200 76810 242374
rect 80197 242371 80263 242374
rect 237014 242336 237074 242782
rect 86453 242298 86519 242301
rect 131349 242298 131415 242301
rect 86453 242296 90028 242298
rect 86453 242240 86458 242296
rect 86514 242240 90028 242296
rect 86453 242238 90028 242240
rect 129772 242296 131415 242298
rect 129772 242240 131354 242296
rect 131410 242240 131415 242296
rect 129772 242238 131415 242240
rect 86453 242235 86519 242238
rect 131349 242235 131415 242238
rect 180293 242298 180359 242301
rect 226385 242298 226451 242301
rect 180293 242296 184052 242298
rect 180293 242240 180298 242296
rect 180354 242240 184052 242296
rect 180293 242238 184052 242240
rect 223796 242296 226451 242298
rect 223796 242240 226390 242296
rect 226446 242240 226451 242296
rect 223796 242238 226451 242240
rect 180293 242235 180359 242238
rect 226385 242235 226451 242238
rect 264657 242298 264723 242301
rect 264798 242298 264858 242812
rect 264657 242296 264858 242298
rect 264657 242240 264662 242296
rect 264718 242240 264858 242296
rect 264657 242238 264858 242240
rect 264657 242235 264723 242238
rect 172841 242162 172907 242165
rect 170804 242160 172907 242162
rect 170804 242104 172846 242160
rect 172902 242104 172907 242160
rect 170804 242102 172907 242104
rect 172841 242099 172907 242102
rect 87373 242026 87439 242029
rect 131349 242026 131415 242029
rect 87373 242024 90028 242026
rect 87373 241968 87378 242024
rect 87434 241968 90028 242024
rect 87373 241966 90028 241968
rect 129772 242024 131415 242026
rect 129772 241968 131354 242024
rect 131410 241968 131415 242024
rect 129772 241966 131415 241968
rect 87373 241963 87439 241966
rect 131349 241963 131415 241966
rect 140549 242026 140615 242029
rect 181581 242026 181647 242029
rect 226017 242026 226083 242029
rect 140549 242024 143020 242026
rect 140549 241968 140554 242024
rect 140610 241968 143020 242024
rect 140549 241966 143020 241968
rect 181581 242024 184052 242026
rect 181581 241968 181586 242024
rect 181642 241968 184052 242024
rect 181581 241966 184052 241968
rect 223796 242024 226083 242026
rect 223796 241968 226022 242024
rect 226078 241968 226083 242024
rect 223796 241966 226083 241968
rect 140549 241963 140615 241966
rect 181581 241963 181647 241966
rect 226017 241963 226083 241966
rect 233469 242026 233535 242029
rect 233469 242024 237074 242026
rect 233469 241968 233474 242024
rect 233530 241968 237074 242024
rect 233469 241966 237074 241968
rect 233469 241963 233535 241966
rect 140181 241890 140247 241893
rect 140181 241888 143050 241890
rect 140181 241832 140186 241888
rect 140242 241832 143050 241888
rect 140181 241830 143050 241832
rect 140181 241827 140247 241830
rect 80197 241754 80263 241757
rect 76750 241752 80263 241754
rect 76750 241696 80202 241752
rect 80258 241696 80263 241752
rect 76750 241694 80263 241696
rect 76750 241520 76810 241694
rect 80197 241691 80263 241694
rect 142990 241384 143050 241830
rect 237014 241656 237074 241966
rect 300169 241618 300235 241621
rect 303416 241618 303896 241648
rect 300169 241616 303896 241618
rect 300169 241560 300174 241616
rect 300230 241560 303896 241616
rect 300169 241558 303896 241560
rect 300169 241555 300235 241558
rect 303416 241528 303896 241558
rect 173577 241482 173643 241485
rect 170804 241480 173643 241482
rect 170804 241424 173582 241480
rect 173638 241424 173643 241480
rect 170804 241422 173643 241424
rect 173577 241419 173643 241422
rect 233653 241482 233719 241485
rect 233653 241480 237074 241482
rect 233653 241424 233658 241480
rect 233714 241424 237074 241480
rect 233653 241422 237074 241424
rect 233653 241419 233719 241422
rect 79093 241346 79159 241349
rect 76750 241344 79159 241346
rect 76750 241288 79098 241344
rect 79154 241288 79159 241344
rect 76750 241286 79159 241288
rect 76750 240840 76810 241286
rect 79093 241283 79159 241286
rect 237014 240976 237074 241422
rect 173669 240802 173735 240805
rect 170804 240800 173735 240802
rect 170804 240744 173674 240800
rect 173730 240744 173735 240800
rect 170804 240742 173735 240744
rect 173669 240739 173735 240742
rect 80105 240666 80171 240669
rect 76750 240664 80171 240666
rect 76750 240608 80110 240664
rect 80166 240608 80171 240664
rect 76750 240606 80171 240608
rect 76750 240160 76810 240606
rect 80105 240603 80171 240606
rect 139537 240666 139603 240669
rect 233745 240666 233811 240669
rect 139537 240664 143020 240666
rect 139537 240608 139542 240664
rect 139598 240608 143020 240664
rect 139537 240606 143020 240608
rect 233745 240664 237074 240666
rect 233745 240608 233750 240664
rect 233806 240608 237074 240664
rect 233745 240606 237074 240608
rect 139537 240603 139603 240606
rect 233745 240603 233811 240606
rect 141009 240530 141075 240533
rect 142246 240530 142252 240532
rect 141009 240528 142252 240530
rect 141009 240472 141014 240528
rect 141070 240472 142252 240528
rect 141009 240470 142252 240472
rect 141009 240467 141075 240470
rect 142246 240468 142252 240470
rect 142316 240468 142322 240532
rect 139353 240394 139419 240397
rect 139353 240392 143050 240394
rect 139353 240336 139358 240392
rect 139414 240336 143050 240392
rect 139353 240334 143050 240336
rect 139353 240331 139419 240334
rect 142990 240024 143050 240334
rect 237014 240296 237074 240606
rect 173485 240122 173551 240125
rect 170804 240120 173551 240122
rect 170804 240064 173490 240120
rect 173546 240064 173551 240120
rect 170804 240062 173551 240064
rect 173485 240059 173551 240062
rect 233837 240122 233903 240125
rect 233837 240120 237074 240122
rect 233837 240064 233842 240120
rect 233898 240064 237074 240120
rect 233837 240062 237074 240064
rect 233837 240059 233903 240062
rect 79921 239986 79987 239989
rect 76750 239984 79987 239986
rect 76750 239928 79926 239984
rect 79982 239928 79987 239984
rect 76750 239926 79987 239928
rect 76750 239480 76810 239926
rect 79921 239923 79987 239926
rect 237014 239616 237074 240062
rect 173853 239442 173919 239445
rect 170804 239440 173919 239442
rect 170804 239384 173858 239440
rect 173914 239384 173919 239440
rect 170804 239382 173919 239384
rect 173853 239379 173919 239382
rect 140549 239306 140615 239309
rect 140549 239304 143020 239306
rect 140549 239248 140554 239304
rect 140610 239248 143020 239304
rect 140549 239246 143020 239248
rect 140549 239243 140615 239246
rect 140641 239170 140707 239173
rect 233469 239170 233535 239173
rect 140641 239168 143050 239170
rect 140641 239112 140646 239168
rect 140702 239112 143050 239168
rect 140641 239110 143050 239112
rect 140641 239107 140707 239110
rect 80197 239034 80263 239037
rect 76750 239032 80263 239034
rect 76750 238976 80202 239032
rect 80258 238976 80263 239032
rect 76750 238974 80263 238976
rect 76750 238800 76810 238974
rect 80197 238971 80263 238974
rect 142990 238800 143050 239110
rect 233469 239168 237074 239170
rect 233469 239112 233474 239168
rect 233530 239112 237074 239168
rect 233469 239110 237074 239112
rect 233469 239107 233535 239110
rect 237014 238936 237074 239110
rect 173669 238762 173735 238765
rect 170804 238760 173735 238762
rect 170804 238704 173674 238760
rect 173730 238704 173735 238760
rect 170804 238702 173735 238704
rect 173669 238699 173735 238702
rect 233561 238762 233627 238765
rect 233561 238760 237074 238762
rect 233561 238704 233566 238760
rect 233622 238704 237074 238760
rect 233561 238702 237074 238704
rect 233561 238699 233627 238702
rect 79277 238626 79343 238629
rect 76750 238624 79343 238626
rect 76750 238568 79282 238624
rect 79338 238568 79343 238624
rect 76750 238566 79343 238568
rect 76750 238120 76810 238566
rect 79277 238563 79343 238566
rect 139445 238626 139511 238629
rect 139445 238624 143050 238626
rect 139445 238568 139450 238624
rect 139506 238568 143050 238624
rect 139445 238566 143050 238568
rect 139445 238563 139511 238566
rect 142990 238120 143050 238566
rect 237014 238256 237074 238702
rect 173761 238082 173827 238085
rect 170804 238080 173827 238082
rect 170804 238024 173766 238080
rect 173822 238024 173827 238080
rect 170804 238022 173827 238024
rect 173761 238019 173827 238022
rect 233469 237810 233535 237813
rect 233469 237808 237074 237810
rect 233469 237752 233474 237808
rect 233530 237752 237074 237808
rect 233469 237750 237074 237752
rect 233469 237747 233535 237750
rect 80197 237674 80263 237677
rect 76750 237672 80263 237674
rect 76750 237616 80202 237672
rect 80258 237616 80263 237672
rect 76750 237614 80263 237616
rect 76750 237440 76810 237614
rect 80197 237611 80263 237614
rect 237014 237576 237074 237750
rect 140549 237402 140615 237405
rect 173577 237402 173643 237405
rect 140549 237400 143020 237402
rect 140549 237344 140554 237400
rect 140610 237344 143020 237400
rect 140549 237342 143020 237344
rect 170804 237400 173643 237402
rect 170804 237344 173582 237400
rect 173638 237344 173643 237400
rect 170804 237342 173643 237344
rect 140549 237339 140615 237342
rect 173577 237339 173643 237342
rect 233561 237402 233627 237405
rect 233561 237400 237074 237402
rect 233561 237344 233566 237400
rect 233622 237344 237074 237400
rect 233561 237342 237074 237344
rect 233561 237339 233627 237342
rect 140273 237266 140339 237269
rect 140273 237264 143050 237266
rect 140273 237208 140278 237264
rect 140334 237208 143050 237264
rect 140273 237206 143050 237208
rect 140273 237203 140339 237206
rect 80197 236994 80263 236997
rect 76750 236992 80263 236994
rect 76750 236936 80202 236992
rect 80258 236936 80263 236992
rect 76750 236934 80263 236936
rect 76750 236760 76810 236934
rect 80197 236931 80263 236934
rect 142990 236760 143050 237206
rect 237014 236896 237074 237342
rect 173393 236722 173459 236725
rect 170804 236720 173459 236722
rect 170804 236664 173398 236720
rect 173454 236664 173459 236720
rect 170804 236662 173459 236664
rect 173393 236659 173459 236662
rect 139261 236450 139327 236453
rect 234113 236450 234179 236453
rect 139261 236448 143050 236450
rect 139261 236392 139266 236448
rect 139322 236392 143050 236448
rect 139261 236390 143050 236392
rect 139261 236387 139327 236390
rect 142990 236216 143050 236390
rect 234113 236448 237074 236450
rect 234113 236392 234118 236448
rect 234174 236392 237074 236448
rect 234113 236390 237074 236392
rect 234113 236387 234179 236390
rect 237014 236216 237074 236390
rect 80197 236178 80263 236181
rect 173577 236178 173643 236181
rect 76780 236176 80263 236178
rect 76780 236120 80202 236176
rect 80258 236120 80263 236176
rect 76780 236118 80263 236120
rect 170804 236176 173643 236178
rect 170804 236120 173582 236176
rect 173638 236120 173643 236176
rect 170804 236118 173643 236120
rect 80197 236115 80263 236118
rect 173577 236115 173643 236118
rect 203109 233730 203175 233733
rect 264197 233730 264263 233733
rect 203109 233728 264263 233730
rect 203109 233672 203114 233728
rect 203170 233672 264202 233728
rect 264258 233672 264263 233728
rect 203109 233670 264263 233672
rect 203109 233667 203175 233670
rect 264197 233667 264263 233670
rect 60693 233050 60759 233053
rect 73665 233050 73731 233053
rect 60693 233048 73731 233050
rect 60693 232992 60698 233048
rect 60754 232992 73670 233048
rect 73726 232992 73731 233048
rect 60693 232990 73731 232992
rect 60693 232987 60759 232990
rect 73665 232987 73731 232990
rect 156005 233050 156071 233053
rect 169989 233050 170055 233053
rect 156005 233048 170055 233050
rect 156005 232992 156010 233048
rect 156066 232992 169994 233048
rect 170050 232992 170055 233048
rect 156005 232990 170055 232992
rect 156005 232987 156071 232990
rect 169989 232987 170055 232990
rect 152969 231010 153035 231013
rect 153153 231010 153219 231013
rect 152969 231008 153219 231010
rect 152969 230952 152974 231008
rect 153030 230952 153158 231008
rect 153214 230952 153219 231008
rect 152969 230950 153219 230952
rect 152969 230947 153035 230950
rect 153153 230947 153219 230950
rect 137697 227066 137763 227069
rect 231997 227066 232063 227069
rect 134740 227064 137763 227066
rect 134740 227008 137702 227064
rect 137758 227008 137763 227064
rect 134740 227006 137763 227008
rect 228764 227064 232063 227066
rect 228764 227008 232002 227064
rect 232058 227008 232063 227064
rect 228764 227006 232063 227008
rect 137697 227003 137763 227006
rect 231997 227003 232063 227006
rect 137513 225570 137579 225573
rect 231905 225570 231971 225573
rect 134740 225568 137579 225570
rect 134740 225512 137518 225568
rect 137574 225512 137579 225568
rect 134740 225510 137579 225512
rect 228764 225568 231971 225570
rect 228764 225512 231910 225568
rect 231966 225512 231971 225568
rect 228764 225510 231971 225512
rect 137513 225507 137579 225510
rect 231905 225507 231971 225510
rect 61153 224346 61219 224349
rect 62901 224346 62967 224349
rect 61153 224344 62967 224346
rect 61153 224288 61158 224344
rect 61214 224288 62906 224344
rect 62962 224288 62967 224344
rect 61153 224286 62967 224288
rect 61153 224283 61219 224286
rect 62901 224283 62967 224286
rect 24169 224210 24235 224213
rect 69750 224210 69756 224212
rect 24169 224208 69756 224210
rect 24169 224152 24174 224208
rect 24230 224152 69756 224208
rect 24169 224150 69756 224152
rect 24169 224147 24235 224150
rect 69750 224148 69756 224150
rect 69820 224148 69826 224212
rect 137697 223938 137763 223941
rect 231997 223938 232063 223941
rect 134740 223936 137763 223938
rect 134740 223880 137702 223936
rect 137758 223880 137763 223936
rect 134740 223878 137763 223880
rect 228764 223936 232063 223938
rect 228764 223880 232002 223936
rect 232058 223880 232063 223936
rect 228764 223878 232063 223880
rect 137697 223875 137763 223878
rect 231997 223875 232063 223878
rect 134710 221762 134770 222344
rect 228734 221898 228794 222344
rect 231077 221898 231143 221901
rect 228734 221896 231143 221898
rect 228734 221840 231082 221896
rect 231138 221840 231143 221896
rect 228734 221838 231143 221840
rect 231077 221835 231143 221838
rect 137697 221762 137763 221765
rect 134710 221760 137763 221762
rect 134710 221704 137702 221760
rect 137758 221704 137763 221760
rect 134710 221702 137763 221704
rect 137697 221699 137763 221702
rect 148737 221626 148803 221629
rect 148737 221624 148938 221626
rect 148737 221568 148742 221624
rect 148798 221568 148938 221624
rect 148737 221566 148938 221568
rect 148737 221563 148803 221566
rect 148878 221460 148938 221566
rect 241606 221564 241612 221628
rect 241676 221626 241682 221628
rect 241676 221566 242962 221626
rect 241676 221564 241682 221566
rect 242902 221460 242962 221566
rect 9896 221218 10376 221248
rect 12945 221218 13011 221221
rect 9896 221216 13011 221218
rect 9896 221160 12950 221216
rect 13006 221160 13011 221216
rect 9896 221158 13011 221160
rect 9896 221128 10376 221158
rect 12945 221155 13011 221158
rect 137605 220810 137671 220813
rect 231721 220810 231787 220813
rect 134740 220808 137671 220810
rect 134740 220752 137610 220808
rect 137666 220752 137671 220808
rect 134740 220750 137671 220752
rect 228764 220808 231787 220810
rect 228764 220752 231726 220808
rect 231782 220752 231787 220808
rect 228764 220750 231787 220752
rect 137605 220747 137671 220750
rect 231721 220747 231787 220750
rect 145609 219314 145675 219317
rect 145609 219312 148938 219314
rect 145609 219256 145614 219312
rect 145670 219256 148938 219312
rect 145609 219254 148938 219256
rect 145609 219251 145675 219254
rect 148878 219216 148938 219254
rect 134710 218906 134770 219216
rect 228734 219042 228794 219216
rect 230985 219042 231051 219045
rect 228734 219040 231051 219042
rect 228734 218984 230990 219040
rect 231046 218984 231051 219040
rect 228734 218982 231051 218984
rect 230985 218979 231051 218982
rect 137605 218906 137671 218909
rect 134710 218904 137671 218906
rect 134710 218848 137610 218904
rect 137666 218848 137671 218904
rect 134710 218846 137671 218848
rect 137605 218843 137671 218846
rect 38102 218770 38108 218772
rect 35748 218710 38108 218770
rect 38102 218708 38108 218710
rect 38172 218708 38178 218772
rect 240921 218770 240987 218773
rect 242902 218770 242962 219148
rect 240921 218768 242962 218770
rect 240921 218712 240926 218768
rect 240982 218712 242962 218768
rect 240921 218710 242962 218712
rect 240921 218707 240987 218710
rect 137789 217682 137855 217685
rect 231813 217682 231879 217685
rect 134740 217680 137855 217682
rect 134740 217624 137794 217680
rect 137850 217624 137855 217680
rect 134740 217622 137855 217624
rect 228764 217680 231879 217682
rect 228764 217624 231818 217680
rect 231874 217624 231879 217680
rect 228764 217622 231879 217624
rect 137789 217619 137855 217622
rect 231813 217619 231879 217622
rect 276157 217682 276223 217685
rect 276157 217680 278076 217682
rect 276157 217624 276162 217680
rect 276218 217624 278076 217680
rect 276157 217622 278076 217624
rect 276157 217619 276223 217622
rect 300169 217138 300235 217141
rect 303416 217138 303896 217168
rect 300169 217136 303896 217138
rect 300169 217080 300174 217136
rect 300230 217080 303896 217136
rect 300169 217078 303896 217080
rect 300169 217075 300235 217078
rect 303416 217048 303896 217078
rect 145609 217002 145675 217005
rect 145609 217000 148938 217002
rect 145609 216944 145614 217000
rect 145670 216944 148938 217000
rect 145609 216942 148938 216944
rect 145609 216939 145675 216942
rect 148878 216904 148938 216942
rect 240461 216322 240527 216325
rect 242902 216322 242962 216836
rect 265209 216596 265275 216597
rect 265158 216532 265164 216596
rect 265228 216594 265275 216596
rect 265228 216592 265320 216594
rect 265270 216536 265320 216592
rect 265228 216534 265320 216536
rect 265228 216532 265275 216534
rect 293678 216532 293684 216596
rect 293748 216532 293754 216596
rect 265209 216531 265275 216532
rect 240461 216320 242962 216322
rect 240461 216264 240466 216320
rect 240522 216264 242962 216320
rect 240461 216262 242962 216264
rect 240461 216259 240527 216262
rect 51953 216186 52019 216189
rect 52270 216186 52276 216188
rect 51953 216184 52276 216186
rect 51953 216128 51958 216184
rect 52014 216128 52276 216184
rect 51953 216126 52276 216128
rect 51953 216123 52019 216126
rect 52270 216124 52276 216126
rect 52340 216186 52346 216188
rect 54486 216186 55068 216242
rect 293686 216224 293746 216532
rect 52340 216182 55068 216186
rect 52340 216126 54546 216182
rect 52340 216124 52346 216126
rect 134710 215914 134770 216088
rect 228734 216050 228794 216088
rect 231997 216050 232063 216053
rect 228734 216048 232063 216050
rect 228734 215992 232002 216048
rect 232058 215992 232063 216048
rect 228734 215990 232063 215992
rect 231997 215987 232063 215990
rect 137789 215914 137855 215917
rect 134710 215912 137855 215914
rect 134710 215856 137794 215912
rect 137850 215856 137855 215912
rect 134710 215854 137855 215856
rect 137789 215851 137855 215854
rect 175509 215778 175575 215781
rect 175509 215776 179114 215778
rect 175509 215720 175514 215776
rect 175570 215720 179114 215776
rect 175509 215718 179114 215720
rect 175509 215715 175575 215718
rect 179054 215476 179114 215718
rect 81710 215172 81716 215236
rect 81780 215234 81786 215236
rect 85030 215234 85090 215408
rect 81780 215174 85090 215234
rect 81780 215172 81786 215174
rect 137881 214554 137947 214557
rect 231629 214554 231695 214557
rect 134740 214552 137947 214554
rect 134740 214496 137886 214552
rect 137942 214496 137947 214552
rect 134740 214494 137947 214496
rect 228764 214552 231695 214554
rect 228764 214496 231634 214552
rect 231690 214496 231695 214552
rect 228764 214494 231695 214496
rect 137881 214491 137947 214494
rect 231629 214491 231695 214494
rect 148694 214426 148908 214486
rect 145609 214418 145675 214421
rect 148694 214418 148754 214426
rect 145609 214416 148754 214418
rect 145609 214360 145614 214416
rect 145670 214360 148754 214416
rect 145609 214358 148754 214360
rect 145609 214355 145675 214358
rect 240921 213874 240987 213877
rect 242902 213874 242962 214388
rect 240921 213872 242962 213874
rect 240921 213816 240926 213872
rect 240982 213816 242962 213872
rect 240921 213814 242962 213816
rect 240921 213811 240987 213814
rect 134710 212378 134770 212960
rect 164732 212782 164946 212842
rect 164886 212652 164946 212782
rect 164878 212588 164884 212652
rect 164948 212588 164954 212652
rect 137881 212378 137947 212381
rect 134710 212376 137947 212378
rect 134710 212320 137886 212376
rect 137942 212320 137947 212376
rect 134710 212318 137947 212320
rect 228734 212378 228794 212960
rect 261161 212786 261227 212789
rect 262357 212786 262423 212789
rect 258756 212784 262423 212786
rect 258756 212728 261166 212784
rect 261222 212728 262362 212784
rect 262418 212728 262423 212784
rect 258756 212726 262423 212728
rect 261161 212723 261227 212726
rect 262357 212723 262423 212726
rect 231997 212378 232063 212381
rect 228734 212376 232063 212378
rect 228734 212320 232002 212376
rect 232058 212320 232063 212376
rect 228734 212318 232063 212320
rect 137881 212315 137947 212318
rect 231997 212315 232063 212318
rect 145609 212242 145675 212245
rect 145609 212240 148938 212242
rect 145609 212184 145614 212240
rect 145670 212184 148938 212240
rect 145609 212182 148938 212184
rect 145609 212179 145675 212182
rect 148878 212144 148938 212182
rect 240921 211970 240987 211973
rect 242902 211970 242962 212076
rect 240921 211968 242962 211970
rect 240921 211912 240926 211968
rect 240982 211912 242962 211968
rect 240921 211910 242962 211912
rect 240921 211907 240987 211910
rect 134569 211834 134635 211837
rect 135254 211834 135260 211836
rect 134569 211832 135260 211834
rect 134569 211776 134574 211832
rect 134630 211776 135260 211832
rect 134569 211774 135260 211776
rect 134569 211771 134635 211774
rect 135254 211772 135260 211774
rect 135324 211772 135330 211836
rect 137973 211426 138039 211429
rect 231537 211426 231603 211429
rect 134740 211424 138039 211426
rect 134740 211368 137978 211424
rect 138034 211368 138039 211424
rect 134740 211366 138039 211368
rect 228764 211424 231603 211426
rect 228764 211368 231542 211424
rect 231598 211368 231603 211424
rect 228764 211366 231603 211368
rect 137973 211363 138039 211366
rect 231537 211363 231603 211366
rect 38245 211290 38311 211293
rect 35718 211288 38311 211290
rect 35718 211232 38250 211288
rect 38306 211232 38311 211288
rect 35718 211230 38311 211232
rect 35718 210784 35778 211230
rect 38245 211227 38311 211230
rect 145609 209930 145675 209933
rect 145609 209928 148938 209930
rect 145609 209872 145614 209928
rect 145670 209872 148938 209928
rect 145609 209870 148938 209872
rect 145609 209867 145675 209870
rect 148878 209832 148938 209870
rect 134710 209386 134770 209832
rect 228734 209522 228794 209832
rect 231997 209522 232063 209525
rect 228734 209520 232063 209522
rect 228734 209464 232002 209520
rect 232058 209464 232063 209520
rect 228734 209462 232063 209464
rect 231997 209459 232063 209462
rect 137973 209386 138039 209389
rect 134710 209384 138039 209386
rect 134710 209328 137978 209384
rect 138034 209328 138039 209384
rect 134710 209326 138039 209328
rect 137973 209323 138039 209326
rect 240461 209250 240527 209253
rect 242902 209250 242962 209764
rect 240461 209248 242962 209250
rect 240461 209192 240466 209248
rect 240522 209192 242962 209248
rect 240461 209190 242962 209192
rect 240461 209187 240527 209190
rect 274869 208434 274935 208437
rect 274869 208432 278106 208434
rect 274869 208376 274874 208432
rect 274930 208376 278106 208432
rect 274869 208374 278106 208376
rect 274869 208371 274935 208374
rect 138065 208298 138131 208301
rect 231445 208298 231511 208301
rect 134740 208296 138131 208298
rect 134740 208240 138070 208296
rect 138126 208240 138131 208296
rect 134740 208238 138131 208240
rect 228764 208296 231511 208298
rect 228764 208240 231450 208296
rect 231506 208240 231511 208296
rect 228764 208238 231511 208240
rect 138065 208235 138131 208238
rect 231445 208235 231511 208238
rect 278046 207792 278106 208374
rect 145793 207482 145859 207485
rect 145793 207480 148938 207482
rect 145793 207424 145798 207480
rect 145854 207424 148938 207480
rect 145793 207422 148938 207424
rect 145793 207419 145859 207422
rect 148878 207384 148938 207422
rect 240645 206802 240711 206805
rect 242902 206802 242962 207316
rect 240645 206800 242962 206802
rect 240645 206744 240650 206800
rect 240706 206744 242962 206800
rect 240645 206742 242962 206744
rect 240645 206739 240711 206742
rect 134710 206258 134770 206704
rect 228734 206530 228794 206704
rect 231997 206530 232063 206533
rect 228734 206528 232063 206530
rect 228734 206472 232002 206528
rect 232058 206472 232063 206528
rect 228734 206470 232063 206472
rect 231997 206467 232063 206470
rect 138065 206258 138131 206261
rect 134710 206256 138131 206258
rect 134710 206200 138070 206256
rect 138126 206200 138131 206256
rect 134710 206198 138131 206200
rect 138065 206195 138131 206198
rect 138157 205170 138223 205173
rect 134740 205168 138223 205170
rect 134740 205112 138162 205168
rect 138218 205112 138223 205168
rect 134740 205110 138223 205112
rect 138157 205107 138223 205110
rect 145609 205170 145675 205173
rect 231353 205170 231419 205173
rect 145609 205168 148938 205170
rect 145609 205112 145614 205168
rect 145670 205112 148938 205168
rect 145609 205110 148938 205112
rect 228764 205168 231419 205170
rect 228764 205112 231358 205168
rect 231414 205112 231419 205168
rect 228764 205110 231419 205112
rect 145609 205107 145675 205110
rect 148878 205072 148938 205110
rect 231353 205107 231419 205110
rect 240921 204898 240987 204901
rect 242902 204898 242962 205004
rect 240921 204896 242962 204898
rect 240921 204840 240926 204896
rect 240982 204840 242962 204896
rect 240921 204838 242962 204840
rect 240921 204835 240987 204838
rect 134710 203538 134770 203576
rect 138157 203538 138223 203541
rect 134710 203536 138223 203538
rect 134710 203480 138162 203536
rect 138218 203480 138223 203536
rect 134710 203478 138223 203480
rect 228734 203538 228794 203576
rect 231353 203538 231419 203541
rect 228734 203536 231419 203538
rect 228734 203480 231358 203536
rect 231414 203480 231419 203536
rect 228734 203478 231419 203480
rect 138157 203475 138223 203478
rect 231353 203475 231419 203478
rect 38153 203402 38219 203405
rect 35718 203400 38219 203402
rect 35718 203344 38158 203400
rect 38214 203344 38219 203400
rect 35718 203342 38219 203344
rect 20078 202316 20138 202828
rect 35718 202760 35778 203342
rect 38153 203339 38219 203342
rect 52454 202932 52460 202996
rect 52524 202994 52530 202996
rect 52524 202934 54546 202994
rect 52524 202932 52530 202934
rect 54486 202926 54546 202934
rect 54486 202866 55068 202926
rect 70892 202866 71474 202926
rect 71414 202858 71474 202866
rect 74033 202858 74099 202861
rect 71414 202856 74099 202858
rect 71414 202800 74038 202856
rect 74094 202800 74099 202856
rect 71414 202798 74099 202800
rect 74033 202795 74099 202798
rect 145517 202858 145583 202861
rect 296213 202858 296279 202861
rect 145517 202856 148938 202858
rect 145517 202800 145522 202856
rect 145578 202800 148938 202856
rect 145517 202798 148938 202800
rect 293716 202856 296279 202858
rect 293716 202800 296218 202856
rect 296274 202800 296279 202856
rect 293716 202798 296279 202800
rect 145517 202795 145583 202798
rect 148878 202760 148938 202798
rect 296213 202795 296279 202798
rect 240369 202450 240435 202453
rect 242902 202450 242962 202692
rect 240369 202448 242962 202450
rect 240369 202392 240374 202448
rect 240430 202392 242962 202448
rect 240369 202390 242962 202392
rect 240369 202387 240435 202390
rect 20070 202252 20076 202316
rect 20140 202252 20146 202316
rect 228910 202252 228916 202316
rect 228980 202314 228986 202316
rect 242894 202314 242900 202316
rect 228980 202254 242900 202314
rect 228980 202252 228986 202254
rect 242894 202252 242900 202254
rect 242964 202252 242970 202316
rect 258902 202252 258908 202316
rect 258972 202314 258978 202316
rect 278038 202314 278044 202316
rect 258972 202254 278044 202314
rect 258972 202252 258978 202254
rect 278038 202252 278044 202254
rect 278108 202252 278114 202316
rect 293678 202252 293684 202316
rect 293748 202314 293754 202316
rect 300445 202314 300511 202317
rect 293748 202312 300511 202314
rect 293748 202256 300450 202312
rect 300506 202256 300511 202312
rect 293748 202254 300511 202256
rect 293748 202252 293754 202254
rect 300445 202251 300511 202254
rect 35894 202116 35900 202180
rect 35964 202178 35970 202180
rect 51953 202178 52019 202181
rect 35964 202176 52019 202178
rect 35964 202120 51958 202176
rect 52014 202120 52019 202176
rect 35964 202118 52019 202120
rect 35964 202116 35970 202118
rect 51953 202115 52019 202118
rect 137421 202042 137487 202045
rect 231721 202042 231787 202045
rect 134740 202040 137487 202042
rect 134740 201984 137426 202040
rect 137482 201984 137487 202040
rect 134740 201982 137487 201984
rect 228764 202040 231787 202042
rect 228764 201984 231726 202040
rect 231782 201984 231787 202040
rect 228764 201982 231787 201984
rect 137421 201979 137487 201982
rect 231721 201979 231787 201982
rect 137329 200546 137395 200549
rect 134740 200544 137395 200546
rect 134740 200488 137334 200544
rect 137390 200488 137395 200544
rect 134740 200486 137395 200488
rect 137329 200483 137395 200486
rect 144413 200546 144479 200549
rect 231813 200546 231879 200549
rect 144413 200544 148938 200546
rect 144413 200488 144418 200544
rect 144474 200488 148938 200544
rect 144413 200486 148938 200488
rect 228764 200544 231879 200546
rect 228764 200488 231818 200544
rect 231874 200488 231879 200544
rect 228764 200486 231879 200488
rect 144413 200483 144479 200486
rect 148878 200448 148938 200486
rect 231813 200483 231879 200486
rect 240461 199866 240527 199869
rect 242902 199866 242962 200380
rect 240461 199864 242962 199866
rect 240461 199808 240466 199864
rect 240522 199808 242962 199864
rect 240461 199806 242962 199808
rect 240461 199803 240527 199806
rect 137145 198914 137211 198917
rect 231905 198914 231971 198917
rect 134740 198912 137211 198914
rect 134740 198856 137150 198912
rect 137206 198856 137211 198912
rect 134740 198854 137211 198856
rect 228764 198912 231971 198914
rect 228764 198856 231910 198912
rect 231966 198856 231971 198912
rect 228764 198854 231971 198856
rect 137145 198851 137211 198854
rect 231905 198851 231971 198854
rect 145609 198098 145675 198101
rect 240921 198098 240987 198101
rect 145609 198096 148938 198098
rect 145609 198040 145614 198096
rect 145670 198040 148938 198096
rect 145609 198038 148938 198040
rect 145609 198035 145675 198038
rect 148878 198000 148938 198038
rect 240921 198096 242962 198098
rect 240921 198040 240926 198096
rect 240982 198040 242962 198096
rect 240921 198038 242962 198040
rect 240921 198035 240987 198038
rect 242902 198000 242962 198038
rect 274869 197690 274935 197693
rect 274869 197688 278076 197690
rect 274869 197632 274874 197688
rect 274930 197632 278076 197688
rect 274869 197630 278076 197632
rect 274869 197627 274935 197630
rect 137237 197418 137303 197421
rect 231629 197418 231695 197421
rect 134740 197416 137303 197418
rect 134740 197360 137242 197416
rect 137298 197360 137303 197416
rect 134740 197358 137303 197360
rect 228764 197416 231695 197418
rect 228764 197360 231634 197416
rect 231690 197360 231695 197416
rect 228764 197358 231695 197360
rect 137237 197355 137303 197358
rect 231629 197355 231695 197358
rect 137053 195786 137119 195789
rect 134740 195784 137119 195786
rect 134740 195728 137058 195784
rect 137114 195728 137119 195784
rect 134740 195726 137119 195728
rect 137053 195723 137119 195726
rect 145609 195786 145675 195789
rect 231537 195786 231603 195789
rect 145609 195784 148938 195786
rect 145609 195728 145614 195784
rect 145670 195728 148938 195784
rect 145609 195726 148938 195728
rect 228764 195784 231603 195786
rect 228764 195728 231542 195784
rect 231598 195728 231603 195784
rect 228764 195726 231603 195728
rect 145609 195723 145675 195726
rect 148878 195688 148938 195726
rect 231537 195723 231603 195726
rect 240921 195242 240987 195245
rect 242902 195242 242962 195620
rect 240921 195240 242962 195242
rect 240921 195184 240926 195240
rect 240982 195184 242962 195240
rect 240921 195182 242962 195184
rect 240921 195179 240987 195182
rect 38153 194698 38219 194701
rect 35748 194696 38219 194698
rect 35748 194640 38158 194696
rect 38214 194640 38219 194696
rect 35748 194638 38219 194640
rect 38153 194635 38219 194638
rect 137421 194290 137487 194293
rect 231997 194290 232063 194293
rect 134740 194288 137487 194290
rect 134740 194232 137426 194288
rect 137482 194232 137487 194288
rect 134740 194230 137487 194232
rect 228764 194288 232063 194290
rect 228764 194232 232002 194288
rect 232058 194232 232063 194288
rect 228764 194230 232063 194232
rect 137421 194227 137487 194230
rect 231997 194227 232063 194230
rect 145793 193474 145859 193477
rect 145793 193472 148938 193474
rect 145793 193416 145798 193472
rect 145854 193416 148938 193472
rect 145793 193414 148938 193416
rect 145793 193411 145859 193414
rect 148878 193376 148938 193414
rect 164732 192794 165314 192850
rect 167873 192794 167939 192797
rect 164732 192792 167939 192794
rect 164732 192790 167878 192792
rect 165254 192736 167878 192790
rect 167934 192736 167939 192792
rect 165254 192734 167939 192736
rect 167873 192731 167939 192734
rect 240461 192794 240527 192797
rect 242902 192794 242962 193308
rect 262357 192794 262423 192797
rect 240461 192792 242962 192794
rect 240461 192736 240466 192792
rect 240522 192736 242962 192792
rect 240461 192734 242962 192736
rect 258756 192792 262423 192794
rect 258756 192736 262362 192792
rect 262418 192736 262423 192792
rect 258756 192734 262423 192736
rect 240461 192731 240527 192734
rect 262357 192731 262423 192734
rect 136961 192658 137027 192661
rect 231445 192658 231511 192661
rect 134740 192656 137027 192658
rect 134740 192600 136966 192656
rect 137022 192600 137027 192656
rect 134740 192598 137027 192600
rect 228764 192656 231511 192658
rect 228764 192600 231450 192656
rect 231506 192600 231511 192656
rect 228764 192598 231511 192600
rect 136961 192595 137027 192598
rect 231445 192595 231511 192598
rect 300445 192658 300511 192661
rect 303416 192658 303896 192688
rect 300445 192656 303896 192658
rect 300445 192600 300450 192656
rect 300506 192600 303896 192656
rect 300445 192598 303896 192600
rect 300445 192595 300511 192598
rect 303416 192568 303896 192598
rect 137421 191162 137487 191165
rect 231261 191162 231327 191165
rect 134740 191160 137487 191162
rect 134740 191104 137426 191160
rect 137482 191104 137487 191160
rect 134740 191102 137487 191104
rect 228764 191160 231327 191162
rect 228764 191104 231266 191160
rect 231322 191104 231327 191160
rect 228764 191102 231327 191104
rect 137421 191099 137487 191102
rect 231261 191099 231327 191102
rect 148326 190898 148908 190958
rect 145149 190890 145215 190893
rect 148326 190890 148386 190898
rect 145149 190888 148386 190890
rect 145149 190832 145154 190888
rect 145210 190832 148386 190888
rect 145149 190830 148386 190832
rect 175509 190890 175575 190893
rect 175509 190888 179114 190890
rect 175509 190832 175514 190888
rect 175570 190832 179114 190888
rect 175509 190830 179114 190832
rect 145149 190827 145215 190830
rect 175509 190827 175575 190830
rect 81669 190482 81735 190485
rect 81669 190480 85060 190482
rect 81669 190424 81674 190480
rect 81730 190424 85060 190480
rect 179054 190452 179114 190830
rect 81669 190422 85060 190424
rect 81669 190419 81735 190422
rect 240645 190346 240711 190349
rect 242902 190346 242962 190860
rect 240645 190344 242962 190346
rect 240645 190288 240650 190344
rect 240706 190288 242962 190344
rect 240645 190286 242962 190288
rect 240645 190283 240711 190286
rect 51309 189530 51375 189533
rect 54486 189530 55068 189586
rect 137421 189530 137487 189533
rect 231721 189530 231787 189533
rect 51309 189528 55068 189530
rect 51309 189472 51314 189528
rect 51370 189526 55068 189528
rect 134740 189528 137487 189530
rect 51370 189472 54546 189526
rect 51309 189470 54546 189472
rect 134740 189472 137426 189528
rect 137482 189472 137487 189528
rect 134740 189470 137487 189472
rect 228764 189528 231787 189530
rect 228764 189472 231726 189528
rect 231782 189472 231787 189528
rect 228764 189470 231787 189472
rect 51309 189467 51375 189470
rect 137421 189467 137487 189470
rect 231721 189467 231787 189470
rect 293502 188989 293562 189500
rect 293502 188984 293611 188989
rect 293502 188928 293550 188984
rect 293606 188928 293611 188984
rect 293502 188926 293611 188928
rect 293545 188923 293611 188926
rect 145609 188714 145675 188717
rect 145609 188712 148938 188714
rect 145609 188656 145614 188712
rect 145670 188656 148938 188712
rect 145609 188654 148938 188656
rect 145609 188651 145675 188654
rect 148878 188616 148938 188654
rect 9896 188578 10376 188608
rect 13497 188578 13563 188581
rect 9896 188576 13563 188578
rect 9896 188520 13502 188576
rect 13558 188520 13563 188576
rect 9896 188518 13563 188520
rect 9896 188488 10376 188518
rect 13497 188515 13563 188518
rect 240737 188306 240803 188309
rect 242902 188306 242962 188548
rect 240737 188304 242962 188306
rect 240737 188248 240742 188304
rect 240798 188248 242962 188304
rect 240737 188246 242962 188248
rect 240737 188243 240803 188246
rect 275513 188170 275579 188173
rect 275513 188168 278106 188170
rect 275513 188112 275518 188168
rect 275574 188112 278106 188168
rect 275513 188110 278106 188112
rect 275513 188107 275579 188110
rect 137421 188034 137487 188037
rect 231813 188034 231879 188037
rect 134740 188032 137487 188034
rect 134740 187976 137426 188032
rect 137482 187976 137487 188032
rect 134740 187974 137487 187976
rect 228764 188032 231879 188034
rect 228764 187976 231818 188032
rect 231874 187976 231879 188032
rect 228764 187974 231879 187976
rect 137421 187971 137487 187974
rect 231813 187971 231879 187974
rect 278046 187800 278106 188110
rect 38797 186810 38863 186813
rect 35748 186808 38863 186810
rect 35748 186752 38802 186808
rect 38858 186752 38863 186808
rect 35748 186750 38863 186752
rect 38797 186747 38863 186750
rect 137421 186402 137487 186405
rect 134740 186400 137487 186402
rect 134740 186344 137426 186400
rect 137482 186344 137487 186400
rect 134740 186342 137487 186344
rect 137421 186339 137487 186342
rect 144781 186402 144847 186405
rect 231813 186402 231879 186405
rect 144781 186400 148938 186402
rect 144781 186344 144786 186400
rect 144842 186344 148938 186400
rect 144781 186342 148938 186344
rect 228764 186400 231879 186402
rect 228764 186344 231818 186400
rect 231874 186344 231879 186400
rect 228764 186342 231879 186344
rect 144781 186339 144847 186342
rect 148878 186304 148938 186342
rect 231813 186339 231879 186342
rect 240921 185858 240987 185861
rect 242902 185858 242962 186236
rect 240921 185856 242962 185858
rect 240921 185800 240926 185856
rect 240982 185800 242962 185856
rect 240921 185798 242962 185800
rect 240921 185795 240987 185798
rect 231813 184906 231879 184909
rect 228764 184904 231879 184906
rect 228764 184848 231818 184904
rect 231874 184848 231879 184904
rect 228764 184846 231879 184848
rect 231813 184843 231879 184846
rect 134710 184634 134770 184808
rect 137421 184634 137487 184637
rect 134710 184632 137487 184634
rect 134710 184576 137426 184632
rect 137482 184576 137487 184632
rect 134710 184574 137487 184576
rect 137421 184571 137487 184574
rect 145793 183410 145859 183413
rect 149062 183410 149122 183924
rect 145793 183408 149122 183410
rect 145793 183352 145798 183408
rect 145854 183352 149122 183408
rect 145793 183350 149122 183352
rect 239633 183410 239699 183413
rect 242902 183410 242962 183924
rect 239633 183408 242962 183410
rect 239633 183352 239638 183408
rect 239694 183352 242962 183408
rect 239633 183350 242962 183352
rect 145793 183347 145859 183350
rect 239633 183347 239699 183350
rect 137053 183274 137119 183277
rect 230801 183274 230867 183277
rect 134740 183272 137119 183274
rect 134740 183216 137058 183272
rect 137114 183216 137119 183272
rect 134740 183214 137119 183216
rect 228764 183272 230867 183274
rect 228764 183216 230806 183272
rect 230862 183216 230867 183272
rect 228764 183214 230867 183216
rect 137053 183211 137119 183214
rect 230801 183211 230867 183214
rect 137329 181778 137395 181781
rect 231261 181778 231327 181781
rect 134740 181776 137395 181778
rect 134740 181720 137334 181776
rect 137390 181720 137395 181776
rect 134740 181718 137395 181720
rect 228764 181776 231327 181778
rect 228764 181720 231266 181776
rect 231322 181720 231327 181776
rect 228764 181718 231327 181720
rect 137329 181715 137395 181718
rect 231261 181715 231327 181718
rect 241606 181172 241612 181236
rect 241676 181234 241682 181236
rect 285909 181234 285975 181237
rect 241676 181232 285975 181234
rect 241676 181176 285914 181232
rect 285970 181176 285975 181232
rect 241676 181174 285975 181176
rect 241676 181172 241682 181174
rect 285909 181171 285975 181174
rect 137421 180146 137487 180149
rect 231629 180146 231695 180149
rect 134740 180144 137487 180146
rect 134740 180088 137426 180144
rect 137482 180088 137487 180144
rect 134740 180086 137487 180088
rect 228764 180144 231695 180146
rect 228764 180088 231634 180144
rect 231690 180088 231695 180144
rect 228764 180086 231695 180088
rect 137421 180083 137487 180086
rect 231629 180083 231695 180086
rect 137421 178650 137487 178653
rect 231629 178650 231695 178653
rect 134740 178648 137487 178650
rect 134740 178592 137426 178648
rect 137482 178592 137487 178648
rect 134740 178590 137487 178592
rect 228764 178648 231695 178650
rect 228764 178592 231634 178648
rect 231690 178592 231695 178648
rect 228764 178590 231695 178592
rect 137421 178587 137487 178590
rect 231629 178587 231695 178590
rect 85022 174644 85028 174708
rect 85092 174706 85098 174708
rect 85533 174706 85599 174709
rect 85092 174704 85599 174706
rect 85092 174648 85538 174704
rect 85594 174648 85599 174704
rect 85092 174646 85599 174648
rect 85092 174644 85098 174646
rect 85533 174643 85599 174646
rect 132729 174706 132795 174709
rect 133230 174706 133236 174708
rect 132729 174704 133236 174706
rect 132729 174648 132734 174704
rect 132790 174648 133236 174704
rect 132729 174646 133236 174648
rect 132729 174643 132795 174646
rect 133230 174644 133236 174646
rect 133300 174644 133306 174708
rect 127301 174570 127367 174573
rect 128446 174570 128452 174572
rect 127301 174568 128452 174570
rect 127301 174512 127306 174568
rect 127362 174512 128452 174568
rect 127301 174510 128452 174512
rect 127301 174507 127367 174510
rect 128446 174508 128452 174510
rect 128516 174508 128522 174572
rect 154625 172938 154691 172941
rect 166309 172938 166375 172941
rect 154625 172936 166375 172938
rect 154625 172880 154630 172936
rect 154686 172880 166314 172936
rect 166370 172880 166375 172936
rect 154625 172878 166375 172880
rect 154625 172875 154691 172878
rect 166309 172875 166375 172878
rect 60877 172802 60943 172805
rect 73021 172802 73087 172805
rect 60877 172800 73087 172802
rect 60877 172744 60882 172800
rect 60938 172744 73026 172800
rect 73082 172744 73087 172800
rect 60877 172742 73087 172744
rect 60877 172739 60943 172742
rect 73021 172739 73087 172742
rect 154257 172802 154323 172805
rect 165849 172802 165915 172805
rect 154257 172800 165915 172802
rect 154257 172744 154262 172800
rect 154318 172744 165854 172800
rect 165910 172744 165915 172800
rect 154257 172742 165915 172744
rect 154257 172739 154323 172742
rect 165849 172739 165915 172742
rect 249937 172802 250003 172805
rect 261069 172802 261135 172805
rect 249937 172800 261135 172802
rect 249937 172744 249942 172800
rect 249998 172744 261074 172800
rect 261130 172744 261135 172800
rect 249937 172742 261135 172744
rect 249937 172739 250003 172742
rect 261069 172739 261135 172742
rect 59497 172666 59563 172669
rect 70997 172666 71063 172669
rect 59497 172664 71063 172666
rect 59497 172608 59502 172664
rect 59558 172608 71002 172664
rect 71058 172608 71063 172664
rect 59497 172606 71063 172608
rect 59497 172603 59563 172606
rect 70997 172603 71063 172606
rect 137697 172666 137763 172669
rect 157569 172666 157635 172669
rect 137697 172664 157635 172666
rect 137697 172608 137702 172664
rect 137758 172608 157574 172664
rect 157630 172608 157635 172664
rect 137697 172606 157635 172608
rect 137697 172603 137763 172606
rect 157569 172603 157635 172606
rect 251041 172666 251107 172669
rect 262541 172666 262607 172669
rect 251041 172664 262607 172666
rect 251041 172608 251046 172664
rect 251102 172608 262546 172664
rect 262602 172608 262607 172664
rect 251041 172606 262607 172608
rect 251041 172603 251107 172606
rect 262541 172603 262607 172606
rect 60693 172530 60759 172533
rect 72377 172530 72443 172533
rect 60693 172528 72443 172530
rect 60693 172472 60698 172528
rect 60754 172472 72382 172528
rect 72438 172472 72443 172528
rect 60693 172470 72443 172472
rect 60693 172467 60759 172470
rect 72377 172467 72443 172470
rect 137513 172530 137579 172533
rect 157937 172530 158003 172533
rect 137513 172528 158003 172530
rect 137513 172472 137518 172528
rect 137574 172472 157942 172528
rect 157998 172472 158003 172528
rect 137513 172470 158003 172472
rect 137513 172467 137579 172470
rect 157937 172467 158003 172470
rect 158305 172530 158371 172533
rect 164469 172530 164535 172533
rect 158305 172528 164535 172530
rect 158305 172472 158310 172528
rect 158366 172472 164474 172528
rect 164530 172472 164535 172528
rect 158305 172470 164535 172472
rect 158305 172467 158371 172470
rect 164469 172467 164535 172470
rect 249477 172530 249543 172533
rect 261437 172530 261503 172533
rect 249477 172528 261503 172530
rect 249477 172472 249482 172528
rect 249538 172472 261442 172528
rect 261498 172472 261503 172528
rect 249477 172470 261503 172472
rect 249477 172467 249543 172470
rect 261437 172467 261503 172470
rect 61889 172394 61955 172397
rect 75781 172394 75847 172397
rect 61889 172392 75847 172394
rect 61889 172336 61894 172392
rect 61950 172336 75786 172392
rect 75842 172336 75847 172392
rect 61889 172334 75847 172336
rect 61889 172331 61955 172334
rect 75781 172331 75847 172334
rect 113869 172394 113935 172397
rect 170173 172394 170239 172397
rect 113869 172392 170239 172394
rect 113869 172336 113874 172392
rect 113930 172336 170178 172392
rect 170234 172336 170239 172392
rect 113869 172334 170239 172336
rect 113869 172331 113935 172334
rect 170173 172331 170239 172334
rect 218657 172394 218723 172397
rect 264197 172394 264263 172397
rect 218657 172392 264263 172394
rect 218657 172336 218662 172392
rect 218718 172336 264202 172392
rect 264258 172336 264263 172392
rect 218657 172334 264263 172336
rect 218657 172331 218723 172334
rect 264197 172331 264263 172334
rect 62165 172258 62231 172261
rect 75045 172258 75111 172261
rect 62165 172256 75111 172258
rect 62165 172200 62170 172256
rect 62226 172200 75050 172256
rect 75106 172200 75111 172256
rect 62165 172198 75111 172200
rect 62165 172195 62231 172198
rect 75045 172195 75111 172198
rect 108441 172258 108507 172261
rect 169989 172258 170055 172261
rect 108441 172256 170055 172258
rect 108441 172200 108446 172256
rect 108502 172200 169994 172256
rect 170050 172200 170055 172256
rect 108441 172198 170055 172200
rect 108441 172195 108507 172198
rect 169989 172195 170055 172198
rect 207893 172258 207959 172261
rect 263829 172258 263895 172261
rect 207893 172256 263895 172258
rect 207893 172200 207898 172256
rect 207954 172200 263834 172256
rect 263890 172200 263895 172256
rect 207893 172198 263895 172200
rect 207893 172195 207959 172198
rect 263829 172195 263895 172198
rect 80013 169538 80079 169541
rect 76780 169536 80079 169538
rect 76780 169480 80018 169536
rect 80074 169480 80079 169536
rect 76780 169478 80079 169480
rect 80013 169475 80079 169478
rect 139629 169538 139695 169541
rect 171369 169538 171435 169541
rect 139629 169536 143020 169538
rect 139629 169480 139634 169536
rect 139690 169480 143020 169536
rect 139629 169478 143020 169480
rect 170804 169536 171435 169538
rect 170804 169480 171374 169536
rect 171430 169480 171435 169536
rect 170804 169478 171435 169480
rect 139629 169475 139695 169478
rect 171369 169475 171435 169478
rect 233469 169538 233535 169541
rect 233469 169536 237044 169538
rect 233469 169480 233474 169536
rect 233530 169480 237044 169536
rect 233469 169478 237044 169480
rect 233469 169475 233535 169478
rect 170725 169266 170791 169269
rect 170725 169264 170834 169266
rect 170725 169208 170730 169264
rect 170786 169208 170834 169264
rect 170725 169203 170834 169208
rect 80197 168994 80263 168997
rect 76780 168992 80263 168994
rect 76780 168936 80202 168992
rect 80258 168936 80263 168992
rect 170774 168964 170834 169203
rect 76780 168934 80263 168936
rect 80197 168931 80263 168934
rect 139629 168858 139695 168861
rect 233469 168858 233535 168861
rect 139629 168856 143020 168858
rect 139629 168800 139634 168856
rect 139690 168800 143020 168856
rect 139629 168798 143020 168800
rect 233469 168856 237044 168858
rect 233469 168800 233474 168856
rect 233530 168800 237044 168856
rect 233469 168798 237044 168800
rect 139629 168795 139695 168798
rect 233469 168795 233535 168798
rect 79921 168450 79987 168453
rect 173301 168450 173367 168453
rect 76780 168448 79987 168450
rect 76780 168392 79926 168448
rect 79982 168392 79987 168448
rect 76780 168390 79987 168392
rect 170804 168448 173367 168450
rect 170804 168392 173306 168448
rect 173362 168392 173367 168448
rect 170804 168390 173367 168392
rect 79921 168387 79987 168390
rect 173301 168387 173367 168390
rect 233653 168178 233719 168181
rect 300169 168178 300235 168181
rect 303416 168178 303896 168208
rect 233653 168176 237044 168178
rect 233653 168120 233658 168176
rect 233714 168120 237044 168176
rect 233653 168118 237044 168120
rect 300169 168176 303896 168178
rect 300169 168120 300174 168176
rect 300230 168120 303896 168176
rect 300169 168118 303896 168120
rect 233653 168115 233719 168118
rect 300169 168115 300235 168118
rect 303416 168088 303896 168118
rect 80105 167770 80171 167773
rect 76780 167768 80171 167770
rect 76780 167712 80110 167768
rect 80166 167712 80171 167768
rect 76780 167710 80171 167712
rect 80105 167707 80171 167710
rect 140825 167770 140891 167773
rect 142990 167770 143050 168080
rect 174037 167906 174103 167909
rect 170804 167904 174103 167906
rect 170804 167848 174042 167904
rect 174098 167848 174103 167904
rect 170804 167846 174103 167848
rect 174037 167843 174103 167846
rect 140825 167768 143050 167770
rect 140825 167712 140830 167768
rect 140886 167712 143050 167768
rect 140825 167710 143050 167712
rect 140825 167707 140891 167710
rect 236689 167566 236755 167569
rect 236689 167564 237044 167566
rect 236689 167508 236694 167564
rect 236750 167508 237044 167564
rect 236689 167506 237044 167508
rect 236689 167503 236755 167506
rect 79829 167226 79895 167229
rect 76780 167224 79895 167226
rect 76780 167168 79834 167224
rect 79890 167168 79895 167224
rect 76780 167166 79895 167168
rect 79829 167163 79895 167166
rect 139721 167090 139787 167093
rect 142990 167090 143050 167400
rect 173301 167362 173367 167365
rect 170804 167360 173367 167362
rect 170804 167304 173306 167360
rect 173362 167304 173367 167360
rect 170804 167302 173367 167304
rect 173301 167299 173367 167302
rect 139721 167088 143050 167090
rect 139721 167032 139726 167088
rect 139782 167032 143050 167088
rect 139721 167030 143050 167032
rect 139721 167027 139787 167030
rect 233469 166954 233535 166957
rect 233469 166952 237044 166954
rect 233469 166896 233474 166952
rect 233530 166896 237044 166952
rect 233469 166894 237044 166896
rect 233469 166891 233535 166894
rect 173117 166818 173183 166821
rect 170804 166816 173183 166818
rect 170804 166760 173122 166816
rect 173178 166760 173183 166816
rect 170804 166758 173183 166760
rect 173117 166755 173183 166758
rect 79645 166682 79711 166685
rect 76780 166680 79711 166682
rect 76780 166624 79650 166680
rect 79706 166624 79711 166680
rect 76780 166622 79711 166624
rect 79645 166619 79711 166622
rect 139629 166546 139695 166549
rect 142990 166546 143050 166720
rect 139629 166544 143050 166546
rect 139629 166488 139634 166544
rect 139690 166488 143050 166544
rect 139629 166486 143050 166488
rect 139629 166483 139695 166486
rect 173117 166274 173183 166277
rect 170804 166272 173183 166274
rect 170804 166216 173122 166272
rect 173178 166216 173183 166272
rect 170804 166214 173183 166216
rect 173117 166211 173183 166214
rect 233469 166274 233535 166277
rect 233469 166272 237044 166274
rect 233469 166216 233474 166272
rect 233530 166216 237044 166272
rect 233469 166214 237044 166216
rect 233469 166211 233535 166214
rect 79553 166002 79619 166005
rect 76780 166000 79619 166002
rect 76780 165944 79558 166000
rect 79614 165944 79619 166000
rect 76780 165942 79619 165944
rect 79553 165939 79619 165942
rect 139077 165730 139143 165733
rect 142990 165730 143050 166040
rect 174037 165730 174103 165733
rect 139077 165728 143050 165730
rect 139077 165672 139082 165728
rect 139138 165672 143050 165728
rect 139077 165670 143050 165672
rect 170804 165728 174103 165730
rect 170804 165672 174042 165728
rect 174098 165672 174103 165728
rect 170804 165670 174103 165672
rect 139077 165667 139143 165670
rect 174037 165667 174103 165670
rect 233561 165730 233627 165733
rect 233561 165728 237044 165730
rect 233561 165672 233566 165728
rect 233622 165672 237044 165728
rect 233561 165670 237044 165672
rect 233561 165667 233627 165670
rect 79737 165458 79803 165461
rect 76780 165456 79803 165458
rect 76780 165400 79742 165456
rect 79798 165400 79803 165456
rect 76780 165398 79803 165400
rect 79737 165395 79803 165398
rect 138985 165050 139051 165053
rect 142990 165050 143050 165360
rect 173945 165050 174011 165053
rect 138985 165048 143050 165050
rect 138985 164992 138990 165048
rect 139046 164992 143050 165048
rect 138985 164990 143050 164992
rect 170804 165048 174011 165050
rect 170804 164992 173950 165048
rect 174006 164992 174011 165048
rect 170804 164990 174011 164992
rect 138985 164987 139051 164990
rect 173945 164987 174011 164990
rect 233469 165050 233535 165053
rect 233469 165048 237044 165050
rect 233469 164992 233474 165048
rect 233530 164992 237044 165048
rect 233469 164990 237044 164992
rect 233469 164987 233535 164990
rect 80197 164914 80263 164917
rect 76780 164912 80263 164914
rect 76780 164856 80202 164912
rect 80258 164856 80263 164912
rect 76780 164854 80263 164856
rect 80197 164851 80263 164854
rect 87189 164370 87255 164373
rect 140365 164370 140431 164373
rect 142990 164370 143050 164680
rect 173025 164506 173091 164509
rect 170804 164504 173091 164506
rect 170804 164448 173030 164504
rect 173086 164448 173091 164504
rect 170804 164446 173091 164448
rect 173025 164443 173091 164446
rect 87189 164368 90058 164370
rect 87189 164312 87194 164368
rect 87250 164312 90058 164368
rect 87189 164310 90058 164312
rect 87189 164307 87255 164310
rect 76750 164098 76810 164272
rect 80197 164098 80263 164101
rect 76750 164096 80263 164098
rect 76750 164040 80202 164096
rect 80258 164040 80263 164096
rect 76750 164038 80263 164040
rect 80197 164035 80263 164038
rect 89998 163728 90058 164310
rect 140365 164368 143050 164370
rect 140365 164312 140370 164368
rect 140426 164312 143050 164368
rect 140365 164310 143050 164312
rect 233745 164370 233811 164373
rect 233745 164368 237044 164370
rect 233745 164312 233750 164368
rect 233806 164312 237044 164368
rect 233745 164310 237044 164312
rect 140365 164307 140431 164310
rect 233745 164307 233811 164310
rect 140549 163826 140615 163829
rect 142990 163826 143050 164000
rect 173209 163962 173275 163965
rect 170804 163960 173275 163962
rect 170804 163904 173214 163960
rect 173270 163904 173275 163960
rect 170804 163902 173275 163904
rect 173209 163899 173275 163902
rect 140549 163824 143050 163826
rect 140549 163768 140554 163824
rect 140610 163768 143050 163824
rect 140549 163766 143050 163768
rect 233837 163826 233903 163829
rect 233837 163824 237044 163826
rect 233837 163768 233842 163824
rect 233898 163768 237044 163824
rect 233837 163766 237044 163768
rect 140549 163763 140615 163766
rect 233837 163763 233903 163766
rect 80197 163690 80263 163693
rect 131993 163690 132059 163693
rect 76780 163688 80263 163690
rect 76780 163632 80202 163688
rect 80258 163632 80263 163688
rect 76780 163630 80263 163632
rect 129772 163688 132059 163690
rect 129772 163632 131998 163688
rect 132054 163632 132059 163688
rect 129772 163630 132059 163632
rect 80197 163627 80263 163630
rect 131993 163627 132059 163630
rect 181765 163690 181831 163693
rect 225925 163690 225991 163693
rect 181765 163688 184052 163690
rect 181765 163632 181770 163688
rect 181826 163632 184052 163688
rect 181765 163630 184052 163632
rect 223796 163688 225991 163690
rect 223796 163632 225930 163688
rect 225986 163632 225991 163688
rect 223796 163630 225991 163632
rect 181765 163627 181831 163630
rect 225925 163627 225991 163630
rect 140641 163418 140707 163421
rect 174037 163418 174103 163421
rect 140641 163416 143020 163418
rect 140641 163360 140646 163416
rect 140702 163360 143020 163416
rect 140641 163358 143020 163360
rect 170804 163416 174103 163418
rect 170804 163360 174042 163416
rect 174098 163360 174103 163416
rect 170804 163358 174103 163360
rect 140641 163355 140707 163358
rect 174037 163355 174103 163358
rect 228685 163418 228751 163421
rect 228869 163418 228935 163421
rect 228685 163416 228935 163418
rect 228685 163360 228690 163416
rect 228746 163360 228874 163416
rect 228930 163360 228935 163416
rect 228685 163358 228935 163360
rect 228685 163355 228751 163358
rect 228869 163355 228935 163358
rect 87281 163282 87347 163285
rect 132453 163282 132519 163285
rect 87281 163280 90028 163282
rect 87281 163224 87286 163280
rect 87342 163224 90028 163280
rect 87281 163222 90028 163224
rect 129772 163280 132519 163282
rect 129772 163224 132458 163280
rect 132514 163224 132519 163280
rect 129772 163222 132519 163224
rect 87281 163219 87347 163222
rect 132453 163219 132519 163222
rect 180937 163282 181003 163285
rect 226385 163282 226451 163285
rect 264841 163282 264907 163285
rect 180937 163280 184052 163282
rect 180937 163224 180942 163280
rect 180998 163224 184052 163280
rect 180937 163222 184052 163224
rect 223796 163280 226451 163282
rect 223796 163224 226390 163280
rect 226446 163224 226451 163280
rect 223796 163222 226451 163224
rect 180937 163219 181003 163222
rect 226385 163219 226451 163222
rect 264798 163280 264907 163282
rect 264798 163224 264846 163280
rect 264902 163224 264907 163280
rect 264798 163219 264907 163224
rect 80105 163146 80171 163149
rect 76780 163144 80171 163146
rect 76780 163088 80110 163144
rect 80166 163088 80171 163144
rect 76780 163086 80171 163088
rect 80105 163083 80171 163086
rect 233561 163146 233627 163149
rect 233561 163144 237044 163146
rect 233561 163088 233566 163144
rect 233622 163088 237044 163144
rect 233561 163086 237044 163088
rect 233561 163083 233627 163086
rect 46985 162874 47051 162877
rect 87189 162874 87255 162877
rect 132545 162874 132611 162877
rect 172933 162874 172999 162877
rect 46985 162872 48996 162874
rect 46985 162816 46990 162872
rect 47046 162816 48996 162872
rect 46985 162814 48996 162816
rect 87189 162872 90028 162874
rect 87189 162816 87194 162872
rect 87250 162816 90028 162872
rect 87189 162814 90028 162816
rect 129772 162872 132611 162874
rect 129772 162816 132550 162872
rect 132606 162816 132611 162872
rect 129772 162814 132611 162816
rect 170804 162872 172999 162874
rect 170804 162816 172938 162872
rect 172994 162816 172999 162872
rect 170804 162814 172999 162816
rect 46985 162811 47051 162814
rect 87189 162811 87255 162814
rect 132545 162811 132611 162814
rect 172933 162811 172999 162814
rect 181121 162874 181187 162877
rect 226477 162874 226543 162877
rect 181121 162872 184052 162874
rect 181121 162816 181126 162872
rect 181182 162816 184052 162872
rect 181121 162814 184052 162816
rect 223796 162872 226543 162874
rect 223796 162816 226482 162872
rect 226538 162816 226543 162872
rect 264798 162844 264858 163219
rect 223796 162814 226543 162816
rect 181121 162811 181187 162814
rect 226477 162811 226543 162814
rect 80197 162602 80263 162605
rect 76780 162600 80263 162602
rect 76780 162544 80202 162600
rect 80258 162544 80263 162600
rect 76780 162542 80263 162544
rect 80197 162539 80263 162542
rect 140457 162602 140523 162605
rect 142990 162602 143050 162776
rect 140457 162600 143050 162602
rect 140457 162544 140462 162600
rect 140518 162544 143050 162600
rect 140457 162542 143050 162544
rect 140457 162539 140523 162542
rect 87189 162466 87255 162469
rect 132637 162466 132703 162469
rect 87189 162464 90028 162466
rect 87189 162408 87194 162464
rect 87250 162408 90028 162464
rect 87189 162406 90028 162408
rect 129772 162464 132703 162466
rect 129772 162408 132642 162464
rect 132698 162408 132703 162464
rect 129772 162406 132703 162408
rect 87189 162403 87255 162406
rect 132637 162403 132703 162406
rect 181213 162466 181279 162469
rect 225557 162466 225623 162469
rect 181213 162464 184052 162466
rect 181213 162408 181218 162464
rect 181274 162408 184052 162464
rect 181213 162406 184052 162408
rect 223796 162464 225623 162466
rect 223796 162408 225562 162464
rect 225618 162408 225623 162464
rect 223796 162406 225623 162408
rect 181213 162403 181279 162406
rect 225557 162403 225623 162406
rect 233469 162466 233535 162469
rect 233469 162464 237044 162466
rect 233469 162408 233474 162464
rect 233530 162408 237044 162464
rect 233469 162406 237044 162408
rect 233469 162403 233535 162406
rect 172933 162330 172999 162333
rect 170804 162328 172999 162330
rect 170804 162272 172938 162328
rect 172994 162272 172999 162328
rect 170804 162270 172999 162272
rect 172933 162267 172999 162270
rect 140549 162194 140615 162197
rect 140549 162192 143020 162194
rect 140549 162136 140554 162192
rect 140610 162136 143020 162192
rect 140549 162134 143020 162136
rect 140549 162131 140615 162134
rect 87281 162058 87347 162061
rect 132637 162058 132703 162061
rect 87281 162056 90028 162058
rect 87281 162000 87286 162056
rect 87342 162000 90028 162056
rect 87281 161998 90028 162000
rect 129772 162056 132703 162058
rect 129772 162000 132642 162056
rect 132698 162000 132703 162056
rect 129772 161998 132703 162000
rect 87281 161995 87347 161998
rect 132637 161995 132703 161998
rect 182317 162058 182383 162061
rect 225925 162058 225991 162061
rect 182317 162056 184052 162058
rect 182317 162000 182322 162056
rect 182378 162000 184052 162056
rect 182317 161998 184052 162000
rect 223796 162056 225991 162058
rect 223796 162000 225930 162056
rect 225986 162000 225991 162056
rect 223796 161998 225991 162000
rect 182317 161995 182383 161998
rect 225925 161995 225991 161998
rect 233653 161922 233719 161925
rect 233653 161920 237044 161922
rect 233653 161864 233658 161920
rect 233714 161864 237044 161920
rect 233653 161862 237044 161864
rect 233653 161859 233719 161862
rect 76750 161650 76810 161824
rect 173945 161786 174011 161789
rect 170804 161784 174011 161786
rect 170804 161728 173950 161784
rect 174006 161728 174011 161784
rect 170804 161726 174011 161728
rect 173945 161723 174011 161726
rect 80013 161650 80079 161653
rect 76750 161648 80079 161650
rect 76750 161592 80018 161648
rect 80074 161592 80079 161648
rect 76750 161590 80079 161592
rect 80013 161587 80079 161590
rect 87281 161650 87347 161653
rect 132637 161650 132703 161653
rect 87281 161648 90028 161650
rect 87281 161592 87286 161648
rect 87342 161592 90028 161648
rect 87281 161590 90028 161592
rect 129772 161648 132703 161650
rect 129772 161592 132642 161648
rect 132698 161592 132703 161648
rect 129772 161590 132703 161592
rect 87281 161587 87347 161590
rect 132637 161587 132703 161590
rect 182317 161650 182383 161653
rect 226477 161650 226543 161653
rect 182317 161648 184052 161650
rect 182317 161592 182322 161648
rect 182378 161592 184052 161648
rect 182317 161590 184052 161592
rect 223796 161648 226543 161650
rect 223796 161592 226482 161648
rect 226538 161592 226543 161648
rect 223796 161590 226543 161592
rect 182317 161587 182383 161590
rect 226477 161587 226543 161590
rect 80197 161378 80263 161381
rect 76780 161376 80263 161378
rect 76780 161320 80202 161376
rect 80258 161320 80263 161376
rect 76780 161318 80263 161320
rect 80197 161315 80263 161318
rect 87189 161242 87255 161245
rect 132545 161242 132611 161245
rect 87189 161240 90028 161242
rect 87189 161184 87194 161240
rect 87250 161184 90028 161240
rect 87189 161182 90028 161184
rect 129772 161240 132611 161242
rect 129772 161184 132550 161240
rect 132606 161184 132611 161240
rect 129772 161182 132611 161184
rect 87189 161179 87255 161182
rect 132545 161179 132611 161182
rect 139813 161106 139879 161109
rect 142990 161106 143050 161416
rect 174037 161242 174103 161245
rect 170804 161240 174103 161242
rect 170804 161184 174042 161240
rect 174098 161184 174103 161240
rect 170804 161182 174103 161184
rect 174037 161179 174103 161182
rect 181397 161242 181463 161245
rect 226477 161242 226543 161245
rect 181397 161240 184052 161242
rect 181397 161184 181402 161240
rect 181458 161184 184052 161240
rect 181397 161182 184052 161184
rect 223796 161240 226543 161242
rect 223796 161184 226482 161240
rect 226538 161184 226543 161240
rect 223796 161182 226543 161184
rect 181397 161179 181463 161182
rect 226477 161179 226543 161182
rect 233469 161242 233535 161245
rect 233469 161240 237044 161242
rect 233469 161184 233474 161240
rect 233530 161184 237044 161240
rect 233469 161182 237044 161184
rect 233469 161179 233535 161182
rect 139813 161104 143050 161106
rect 139813 161048 139818 161104
rect 139874 161048 143050 161104
rect 139813 161046 143050 161048
rect 139813 161043 139879 161046
rect 80105 160834 80171 160837
rect 76780 160832 80171 160834
rect 76780 160776 80110 160832
rect 80166 160776 80171 160832
rect 76780 160774 80171 160776
rect 80105 160771 80171 160774
rect 87373 160834 87439 160837
rect 133373 160834 133439 160837
rect 87373 160832 90028 160834
rect 87373 160776 87378 160832
rect 87434 160776 90028 160832
rect 87373 160774 90028 160776
rect 129772 160832 133439 160834
rect 129772 160776 133378 160832
rect 133434 160776 133439 160832
rect 129772 160774 133439 160776
rect 87373 160771 87439 160774
rect 133373 160771 133439 160774
rect 140457 160834 140523 160837
rect 182133 160834 182199 160837
rect 225925 160834 225991 160837
rect 140457 160832 143020 160834
rect 140457 160776 140462 160832
rect 140518 160776 143020 160832
rect 140457 160774 143020 160776
rect 182133 160832 184052 160834
rect 182133 160776 182138 160832
rect 182194 160776 184052 160832
rect 182133 160774 184052 160776
rect 223796 160832 225991 160834
rect 223796 160776 225930 160832
rect 225986 160776 225991 160832
rect 223796 160774 225991 160776
rect 140457 160771 140523 160774
rect 182133 160771 182199 160774
rect 225925 160771 225991 160774
rect 132453 160562 132519 160565
rect 172749 160562 172815 160565
rect 226477 160562 226543 160565
rect 129772 160560 132519 160562
rect 129772 160504 132458 160560
rect 132514 160504 132519 160560
rect 129772 160502 132519 160504
rect 170804 160560 172815 160562
rect 170804 160504 172754 160560
rect 172810 160504 172815 160560
rect 170804 160502 172815 160504
rect 223796 160560 226543 160562
rect 223796 160504 226482 160560
rect 226538 160504 226543 160560
rect 223796 160502 226543 160504
rect 132453 160499 132519 160502
rect 172749 160499 172815 160502
rect 226477 160499 226543 160502
rect 233561 160562 233627 160565
rect 233561 160560 237044 160562
rect 233561 160504 233566 160560
rect 233622 160504 237044 160560
rect 233561 160502 237044 160504
rect 233561 160499 233627 160502
rect 87281 160426 87347 160429
rect 181397 160426 181463 160429
rect 87281 160424 90028 160426
rect 87281 160368 87286 160424
rect 87342 160368 90028 160424
rect 87281 160366 90028 160368
rect 181397 160424 184052 160426
rect 181397 160368 181402 160424
rect 181458 160368 184052 160424
rect 181397 160366 184052 160368
rect 87281 160363 87347 160366
rect 181397 160363 181463 160366
rect 80197 160290 80263 160293
rect 76780 160288 80263 160290
rect 76780 160232 80202 160288
rect 80258 160232 80263 160288
rect 76780 160230 80263 160232
rect 80197 160227 80263 160230
rect 132637 160154 132703 160157
rect 225557 160154 225623 160157
rect 129772 160152 132703 160154
rect 129772 160096 132642 160152
rect 132698 160096 132703 160152
rect 129772 160094 132703 160096
rect 223796 160152 225623 160154
rect 223796 160096 225562 160152
rect 225618 160096 225623 160152
rect 223796 160094 225623 160096
rect 132637 160091 132703 160094
rect 225557 160091 225623 160094
rect 87189 160018 87255 160021
rect 87189 160016 90028 160018
rect 87189 159960 87194 160016
rect 87250 159960 90028 160016
rect 87189 159958 90028 159960
rect 87189 159955 87255 159958
rect 132545 159746 132611 159749
rect 129772 159744 132611 159746
rect 129772 159688 132550 159744
rect 132606 159688 132611 159744
rect 129772 159686 132611 159688
rect 132545 159683 132611 159686
rect 139353 159746 139419 159749
rect 142990 159746 143050 160056
rect 173301 160018 173367 160021
rect 170804 160016 173367 160018
rect 170804 159960 173306 160016
rect 173362 159960 173367 160016
rect 170804 159958 173367 159960
rect 173301 159955 173367 159958
rect 181305 160018 181371 160021
rect 233469 160018 233535 160021
rect 181305 160016 184052 160018
rect 181305 159960 181310 160016
rect 181366 159960 184052 160016
rect 181305 159958 184052 159960
rect 233469 160016 237044 160018
rect 233469 159960 233474 160016
rect 233530 159960 237044 160016
rect 233469 159958 237044 159960
rect 181305 159955 181371 159958
rect 233469 159955 233535 159958
rect 225925 159746 225991 159749
rect 139353 159744 143050 159746
rect 139353 159688 139358 159744
rect 139414 159688 143050 159744
rect 139353 159686 143050 159688
rect 223796 159744 225991 159746
rect 223796 159688 225930 159744
rect 225986 159688 225991 159744
rect 223796 159686 225991 159688
rect 139353 159683 139419 159686
rect 225925 159683 225991 159686
rect 80105 159610 80171 159613
rect 76780 159608 80171 159610
rect 76780 159552 80110 159608
rect 80166 159552 80171 159608
rect 76780 159550 80171 159552
rect 80105 159547 80171 159550
rect 87189 159610 87255 159613
rect 181029 159610 181095 159613
rect 87189 159608 90028 159610
rect 87189 159552 87194 159608
rect 87250 159552 90028 159608
rect 87189 159550 90028 159552
rect 181029 159608 184052 159610
rect 181029 159552 181034 159608
rect 181090 159552 184052 159608
rect 181029 159550 184052 159552
rect 87189 159547 87255 159550
rect 181029 159547 181095 159550
rect 139445 159474 139511 159477
rect 174037 159474 174103 159477
rect 139445 159472 143020 159474
rect 139445 159416 139450 159472
rect 139506 159416 143020 159472
rect 139445 159414 143020 159416
rect 170804 159472 174103 159474
rect 170804 159416 174042 159472
rect 174098 159416 174103 159472
rect 170804 159414 174103 159416
rect 139445 159411 139511 159414
rect 174037 159411 174103 159414
rect 132637 159338 132703 159341
rect 226477 159338 226543 159341
rect 129772 159336 132703 159338
rect 129772 159280 132642 159336
rect 132698 159280 132703 159336
rect 129772 159278 132703 159280
rect 223796 159336 226543 159338
rect 223796 159280 226482 159336
rect 226538 159280 226543 159336
rect 223796 159278 226543 159280
rect 132637 159275 132703 159278
rect 226477 159275 226543 159278
rect 233561 159338 233627 159341
rect 233561 159336 237044 159338
rect 233561 159280 233566 159336
rect 233622 159280 237044 159336
rect 233561 159278 237044 159280
rect 233561 159275 233627 159278
rect 87281 159202 87347 159205
rect 181489 159202 181555 159205
rect 87281 159200 90028 159202
rect 87281 159144 87286 159200
rect 87342 159144 90028 159200
rect 87281 159142 90028 159144
rect 181489 159200 184052 159202
rect 181489 159144 181494 159200
rect 181550 159144 184052 159200
rect 181489 159142 184052 159144
rect 87281 159139 87347 159142
rect 181489 159139 181555 159142
rect 80197 159066 80263 159069
rect 76780 159064 80263 159066
rect 76780 159008 80202 159064
rect 80258 159008 80263 159064
rect 76780 159006 80263 159008
rect 80197 159003 80263 159006
rect 132545 158930 132611 158933
rect 173117 158930 173183 158933
rect 226477 158930 226543 158933
rect 129772 158928 132611 158930
rect 129772 158872 132550 158928
rect 132606 158872 132611 158928
rect 129772 158870 132611 158872
rect 170804 158928 173183 158930
rect 170804 158872 173122 158928
rect 173178 158872 173183 158928
rect 170804 158870 173183 158872
rect 223796 158928 226543 158930
rect 223796 158872 226482 158928
rect 226538 158872 226543 158928
rect 223796 158870 226543 158872
rect 132545 158867 132611 158870
rect 173117 158867 173183 158870
rect 226477 158867 226543 158870
rect 87373 158794 87439 158797
rect 182133 158794 182199 158797
rect 87373 158792 90028 158794
rect 87373 158736 87378 158792
rect 87434 158736 90028 158792
rect 87373 158734 90028 158736
rect 182133 158792 184052 158794
rect 182133 158736 182138 158792
rect 182194 158736 184052 158792
rect 182133 158734 184052 158736
rect 87373 158731 87439 158734
rect 182133 158731 182199 158734
rect 80197 158522 80263 158525
rect 132453 158522 132519 158525
rect 76780 158520 80263 158522
rect 76780 158464 80202 158520
rect 80258 158464 80263 158520
rect 76780 158462 80263 158464
rect 129772 158520 132519 158522
rect 129772 158464 132458 158520
rect 132514 158464 132519 158520
rect 129772 158462 132519 158464
rect 80197 158459 80263 158462
rect 132453 158459 132519 158462
rect 87281 158386 87347 158389
rect 140365 158386 140431 158389
rect 142990 158386 143050 158696
rect 233469 158658 233535 158661
rect 233469 158656 237044 158658
rect 233469 158600 233474 158656
rect 233530 158600 237044 158656
rect 233469 158598 237044 158600
rect 233469 158595 233535 158598
rect 225557 158522 225623 158525
rect 223796 158520 225623 158522
rect 223796 158464 225562 158520
rect 225618 158464 225623 158520
rect 223796 158462 225623 158464
rect 225557 158459 225623 158462
rect 173301 158386 173367 158389
rect 87281 158384 90028 158386
rect 87281 158328 87286 158384
rect 87342 158328 90028 158384
rect 87281 158326 90028 158328
rect 140365 158384 143050 158386
rect 140365 158328 140370 158384
rect 140426 158328 143050 158384
rect 140365 158326 143050 158328
rect 170804 158384 173367 158386
rect 170804 158328 173306 158384
rect 173362 158328 173367 158384
rect 170804 158326 173367 158328
rect 87281 158323 87347 158326
rect 140365 158323 140431 158326
rect 173301 158323 173367 158326
rect 182317 158386 182383 158389
rect 182317 158384 184052 158386
rect 182317 158328 182322 158384
rect 182378 158328 184052 158384
rect 182317 158326 184052 158328
rect 182317 158323 182383 158326
rect 132637 158114 132703 158117
rect 129772 158112 132703 158114
rect 129772 158056 132642 158112
rect 132698 158056 132703 158112
rect 129772 158054 132703 158056
rect 132637 158051 132703 158054
rect 139169 158114 139235 158117
rect 226385 158114 226451 158117
rect 139169 158112 143020 158114
rect 139169 158056 139174 158112
rect 139230 158056 143020 158112
rect 139169 158054 143020 158056
rect 223796 158112 226451 158114
rect 223796 158056 226390 158112
rect 226446 158056 226451 158112
rect 223796 158054 226451 158056
rect 139169 158051 139235 158054
rect 226385 158051 226451 158054
rect 233469 158114 233535 158117
rect 233469 158112 237044 158114
rect 233469 158056 233474 158112
rect 233530 158056 237044 158112
rect 233469 158054 237044 158056
rect 233469 158051 233535 158054
rect 87189 157978 87255 157981
rect 180753 157978 180819 157981
rect 87189 157976 90028 157978
rect 87189 157920 87194 157976
rect 87250 157920 90028 157976
rect 87189 157918 90028 157920
rect 180753 157976 184052 157978
rect 180753 157920 180758 157976
rect 180814 157920 184052 157976
rect 180753 157918 184052 157920
rect 87189 157915 87255 157918
rect 180753 157915 180819 157918
rect 79461 157842 79527 157845
rect 172933 157842 172999 157845
rect 76780 157840 79527 157842
rect 76780 157784 79466 157840
rect 79522 157784 79527 157840
rect 76780 157782 79527 157784
rect 170804 157840 172999 157842
rect 170804 157784 172938 157840
rect 172994 157784 172999 157840
rect 170804 157782 172999 157784
rect 79461 157779 79527 157782
rect 172933 157779 172999 157782
rect 132545 157706 132611 157709
rect 226293 157706 226359 157709
rect 129772 157704 132611 157706
rect 129772 157648 132550 157704
rect 132606 157648 132611 157704
rect 129772 157646 132611 157648
rect 223796 157704 226359 157706
rect 223796 157648 226298 157704
rect 226354 157648 226359 157704
rect 223796 157646 226359 157648
rect 132545 157643 132611 157646
rect 226293 157643 226359 157646
rect 87281 157570 87347 157573
rect 180937 157570 181003 157573
rect 87281 157568 90028 157570
rect 87281 157512 87286 157568
rect 87342 157512 90028 157568
rect 87281 157510 90028 157512
rect 180937 157568 184052 157570
rect 180937 157512 180942 157568
rect 180998 157512 184052 157568
rect 180937 157510 184052 157512
rect 87281 157507 87347 157510
rect 180937 157507 181003 157510
rect 132637 157434 132703 157437
rect 226477 157434 226543 157437
rect 129772 157432 132703 157434
rect 129772 157376 132642 157432
rect 132698 157376 132703 157432
rect 129772 157374 132703 157376
rect 223796 157432 226543 157434
rect 223796 157376 226482 157432
rect 226538 157376 226543 157432
rect 223796 157374 226543 157376
rect 132637 157371 132703 157374
rect 226477 157371 226543 157374
rect 233469 157434 233535 157437
rect 233469 157432 237044 157434
rect 233469 157376 233474 157432
rect 233530 157376 237044 157432
rect 233469 157374 237044 157376
rect 233469 157371 233535 157374
rect 80197 157298 80263 157301
rect 76780 157296 80263 157298
rect 76780 157240 80202 157296
rect 80258 157240 80263 157296
rect 76780 157238 80263 157240
rect 80197 157235 80263 157238
rect 87189 157162 87255 157165
rect 87189 157160 90028 157162
rect 87189 157104 87194 157160
rect 87250 157104 90028 157160
rect 87189 157102 90028 157104
rect 87189 157099 87255 157102
rect 132545 157026 132611 157029
rect 129772 157024 132611 157026
rect 129772 156968 132550 157024
rect 132606 156968 132611 157024
rect 129772 156966 132611 156968
rect 132545 156963 132611 156966
rect 140181 157026 140247 157029
rect 142990 157026 143050 157336
rect 173209 157298 173275 157301
rect 170804 157296 173275 157298
rect 170804 157240 173214 157296
rect 173270 157240 173275 157296
rect 170804 157238 173275 157240
rect 173209 157235 173275 157238
rect 182041 157162 182107 157165
rect 182041 157160 184052 157162
rect 182041 157104 182046 157160
rect 182102 157104 184052 157160
rect 182041 157102 184052 157104
rect 182041 157099 182107 157102
rect 226477 157026 226543 157029
rect 140181 157024 143050 157026
rect 140181 156968 140186 157024
rect 140242 156968 143050 157024
rect 140181 156966 143050 156968
rect 223796 157024 226543 157026
rect 223796 156968 226482 157024
rect 226538 156968 226543 157024
rect 223796 156966 226543 156968
rect 140181 156963 140247 156966
rect 226477 156963 226543 156966
rect 80105 156754 80171 156757
rect 76780 156752 80171 156754
rect 76780 156696 80110 156752
rect 80166 156696 80171 156752
rect 76780 156694 80171 156696
rect 80105 156691 80171 156694
rect 87097 156754 87163 156757
rect 139537 156754 139603 156757
rect 173117 156754 173183 156757
rect 87097 156752 90028 156754
rect 87097 156696 87102 156752
rect 87158 156696 90028 156752
rect 87097 156694 90028 156696
rect 139537 156752 143020 156754
rect 139537 156696 139542 156752
rect 139598 156696 143020 156752
rect 139537 156694 143020 156696
rect 170804 156752 173183 156754
rect 170804 156696 173122 156752
rect 173178 156696 173183 156752
rect 170804 156694 173183 156696
rect 87097 156691 87163 156694
rect 139537 156691 139603 156694
rect 173117 156691 173183 156694
rect 180569 156754 180635 156757
rect 233469 156754 233535 156757
rect 180569 156752 184052 156754
rect 180569 156696 180574 156752
rect 180630 156696 184052 156752
rect 180569 156694 184052 156696
rect 233469 156752 237044 156754
rect 233469 156696 233474 156752
rect 233530 156696 237044 156752
rect 233469 156694 237044 156696
rect 180569 156691 180635 156694
rect 233469 156691 233535 156694
rect 132637 156618 132703 156621
rect 225373 156618 225439 156621
rect 129772 156616 132703 156618
rect 129772 156560 132642 156616
rect 132698 156560 132703 156616
rect 129772 156558 132703 156560
rect 223796 156616 225439 156618
rect 223796 156560 225378 156616
rect 225434 156560 225439 156616
rect 223796 156558 225439 156560
rect 132637 156555 132703 156558
rect 225373 156555 225439 156558
rect 87373 156346 87439 156349
rect 180845 156346 180911 156349
rect 87373 156344 90028 156346
rect 87373 156288 87378 156344
rect 87434 156288 90028 156344
rect 87373 156286 90028 156288
rect 180845 156344 184052 156346
rect 180845 156288 180850 156344
rect 180906 156288 184052 156344
rect 180845 156286 184052 156288
rect 87373 156283 87439 156286
rect 180845 156283 180911 156286
rect 80197 156210 80263 156213
rect 131809 156210 131875 156213
rect 174037 156210 174103 156213
rect 226477 156210 226543 156213
rect 76780 156208 80263 156210
rect 76780 156152 80202 156208
rect 80258 156152 80263 156208
rect 76780 156150 80263 156152
rect 129772 156208 131875 156210
rect 129772 156152 131814 156208
rect 131870 156152 131875 156208
rect 129772 156150 131875 156152
rect 170804 156208 174103 156210
rect 170804 156152 174042 156208
rect 174098 156152 174103 156208
rect 170804 156150 174103 156152
rect 223796 156208 226543 156210
rect 223796 156152 226482 156208
rect 226538 156152 226543 156208
rect 223796 156150 226543 156152
rect 80197 156147 80263 156150
rect 131809 156147 131875 156150
rect 174037 156147 174103 156150
rect 226477 156147 226543 156150
rect 233469 156210 233535 156213
rect 233469 156208 237044 156210
rect 233469 156152 233474 156208
rect 233530 156152 237044 156208
rect 233469 156150 237044 156152
rect 233469 156147 233535 156150
rect 87189 156074 87255 156077
rect 87189 156072 90028 156074
rect 87189 156016 87194 156072
rect 87250 156016 90028 156072
rect 87189 156014 90028 156016
rect 87189 156011 87255 156014
rect 9896 155802 10376 155832
rect 13589 155802 13655 155805
rect 132269 155802 132335 155805
rect 9896 155800 13655 155802
rect 9896 155744 13594 155800
rect 13650 155744 13655 155800
rect 9896 155742 13655 155744
rect 129772 155800 132335 155802
rect 129772 155744 132274 155800
rect 132330 155744 132335 155800
rect 129772 155742 132335 155744
rect 9896 155712 10376 155742
rect 13589 155739 13655 155742
rect 132269 155739 132335 155742
rect 139813 155802 139879 155805
rect 142990 155802 143050 156112
rect 181949 156074 182015 156077
rect 181949 156072 184052 156074
rect 181949 156016 181954 156072
rect 182010 156016 184052 156072
rect 181949 156014 184052 156016
rect 181949 156011 182015 156014
rect 226477 155802 226543 155805
rect 139813 155800 143050 155802
rect 139813 155744 139818 155800
rect 139874 155744 143050 155800
rect 139813 155742 143050 155744
rect 223796 155800 226543 155802
rect 223796 155744 226482 155800
rect 226538 155744 226543 155800
rect 223796 155742 226543 155744
rect 139813 155739 139879 155742
rect 226477 155739 226543 155742
rect 87005 155666 87071 155669
rect 180293 155666 180359 155669
rect 87005 155664 90028 155666
rect 87005 155608 87010 155664
rect 87066 155608 90028 155664
rect 87005 155606 90028 155608
rect 180293 155664 184052 155666
rect 180293 155608 180298 155664
rect 180354 155608 184052 155664
rect 180293 155606 184052 155608
rect 87005 155603 87071 155606
rect 180293 155603 180359 155606
rect 80105 155530 80171 155533
rect 173945 155530 174011 155533
rect 76780 155528 80171 155530
rect 76780 155472 80110 155528
rect 80166 155472 80171 155528
rect 76780 155470 80171 155472
rect 170804 155528 174011 155530
rect 170804 155472 173950 155528
rect 174006 155472 174011 155528
rect 170804 155470 174011 155472
rect 80105 155467 80171 155470
rect 173945 155467 174011 155470
rect 233469 155530 233535 155533
rect 233469 155528 237044 155530
rect 233469 155472 233474 155528
rect 233530 155472 237044 155528
rect 233469 155470 237044 155472
rect 233469 155467 233535 155470
rect 131533 155394 131599 155397
rect 129772 155392 131599 155394
rect 129772 155336 131538 155392
rect 131594 155336 131599 155392
rect 129772 155334 131599 155336
rect 131533 155331 131599 155334
rect 86913 155258 86979 155261
rect 139721 155258 139787 155261
rect 142990 155258 143050 155432
rect 225557 155394 225623 155397
rect 223796 155392 225623 155394
rect 223796 155336 225562 155392
rect 225618 155336 225623 155392
rect 223796 155334 225623 155336
rect 225557 155331 225623 155334
rect 86913 155256 90028 155258
rect 86913 155200 86918 155256
rect 86974 155200 90028 155256
rect 86913 155198 90028 155200
rect 139721 155256 143050 155258
rect 139721 155200 139726 155256
rect 139782 155200 143050 155256
rect 139721 155198 143050 155200
rect 181029 155258 181095 155261
rect 181029 155256 184052 155258
rect 181029 155200 181034 155256
rect 181090 155200 184052 155256
rect 181029 155198 184052 155200
rect 86913 155195 86979 155198
rect 139721 155195 139787 155198
rect 181029 155195 181095 155198
rect 80197 154986 80263 154989
rect 131349 154986 131415 154989
rect 173945 154986 174011 154989
rect 225741 154986 225807 154989
rect 76780 154984 80263 154986
rect 76780 154928 80202 154984
rect 80258 154928 80263 154984
rect 76780 154926 80263 154928
rect 129772 154984 131415 154986
rect 129772 154928 131354 154984
rect 131410 154928 131415 154984
rect 129772 154926 131415 154928
rect 170804 154984 174011 154986
rect 170804 154928 173950 154984
rect 174006 154928 174011 154984
rect 170804 154926 174011 154928
rect 223796 154984 225807 154986
rect 223796 154928 225746 154984
rect 225802 154928 225807 154984
rect 223796 154926 225807 154928
rect 80197 154923 80263 154926
rect 131349 154923 131415 154926
rect 173945 154923 174011 154926
rect 225741 154923 225807 154926
rect 86821 154850 86887 154853
rect 139629 154850 139695 154853
rect 181029 154850 181095 154853
rect 233561 154850 233627 154853
rect 86821 154848 90028 154850
rect 86821 154792 86826 154848
rect 86882 154792 90028 154848
rect 86821 154790 90028 154792
rect 139629 154848 143020 154850
rect 139629 154792 139634 154848
rect 139690 154792 143020 154848
rect 139629 154790 143020 154792
rect 181029 154848 184052 154850
rect 181029 154792 181034 154848
rect 181090 154792 184052 154848
rect 181029 154790 184052 154792
rect 233561 154848 237044 154850
rect 233561 154792 233566 154848
rect 233622 154792 237044 154848
rect 233561 154790 237044 154792
rect 86821 154787 86887 154790
rect 139629 154787 139695 154790
rect 181029 154787 181095 154790
rect 233561 154787 233627 154790
rect 132085 154578 132151 154581
rect 226109 154578 226175 154581
rect 129772 154576 132151 154578
rect 129772 154520 132090 154576
rect 132146 154520 132151 154576
rect 129772 154518 132151 154520
rect 223796 154576 226175 154578
rect 223796 154520 226114 154576
rect 226170 154520 226175 154576
rect 223796 154518 226175 154520
rect 132085 154515 132151 154518
rect 226109 154515 226175 154518
rect 80105 154442 80171 154445
rect 76780 154440 80171 154442
rect 76780 154384 80110 154440
rect 80166 154384 80171 154440
rect 76780 154382 80171 154384
rect 80105 154379 80171 154382
rect 87097 154442 87163 154445
rect 173117 154442 173183 154445
rect 87097 154440 90028 154442
rect 87097 154384 87102 154440
rect 87158 154384 90028 154440
rect 87097 154382 90028 154384
rect 170804 154440 173183 154442
rect 170804 154384 173122 154440
rect 173178 154384 173183 154440
rect 170804 154382 173183 154384
rect 87097 154379 87163 154382
rect 173117 154379 173183 154382
rect 181213 154442 181279 154445
rect 181213 154440 184052 154442
rect 181213 154384 181218 154440
rect 181274 154384 184052 154440
rect 181213 154382 184052 154384
rect 181213 154379 181279 154382
rect 131441 154306 131507 154309
rect 225833 154306 225899 154309
rect 129772 154304 131507 154306
rect 129772 154248 131446 154304
rect 131502 154248 131507 154304
rect 129772 154246 131507 154248
rect 223796 154304 225899 154306
rect 223796 154248 225838 154304
rect 225894 154248 225899 154304
rect 223796 154246 225899 154248
rect 131441 154243 131507 154246
rect 225833 154243 225899 154246
rect 139721 154170 139787 154173
rect 233469 154170 233535 154173
rect 139721 154168 143020 154170
rect 139721 154112 139726 154168
rect 139782 154112 143020 154168
rect 139721 154110 143020 154112
rect 233469 154168 237044 154170
rect 233469 154112 233474 154168
rect 233530 154112 237044 154168
rect 233469 154110 237044 154112
rect 139721 154107 139787 154110
rect 233469 154107 233535 154110
rect 87189 154034 87255 154037
rect 181121 154034 181187 154037
rect 87189 154032 90028 154034
rect 87189 153976 87194 154032
rect 87250 153976 90028 154032
rect 87189 153974 90028 153976
rect 181121 154032 184052 154034
rect 181121 153976 181126 154032
rect 181182 153976 184052 154032
rect 181121 153974 184052 153976
rect 87189 153971 87255 153974
rect 181121 153971 181187 153974
rect 131349 153898 131415 153901
rect 172933 153898 172999 153901
rect 226477 153898 226543 153901
rect 129772 153896 131415 153898
rect 129772 153840 131354 153896
rect 131410 153840 131415 153896
rect 129772 153838 131415 153840
rect 170804 153896 172999 153898
rect 170804 153840 172938 153896
rect 172994 153840 172999 153896
rect 170804 153838 172999 153840
rect 223796 153896 226543 153898
rect 223796 153840 226482 153896
rect 226538 153840 226543 153896
rect 223796 153838 226543 153840
rect 131349 153835 131415 153838
rect 172933 153835 172999 153838
rect 226477 153835 226543 153838
rect 80013 153762 80079 153765
rect 76780 153760 80079 153762
rect 76780 153704 80018 153760
rect 80074 153704 80079 153760
rect 76780 153702 80079 153704
rect 80013 153699 80079 153702
rect 228409 153762 228475 153765
rect 228685 153762 228751 153765
rect 228409 153760 228751 153762
rect 228409 153704 228414 153760
rect 228470 153704 228690 153760
rect 228746 153704 228751 153760
rect 228409 153702 228751 153704
rect 228409 153699 228475 153702
rect 228685 153699 228751 153702
rect 87925 153626 87991 153629
rect 181673 153626 181739 153629
rect 233561 153626 233627 153629
rect 87925 153624 90028 153626
rect 87925 153568 87930 153624
rect 87986 153568 90028 153624
rect 87925 153566 90028 153568
rect 181673 153624 184052 153626
rect 181673 153568 181678 153624
rect 181734 153568 184052 153624
rect 181673 153566 184052 153568
rect 233561 153624 237044 153626
rect 233561 153568 233566 153624
rect 233622 153568 237044 153624
rect 233561 153566 237044 153568
rect 87925 153563 87991 153566
rect 181673 153563 181739 153566
rect 233561 153563 233627 153566
rect 132177 153490 132243 153493
rect 129772 153488 132243 153490
rect 129772 153432 132182 153488
rect 132238 153432 132243 153488
rect 129772 153430 132243 153432
rect 132177 153427 132243 153430
rect 140089 153490 140155 153493
rect 226109 153490 226175 153493
rect 140089 153488 143020 153490
rect 140089 153432 140094 153488
rect 140150 153432 143020 153488
rect 140089 153430 143020 153432
rect 223796 153488 226175 153490
rect 223796 153432 226114 153488
rect 226170 153432 226175 153488
rect 223796 153430 226175 153432
rect 140089 153427 140155 153430
rect 226109 153427 226175 153430
rect 174037 153354 174103 153357
rect 170804 153352 174103 153354
rect 170804 153296 174042 153352
rect 174098 153296 174103 153352
rect 170804 153294 174103 153296
rect 174037 153291 174103 153294
rect 80197 153218 80263 153221
rect 76780 153216 80263 153218
rect 76780 153160 80202 153216
rect 80258 153160 80263 153216
rect 76780 153158 80263 153160
rect 80197 153155 80263 153158
rect 87557 153218 87623 153221
rect 181029 153218 181095 153221
rect 87557 153216 90028 153218
rect 87557 153160 87562 153216
rect 87618 153160 90028 153216
rect 87557 153158 90028 153160
rect 181029 153216 184052 153218
rect 181029 153160 181034 153216
rect 181090 153160 184052 153216
rect 181029 153158 184052 153160
rect 87557 153155 87623 153158
rect 181029 153155 181095 153158
rect 132545 153082 132611 153085
rect 225741 153082 225807 153085
rect 129772 153080 132611 153082
rect 129772 153024 132550 153080
rect 132606 153024 132611 153080
rect 129772 153022 132611 153024
rect 223796 153080 225807 153082
rect 223796 153024 225746 153080
rect 225802 153024 225807 153080
rect 223796 153022 225807 153024
rect 132545 153019 132611 153022
rect 225741 153019 225807 153022
rect 233469 152946 233535 152949
rect 233469 152944 237044 152946
rect 233469 152888 233474 152944
rect 233530 152888 237044 152944
rect 233469 152886 237044 152888
rect 233469 152883 233535 152886
rect 87741 152810 87807 152813
rect 139905 152810 139971 152813
rect 173301 152810 173367 152813
rect 87741 152808 90028 152810
rect 87741 152752 87746 152808
rect 87802 152752 90028 152808
rect 87741 152750 90028 152752
rect 139905 152808 143020 152810
rect 139905 152752 139910 152808
rect 139966 152752 143020 152808
rect 139905 152750 143020 152752
rect 170804 152808 173367 152810
rect 170804 152752 173306 152808
rect 173362 152752 173367 152808
rect 170804 152750 173367 152752
rect 87741 152747 87807 152750
rect 139905 152747 139971 152750
rect 173301 152747 173367 152750
rect 181213 152810 181279 152813
rect 181213 152808 184052 152810
rect 181213 152752 181218 152808
rect 181274 152752 184052 152808
rect 181213 152750 184052 152752
rect 181213 152747 181279 152750
rect 80197 152674 80263 152677
rect 132453 152674 132519 152677
rect 225373 152674 225439 152677
rect 76780 152672 80263 152674
rect 76780 152616 80202 152672
rect 80258 152616 80263 152672
rect 76780 152614 80263 152616
rect 129772 152672 132519 152674
rect 129772 152616 132458 152672
rect 132514 152616 132519 152672
rect 129772 152614 132519 152616
rect 223796 152672 225439 152674
rect 223796 152616 225378 152672
rect 225434 152616 225439 152672
rect 223796 152614 225439 152616
rect 80197 152611 80263 152614
rect 132453 152611 132519 152614
rect 225373 152611 225439 152614
rect 88109 152402 88175 152405
rect 181121 152402 181187 152405
rect 88109 152400 90028 152402
rect 88109 152344 88114 152400
rect 88170 152344 90028 152400
rect 88109 152342 90028 152344
rect 181121 152400 184052 152402
rect 181121 152344 181126 152400
rect 181182 152344 184052 152400
rect 181121 152342 184052 152344
rect 88109 152339 88175 152342
rect 181121 152339 181187 152342
rect 131349 152266 131415 152269
rect 174037 152266 174103 152269
rect 225925 152266 225991 152269
rect 129772 152264 131415 152266
rect 129772 152208 131354 152264
rect 131410 152208 131415 152264
rect 129772 152206 131415 152208
rect 170804 152264 174103 152266
rect 170804 152208 174042 152264
rect 174098 152208 174103 152264
rect 170804 152206 174103 152208
rect 223796 152264 225991 152266
rect 223796 152208 225930 152264
rect 225986 152208 225991 152264
rect 223796 152206 225991 152208
rect 131349 152203 131415 152206
rect 174037 152203 174103 152206
rect 225925 152203 225991 152206
rect 233653 152266 233719 152269
rect 233653 152264 237044 152266
rect 233653 152208 233658 152264
rect 233714 152208 237044 152264
rect 233653 152206 237044 152208
rect 233653 152203 233719 152206
rect 139997 152130 140063 152133
rect 139997 152128 143020 152130
rect 139997 152072 140002 152128
rect 140058 152072 143020 152128
rect 139997 152070 143020 152072
rect 139997 152067 140063 152070
rect 87373 151994 87439 151997
rect 181765 151994 181831 151997
rect 87373 151992 90028 151994
rect 87373 151936 87378 151992
rect 87434 151936 90028 151992
rect 87373 151934 90028 151936
rect 181765 151992 184052 151994
rect 181765 151936 181770 151992
rect 181826 151936 184052 151992
rect 181765 151934 184052 151936
rect 87373 151931 87439 151934
rect 181765 151931 181831 151934
rect 76750 151722 76810 151896
rect 131349 151858 131415 151861
rect 226109 151858 226175 151861
rect 129772 151856 131415 151858
rect 129772 151800 131354 151856
rect 131410 151800 131415 151856
rect 129772 151798 131415 151800
rect 223796 151856 226175 151858
rect 223796 151800 226114 151856
rect 226170 151800 226175 151856
rect 223796 151798 226175 151800
rect 131349 151795 131415 151798
rect 226109 151795 226175 151798
rect 80197 151722 80263 151725
rect 173301 151722 173367 151725
rect 76750 151720 80263 151722
rect 76750 151664 80202 151720
rect 80258 151664 80263 151720
rect 76750 151662 80263 151664
rect 170804 151720 173367 151722
rect 170804 151664 173306 151720
rect 173362 151664 173367 151720
rect 170804 151662 173367 151664
rect 80197 151659 80263 151662
rect 173301 151659 173367 151662
rect 233745 151722 233811 151725
rect 233745 151720 237044 151722
rect 233745 151664 233750 151720
rect 233806 151664 237044 151720
rect 233745 151662 237044 151664
rect 233745 151659 233811 151662
rect 87281 151586 87347 151589
rect 181029 151586 181095 151589
rect 87281 151584 90028 151586
rect 87281 151528 87286 151584
rect 87342 151528 90028 151584
rect 87281 151526 90028 151528
rect 181029 151584 184052 151586
rect 181029 151528 181034 151584
rect 181090 151528 184052 151584
rect 181029 151526 184052 151528
rect 87281 151523 87347 151526
rect 181029 151523 181095 151526
rect 80105 151450 80171 151453
rect 131441 151450 131507 151453
rect 76780 151448 80171 151450
rect 76780 151392 80110 151448
rect 80166 151392 80171 151448
rect 76780 151390 80171 151392
rect 129772 151448 131507 151450
rect 129772 151392 131446 151448
rect 131502 151392 131507 151448
rect 129772 151390 131507 151392
rect 80105 151387 80171 151390
rect 131441 151387 131507 151390
rect 140181 151450 140247 151453
rect 225373 151450 225439 151453
rect 140181 151448 143020 151450
rect 140181 151392 140186 151448
rect 140242 151392 143020 151448
rect 140181 151390 143020 151392
rect 223796 151448 225439 151450
rect 223796 151392 225378 151448
rect 225434 151392 225439 151448
rect 223796 151390 225439 151392
rect 140181 151387 140247 151390
rect 225373 151387 225439 151390
rect 87189 151178 87255 151181
rect 131533 151178 131599 151181
rect 87189 151176 90028 151178
rect 87189 151120 87194 151176
rect 87250 151120 90028 151176
rect 87189 151118 90028 151120
rect 129772 151176 131599 151178
rect 129772 151120 131538 151176
rect 131594 151120 131599 151176
rect 129772 151118 131599 151120
rect 87189 151115 87255 151118
rect 131533 151115 131599 151118
rect 181121 151178 181187 151181
rect 226477 151178 226543 151181
rect 181121 151176 184052 151178
rect 181121 151120 181126 151176
rect 181182 151120 184052 151176
rect 181121 151118 184052 151120
rect 223796 151176 226543 151178
rect 223796 151120 226482 151176
rect 226538 151120 226543 151176
rect 223796 151118 226543 151120
rect 181121 151115 181187 151118
rect 226477 151115 226543 151118
rect 173945 151042 174011 151045
rect 170804 151040 174011 151042
rect 170804 150984 173950 151040
rect 174006 150984 174011 151040
rect 170804 150982 174011 150984
rect 173945 150979 174011 150982
rect 233561 151042 233627 151045
rect 233561 151040 237044 151042
rect 233561 150984 233566 151040
rect 233622 150984 237044 151040
rect 233561 150982 237044 150984
rect 233561 150979 233627 150982
rect 80105 150906 80171 150909
rect 76780 150904 80171 150906
rect 76780 150848 80110 150904
rect 80166 150848 80171 150904
rect 76780 150846 80171 150848
rect 80105 150843 80171 150846
rect 87373 150770 87439 150773
rect 131349 150770 131415 150773
rect 87373 150768 90028 150770
rect 87373 150712 87378 150768
rect 87434 150712 90028 150768
rect 87373 150710 90028 150712
rect 129772 150768 131415 150770
rect 129772 150712 131354 150768
rect 131410 150712 131415 150768
rect 129772 150710 131415 150712
rect 87373 150707 87439 150710
rect 131349 150707 131415 150710
rect 139629 150770 139695 150773
rect 182041 150770 182107 150773
rect 225557 150770 225623 150773
rect 139629 150768 143020 150770
rect 139629 150712 139634 150768
rect 139690 150712 143020 150768
rect 139629 150710 143020 150712
rect 182041 150768 184052 150770
rect 182041 150712 182046 150768
rect 182102 150712 184052 150768
rect 182041 150710 184052 150712
rect 223796 150768 225623 150770
rect 223796 150712 225562 150768
rect 225618 150712 225623 150768
rect 223796 150710 225623 150712
rect 139629 150707 139695 150710
rect 182041 150707 182107 150710
rect 225557 150707 225623 150710
rect 174037 150498 174103 150501
rect 170804 150496 174103 150498
rect 170804 150440 174042 150496
rect 174098 150440 174103 150496
rect 170804 150438 174103 150440
rect 174037 150435 174103 150438
rect 80197 150362 80263 150365
rect 76780 150360 80263 150362
rect 76780 150304 80202 150360
rect 80258 150304 80263 150360
rect 76780 150302 80263 150304
rect 80197 150299 80263 150302
rect 87281 150362 87347 150365
rect 131441 150362 131507 150365
rect 87281 150360 90028 150362
rect 87281 150304 87286 150360
rect 87342 150304 90028 150360
rect 87281 150302 90028 150304
rect 129772 150360 131507 150362
rect 129772 150304 131446 150360
rect 131502 150304 131507 150360
rect 129772 150302 131507 150304
rect 87281 150299 87347 150302
rect 131441 150299 131507 150302
rect 181857 150362 181923 150365
rect 225741 150362 225807 150365
rect 181857 150360 184052 150362
rect 181857 150304 181862 150360
rect 181918 150304 184052 150360
rect 181857 150302 184052 150304
rect 223796 150360 225807 150362
rect 223796 150304 225746 150360
rect 225802 150304 225807 150360
rect 223796 150302 225807 150304
rect 181857 150299 181923 150302
rect 225741 150299 225807 150302
rect 233469 150362 233535 150365
rect 233469 150360 237044 150362
rect 233469 150304 233474 150360
rect 233530 150304 237044 150360
rect 233469 150302 237044 150304
rect 233469 150299 233535 150302
rect 139261 150090 139327 150093
rect 139261 150088 143020 150090
rect 139261 150032 139266 150088
rect 139322 150032 143020 150088
rect 139261 150030 143020 150032
rect 139261 150027 139327 150030
rect 87189 149954 87255 149957
rect 131349 149954 131415 149957
rect 172933 149954 172999 149957
rect 87189 149952 90028 149954
rect 87189 149896 87194 149952
rect 87250 149896 90028 149952
rect 87189 149894 90028 149896
rect 129772 149952 131415 149954
rect 129772 149896 131354 149952
rect 131410 149896 131415 149952
rect 129772 149894 131415 149896
rect 170804 149952 172999 149954
rect 170804 149896 172938 149952
rect 172994 149896 172999 149952
rect 170804 149894 172999 149896
rect 87189 149891 87255 149894
rect 131349 149891 131415 149894
rect 172933 149891 172999 149894
rect 180661 149954 180727 149957
rect 226477 149954 226543 149957
rect 180661 149952 184052 149954
rect 180661 149896 180666 149952
rect 180722 149896 184052 149952
rect 180661 149894 184052 149896
rect 223796 149952 226543 149954
rect 223796 149896 226482 149952
rect 226538 149896 226543 149952
rect 223796 149894 226543 149896
rect 180661 149891 180727 149894
rect 226477 149891 226543 149894
rect 233837 149818 233903 149821
rect 233837 149816 237044 149818
rect 233837 149760 233842 149816
rect 233898 149760 237044 149816
rect 233837 149758 237044 149760
rect 233837 149755 233903 149758
rect 80105 149682 80171 149685
rect 76780 149680 80171 149682
rect 76780 149624 80110 149680
rect 80166 149624 80171 149680
rect 76780 149622 80171 149624
rect 80105 149619 80171 149622
rect 87465 149546 87531 149549
rect 131441 149546 131507 149549
rect 87465 149544 90028 149546
rect 87465 149488 87470 149544
rect 87526 149488 90028 149544
rect 87465 149486 90028 149488
rect 129772 149544 131507 149546
rect 129772 149488 131446 149544
rect 131502 149488 131507 149544
rect 129772 149486 131507 149488
rect 87465 149483 87531 149486
rect 131441 149483 131507 149486
rect 180477 149546 180543 149549
rect 225557 149546 225623 149549
rect 180477 149544 184052 149546
rect 180477 149488 180482 149544
rect 180538 149488 184052 149544
rect 180477 149486 184052 149488
rect 223796 149544 225623 149546
rect 223796 149488 225562 149544
rect 225618 149488 225623 149544
rect 223796 149486 225623 149488
rect 180477 149483 180543 149486
rect 225557 149483 225623 149486
rect 140917 149410 140983 149413
rect 174037 149410 174103 149413
rect 140917 149408 143020 149410
rect 140917 149352 140922 149408
rect 140978 149352 143020 149408
rect 140917 149350 143020 149352
rect 170804 149408 174103 149410
rect 170804 149352 174042 149408
rect 174098 149352 174103 149408
rect 170804 149350 174103 149352
rect 140917 149347 140983 149350
rect 174037 149347 174103 149350
rect 264749 149410 264815 149413
rect 264749 149408 264858 149410
rect 264749 149352 264754 149408
rect 264810 149352 264858 149408
rect 264749 149347 264858 149352
rect 80197 149138 80263 149141
rect 76780 149136 80263 149138
rect 76780 149080 80202 149136
rect 80258 149080 80263 149136
rect 76780 149078 80263 149080
rect 80197 149075 80263 149078
rect 87557 149138 87623 149141
rect 131349 149138 131415 149141
rect 87557 149136 90028 149138
rect 87557 149080 87562 149136
rect 87618 149080 90028 149136
rect 87557 149078 90028 149080
rect 129772 149136 131415 149138
rect 129772 149080 131354 149136
rect 131410 149080 131415 149136
rect 129772 149078 131415 149080
rect 87557 149075 87623 149078
rect 131349 149075 131415 149078
rect 180385 149138 180451 149141
rect 225373 149138 225439 149141
rect 180385 149136 184052 149138
rect 180385 149080 180390 149136
rect 180446 149080 184052 149136
rect 180385 149078 184052 149080
rect 223796 149136 225439 149138
rect 223796 149080 225378 149136
rect 225434 149080 225439 149136
rect 223796 149078 225439 149080
rect 180385 149075 180451 149078
rect 225373 149075 225439 149078
rect 233469 149138 233535 149141
rect 233469 149136 237044 149138
rect 233469 149080 233474 149136
rect 233530 149080 237044 149136
rect 233469 149078 237044 149080
rect 233469 149075 233535 149078
rect 47077 148866 47143 148869
rect 140733 148866 140799 148869
rect 174037 148866 174103 148869
rect 47077 148864 48996 148866
rect 47077 148808 47082 148864
rect 47138 148808 48996 148864
rect 47077 148806 48996 148808
rect 140733 148864 143020 148866
rect 140733 148808 140738 148864
rect 140794 148808 143020 148864
rect 140733 148806 143020 148808
rect 170804 148864 174103 148866
rect 170804 148808 174042 148864
rect 174098 148808 174103 148864
rect 264798 148836 264858 149347
rect 170804 148806 174103 148808
rect 47077 148803 47143 148806
rect 140733 148803 140799 148806
rect 174037 148803 174103 148806
rect 87189 148730 87255 148733
rect 131625 148730 131691 148733
rect 87189 148728 90028 148730
rect 87189 148672 87194 148728
rect 87250 148672 90028 148728
rect 87189 148670 90028 148672
rect 129772 148728 131691 148730
rect 129772 148672 131630 148728
rect 131686 148672 131691 148728
rect 129772 148670 131691 148672
rect 87189 148667 87255 148670
rect 131625 148667 131691 148670
rect 182317 148730 182383 148733
rect 226477 148730 226543 148733
rect 182317 148728 184052 148730
rect 182317 148672 182322 148728
rect 182378 148672 184052 148728
rect 182317 148670 184052 148672
rect 223796 148728 226543 148730
rect 223796 148672 226482 148728
rect 226538 148672 226543 148728
rect 223796 148670 226543 148672
rect 182317 148667 182383 148670
rect 226477 148667 226543 148670
rect 80105 148594 80171 148597
rect 76780 148592 80171 148594
rect 76780 148536 80110 148592
rect 80166 148536 80171 148592
rect 76780 148534 80171 148536
rect 80105 148531 80171 148534
rect 233561 148458 233627 148461
rect 233561 148456 237044 148458
rect 233561 148400 233566 148456
rect 233622 148400 237044 148456
rect 233561 148398 237044 148400
rect 233561 148395 233627 148398
rect 87281 148322 87347 148325
rect 131533 148322 131599 148325
rect 173853 148322 173919 148325
rect 87281 148320 90028 148322
rect 87281 148264 87286 148320
rect 87342 148264 90028 148320
rect 87281 148262 90028 148264
rect 129772 148320 131599 148322
rect 129772 148264 131538 148320
rect 131594 148264 131599 148320
rect 129772 148262 131599 148264
rect 170804 148320 173919 148322
rect 170804 148264 173858 148320
rect 173914 148264 173919 148320
rect 170804 148262 173919 148264
rect 87281 148259 87347 148262
rect 131533 148259 131599 148262
rect 173853 148259 173919 148262
rect 181765 148322 181831 148325
rect 226477 148322 226543 148325
rect 181765 148320 184052 148322
rect 181765 148264 181770 148320
rect 181826 148264 184052 148320
rect 181765 148262 184052 148264
rect 223796 148320 226543 148322
rect 223796 148264 226482 148320
rect 226538 148264 226543 148320
rect 223796 148262 226543 148264
rect 181765 148259 181831 148262
rect 226477 148259 226543 148262
rect 139721 148186 139787 148189
rect 139721 148184 143020 148186
rect 139721 148128 139726 148184
rect 139782 148128 143020 148184
rect 139721 148126 143020 148128
rect 139721 148123 139787 148126
rect 87373 148050 87439 148053
rect 131349 148050 131415 148053
rect 87373 148048 90028 148050
rect 87373 147992 87378 148048
rect 87434 147992 90028 148048
rect 87373 147990 90028 147992
rect 129772 148048 131415 148050
rect 129772 147992 131354 148048
rect 131410 147992 131415 148048
rect 129772 147990 131415 147992
rect 87373 147987 87439 147990
rect 131349 147987 131415 147990
rect 182317 148050 182383 148053
rect 225557 148050 225623 148053
rect 182317 148048 184052 148050
rect 182317 147992 182322 148048
rect 182378 147992 184052 148048
rect 182317 147990 184052 147992
rect 223796 148048 225623 148050
rect 223796 147992 225562 148048
rect 225618 147992 225623 148048
rect 223796 147990 225623 147992
rect 182317 147987 182383 147990
rect 225557 147987 225623 147990
rect 79737 147914 79803 147917
rect 76780 147912 79803 147914
rect 76780 147856 79742 147912
rect 79798 147856 79803 147912
rect 76780 147854 79803 147856
rect 79737 147851 79803 147854
rect 233469 147914 233535 147917
rect 233469 147912 237044 147914
rect 233469 147856 233474 147912
rect 233530 147856 237044 147912
rect 233469 147854 237044 147856
rect 233469 147851 233535 147854
rect 174037 147778 174103 147781
rect 170804 147776 174103 147778
rect 170804 147720 174042 147776
rect 174098 147720 174103 147776
rect 170804 147718 174103 147720
rect 174037 147715 174103 147718
rect 140641 147506 140707 147509
rect 140641 147504 143020 147506
rect 140641 147448 140646 147504
rect 140702 147448 143020 147504
rect 140641 147446 143020 147448
rect 140641 147443 140707 147446
rect 79369 147370 79435 147373
rect 76780 147368 79435 147370
rect 76780 147312 79374 147368
rect 79430 147312 79435 147368
rect 76780 147310 79435 147312
rect 79369 147307 79435 147310
rect 172749 147234 172815 147237
rect 170804 147232 172815 147234
rect 170804 147176 172754 147232
rect 172810 147176 172815 147232
rect 170804 147174 172815 147176
rect 172749 147171 172815 147174
rect 233561 147234 233627 147237
rect 233561 147232 237044 147234
rect 233561 147176 233566 147232
rect 233622 147176 237044 147232
rect 233561 147174 237044 147176
rect 233561 147171 233627 147174
rect 79277 146826 79343 146829
rect 76780 146824 79343 146826
rect 76780 146768 79282 146824
rect 79338 146768 79343 146824
rect 76780 146766 79343 146768
rect 79277 146763 79343 146766
rect 139721 146826 139787 146829
rect 139721 146824 143020 146826
rect 139721 146768 139726 146824
rect 139782 146768 143020 146824
rect 139721 146766 143020 146768
rect 139721 146763 139787 146766
rect 174037 146554 174103 146557
rect 170804 146552 174103 146554
rect 170804 146496 174042 146552
rect 174098 146496 174103 146552
rect 170804 146494 174103 146496
rect 174037 146491 174103 146494
rect 233469 146554 233535 146557
rect 233469 146552 237044 146554
rect 233469 146496 233474 146552
rect 233530 146496 237044 146552
rect 233469 146494 237044 146496
rect 233469 146491 233535 146494
rect 80013 146282 80079 146285
rect 76780 146280 80079 146282
rect 76780 146224 80018 146280
rect 80074 146224 80079 146280
rect 76780 146222 80079 146224
rect 80013 146219 80079 146222
rect 140549 146146 140615 146149
rect 140549 146144 143020 146146
rect 140549 146088 140554 146144
rect 140610 146088 143020 146144
rect 140549 146086 143020 146088
rect 140549 146083 140615 146086
rect 172749 146010 172815 146013
rect 170804 146008 172815 146010
rect 170804 145952 172754 146008
rect 172810 145952 172815 146008
rect 170804 145950 172815 145952
rect 172749 145947 172815 145950
rect 233469 146010 233535 146013
rect 233469 146008 237044 146010
rect 233469 145952 233474 146008
rect 233530 145952 237044 146008
rect 233469 145950 237044 145952
rect 233469 145947 233535 145950
rect 79921 145602 79987 145605
rect 76780 145600 79987 145602
rect 76780 145544 79926 145600
rect 79982 145544 79987 145600
rect 76780 145542 79987 145544
rect 79921 145539 79987 145542
rect 139905 145466 139971 145469
rect 173669 145466 173735 145469
rect 139905 145464 143020 145466
rect 139905 145408 139910 145464
rect 139966 145408 143020 145464
rect 139905 145406 143020 145408
rect 170804 145464 173735 145466
rect 170804 145408 173674 145464
rect 173730 145408 173735 145464
rect 170804 145406 173735 145408
rect 139905 145403 139971 145406
rect 173669 145403 173735 145406
rect 233469 145330 233535 145333
rect 233469 145328 237044 145330
rect 233469 145272 233474 145328
rect 233530 145272 237044 145328
rect 233469 145270 237044 145272
rect 233469 145267 233535 145270
rect 79829 145058 79895 145061
rect 76780 145056 79895 145058
rect 76780 145000 79834 145056
rect 79890 145000 79895 145056
rect 76780 144998 79895 145000
rect 79829 144995 79895 144998
rect 173577 144922 173643 144925
rect 170804 144920 173643 144922
rect 170804 144864 173582 144920
rect 173638 144864 173643 144920
rect 170804 144862 173643 144864
rect 173577 144859 173643 144862
rect 140457 144786 140523 144789
rect 140457 144784 143020 144786
rect 140457 144728 140462 144784
rect 140518 144728 143020 144784
rect 140457 144726 143020 144728
rect 140457 144723 140523 144726
rect 233653 144650 233719 144653
rect 233653 144648 237044 144650
rect 233653 144592 233658 144648
rect 233714 144592 237044 144648
rect 233653 144590 237044 144592
rect 233653 144587 233719 144590
rect 80197 144514 80263 144517
rect 76780 144512 80263 144514
rect 76780 144456 80202 144512
rect 80258 144456 80263 144512
rect 76780 144454 80263 144456
rect 80197 144451 80263 144454
rect 173945 144378 174011 144381
rect 170804 144376 174011 144378
rect 170804 144320 173950 144376
rect 174006 144320 174011 144376
rect 170804 144318 174011 144320
rect 173945 144315 174011 144318
rect 46985 144106 47051 144109
rect 48222 144106 48228 144108
rect 46985 144104 48228 144106
rect 46985 144048 46990 144104
rect 47046 144048 48228 144104
rect 46985 144046 48228 144048
rect 46985 144043 47051 144046
rect 48222 144044 48228 144046
rect 48292 144044 48298 144108
rect 138893 144106 138959 144109
rect 233745 144106 233811 144109
rect 138893 144104 143020 144106
rect 138893 144048 138898 144104
rect 138954 144048 143020 144104
rect 138893 144046 143020 144048
rect 233745 144104 237044 144106
rect 233745 144048 233750 144104
rect 233806 144048 237044 144104
rect 233745 144046 237044 144048
rect 138893 144043 138959 144046
rect 233745 144043 233811 144046
rect 109545 143972 109611 143973
rect 109494 143908 109500 143972
rect 109564 143970 109611 143972
rect 109564 143968 109656 143970
rect 109606 143912 109656 143968
rect 109564 143910 109656 143912
rect 109564 143908 109611 143910
rect 109545 143907 109611 143908
rect 80197 143834 80263 143837
rect 173485 143834 173551 143837
rect 76780 143832 80263 143834
rect 76780 143776 80202 143832
rect 80258 143776 80263 143832
rect 76780 143774 80263 143776
rect 170804 143832 173551 143834
rect 170804 143776 173490 143832
rect 173546 143776 173551 143832
rect 170804 143774 173551 143776
rect 80197 143771 80263 143774
rect 173485 143771 173551 143774
rect 300169 143562 300235 143565
rect 303416 143562 303896 143592
rect 300169 143560 303896 143562
rect 300169 143504 300174 143560
rect 300230 143504 303896 143560
rect 300169 143502 303896 143504
rect 300169 143499 300235 143502
rect 303416 143472 303896 143502
rect 140365 143426 140431 143429
rect 233929 143426 233995 143429
rect 140365 143424 143020 143426
rect 140365 143368 140370 143424
rect 140426 143368 143020 143424
rect 140365 143366 143020 143368
rect 233929 143424 237044 143426
rect 233929 143368 233934 143424
rect 233990 143368 237044 143424
rect 233929 143366 237044 143368
rect 140365 143363 140431 143366
rect 233929 143363 233995 143366
rect 80013 143290 80079 143293
rect 173853 143290 173919 143293
rect 76780 143288 80079 143290
rect 76780 143232 80018 143288
rect 80074 143232 80079 143288
rect 76780 143230 80079 143232
rect 170804 143288 173919 143290
rect 170804 143232 173858 143288
rect 173914 143232 173919 143288
rect 170804 143230 173919 143232
rect 80013 143227 80079 143230
rect 173853 143227 173919 143230
rect 80105 142746 80171 142749
rect 76780 142744 80171 142746
rect 76780 142688 80110 142744
rect 80166 142688 80171 142744
rect 76780 142686 80171 142688
rect 80105 142683 80171 142686
rect 139721 142746 139787 142749
rect 173301 142746 173367 142749
rect 139721 142744 143020 142746
rect 139721 142688 139726 142744
rect 139782 142688 143020 142744
rect 139721 142686 143020 142688
rect 170804 142744 173367 142746
rect 170804 142688 173306 142744
rect 173362 142688 173367 142744
rect 170804 142686 173367 142688
rect 139721 142683 139787 142686
rect 173301 142683 173367 142686
rect 233837 142746 233903 142749
rect 233837 142744 237044 142746
rect 233837 142688 233842 142744
rect 233898 142688 237044 142744
rect 233837 142686 237044 142688
rect 233837 142683 233903 142686
rect 80197 142202 80263 142205
rect 76780 142200 80263 142202
rect 76780 142144 80202 142200
rect 80258 142144 80263 142200
rect 76780 142142 80263 142144
rect 80197 142139 80263 142142
rect 139629 142202 139695 142205
rect 173393 142202 173459 142205
rect 139629 142200 143020 142202
rect 139629 142144 139634 142200
rect 139690 142144 143020 142200
rect 139629 142142 143020 142144
rect 170804 142200 173459 142202
rect 170804 142144 173398 142200
rect 173454 142144 173459 142200
rect 170804 142142 173459 142144
rect 139629 142139 139695 142142
rect 173393 142139 173459 142142
rect 233469 142202 233535 142205
rect 233469 142200 237044 142202
rect 233469 142144 233474 142200
rect 233530 142144 237044 142200
rect 233469 142142 237044 142144
rect 233469 142139 233535 142142
rect 128446 139828 128452 139892
rect 128516 139890 128522 139892
rect 170541 139890 170607 139893
rect 128516 139888 170607 139890
rect 128516 139832 170546 139888
rect 170602 139832 170607 139888
rect 128516 139830 170607 139832
rect 128516 139828 128522 139830
rect 170541 139827 170607 139830
rect 232825 139890 232891 139893
rect 263277 139890 263343 139893
rect 232825 139888 263343 139890
rect 232825 139832 232830 139888
rect 232886 139832 263282 139888
rect 263338 139832 263343 139888
rect 232825 139830 263343 139832
rect 232825 139827 232891 139830
rect 263277 139827 263343 139830
rect 264565 138666 264631 138669
rect 264974 138666 264980 138668
rect 264565 138664 264980 138666
rect 264565 138608 264570 138664
rect 264626 138608 264980 138664
rect 264565 138606 264980 138608
rect 264565 138603 264631 138606
rect 264974 138604 264980 138606
rect 265044 138604 265050 138668
rect 134710 132954 134770 132988
rect 136869 132954 136935 132957
rect 134710 132952 136935 132954
rect 134710 132896 136874 132952
rect 136930 132896 136935 132952
rect 134710 132894 136935 132896
rect 228734 132954 228794 132988
rect 231905 132954 231971 132957
rect 228734 132952 231971 132954
rect 228734 132896 231910 132952
rect 231966 132896 231971 132952
rect 228734 132894 231971 132896
rect 136869 132891 136935 132894
rect 231905 132891 231971 132894
rect 13681 131594 13747 131597
rect 20806 131594 20812 131596
rect 13681 131592 20812 131594
rect 13681 131536 13686 131592
rect 13742 131536 20812 131592
rect 13681 131534 20812 131536
rect 13681 131531 13747 131534
rect 20806 131532 20812 131534
rect 20876 131532 20882 131596
rect 60509 131458 60575 131461
rect 61613 131458 61679 131461
rect 60509 131456 61679 131458
rect 60509 131400 60514 131456
rect 60570 131400 61618 131456
rect 61674 131400 61679 131456
rect 60509 131398 61679 131400
rect 60509 131395 60575 131398
rect 61613 131395 61679 131398
rect 58761 131186 58827 131189
rect 60877 131186 60943 131189
rect 58761 131184 60943 131186
rect 58761 131128 58766 131184
rect 58822 131128 60882 131184
rect 60938 131128 60943 131184
rect 58761 131126 60943 131128
rect 58761 131123 58827 131126
rect 60877 131123 60943 131126
rect 134710 130914 134770 131492
rect 138893 130914 138959 130917
rect 134710 130912 138959 130914
rect 134710 130856 138898 130912
rect 138954 130856 138959 130912
rect 134710 130854 138959 130856
rect 228734 130914 228794 131492
rect 232733 130914 232799 130917
rect 228734 130912 232799 130914
rect 228734 130856 232738 130912
rect 232794 130856 232799 130912
rect 228734 130854 232799 130856
rect 138893 130851 138959 130854
rect 232733 130851 232799 130854
rect 23893 130370 23959 130373
rect 69750 130370 69756 130372
rect 23893 130368 69756 130370
rect 23893 130312 23898 130368
rect 23954 130312 69756 130368
rect 23893 130310 69756 130312
rect 23893 130307 23959 130310
rect 69750 130308 69756 130310
rect 69820 130308 69826 130372
rect 288710 130308 288716 130372
rect 288780 130370 288786 130372
rect 289865 130370 289931 130373
rect 288780 130368 289931 130370
rect 288780 130312 289870 130368
rect 289926 130312 289931 130368
rect 288780 130310 289931 130312
rect 288780 130308 288786 130310
rect 289865 130307 289931 130310
rect 58158 130172 58164 130236
rect 58228 130234 58234 130236
rect 61470 130234 61476 130236
rect 58228 130174 61476 130234
rect 58228 130172 58234 130174
rect 61470 130172 61476 130174
rect 61540 130172 61546 130236
rect 135438 130172 135444 130236
rect 135508 130234 135514 130236
rect 138750 130234 138756 130236
rect 135508 130174 138756 130234
rect 135508 130172 135514 130174
rect 138750 130172 138756 130174
rect 138820 130172 138826 130236
rect 231997 130234 232063 130237
rect 228734 130232 232063 130234
rect 228734 130176 232002 130232
rect 232058 130176 232063 130232
rect 228734 130174 232063 130176
rect 136869 130098 136935 130101
rect 134710 130096 136935 130098
rect 134710 130040 136874 130096
rect 136930 130040 136935 130096
rect 134710 130038 136935 130040
rect 134710 129864 134770 130038
rect 136869 130035 136935 130038
rect 228734 129864 228794 130174
rect 231997 130171 232063 130174
rect 243998 130172 244004 130236
rect 244068 130234 244074 130236
rect 245102 130234 245108 130236
rect 244068 130174 245108 130234
rect 244068 130172 244074 130174
rect 245102 130172 245108 130174
rect 245172 130172 245178 130236
rect 48590 129492 48596 129556
rect 48660 129554 48666 129556
rect 57790 129554 57796 129556
rect 48660 129494 57796 129554
rect 48660 129492 48666 129494
rect 57790 129492 57796 129494
rect 57860 129492 57866 129556
rect 251358 129492 251364 129556
rect 251428 129554 251434 129556
rect 269206 129554 269212 129556
rect 251428 129494 269212 129554
rect 251428 129492 251434 129494
rect 269206 129492 269212 129494
rect 269276 129492 269282 129556
rect 134710 127922 134770 128364
rect 136869 127922 136935 127925
rect 134710 127920 136935 127922
rect 134710 127864 136874 127920
rect 136930 127864 136935 127920
rect 134710 127862 136935 127864
rect 228734 127922 228794 128364
rect 230709 127922 230775 127925
rect 228734 127920 230775 127922
rect 228734 127864 230714 127920
rect 230770 127864 230775 127920
rect 228734 127862 230775 127864
rect 136869 127859 136935 127862
rect 230709 127859 230775 127862
rect 148694 127590 148938 127650
rect 148694 127517 148754 127590
rect 148694 127512 148803 127517
rect 148694 127456 148742 127512
rect 148798 127456 148803 127512
rect 148878 127484 148938 127590
rect 148694 127454 148803 127456
rect 148737 127451 148803 127454
rect 241606 127452 241612 127516
rect 241676 127514 241682 127516
rect 241676 127454 242932 127514
rect 241676 127452 241682 127454
rect 137881 127378 137947 127381
rect 134710 127376 137947 127378
rect 134710 127320 137886 127376
rect 137942 127320 137947 127376
rect 134710 127318 137947 127320
rect 134710 126736 134770 127318
rect 137881 127315 137947 127318
rect 231721 127106 231787 127109
rect 228734 127104 231787 127106
rect 228734 127048 231726 127104
rect 231782 127048 231787 127104
rect 228734 127046 231787 127048
rect 228734 126736 228794 127046
rect 231721 127043 231787 127046
rect 145609 125338 145675 125341
rect 145609 125336 148938 125338
rect 145609 125280 145614 125336
rect 145670 125280 148938 125336
rect 145609 125278 148938 125280
rect 145609 125275 145675 125278
rect 134710 125066 134770 125236
rect 148878 125172 148938 125278
rect 228734 125202 228794 125236
rect 231629 125202 231695 125205
rect 228734 125200 231695 125202
rect 228734 125144 231634 125200
rect 231690 125144 231695 125200
rect 228734 125142 231695 125144
rect 231629 125139 231695 125142
rect 240921 125202 240987 125205
rect 240921 125200 242932 125202
rect 240921 125144 240926 125200
rect 240982 125144 242932 125200
rect 240921 125142 242932 125144
rect 240921 125139 240987 125142
rect 138157 125066 138223 125069
rect 134710 125064 138223 125066
rect 134710 125008 138162 125064
rect 138218 125008 138223 125064
rect 134710 125006 138223 125008
rect 138157 125003 138223 125006
rect 38153 124794 38219 124797
rect 35748 124792 38219 124794
rect 35748 124736 38158 124792
rect 38214 124736 38219 124792
rect 35748 124734 38219 124736
rect 38153 124731 38219 124734
rect 137973 124250 138039 124253
rect 231813 124250 231879 124253
rect 134710 124248 138039 124250
rect 134710 124192 137978 124248
rect 138034 124192 138039 124248
rect 134710 124190 138039 124192
rect 134710 123608 134770 124190
rect 137973 124187 138039 124190
rect 228734 124248 231879 124250
rect 228734 124192 231818 124248
rect 231874 124192 231879 124248
rect 228734 124190 231879 124192
rect 228734 123608 228794 124190
rect 231813 124187 231879 124190
rect 276065 123706 276131 123709
rect 276065 123704 278076 123706
rect 276065 123648 276070 123704
rect 276126 123648 278076 123704
rect 276065 123646 278076 123648
rect 276065 123643 276131 123646
rect 47813 123298 47879 123301
rect 48222 123298 48228 123300
rect 47813 123296 48228 123298
rect 47813 123240 47818 123296
rect 47874 123240 48228 123296
rect 47813 123238 48228 123240
rect 47813 123235 47879 123238
rect 48222 123236 48228 123238
rect 48292 123236 48298 123300
rect 9896 123162 10376 123192
rect 13405 123162 13471 123165
rect 9896 123160 13471 123162
rect 9896 123104 13410 123160
rect 13466 123104 13471 123160
rect 9896 123102 13471 123104
rect 9896 123072 10376 123102
rect 13405 123099 13471 123102
rect 145609 123026 145675 123029
rect 145609 123024 148938 123026
rect 145609 122968 145614 123024
rect 145670 122968 148938 123024
rect 145609 122966 148938 122968
rect 145609 122963 145675 122966
rect 148878 122860 148938 122966
rect 240921 122890 240987 122893
rect 240921 122888 242932 122890
rect 240921 122832 240926 122888
rect 240982 122832 242932 122888
rect 240921 122830 242932 122832
rect 240921 122827 240987 122830
rect 51309 122210 51375 122213
rect 51309 122208 55068 122210
rect 51309 122152 51314 122208
rect 51370 122152 55068 122208
rect 51309 122150 55068 122152
rect 51309 122147 51375 122150
rect 134710 122074 134770 122108
rect 138157 122074 138223 122077
rect 134710 122072 138223 122074
rect 134710 122016 138162 122072
rect 138218 122016 138223 122072
rect 134710 122014 138223 122016
rect 228734 122074 228794 122108
rect 231629 122074 231695 122077
rect 293686 122076 293746 122180
rect 228734 122072 231695 122074
rect 228734 122016 231634 122072
rect 231690 122016 231695 122072
rect 228734 122014 231695 122016
rect 138157 122011 138223 122014
rect 231629 122011 231695 122014
rect 293678 122012 293684 122076
rect 293748 122012 293754 122076
rect 175509 121938 175575 121941
rect 175509 121936 178930 121938
rect 175509 121880 175514 121936
rect 175570 121880 178930 121936
rect 175509 121878 178930 121880
rect 175509 121875 175575 121878
rect 178870 121432 178930 121878
rect 81710 121332 81716 121396
rect 81780 121394 81786 121396
rect 85030 121394 85090 121428
rect 81780 121334 85090 121394
rect 81780 121332 81786 121334
rect 261069 120716 261135 120717
rect 261069 120714 261116 120716
rect 260988 120712 261116 120714
rect 261180 120714 261186 120716
rect 264974 120714 264980 120716
rect 260988 120656 261074 120712
rect 260988 120654 261116 120656
rect 261069 120652 261116 120654
rect 261180 120654 264980 120714
rect 261180 120652 261186 120654
rect 264974 120652 264980 120654
rect 265044 120652 265050 120716
rect 261069 120651 261135 120652
rect 137789 120578 137855 120581
rect 134710 120576 137855 120578
rect 134710 120520 137794 120576
rect 137850 120520 137855 120576
rect 134710 120518 137855 120520
rect 134710 120480 134770 120518
rect 137789 120515 137855 120518
rect 145609 120578 145675 120581
rect 231721 120578 231787 120581
rect 145609 120576 148938 120578
rect 145609 120520 145614 120576
rect 145670 120520 148938 120576
rect 145609 120518 148938 120520
rect 145609 120515 145675 120518
rect 148878 120412 148938 120518
rect 228734 120576 231787 120578
rect 228734 120520 231726 120576
rect 231782 120520 231787 120576
rect 228734 120518 231787 120520
rect 228734 120480 228794 120518
rect 231721 120515 231787 120518
rect 240921 120442 240987 120445
rect 240921 120440 242932 120442
rect 240921 120384 240926 120440
rect 240982 120384 242932 120440
rect 240921 120382 242932 120384
rect 240921 120379 240987 120382
rect 228501 120306 228567 120309
rect 229646 120306 229652 120308
rect 228501 120304 229652 120306
rect 228501 120248 228506 120304
rect 228562 120248 229652 120304
rect 228501 120246 229652 120248
rect 228501 120243 228567 120246
rect 229646 120244 229652 120246
rect 229716 120244 229722 120308
rect 300169 119082 300235 119085
rect 303416 119082 303896 119112
rect 300169 119080 303896 119082
rect 300169 119024 300174 119080
rect 300230 119024 303896 119080
rect 300169 119022 303896 119024
rect 300169 119019 300235 119022
rect 303416 118992 303896 119022
rect 134710 118402 134770 118980
rect 167229 118810 167295 118813
rect 167873 118810 167939 118813
rect 164732 118808 167939 118810
rect 164732 118752 167234 118808
rect 167290 118752 167878 118808
rect 167934 118752 167939 118808
rect 164732 118750 167939 118752
rect 228734 118810 228794 118980
rect 231629 118810 231695 118813
rect 261069 118810 261135 118813
rect 228734 118808 231695 118810
rect 228734 118752 231634 118808
rect 231690 118752 231695 118808
rect 228734 118750 231695 118752
rect 258756 118808 261135 118810
rect 258756 118752 261074 118808
rect 261130 118752 261135 118808
rect 258756 118750 261135 118752
rect 167229 118747 167295 118750
rect 167873 118747 167939 118750
rect 231629 118747 231695 118750
rect 261069 118747 261135 118750
rect 138157 118402 138223 118405
rect 134710 118400 138223 118402
rect 134710 118344 138162 118400
rect 138218 118344 138223 118400
rect 134710 118342 138223 118344
rect 138157 118339 138223 118342
rect 145609 118266 145675 118269
rect 145609 118264 148938 118266
rect 145609 118208 145614 118264
rect 145670 118208 148938 118264
rect 145609 118206 148938 118208
rect 145609 118203 145675 118206
rect 148878 118100 148938 118206
rect 240921 118130 240987 118133
rect 240921 118128 242932 118130
rect 240921 118072 240926 118128
rect 240982 118072 242932 118128
rect 240921 118070 242932 118072
rect 240921 118067 240987 118070
rect 137697 117858 137763 117861
rect 134710 117856 137763 117858
rect 134710 117800 137702 117856
rect 137758 117800 137763 117856
rect 134710 117798 137763 117800
rect 38337 117450 38403 117453
rect 35718 117448 38403 117450
rect 35718 117392 38342 117448
rect 38398 117392 38403 117448
rect 35718 117390 38403 117392
rect 35718 116808 35778 117390
rect 38337 117387 38403 117390
rect 134710 117352 134770 117798
rect 137697 117795 137763 117798
rect 231537 117586 231603 117589
rect 228734 117584 231603 117586
rect 228734 117528 231542 117584
rect 231598 117528 231603 117584
rect 228734 117526 231603 117528
rect 228734 117352 228794 117526
rect 231537 117523 231603 117526
rect 145609 115954 145675 115957
rect 145609 115952 148938 115954
rect 145609 115896 145614 115952
rect 145670 115896 148938 115952
rect 145609 115894 148938 115896
rect 145609 115891 145675 115894
rect 134710 115274 134770 115852
rect 148878 115788 148938 115894
rect 137329 115274 137395 115277
rect 134710 115272 137395 115274
rect 134710 115216 137334 115272
rect 137390 115216 137395 115272
rect 134710 115214 137395 115216
rect 228734 115274 228794 115852
rect 240921 115818 240987 115821
rect 240921 115816 242932 115818
rect 240921 115760 240926 115816
rect 240982 115760 242932 115816
rect 240921 115758 242932 115760
rect 240921 115755 240987 115758
rect 231261 115274 231327 115277
rect 228734 115272 231327 115274
rect 228734 115216 231266 115272
rect 231322 115216 231327 115272
rect 228734 115214 231327 115216
rect 137329 115211 137395 115214
rect 231261 115211 231327 115214
rect 137605 114866 137671 114869
rect 231353 114866 231419 114869
rect 134710 114864 137671 114866
rect 134710 114808 137610 114864
rect 137666 114808 137671 114864
rect 134710 114806 137671 114808
rect 134710 114224 134770 114806
rect 137605 114803 137671 114806
rect 228734 114864 231419 114866
rect 228734 114808 231358 114864
rect 231414 114808 231419 114864
rect 228734 114806 231419 114808
rect 228734 114224 228794 114806
rect 231353 114803 231419 114806
rect 274869 114458 274935 114461
rect 274869 114456 278106 114458
rect 274869 114400 274874 114456
rect 274930 114400 278106 114456
rect 274869 114398 278106 114400
rect 274869 114395 274935 114398
rect 278046 113816 278106 114398
rect 145609 113506 145675 113509
rect 145609 113504 148938 113506
rect 145609 113448 145614 113504
rect 145670 113448 148938 113504
rect 145609 113446 148938 113448
rect 145609 113443 145675 113446
rect 148878 113340 148938 113446
rect 240737 113370 240803 113373
rect 240737 113368 242932 113370
rect 240737 113312 240742 113368
rect 240798 113312 242932 113368
rect 240737 113310 242932 113312
rect 240737 113307 240803 113310
rect 134710 112690 134770 112724
rect 138157 112690 138223 112693
rect 134710 112688 138223 112690
rect 134710 112632 138162 112688
rect 138218 112632 138223 112688
rect 134710 112630 138223 112632
rect 138157 112627 138223 112630
rect 228734 112418 228794 112724
rect 231353 112418 231419 112421
rect 228734 112416 231419 112418
rect 228734 112360 231358 112416
rect 231414 112360 231419 112416
rect 228734 112358 231419 112360
rect 231353 112355 231419 112358
rect 137513 111738 137579 111741
rect 231445 111738 231511 111741
rect 134710 111736 137579 111738
rect 134710 111680 137518 111736
rect 137574 111680 137579 111736
rect 134710 111678 137579 111680
rect 134710 111096 134770 111678
rect 137513 111675 137579 111678
rect 228734 111736 231511 111738
rect 228734 111680 231450 111736
rect 231506 111680 231511 111736
rect 228734 111678 231511 111680
rect 145609 111194 145675 111197
rect 145609 111192 148938 111194
rect 145609 111136 145614 111192
rect 145670 111136 148938 111192
rect 145609 111134 148938 111136
rect 145609 111131 145675 111134
rect 148878 111028 148938 111134
rect 228734 111096 228794 111678
rect 231445 111675 231511 111678
rect 240921 111058 240987 111061
rect 240921 111056 242932 111058
rect 240921 111000 240926 111056
rect 240982 111000 242932 111056
rect 240921 110998 242932 111000
rect 240921 110995 240987 110998
rect 137513 109698 137579 109701
rect 231537 109698 231603 109701
rect 134710 109696 137579 109698
rect 134710 109640 137518 109696
rect 137574 109640 137579 109696
rect 134710 109638 137579 109640
rect 134710 109600 134770 109638
rect 137513 109635 137579 109638
rect 228734 109696 231603 109698
rect 228734 109640 231542 109696
rect 231598 109640 231603 109696
rect 228734 109638 231603 109640
rect 228734 109600 228794 109638
rect 231537 109635 231603 109638
rect 293545 109562 293611 109565
rect 293502 109560 293611 109562
rect 293502 109504 293550 109560
rect 293606 109504 293611 109560
rect 293502 109499 293611 109504
rect 38245 109426 38311 109429
rect 35718 109424 38311 109426
rect 35718 109368 38250 109424
rect 38306 109368 38311 109424
rect 35718 109366 38311 109368
rect 20078 108476 20138 108852
rect 35718 108784 35778 109366
rect 38245 109363 38311 109366
rect 74033 109018 74099 109021
rect 70862 109016 74099 109018
rect 70862 108960 74038 109016
rect 74094 108960 74099 109016
rect 70862 108958 74099 108960
rect 51309 108882 51375 108885
rect 51309 108880 55068 108882
rect 51309 108824 51314 108880
rect 51370 108824 55068 108880
rect 70862 108852 70922 108958
rect 74033 108955 74099 108958
rect 293502 108920 293562 109499
rect 145609 108882 145675 108885
rect 145609 108880 148938 108882
rect 51309 108822 55068 108824
rect 145609 108824 145614 108880
rect 145670 108824 148938 108880
rect 145609 108822 148938 108824
rect 51309 108819 51375 108822
rect 145609 108819 145675 108822
rect 148878 108716 148938 108822
rect 240829 108746 240895 108749
rect 240829 108744 242932 108746
rect 240829 108688 240834 108744
rect 240890 108688 242932 108744
rect 240829 108686 242932 108688
rect 240829 108683 240895 108686
rect 20070 108412 20076 108476
rect 20140 108412 20146 108476
rect 35894 108276 35900 108340
rect 35964 108338 35970 108340
rect 47077 108338 47143 108341
rect 47813 108338 47879 108341
rect 35964 108336 47879 108338
rect 35964 108280 47082 108336
rect 47138 108280 47818 108336
rect 47874 108280 47879 108336
rect 35964 108278 47879 108280
rect 35964 108276 35970 108278
rect 47077 108275 47143 108278
rect 47813 108275 47879 108278
rect 137881 108202 137947 108205
rect 134710 108200 137947 108202
rect 134710 108144 137886 108200
rect 137942 108144 137947 108200
rect 134710 108142 137947 108144
rect 134710 107968 134770 108142
rect 137881 108139 137947 108142
rect 231721 108066 231787 108069
rect 228734 108064 231787 108066
rect 228734 108008 231726 108064
rect 231782 108008 231787 108064
rect 228734 108006 231787 108008
rect 228734 107968 228794 108006
rect 231721 108003 231787 108006
rect 137973 106706 138039 106709
rect 231813 106706 231879 106709
rect 134710 106704 138039 106706
rect 134710 106648 137978 106704
rect 138034 106648 138039 106704
rect 134710 106646 138039 106648
rect 134710 106472 134770 106646
rect 137973 106643 138039 106646
rect 228734 106704 231879 106706
rect 228734 106648 231818 106704
rect 231874 106648 231879 106704
rect 228734 106646 231879 106648
rect 145609 106570 145675 106573
rect 145609 106568 148938 106570
rect 145609 106512 145614 106568
rect 145670 106512 148938 106568
rect 145609 106510 148938 106512
rect 145609 106507 145675 106510
rect 148878 106404 148938 106510
rect 228734 106472 228794 106646
rect 231813 106643 231879 106646
rect 240921 106434 240987 106437
rect 240921 106432 242932 106434
rect 240921 106376 240926 106432
rect 240982 106376 242932 106432
rect 240921 106374 242932 106376
rect 240921 106371 240987 106374
rect 138065 105346 138131 105349
rect 231905 105346 231971 105349
rect 134710 105344 138131 105346
rect 134710 105288 138070 105344
rect 138126 105288 138131 105344
rect 134710 105286 138131 105288
rect 134710 104840 134770 105286
rect 138065 105283 138131 105286
rect 228734 105344 231971 105346
rect 228734 105288 231910 105344
rect 231966 105288 231971 105344
rect 228734 105286 231971 105288
rect 228734 104840 228794 105286
rect 231905 105283 231971 105286
rect 148694 104062 148938 104122
rect 137789 103986 137855 103989
rect 134710 103984 137855 103986
rect 134710 103928 137794 103984
rect 137850 103928 137855 103984
rect 134710 103926 137855 103928
rect 134710 103344 134770 103926
rect 137789 103923 137855 103926
rect 145425 103986 145491 103989
rect 148694 103986 148754 104062
rect 145425 103984 148754 103986
rect 145425 103928 145430 103984
rect 145486 103928 148754 103984
rect 148878 103956 148938 104062
rect 231629 103986 231695 103989
rect 228734 103984 231695 103986
rect 145425 103926 148754 103928
rect 228734 103928 231634 103984
rect 231690 103928 231695 103984
rect 228734 103926 231695 103928
rect 145425 103923 145491 103926
rect 228734 103344 228794 103926
rect 231629 103923 231695 103926
rect 240737 103986 240803 103989
rect 240737 103984 242932 103986
rect 240737 103928 240742 103984
rect 240798 103928 242932 103984
rect 240737 103926 242932 103928
rect 240737 103923 240803 103926
rect 274869 103714 274935 103717
rect 274869 103712 278076 103714
rect 274869 103656 274874 103712
rect 274930 103656 278076 103712
rect 274869 103654 278076 103656
rect 274869 103651 274935 103654
rect 231537 102354 231603 102357
rect 228734 102352 231603 102354
rect 228734 102296 231542 102352
rect 231598 102296 231603 102352
rect 228734 102294 231603 102296
rect 137697 102218 137763 102221
rect 134710 102216 137763 102218
rect 134710 102160 137702 102216
rect 137758 102160 137763 102216
rect 134710 102158 137763 102160
rect 134710 101712 134770 102158
rect 137697 102155 137763 102158
rect 145609 101810 145675 101813
rect 145609 101808 148938 101810
rect 145609 101752 145614 101808
rect 145670 101752 148938 101808
rect 145609 101750 148938 101752
rect 145609 101747 145675 101750
rect 148878 101644 148938 101750
rect 228734 101712 228794 102294
rect 231537 102291 231603 102294
rect 240369 101674 240435 101677
rect 240369 101672 242932 101674
rect 240369 101616 240374 101672
rect 240430 101616 242932 101672
rect 240369 101614 242932 101616
rect 240369 101611 240435 101614
rect 137421 100858 137487 100861
rect 231261 100858 231327 100861
rect 134710 100856 137487 100858
rect 134710 100800 137426 100856
rect 137482 100800 137487 100856
rect 134710 100798 137487 100800
rect 38245 100722 38311 100725
rect 35748 100720 38311 100722
rect 35748 100664 38250 100720
rect 38306 100664 38311 100720
rect 35748 100662 38311 100664
rect 38245 100659 38311 100662
rect 134710 100216 134770 100798
rect 137421 100795 137487 100798
rect 228734 100856 231327 100858
rect 228734 100800 231266 100856
rect 231322 100800 231327 100856
rect 228734 100798 231327 100800
rect 228734 100216 228794 100798
rect 231261 100795 231327 100798
rect 145609 99498 145675 99501
rect 145609 99496 148938 99498
rect 145609 99440 145614 99496
rect 145670 99440 148938 99496
rect 145609 99438 148938 99440
rect 145609 99435 145675 99438
rect 148878 99332 148938 99438
rect 240829 99362 240895 99365
rect 240829 99360 242932 99362
rect 240829 99304 240834 99360
rect 240890 99304 242932 99360
rect 240829 99302 242932 99304
rect 240829 99299 240895 99302
rect 138157 99226 138223 99229
rect 231997 99226 232063 99229
rect 134710 99224 138223 99226
rect 134710 99168 138162 99224
rect 138218 99168 138223 99224
rect 134710 99166 138223 99168
rect 134710 98584 134770 99166
rect 138157 99163 138223 99166
rect 228734 99224 232063 99226
rect 228734 99168 232002 99224
rect 232058 99168 232063 99224
rect 228734 99166 232063 99168
rect 167873 98818 167939 98821
rect 164732 98816 167939 98818
rect 164732 98760 167878 98816
rect 167934 98760 167939 98816
rect 164732 98758 167939 98760
rect 167873 98755 167939 98758
rect 228734 98584 228794 99166
rect 231997 99163 232063 99166
rect 262357 98818 262423 98821
rect 258756 98816 262423 98818
rect 258756 98760 262362 98816
rect 262418 98760 262423 98816
rect 258756 98758 262423 98760
rect 262357 98755 262423 98758
rect 134710 97050 134770 97084
rect 137329 97050 137395 97053
rect 134710 97048 137395 97050
rect 134710 96992 137334 97048
rect 137390 96992 137395 97048
rect 134710 96990 137395 96992
rect 137329 96987 137395 96990
rect 144597 97050 144663 97053
rect 175509 97050 175575 97053
rect 228734 97050 228794 97084
rect 231445 97050 231511 97053
rect 144597 97048 148938 97050
rect 144597 96992 144602 97048
rect 144658 96992 148938 97048
rect 144597 96990 148938 96992
rect 144597 96987 144663 96990
rect 81669 96914 81735 96917
rect 81669 96912 85090 96914
rect 81669 96856 81674 96912
rect 81730 96856 85090 96912
rect 148878 96884 148938 96990
rect 175509 97048 178930 97050
rect 175509 96992 175514 97048
rect 175570 96992 178930 97048
rect 175509 96990 178930 96992
rect 228734 97048 231511 97050
rect 228734 96992 231450 97048
rect 231506 96992 231511 97048
rect 228734 96990 231511 96992
rect 175509 96987 175575 96990
rect 81669 96854 85090 96856
rect 81669 96851 81735 96854
rect 85030 96408 85090 96854
rect 178870 96408 178930 96990
rect 231445 96987 231511 96990
rect 240921 96914 240987 96917
rect 240921 96912 242932 96914
rect 240921 96856 240926 96912
rect 240982 96856 242932 96912
rect 240921 96854 242932 96856
rect 240921 96851 240987 96854
rect 138157 95690 138223 95693
rect 231721 95690 231787 95693
rect 134710 95688 138223 95690
rect 134710 95632 138162 95688
rect 138218 95632 138223 95688
rect 134710 95630 138223 95632
rect 51309 95554 51375 95557
rect 51309 95552 55068 95554
rect 51309 95496 51314 95552
rect 51370 95496 55068 95552
rect 51309 95494 55068 95496
rect 51309 95491 51375 95494
rect 134710 95456 134770 95630
rect 138157 95627 138223 95630
rect 228734 95688 231787 95690
rect 228734 95632 231726 95688
rect 231782 95632 231787 95688
rect 228734 95630 231787 95632
rect 228734 95456 228794 95630
rect 231721 95627 231787 95630
rect 295569 95554 295635 95557
rect 293716 95552 295635 95554
rect 293716 95496 295574 95552
rect 295630 95496 295635 95552
rect 293716 95494 295635 95496
rect 295569 95491 295635 95494
rect 146345 94738 146411 94741
rect 146345 94736 148938 94738
rect 146345 94680 146350 94736
rect 146406 94680 148938 94736
rect 146345 94678 148938 94680
rect 146345 94675 146411 94678
rect 148878 94572 148938 94678
rect 240921 94602 240987 94605
rect 299709 94602 299775 94605
rect 303416 94602 303896 94632
rect 240921 94600 242932 94602
rect 240921 94544 240926 94600
rect 240982 94544 242932 94600
rect 240921 94542 242932 94544
rect 299709 94600 303896 94602
rect 299709 94544 299714 94600
rect 299770 94544 303896 94600
rect 299709 94542 303896 94544
rect 240921 94539 240987 94542
rect 299709 94539 299775 94542
rect 303416 94512 303896 94542
rect 274869 94330 274935 94333
rect 274869 94328 278106 94330
rect 274869 94272 274874 94328
rect 274930 94272 278106 94328
rect 274869 94270 278106 94272
rect 274869 94267 274935 94270
rect 231813 94194 231879 94197
rect 228734 94192 231879 94194
rect 228734 94136 231818 94192
rect 231874 94136 231879 94192
rect 228734 94134 231879 94136
rect 228734 93960 228794 94134
rect 231813 94131 231879 94134
rect 134710 93922 134770 93956
rect 138157 93922 138223 93925
rect 134710 93920 138223 93922
rect 134710 93864 138162 93920
rect 138218 93864 138223 93920
rect 134710 93862 138223 93864
rect 138157 93859 138223 93862
rect 278046 93824 278106 94270
rect 38797 92970 38863 92973
rect 231445 92970 231511 92973
rect 35902 92968 38863 92970
rect 35902 92912 38802 92968
rect 38858 92912 38863 92968
rect 35902 92910 38863 92912
rect 35902 92902 35962 92910
rect 38797 92907 38863 92910
rect 228734 92968 231511 92970
rect 228734 92912 231450 92968
rect 231506 92912 231511 92968
rect 228734 92910 231511 92912
rect 35748 92842 35962 92902
rect 137789 92698 137855 92701
rect 134710 92696 137855 92698
rect 134710 92640 137794 92696
rect 137850 92640 137855 92696
rect 134710 92638 137855 92640
rect 134710 92328 134770 92638
rect 137789 92635 137855 92638
rect 145241 92426 145307 92429
rect 145241 92424 148938 92426
rect 145241 92368 145246 92424
rect 145302 92368 148938 92424
rect 145241 92366 148938 92368
rect 145241 92363 145307 92366
rect 148878 92260 148938 92366
rect 228734 92328 228794 92910
rect 231445 92907 231511 92910
rect 240921 92290 240987 92293
rect 240921 92288 242932 92290
rect 240921 92232 240926 92288
rect 240982 92232 242932 92288
rect 240921 92230 242932 92232
rect 240921 92227 240987 92230
rect 137605 91474 137671 91477
rect 231445 91474 231511 91477
rect 134710 91472 137671 91474
rect 134710 91416 137610 91472
rect 137666 91416 137671 91472
rect 134710 91414 137671 91416
rect 134710 90832 134770 91414
rect 137605 91411 137671 91414
rect 228734 91472 231511 91474
rect 228734 91416 231450 91472
rect 231506 91416 231511 91472
rect 228734 91414 231511 91416
rect 228734 90832 228794 91414
rect 231445 91411 231511 91414
rect 9896 90522 10376 90552
rect 13773 90522 13839 90525
rect 9896 90520 13839 90522
rect 9896 90464 13778 90520
rect 13834 90464 13839 90520
rect 9896 90462 13839 90464
rect 9896 90432 10376 90462
rect 13773 90459 13839 90462
rect 240921 89978 240987 89981
rect 240921 89976 242932 89978
rect 145241 89434 145307 89437
rect 149062 89434 149122 89948
rect 240921 89920 240926 89976
rect 240982 89920 242932 89976
rect 240921 89918 242932 89920
rect 240921 89915 240987 89918
rect 231629 89842 231695 89845
rect 145241 89432 149122 89434
rect 145241 89376 145246 89432
rect 145302 89376 149122 89432
rect 145241 89374 149122 89376
rect 228734 89840 231695 89842
rect 228734 89784 231634 89840
rect 231690 89784 231695 89840
rect 228734 89782 231695 89784
rect 145241 89371 145307 89374
rect 228734 89200 228794 89782
rect 231629 89779 231695 89782
rect 134710 89162 134770 89196
rect 138157 89162 138223 89165
rect 134710 89160 138223 89162
rect 134710 89104 138162 89160
rect 138218 89104 138223 89160
rect 134710 89102 138223 89104
rect 138157 89099 138223 89102
rect 231629 88346 231695 88349
rect 228734 88344 231695 88346
rect 228734 88288 231634 88344
rect 231690 88288 231695 88344
rect 228734 88286 231695 88288
rect 137605 88210 137671 88213
rect 134710 88208 137671 88210
rect 134710 88152 137610 88208
rect 137666 88152 137671 88208
rect 134710 88150 137671 88152
rect 134710 87704 134770 88150
rect 137605 88147 137671 88150
rect 228734 87704 228794 88286
rect 231629 88283 231695 88286
rect 241606 87332 241612 87396
rect 241676 87394 241682 87396
rect 285909 87394 285975 87397
rect 241676 87392 285975 87394
rect 241676 87336 285914 87392
rect 285970 87336 285975 87392
rect 241676 87334 285975 87336
rect 241676 87332 241682 87334
rect 285909 87331 285975 87334
rect 251409 86442 251475 86445
rect 256561 86442 256627 86445
rect 251409 86440 256627 86442
rect 251409 86384 251414 86440
rect 251470 86384 256566 86440
rect 256622 86384 256627 86440
rect 251409 86382 256627 86384
rect 251409 86379 251475 86382
rect 256561 86379 256627 86382
rect 134710 85626 134770 86068
rect 228734 86034 228794 86068
rect 231629 86034 231695 86037
rect 228734 86032 231695 86034
rect 228734 85976 231634 86032
rect 231690 85976 231695 86032
rect 228734 85974 231695 85976
rect 231629 85971 231695 85974
rect 136869 85626 136935 85629
rect 134710 85624 136935 85626
rect 134710 85568 136874 85624
rect 136930 85568 136935 85624
rect 134710 85566 136935 85568
rect 136869 85563 136935 85566
rect 136869 84674 136935 84677
rect 231629 84674 231695 84677
rect 134710 84672 136935 84674
rect 134710 84616 136874 84672
rect 136930 84616 136935 84672
rect 134710 84614 136935 84616
rect 134710 84576 134770 84614
rect 136869 84611 136935 84614
rect 228734 84672 231695 84674
rect 228734 84616 231634 84672
rect 231690 84616 231695 84672
rect 228734 84614 231695 84616
rect 228734 84576 228794 84614
rect 231629 84611 231695 84614
rect 85022 84068 85028 84132
rect 85092 84130 85098 84132
rect 85165 84130 85231 84133
rect 85092 84128 85231 84130
rect 85092 84072 85170 84128
rect 85226 84072 85231 84128
rect 85092 84070 85231 84072
rect 85092 84068 85098 84070
rect 85165 84067 85231 84070
rect 133230 83660 133236 83724
rect 133300 83722 133306 83724
rect 133373 83722 133439 83725
rect 133300 83720 133439 83722
rect 133300 83664 133378 83720
rect 133434 83664 133439 83720
rect 133300 83662 133439 83664
rect 133300 83660 133306 83662
rect 133373 83659 133439 83662
rect 182133 83724 182199 83725
rect 182133 83720 182180 83724
rect 182244 83722 182250 83724
rect 182133 83664 182138 83720
rect 182133 83660 182180 83664
rect 182244 83662 182290 83722
rect 182244 83660 182250 83662
rect 182133 83659 182199 83660
rect 210561 81410 210627 81413
rect 237006 81410 237012 81412
rect 210561 81408 237012 81410
rect 210561 81352 210566 81408
rect 210622 81352 237012 81408
rect 210561 81350 237012 81352
rect 210561 81347 210627 81350
rect 237006 81348 237012 81350
rect 237076 81348 237082 81412
rect 125553 81274 125619 81277
rect 144270 81274 144276 81276
rect 125553 81272 144276 81274
rect 125553 81216 125558 81272
rect 125614 81216 144276 81272
rect 125553 81214 144276 81216
rect 125553 81211 125619 81214
rect 144270 81212 144276 81214
rect 144340 81212 144346 81276
rect 202465 81274 202531 81277
rect 236822 81274 236828 81276
rect 202465 81272 236828 81274
rect 202465 81216 202470 81272
rect 202526 81216 236828 81272
rect 202465 81214 236828 81216
rect 202465 81211 202531 81214
rect 236822 81212 236828 81214
rect 236892 81212 236898 81276
rect 156005 79370 156071 79373
rect 155502 79368 156071 79370
rect 155502 79312 156010 79368
rect 156066 79312 156071 79368
rect 155502 79310 156071 79312
rect 155361 79234 155427 79237
rect 155502 79234 155562 79310
rect 156005 79307 156071 79310
rect 155361 79232 155562 79234
rect 155361 79176 155366 79232
rect 155422 79176 155562 79232
rect 155361 79174 155562 79176
rect 155361 79171 155427 79174
rect 248557 78962 248623 78965
rect 259781 78962 259847 78965
rect 248557 78960 259847 78962
rect 248557 78904 248562 78960
rect 248618 78904 259786 78960
rect 259842 78904 259847 78960
rect 248557 78902 259847 78904
rect 248557 78899 248623 78902
rect 259781 78899 259847 78902
rect 60785 78826 60851 78829
rect 72469 78826 72535 78829
rect 60785 78824 72535 78826
rect 60785 78768 60790 78824
rect 60846 78768 72474 78824
rect 72530 78768 72535 78824
rect 60785 78766 72535 78768
rect 60785 78763 60851 78766
rect 72469 78763 72535 78766
rect 249845 78826 249911 78829
rect 261069 78826 261135 78829
rect 249845 78824 261135 78826
rect 249845 78768 249850 78824
rect 249906 78768 261074 78824
rect 261130 78768 261135 78824
rect 249845 78766 261135 78768
rect 249845 78763 249911 78766
rect 261069 78763 261135 78766
rect 61521 78690 61587 78693
rect 73757 78690 73823 78693
rect 61521 78688 73823 78690
rect 61521 78632 61526 78688
rect 61582 78632 73762 78688
rect 73818 78632 73823 78688
rect 61521 78630 73823 78632
rect 61521 78627 61587 78630
rect 73757 78627 73823 78630
rect 155269 78690 155335 78693
rect 167321 78690 167387 78693
rect 155269 78688 167387 78690
rect 155269 78632 155274 78688
rect 155330 78632 167326 78688
rect 167382 78632 167387 78688
rect 155269 78630 167387 78632
rect 155269 78627 155335 78630
rect 167321 78627 167387 78630
rect 247085 78690 247151 78693
rect 258309 78690 258375 78693
rect 247085 78688 258375 78690
rect 247085 78632 247090 78688
rect 247146 78632 258314 78688
rect 258370 78632 258375 78688
rect 247085 78630 258375 78632
rect 247085 78627 247151 78630
rect 258309 78627 258375 78630
rect 62073 78554 62139 78557
rect 74493 78554 74559 78557
rect 62073 78552 74559 78554
rect 62073 78496 62078 78552
rect 62134 78496 74498 78552
rect 74554 78496 74559 78552
rect 62073 78494 74559 78496
rect 62073 78491 62139 78494
rect 74493 78491 74559 78494
rect 134845 78554 134911 78557
rect 170081 78554 170147 78557
rect 134845 78552 170147 78554
rect 134845 78496 134850 78552
rect 134906 78496 170086 78552
rect 170142 78496 170147 78552
rect 134845 78494 170147 78496
rect 134845 78491 134911 78494
rect 170081 78491 170147 78494
rect 249661 78554 249727 78557
rect 261437 78554 261503 78557
rect 249661 78552 261503 78554
rect 249661 78496 249666 78552
rect 249722 78496 261442 78552
rect 261498 78496 261503 78552
rect 249661 78494 261503 78496
rect 249661 78491 249727 78494
rect 261437 78491 261503 78494
rect 62165 78418 62231 78421
rect 75137 78418 75203 78421
rect 62165 78416 75203 78418
rect 62165 78360 62170 78416
rect 62226 78360 75142 78416
rect 75198 78360 75203 78416
rect 62165 78358 75203 78360
rect 62165 78355 62231 78358
rect 75137 78355 75203 78358
rect 112949 78418 113015 78421
rect 169069 78418 169135 78421
rect 112949 78416 169135 78418
rect 112949 78360 112954 78416
rect 113010 78360 169074 78416
rect 169130 78360 169135 78416
rect 112949 78358 169135 78360
rect 112949 78355 113015 78358
rect 169069 78355 169135 78358
rect 249109 78418 249175 78421
rect 261989 78418 262055 78421
rect 249109 78416 262055 78418
rect 249109 78360 249114 78416
rect 249170 78360 261994 78416
rect 262050 78360 262055 78416
rect 249109 78358 262055 78360
rect 249109 78355 249175 78358
rect 261989 78355 262055 78358
rect 103974 77812 103980 77876
rect 104044 77874 104050 77876
rect 168609 77874 168675 77877
rect 104044 77872 168675 77874
rect 104044 77816 168614 77872
rect 168670 77816 168675 77872
rect 104044 77814 168675 77816
rect 104044 77812 104050 77814
rect 168609 77811 168675 77814
rect 169989 76106 170055 76109
rect 169989 76104 170650 76106
rect 169989 76048 169994 76104
rect 170050 76048 170650 76104
rect 169989 76046 170650 76048
rect 169989 76043 170055 76046
rect 80197 75562 80263 75565
rect 76780 75560 80263 75562
rect 76780 75504 80202 75560
rect 80258 75504 80263 75560
rect 76780 75502 80263 75504
rect 80197 75499 80263 75502
rect 139629 75562 139695 75565
rect 139629 75560 143020 75562
rect 139629 75504 139634 75560
rect 139690 75504 143020 75560
rect 170590 75532 170650 76046
rect 233469 75562 233535 75565
rect 233469 75560 237044 75562
rect 139629 75502 143020 75504
rect 233469 75504 233474 75560
rect 233530 75504 237044 75560
rect 233469 75502 237044 75504
rect 139629 75499 139695 75502
rect 233469 75499 233535 75502
rect 80105 75018 80171 75021
rect 76780 75016 80171 75018
rect 76780 74960 80110 75016
rect 80166 74960 80171 75016
rect 233469 75018 233535 75021
rect 233469 75016 237044 75018
rect 76780 74958 80171 74960
rect 80105 74955 80171 74958
rect 140917 74882 140983 74885
rect 140917 74880 143020 74882
rect 140917 74824 140922 74880
rect 140978 74824 143020 74880
rect 140917 74822 143020 74824
rect 140917 74819 140983 74822
rect 170590 74749 170650 74988
rect 233469 74960 233474 75016
rect 233530 74960 237044 75016
rect 233469 74958 237044 74960
rect 233469 74955 233535 74958
rect 170590 74744 170699 74749
rect 170817 74746 170883 74749
rect 170590 74688 170638 74744
rect 170694 74688 170699 74744
rect 170590 74686 170699 74688
rect 170633 74683 170699 74686
rect 170774 74744 170883 74746
rect 170774 74688 170822 74744
rect 170878 74688 170883 74744
rect 170774 74683 170883 74688
rect 80013 74474 80079 74477
rect 76780 74472 80079 74474
rect 76780 74416 80018 74472
rect 80074 74416 80079 74472
rect 170774 74444 170834 74683
rect 76780 74414 80079 74416
rect 80013 74411 80079 74414
rect 233561 74338 233627 74341
rect 233561 74336 237044 74338
rect 233561 74280 233566 74336
rect 233622 74280 237044 74336
rect 233561 74278 237044 74280
rect 233561 74275 233627 74278
rect 139629 74202 139695 74205
rect 170725 74202 170791 74205
rect 139629 74200 143020 74202
rect 139629 74144 139634 74200
rect 139690 74144 143020 74200
rect 139629 74142 143020 74144
rect 170725 74200 170834 74202
rect 170725 74144 170730 74200
rect 170786 74144 170834 74200
rect 139629 74139 139695 74142
rect 170725 74139 170834 74144
rect 79921 73930 79987 73933
rect 76780 73928 79987 73930
rect 76780 73872 79926 73928
rect 79982 73872 79987 73928
rect 170774 73900 170834 74139
rect 76780 73870 79987 73872
rect 79921 73867 79987 73870
rect 233653 73794 233719 73797
rect 233653 73792 237044 73794
rect 233653 73736 233658 73792
rect 233714 73736 237044 73792
rect 233653 73734 237044 73736
rect 233653 73731 233719 73734
rect 139721 73522 139787 73525
rect 139721 73520 143020 73522
rect 139721 73464 139726 73520
rect 139782 73464 143020 73520
rect 139721 73462 143020 73464
rect 139721 73459 139787 73462
rect 173301 73386 173367 73389
rect 170804 73384 173367 73386
rect 170804 73328 173306 73384
rect 173362 73328 173367 73384
rect 170804 73326 173367 73328
rect 173301 73323 173367 73326
rect 79645 73250 79711 73253
rect 76780 73248 79711 73250
rect 76780 73192 79650 73248
rect 79706 73192 79711 73248
rect 76780 73190 79711 73192
rect 79645 73187 79711 73190
rect 139629 72978 139695 72981
rect 139629 72976 143020 72978
rect 139629 72920 139634 72976
rect 139690 72920 143020 72976
rect 139629 72918 143020 72920
rect 139629 72915 139695 72918
rect 173945 72842 174011 72845
rect 170804 72840 174011 72842
rect 170804 72784 173950 72840
rect 174006 72784 174011 72840
rect 170804 72782 174011 72784
rect 173945 72779 174011 72782
rect 79829 72706 79895 72709
rect 76780 72704 79895 72706
rect 76780 72648 79834 72704
rect 79890 72648 79895 72704
rect 76780 72646 79895 72648
rect 79829 72643 79895 72646
rect 234113 72706 234179 72709
rect 237014 72706 237074 73016
rect 234113 72704 237074 72706
rect 234113 72648 234118 72704
rect 234174 72648 237074 72704
rect 234113 72646 237074 72648
rect 234113 72643 234179 72646
rect 233469 72570 233535 72573
rect 233469 72568 237044 72570
rect 233469 72512 233474 72568
rect 233530 72512 237044 72568
rect 233469 72510 237044 72512
rect 233469 72507 233535 72510
rect 139629 72298 139695 72301
rect 173669 72298 173735 72301
rect 139629 72296 143020 72298
rect 139629 72240 139634 72296
rect 139690 72240 143020 72296
rect 139629 72238 143020 72240
rect 170804 72296 173735 72298
rect 170804 72240 173674 72296
rect 173730 72240 173735 72296
rect 170804 72238 173735 72240
rect 139629 72235 139695 72238
rect 173669 72235 173735 72238
rect 79737 72162 79803 72165
rect 76780 72160 79803 72162
rect 76780 72104 79742 72160
rect 79798 72104 79803 72160
rect 76780 72102 79803 72104
rect 79737 72099 79803 72102
rect 173853 71754 173919 71757
rect 170804 71752 173919 71754
rect 170804 71696 173858 71752
rect 173914 71696 173919 71752
rect 170804 71694 173919 71696
rect 173853 71691 173919 71694
rect 79553 71618 79619 71621
rect 76780 71616 79619 71618
rect 76780 71560 79558 71616
rect 79614 71560 79619 71616
rect 76780 71558 79619 71560
rect 79553 71555 79619 71558
rect 139905 71618 139971 71621
rect 139905 71616 143020 71618
rect 139905 71560 139910 71616
rect 139966 71560 143020 71616
rect 139905 71558 143020 71560
rect 139905 71555 139971 71558
rect 233561 71482 233627 71485
rect 237014 71482 237074 71792
rect 233561 71480 237074 71482
rect 233561 71424 233566 71480
rect 233622 71424 237074 71480
rect 233561 71422 237074 71424
rect 233561 71419 233627 71422
rect 173485 71346 173551 71349
rect 170804 71344 173551 71346
rect 170804 71288 173490 71344
rect 173546 71288 173551 71344
rect 170804 71286 173551 71288
rect 173485 71283 173551 71286
rect 80197 71074 80263 71077
rect 76780 71072 80263 71074
rect 76780 71016 80202 71072
rect 80258 71016 80263 71072
rect 76780 71014 80263 71016
rect 80197 71011 80263 71014
rect 233469 71074 233535 71077
rect 237014 71074 237074 71248
rect 233469 71072 237074 71074
rect 233469 71016 233474 71072
rect 233530 71016 237074 71072
rect 233469 71014 237074 71016
rect 233469 71011 233535 71014
rect 139813 70938 139879 70941
rect 139813 70936 143020 70938
rect 139813 70880 139818 70936
rect 139874 70880 143020 70936
rect 139813 70878 143020 70880
rect 139813 70875 139879 70878
rect 173761 70802 173827 70805
rect 170804 70800 173827 70802
rect 170804 70744 173766 70800
rect 173822 70744 173827 70800
rect 170804 70742 173827 70744
rect 173761 70739 173827 70742
rect 76750 69986 76810 70296
rect 139721 70258 139787 70261
rect 173577 70258 173643 70261
rect 139721 70256 143020 70258
rect 139721 70200 139726 70256
rect 139782 70200 143020 70256
rect 139721 70198 143020 70200
rect 170804 70256 173643 70258
rect 170804 70200 173582 70256
rect 173638 70200 173643 70256
rect 170804 70198 173643 70200
rect 139721 70195 139787 70198
rect 173577 70195 173643 70198
rect 233653 70258 233719 70261
rect 237014 70258 237074 70568
rect 233653 70256 237074 70258
rect 233653 70200 233658 70256
rect 233714 70200 237074 70256
rect 233653 70198 237074 70200
rect 233653 70195 233719 70198
rect 300169 70122 300235 70125
rect 303416 70122 303896 70152
rect 300169 70120 303896 70122
rect 300169 70064 300174 70120
rect 300230 70064 303896 70120
rect 300169 70062 303896 70064
rect 300169 70059 300235 70062
rect 303416 70032 303896 70062
rect 79461 69986 79527 69989
rect 76750 69984 79527 69986
rect 76750 69928 79466 69984
rect 79522 69928 79527 69984
rect 76750 69926 79527 69928
rect 79461 69923 79527 69926
rect 80197 69850 80263 69853
rect 76780 69848 80263 69850
rect 76780 69792 80202 69848
rect 80258 69792 80263 69848
rect 76780 69790 80263 69792
rect 80197 69787 80263 69790
rect 87189 69714 87255 69717
rect 131349 69714 131415 69717
rect 87189 69712 90028 69714
rect 87189 69656 87194 69712
rect 87250 69656 90028 69712
rect 87189 69654 90028 69656
rect 129772 69712 131415 69714
rect 129772 69656 131354 69712
rect 131410 69656 131415 69712
rect 129772 69654 131415 69656
rect 87189 69651 87255 69654
rect 131349 69651 131415 69654
rect 139629 69714 139695 69717
rect 174037 69714 174103 69717
rect 139629 69712 143020 69714
rect 139629 69656 139634 69712
rect 139690 69656 143020 69712
rect 139629 69654 143020 69656
rect 170804 69712 174103 69714
rect 170804 69656 174042 69712
rect 174098 69656 174103 69712
rect 170804 69654 174103 69656
rect 139629 69651 139695 69654
rect 174037 69651 174103 69654
rect 181765 69714 181831 69717
rect 226017 69714 226083 69717
rect 181765 69712 184052 69714
rect 181765 69656 181770 69712
rect 181826 69656 184052 69712
rect 181765 69654 184052 69656
rect 223796 69712 226083 69714
rect 223796 69656 226022 69712
rect 226078 69656 226083 69712
rect 223796 69654 226083 69656
rect 181765 69651 181831 69654
rect 226017 69651 226083 69654
rect 233745 69578 233811 69581
rect 237014 69578 237074 70024
rect 233745 69576 237074 69578
rect 233745 69520 233750 69576
rect 233806 69520 237074 69576
rect 233745 69518 237074 69520
rect 233745 69515 233811 69518
rect 264841 69442 264907 69445
rect 264798 69440 264907 69442
rect 264798 69384 264846 69440
rect 264902 69384 264907 69440
rect 264798 69379 264907 69384
rect 87189 69306 87255 69309
rect 131349 69306 131415 69309
rect 226017 69306 226083 69309
rect 87189 69304 90028 69306
rect 87189 69248 87194 69304
rect 87250 69248 90028 69304
rect 87189 69246 90028 69248
rect 129772 69304 131415 69306
rect 129772 69248 131354 69304
rect 131410 69248 131415 69304
rect 129772 69246 131415 69248
rect 223796 69304 226083 69306
rect 223796 69248 226022 69304
rect 226078 69248 226083 69304
rect 223796 69246 226083 69248
rect 87189 69243 87255 69246
rect 131349 69243 131415 69246
rect 226017 69243 226083 69246
rect 76750 69034 76810 69208
rect 173301 69170 173367 69173
rect 170804 69168 173367 69170
rect 170804 69112 173306 69168
rect 173362 69112 173367 69168
rect 170804 69110 173367 69112
rect 173301 69107 173367 69110
rect 80197 69034 80263 69037
rect 76750 69032 80263 69034
rect 76750 68976 80202 69032
rect 80258 68976 80263 69032
rect 76750 68974 80263 68976
rect 80197 68971 80263 68974
rect 139721 69034 139787 69037
rect 182317 69034 182383 69037
rect 184022 69034 184082 69208
rect 139721 69032 143020 69034
rect 139721 68976 139726 69032
rect 139782 68976 143020 69032
rect 139721 68974 143020 68976
rect 182317 69032 184082 69034
rect 182317 68976 182322 69032
rect 182378 68976 184082 69032
rect 182317 68974 184082 68976
rect 233653 69034 233719 69037
rect 237014 69034 237074 69344
rect 233653 69032 237074 69034
rect 233653 68976 233658 69032
rect 233714 68976 237074 69032
rect 233653 68974 237074 68976
rect 139721 68971 139787 68974
rect 182317 68971 182383 68974
rect 233653 68971 233719 68974
rect 87281 68898 87347 68901
rect 131441 68898 131507 68901
rect 225741 68898 225807 68901
rect 87281 68896 90028 68898
rect 87281 68840 87286 68896
rect 87342 68840 90028 68896
rect 87281 68838 90028 68840
rect 129772 68896 131507 68898
rect 129772 68840 131446 68896
rect 131502 68840 131507 68896
rect 129772 68838 131507 68840
rect 223796 68896 225807 68898
rect 223796 68840 225746 68896
rect 225802 68840 225807 68896
rect 264798 68868 264858 69379
rect 223796 68838 225807 68840
rect 87281 68835 87347 68838
rect 131441 68835 131507 68838
rect 225741 68835 225807 68838
rect 76750 68490 76810 68664
rect 172841 68626 172907 68629
rect 170804 68624 172907 68626
rect 170804 68568 172846 68624
rect 172902 68568 172907 68624
rect 170804 68566 172907 68568
rect 172841 68563 172907 68566
rect 181765 68626 181831 68629
rect 184022 68626 184082 68800
rect 181765 68624 184082 68626
rect 181765 68568 181770 68624
rect 181826 68568 184082 68624
rect 181765 68566 184082 68568
rect 181765 68563 181831 68566
rect 80105 68490 80171 68493
rect 76750 68488 80171 68490
rect 76750 68432 80110 68488
rect 80166 68432 80171 68488
rect 76750 68430 80171 68432
rect 80105 68427 80171 68430
rect 87189 68490 87255 68493
rect 131533 68490 131599 68493
rect 226293 68490 226359 68493
rect 87189 68488 90028 68490
rect 87189 68432 87194 68488
rect 87250 68432 90028 68488
rect 87189 68430 90028 68432
rect 129772 68488 131599 68490
rect 129772 68432 131538 68488
rect 131594 68432 131599 68488
rect 129772 68430 131599 68432
rect 223796 68488 226359 68490
rect 223796 68432 226298 68488
rect 226354 68432 226359 68488
rect 223796 68430 226359 68432
rect 87189 68427 87255 68430
rect 131533 68427 131599 68430
rect 226293 68427 226359 68430
rect 139629 68354 139695 68357
rect 139629 68352 143020 68354
rect 139629 68296 139634 68352
rect 139690 68296 143020 68352
rect 139629 68294 143020 68296
rect 139629 68291 139695 68294
rect 80197 68218 80263 68221
rect 76780 68216 80263 68218
rect 76780 68160 80202 68216
rect 80258 68160 80263 68216
rect 76780 68158 80263 68160
rect 80197 68155 80263 68158
rect 181581 68218 181647 68221
rect 184022 68218 184082 68392
rect 233561 68354 233627 68357
rect 237014 68354 237074 68800
rect 233561 68352 237074 68354
rect 233561 68296 233566 68352
rect 233622 68296 237074 68352
rect 233561 68294 237074 68296
rect 233561 68291 233627 68294
rect 181581 68216 184082 68218
rect 181581 68160 181586 68216
rect 181642 68160 184082 68216
rect 181581 68158 184082 68160
rect 233469 68218 233535 68221
rect 233469 68216 237044 68218
rect 233469 68160 233474 68216
rect 233530 68160 237044 68216
rect 233469 68158 237044 68160
rect 181581 68155 181647 68158
rect 233469 68155 233535 68158
rect 87189 68082 87255 68085
rect 131993 68082 132059 68085
rect 174037 68082 174103 68085
rect 226293 68082 226359 68085
rect 87189 68080 90028 68082
rect 87189 68024 87194 68080
rect 87250 68024 90028 68080
rect 87189 68022 90028 68024
rect 129772 68080 132059 68082
rect 129772 68024 131998 68080
rect 132054 68024 132059 68080
rect 129772 68022 132059 68024
rect 170804 68080 174103 68082
rect 170804 68024 174042 68080
rect 174098 68024 174103 68080
rect 170804 68022 174103 68024
rect 223796 68080 226359 68082
rect 223796 68024 226298 68080
rect 226354 68024 226359 68080
rect 223796 68022 226359 68024
rect 87189 68019 87255 68022
rect 131993 68019 132059 68022
rect 174037 68019 174103 68022
rect 226293 68019 226359 68022
rect 182317 67810 182383 67813
rect 184022 67810 184082 67984
rect 182317 67808 184082 67810
rect 182317 67752 182322 67808
rect 182378 67752 184082 67808
rect 182317 67750 184082 67752
rect 182317 67747 182383 67750
rect 87281 67674 87347 67677
rect 132545 67674 132611 67677
rect 87281 67672 90028 67674
rect 87281 67616 87286 67672
rect 87342 67616 90028 67672
rect 87281 67614 90028 67616
rect 129772 67672 132611 67674
rect 129772 67616 132550 67672
rect 132606 67616 132611 67672
rect 129772 67614 132611 67616
rect 87281 67611 87347 67614
rect 132545 67611 132611 67614
rect 139629 67674 139695 67677
rect 225557 67674 225623 67677
rect 139629 67672 143020 67674
rect 139629 67616 139634 67672
rect 139690 67616 143020 67672
rect 139629 67614 143020 67616
rect 223796 67672 225623 67674
rect 223796 67616 225562 67672
rect 225618 67616 225623 67672
rect 223796 67614 225623 67616
rect 139629 67611 139695 67614
rect 225557 67611 225623 67614
rect 80197 67538 80263 67541
rect 173945 67538 174011 67541
rect 76780 67536 80263 67538
rect 76780 67480 80202 67536
rect 80258 67480 80263 67536
rect 76780 67478 80263 67480
rect 170804 67536 174011 67538
rect 170804 67480 173950 67536
rect 174006 67480 174011 67536
rect 170804 67478 174011 67480
rect 80197 67475 80263 67478
rect 173945 67475 174011 67478
rect 182225 67402 182291 67405
rect 184022 67402 184082 67576
rect 182225 67400 184082 67402
rect 182225 67344 182230 67400
rect 182286 67344 184082 67400
rect 182225 67342 184082 67344
rect 182225 67339 182291 67342
rect 87189 67266 87255 67269
rect 131809 67266 131875 67269
rect 225465 67266 225531 67269
rect 87189 67264 90028 67266
rect 87189 67208 87194 67264
rect 87250 67208 90028 67264
rect 87189 67206 90028 67208
rect 129772 67264 131875 67266
rect 129772 67208 131814 67264
rect 131870 67208 131875 67264
rect 129772 67206 131875 67208
rect 223796 67264 225531 67266
rect 223796 67208 225470 67264
rect 225526 67208 225531 67264
rect 223796 67206 225531 67208
rect 87189 67203 87255 67206
rect 131809 67203 131875 67206
rect 225465 67203 225531 67206
rect 80105 66994 80171 66997
rect 76780 66992 80171 66994
rect 76780 66936 80110 66992
rect 80166 66936 80171 66992
rect 76780 66934 80171 66936
rect 80105 66931 80171 66934
rect 139721 66994 139787 66997
rect 173485 66994 173551 66997
rect 139721 66992 143020 66994
rect 139721 66936 139726 66992
rect 139782 66936 143020 66992
rect 139721 66934 143020 66936
rect 170804 66992 173551 66994
rect 170804 66936 173490 66992
rect 173546 66936 173551 66992
rect 170804 66934 173551 66936
rect 139721 66931 139787 66934
rect 173485 66931 173551 66934
rect 182317 66994 182383 66997
rect 184022 66994 184082 67168
rect 233561 67130 233627 67133
rect 237014 67130 237074 67576
rect 233561 67128 237074 67130
rect 233561 67072 233566 67128
rect 233622 67072 237074 67128
rect 233561 67070 237074 67072
rect 233561 67067 233627 67070
rect 182317 66992 184082 66994
rect 182317 66936 182322 66992
rect 182378 66936 184082 66992
rect 182317 66934 184082 66936
rect 233469 66994 233535 66997
rect 233469 66992 237044 66994
rect 233469 66936 233474 66992
rect 233530 66936 237044 66992
rect 233469 66934 237044 66936
rect 182317 66931 182383 66934
rect 233469 66931 233535 66934
rect 87281 66858 87347 66861
rect 131349 66858 131415 66861
rect 87281 66856 90028 66858
rect 87281 66800 87286 66856
rect 87342 66800 90028 66856
rect 87281 66798 90028 66800
rect 129772 66856 131415 66858
rect 129772 66800 131354 66856
rect 131410 66800 131415 66856
rect 129772 66798 131415 66800
rect 87281 66795 87347 66798
rect 131349 66795 131415 66798
rect 181397 66858 181463 66861
rect 225833 66858 225899 66861
rect 181397 66856 184052 66858
rect 181397 66800 181402 66856
rect 181458 66800 184052 66856
rect 181397 66798 184052 66800
rect 223796 66856 225899 66858
rect 223796 66800 225838 66856
rect 225894 66800 225899 66856
rect 223796 66798 225899 66800
rect 181397 66795 181463 66798
rect 225833 66795 225899 66798
rect 174037 66586 174103 66589
rect 170804 66584 174103 66586
rect 170804 66528 174042 66584
rect 174098 66528 174103 66584
rect 170804 66526 174103 66528
rect 174037 66523 174103 66526
rect 80105 66450 80171 66453
rect 131349 66450 131415 66453
rect 76780 66448 80171 66450
rect 76780 66392 80110 66448
rect 80166 66392 80171 66448
rect 76780 66390 80171 66392
rect 129772 66448 131415 66450
rect 129772 66392 131354 66448
rect 131410 66392 131415 66448
rect 129772 66390 131415 66392
rect 80105 66387 80171 66390
rect 131349 66387 131415 66390
rect 139721 66450 139787 66453
rect 226017 66450 226083 66453
rect 139721 66448 143020 66450
rect 139721 66392 139726 66448
rect 139782 66392 143020 66448
rect 139721 66390 143020 66392
rect 223796 66448 226083 66450
rect 223796 66392 226022 66448
rect 226078 66392 226083 66448
rect 223796 66390 226083 66392
rect 139721 66387 139787 66390
rect 226017 66387 226083 66390
rect 87281 66178 87347 66181
rect 89998 66178 90058 66352
rect 87281 66176 90058 66178
rect 87281 66120 87286 66176
rect 87342 66120 90058 66176
rect 87281 66118 90058 66120
rect 182317 66178 182383 66181
rect 184022 66178 184082 66352
rect 182317 66176 184082 66178
rect 182317 66120 182322 66176
rect 182378 66120 184082 66176
rect 182317 66118 184082 66120
rect 233469 66178 233535 66181
rect 237014 66178 237074 66352
rect 233469 66176 237074 66178
rect 233469 66120 233474 66176
rect 233530 66120 237074 66176
rect 233469 66118 237074 66120
rect 87281 66115 87347 66118
rect 182317 66115 182383 66118
rect 233469 66115 233535 66118
rect 87189 66042 87255 66045
rect 132177 66042 132243 66045
rect 173577 66042 173643 66045
rect 226293 66042 226359 66045
rect 87189 66040 90028 66042
rect 87189 65984 87194 66040
rect 87250 65984 90028 66040
rect 87189 65982 90028 65984
rect 129772 66040 132243 66042
rect 129772 65984 132182 66040
rect 132238 65984 132243 66040
rect 129772 65982 132243 65984
rect 170804 66040 173643 66042
rect 170804 65984 173582 66040
rect 173638 65984 173643 66040
rect 170804 65982 173643 65984
rect 223796 66040 226359 66042
rect 223796 65984 226298 66040
rect 226354 65984 226359 66040
rect 223796 65982 226359 65984
rect 87189 65979 87255 65982
rect 132177 65979 132243 65982
rect 173577 65979 173643 65982
rect 226293 65979 226359 65982
rect 80197 65906 80263 65909
rect 76780 65904 80263 65906
rect 76780 65848 80202 65904
rect 80258 65848 80263 65904
rect 76780 65846 80263 65848
rect 80197 65843 80263 65846
rect 139629 65770 139695 65773
rect 181397 65770 181463 65773
rect 184022 65770 184082 65944
rect 139629 65768 143020 65770
rect 139629 65712 139634 65768
rect 139690 65712 143020 65768
rect 139629 65710 143020 65712
rect 181397 65768 184082 65770
rect 181397 65712 181402 65768
rect 181458 65712 184082 65768
rect 181397 65710 184082 65712
rect 139629 65707 139695 65710
rect 181397 65707 181463 65710
rect 87189 65634 87255 65637
rect 131349 65634 131415 65637
rect 87189 65632 90028 65634
rect 87189 65576 87194 65632
rect 87250 65576 90028 65632
rect 87189 65574 90028 65576
rect 129772 65632 131415 65634
rect 129772 65576 131354 65632
rect 131410 65576 131415 65632
rect 129772 65574 131415 65576
rect 87189 65571 87255 65574
rect 131349 65571 131415 65574
rect 181305 65634 181371 65637
rect 226385 65634 226451 65637
rect 181305 65632 184052 65634
rect 181305 65576 181310 65632
rect 181366 65576 184052 65632
rect 181305 65574 184052 65576
rect 223796 65632 226451 65634
rect 223796 65576 226390 65632
rect 226446 65576 226451 65632
rect 223796 65574 226451 65576
rect 181305 65571 181371 65574
rect 226385 65571 226451 65574
rect 173853 65498 173919 65501
rect 170804 65496 173919 65498
rect 170804 65440 173858 65496
rect 173914 65440 173919 65496
rect 170804 65438 173919 65440
rect 173853 65435 173919 65438
rect 233469 65498 233535 65501
rect 237014 65498 237074 65672
rect 233469 65496 237074 65498
rect 233469 65440 233474 65496
rect 233530 65440 237074 65496
rect 233469 65438 237074 65440
rect 233469 65435 233535 65438
rect 80197 65362 80263 65365
rect 76780 65360 80263 65362
rect 76780 65304 80202 65360
rect 80258 65304 80263 65360
rect 76780 65302 80263 65304
rect 80197 65299 80263 65302
rect 131349 65226 131415 65229
rect 226293 65226 226359 65229
rect 129772 65224 131415 65226
rect 129772 65168 131354 65224
rect 131410 65168 131415 65224
rect 129772 65166 131415 65168
rect 223796 65224 226359 65226
rect 223796 65168 226298 65224
rect 226354 65168 226359 65224
rect 223796 65166 226359 65168
rect 131349 65163 131415 65166
rect 226293 65163 226359 65166
rect 87281 64954 87347 64957
rect 89998 64954 90058 65128
rect 139721 65090 139787 65093
rect 139721 65088 143020 65090
rect 139721 65032 139726 65088
rect 139782 65032 143020 65088
rect 139721 65030 143020 65032
rect 139721 65027 139787 65030
rect 173485 64954 173551 64957
rect 87281 64952 90058 64954
rect 87281 64896 87286 64952
rect 87342 64896 90058 64952
rect 87281 64894 90058 64896
rect 170804 64952 173551 64954
rect 170804 64896 173490 64952
rect 173546 64896 173551 64952
rect 170804 64894 173551 64896
rect 87281 64891 87347 64894
rect 173485 64891 173551 64894
rect 181029 64954 181095 64957
rect 184022 64954 184082 65128
rect 181029 64952 184082 64954
rect 181029 64896 181034 64952
rect 181090 64896 184082 64952
rect 181029 64894 184082 64896
rect 181029 64891 181095 64894
rect 87189 64818 87255 64821
rect 131441 64818 131507 64821
rect 226293 64818 226359 64821
rect 87189 64816 90028 64818
rect 87189 64760 87194 64816
rect 87250 64760 90028 64816
rect 87189 64758 90028 64760
rect 129772 64816 131507 64818
rect 129772 64760 131446 64816
rect 131502 64760 131507 64816
rect 129772 64758 131507 64760
rect 223796 64816 226359 64818
rect 223796 64760 226298 64816
rect 226354 64760 226359 64816
rect 223796 64758 226359 64760
rect 87189 64755 87255 64758
rect 131441 64755 131507 64758
rect 226293 64755 226359 64758
rect 233561 64818 233627 64821
rect 237014 64818 237074 65128
rect 233561 64816 237074 64818
rect 233561 64760 233566 64816
rect 233622 64760 237074 64816
rect 233561 64758 237074 64760
rect 233561 64755 233627 64758
rect 80197 64682 80263 64685
rect 76780 64680 80263 64682
rect 76780 64624 80202 64680
rect 80258 64624 80263 64680
rect 76780 64622 80263 64624
rect 80197 64619 80263 64622
rect 181121 64546 181187 64549
rect 184022 64546 184082 64720
rect 181121 64544 184082 64546
rect 181121 64488 181126 64544
rect 181182 64488 184082 64544
rect 181121 64486 184082 64488
rect 233469 64546 233535 64549
rect 233469 64544 237044 64546
rect 233469 64488 233474 64544
rect 233530 64488 237044 64544
rect 233469 64486 237044 64488
rect 181121 64483 181187 64486
rect 233469 64483 233535 64486
rect 87649 64410 87715 64413
rect 131809 64410 131875 64413
rect 87649 64408 90028 64410
rect 87649 64352 87654 64408
rect 87710 64352 90028 64408
rect 87649 64350 90028 64352
rect 129772 64408 131875 64410
rect 129772 64352 131814 64408
rect 131870 64352 131875 64408
rect 129772 64350 131875 64352
rect 87649 64347 87715 64350
rect 131809 64347 131875 64350
rect 139629 64410 139695 64413
rect 173761 64410 173827 64413
rect 139629 64408 143020 64410
rect 139629 64352 139634 64408
rect 139690 64352 143020 64408
rect 139629 64350 143020 64352
rect 170804 64408 173827 64410
rect 170804 64352 173766 64408
rect 173822 64352 173827 64408
rect 170804 64350 173827 64352
rect 139629 64347 139695 64350
rect 173761 64347 173827 64350
rect 181397 64410 181463 64413
rect 226385 64410 226451 64413
rect 181397 64408 184052 64410
rect 181397 64352 181402 64408
rect 181458 64352 184052 64408
rect 181397 64350 184052 64352
rect 223796 64408 226451 64410
rect 223796 64352 226390 64408
rect 226446 64352 226451 64408
rect 223796 64350 226451 64352
rect 181397 64347 181463 64350
rect 226385 64347 226451 64350
rect 80105 64138 80171 64141
rect 76780 64136 80171 64138
rect 76780 64080 80110 64136
rect 80166 64080 80171 64136
rect 76780 64078 80171 64080
rect 80105 64075 80171 64078
rect 131809 64002 131875 64005
rect 226385 64002 226451 64005
rect 129772 64000 131875 64002
rect 129772 63944 131814 64000
rect 131870 63944 131875 64000
rect 129772 63942 131875 63944
rect 223796 64000 226451 64002
rect 223796 63944 226390 64000
rect 226446 63944 226451 64000
rect 223796 63942 226451 63944
rect 131809 63939 131875 63942
rect 226385 63939 226451 63942
rect 87189 63730 87255 63733
rect 89998 63730 90058 63904
rect 174037 63866 174103 63869
rect 170804 63864 174103 63866
rect 170804 63808 174042 63864
rect 174098 63808 174103 63864
rect 170804 63806 174103 63808
rect 174037 63803 174103 63806
rect 87189 63728 90058 63730
rect 87189 63672 87194 63728
rect 87250 63672 90058 63728
rect 87189 63670 90058 63672
rect 139721 63730 139787 63733
rect 182317 63730 182383 63733
rect 184022 63730 184082 63904
rect 139721 63728 143020 63730
rect 139721 63672 139726 63728
rect 139782 63672 143020 63728
rect 139721 63670 143020 63672
rect 182317 63728 184082 63730
rect 182317 63672 182322 63728
rect 182378 63672 184082 63728
rect 182317 63670 184082 63672
rect 87189 63667 87255 63670
rect 139721 63667 139787 63670
rect 182317 63667 182383 63670
rect 80197 63594 80263 63597
rect 131349 63594 131415 63597
rect 226293 63594 226359 63597
rect 76780 63592 80263 63594
rect 76780 63536 80202 63592
rect 80258 63536 80263 63592
rect 76780 63534 80263 63536
rect 129772 63592 131415 63594
rect 129772 63536 131354 63592
rect 131410 63536 131415 63592
rect 129772 63534 131415 63536
rect 223796 63592 226359 63594
rect 223796 63536 226298 63592
rect 226354 63536 226359 63592
rect 223796 63534 226359 63536
rect 80197 63531 80263 63534
rect 131349 63531 131415 63534
rect 226293 63531 226359 63534
rect 87281 63322 87347 63325
rect 89998 63322 90058 63496
rect 173853 63322 173919 63325
rect 87281 63320 90058 63322
rect 87281 63264 87286 63320
rect 87342 63264 90058 63320
rect 87281 63262 90058 63264
rect 170804 63320 173919 63322
rect 170804 63264 173858 63320
rect 173914 63264 173919 63320
rect 170804 63262 173919 63264
rect 87281 63259 87347 63262
rect 173853 63259 173919 63262
rect 182041 63322 182107 63325
rect 184022 63322 184082 63496
rect 233469 63458 233535 63461
rect 237014 63458 237074 63904
rect 233469 63456 237074 63458
rect 233469 63400 233474 63456
rect 233530 63400 237074 63456
rect 233469 63398 237074 63400
rect 233469 63395 233535 63398
rect 182041 63320 184082 63322
rect 182041 63264 182046 63320
rect 182102 63264 184082 63320
rect 182041 63262 184082 63264
rect 233653 63322 233719 63325
rect 233653 63320 237044 63322
rect 233653 63264 233658 63320
rect 233714 63264 237044 63320
rect 233653 63262 237044 63264
rect 182041 63259 182107 63262
rect 233653 63259 233719 63262
rect 131349 63186 131415 63189
rect 129772 63184 131415 63186
rect 129772 63128 131354 63184
rect 131410 63128 131415 63184
rect 129772 63126 131415 63128
rect 131349 63123 131415 63126
rect 139629 63186 139695 63189
rect 226293 63186 226359 63189
rect 139629 63184 143020 63186
rect 139629 63128 139634 63184
rect 139690 63128 143020 63184
rect 139629 63126 143020 63128
rect 223796 63184 226359 63186
rect 223796 63128 226298 63184
rect 226354 63128 226359 63184
rect 223796 63126 226359 63128
rect 139629 63123 139695 63126
rect 226293 63123 226359 63126
rect 80197 63050 80263 63053
rect 76780 63048 80263 63050
rect 76780 62992 80202 63048
rect 80258 62992 80263 63048
rect 76780 62990 80263 62992
rect 80197 62987 80263 62990
rect 87189 62914 87255 62917
rect 89998 62914 90058 63088
rect 87189 62912 90058 62914
rect 87189 62856 87194 62912
rect 87250 62856 90058 62912
rect 87189 62854 90058 62856
rect 182133 62914 182199 62917
rect 184022 62914 184082 63088
rect 182133 62912 184082 62914
rect 182133 62856 182138 62912
rect 182194 62856 184082 62912
rect 182133 62854 184082 62856
rect 87189 62851 87255 62854
rect 182133 62851 182199 62854
rect 87005 62778 87071 62781
rect 131993 62778 132059 62781
rect 173945 62778 174011 62781
rect 87005 62776 90028 62778
rect 87005 62720 87010 62776
rect 87066 62720 90028 62776
rect 87005 62718 90028 62720
rect 129772 62776 132059 62778
rect 129772 62720 131998 62776
rect 132054 62720 132059 62776
rect 129772 62718 132059 62720
rect 170804 62776 174011 62778
rect 170804 62720 173950 62776
rect 174006 62720 174011 62776
rect 170804 62718 174011 62720
rect 87005 62715 87071 62718
rect 131993 62715 132059 62718
rect 173945 62715 174011 62718
rect 182225 62778 182291 62781
rect 226293 62778 226359 62781
rect 182225 62776 184052 62778
rect 182225 62720 182230 62776
rect 182286 62720 184052 62776
rect 182225 62718 184052 62720
rect 223796 62776 226359 62778
rect 223796 62720 226298 62776
rect 226354 62720 226359 62776
rect 223796 62718 226359 62720
rect 182225 62715 182291 62718
rect 226293 62715 226359 62718
rect 233561 62778 233627 62781
rect 233561 62776 237044 62778
rect 233561 62720 233566 62776
rect 233622 62720 237044 62776
rect 233561 62718 237044 62720
rect 233561 62715 233627 62718
rect 80197 62506 80263 62509
rect 76780 62504 80263 62506
rect 76780 62448 80202 62504
rect 80258 62448 80263 62504
rect 76780 62446 80263 62448
rect 80197 62443 80263 62446
rect 139721 62506 139787 62509
rect 139721 62504 143020 62506
rect 139721 62448 139726 62504
rect 139782 62448 143020 62504
rect 139721 62446 143020 62448
rect 139721 62443 139787 62446
rect 87281 62370 87347 62373
rect 131441 62370 131507 62373
rect 87281 62368 90028 62370
rect 87281 62312 87286 62368
rect 87342 62312 90028 62368
rect 87281 62310 90028 62312
rect 129772 62368 131507 62370
rect 129772 62312 131446 62368
rect 131502 62312 131507 62368
rect 129772 62310 131507 62312
rect 87281 62307 87347 62310
rect 131441 62307 131507 62310
rect 181765 62370 181831 62373
rect 226385 62370 226451 62373
rect 181765 62368 184052 62370
rect 181765 62312 181770 62368
rect 181826 62312 184052 62368
rect 181765 62310 184052 62312
rect 223796 62368 226451 62370
rect 223796 62312 226390 62368
rect 226446 62312 226451 62368
rect 223796 62310 226451 62312
rect 181765 62307 181831 62310
rect 226385 62307 226451 62310
rect 173301 62234 173367 62237
rect 170804 62232 173367 62234
rect 170804 62176 173306 62232
rect 173362 62176 173367 62232
rect 170804 62174 173367 62176
rect 173301 62171 173367 62174
rect 233469 62234 233535 62237
rect 233469 62232 237044 62234
rect 233469 62176 233474 62232
rect 233530 62176 237044 62232
rect 233469 62174 237044 62176
rect 233469 62171 233535 62174
rect 131349 62098 131415 62101
rect 226201 62098 226267 62101
rect 129772 62096 131415 62098
rect 129772 62040 131354 62096
rect 131410 62040 131415 62096
rect 129772 62038 131415 62040
rect 223796 62096 226267 62098
rect 223796 62040 226206 62096
rect 226262 62040 226267 62096
rect 223796 62038 226267 62040
rect 131349 62035 131415 62038
rect 226201 62035 226267 62038
rect 47077 61962 47143 61965
rect 47077 61960 48996 61962
rect 47077 61904 47082 61960
rect 47138 61904 48996 61960
rect 47077 61902 48996 61904
rect 47077 61899 47143 61902
rect 80105 61826 80171 61829
rect 76780 61824 80171 61826
rect 76780 61768 80110 61824
rect 80166 61768 80171 61824
rect 76780 61766 80171 61768
rect 80105 61763 80171 61766
rect 87189 61826 87255 61829
rect 89998 61826 90058 62000
rect 87189 61824 90058 61826
rect 87189 61768 87194 61824
rect 87250 61768 90058 61824
rect 87189 61766 90058 61768
rect 139629 61826 139695 61829
rect 173761 61826 173827 61829
rect 139629 61824 143020 61826
rect 139629 61768 139634 61824
rect 139690 61768 143020 61824
rect 139629 61766 143020 61768
rect 170804 61824 173827 61826
rect 170804 61768 173766 61824
rect 173822 61768 173827 61824
rect 170804 61766 173827 61768
rect 87189 61763 87255 61766
rect 139629 61763 139695 61766
rect 173761 61763 173827 61766
rect 181857 61826 181923 61829
rect 184022 61826 184082 62000
rect 181857 61824 184082 61826
rect 181857 61768 181862 61824
rect 181918 61768 184082 61824
rect 181857 61766 184082 61768
rect 181857 61763 181923 61766
rect 131349 61690 131415 61693
rect 226293 61690 226359 61693
rect 129772 61688 131415 61690
rect 129772 61632 131354 61688
rect 131410 61632 131415 61688
rect 129772 61630 131415 61632
rect 223796 61688 226359 61690
rect 223796 61632 226298 61688
rect 226354 61632 226359 61688
rect 223796 61630 226359 61632
rect 131349 61627 131415 61630
rect 226293 61627 226359 61630
rect 87097 61418 87163 61421
rect 89998 61418 90058 61592
rect 87097 61416 90058 61418
rect 87097 61360 87102 61416
rect 87158 61360 90058 61416
rect 87097 61358 90058 61360
rect 181949 61418 182015 61421
rect 184022 61418 184082 61592
rect 233469 61554 233535 61557
rect 233469 61552 237044 61554
rect 233469 61496 233474 61552
rect 233530 61496 237044 61552
rect 233469 61494 237044 61496
rect 233469 61491 233535 61494
rect 181949 61416 184082 61418
rect 181949 61360 181954 61416
rect 182010 61360 184082 61416
rect 181949 61358 184082 61360
rect 87097 61355 87163 61358
rect 181949 61355 182015 61358
rect 173945 61282 174011 61285
rect 225741 61282 225807 61285
rect 170804 61280 174011 61282
rect 170804 61224 173950 61280
rect 174006 61224 174011 61280
rect 170804 61222 174011 61224
rect 223796 61280 225807 61282
rect 223796 61224 225746 61280
rect 225802 61224 225807 61280
rect 223796 61222 225807 61224
rect 173945 61219 174011 61222
rect 225741 61219 225807 61222
rect 76750 60874 76810 61184
rect 87189 61010 87255 61013
rect 89998 61010 90058 61184
rect 87189 61008 90058 61010
rect 87189 60952 87194 61008
rect 87250 60952 90058 61008
rect 87189 60950 90058 60952
rect 129742 61010 129802 61184
rect 139629 61146 139695 61149
rect 139629 61144 143020 61146
rect 139629 61088 139634 61144
rect 139690 61088 143020 61144
rect 139629 61086 143020 61088
rect 139629 61083 139695 61086
rect 131441 61010 131507 61013
rect 129742 61008 131507 61010
rect 129742 60952 131446 61008
rect 131502 60952 131507 61008
rect 129742 60950 131507 60952
rect 87189 60947 87255 60950
rect 131441 60947 131507 60950
rect 181673 61010 181739 61013
rect 184022 61010 184082 61184
rect 181673 61008 184082 61010
rect 181673 60952 181678 61008
rect 181734 60952 184082 61008
rect 181673 60950 184082 60952
rect 233469 61010 233535 61013
rect 233469 61008 237044 61010
rect 233469 60952 233474 61008
rect 233530 60952 237044 61008
rect 233469 60950 237044 60952
rect 181673 60947 181739 60950
rect 233469 60947 233535 60950
rect 79093 60874 79159 60877
rect 131349 60874 131415 60877
rect 225925 60874 225991 60877
rect 76750 60872 79159 60874
rect 76750 60816 79098 60872
rect 79154 60816 79159 60872
rect 76750 60814 79159 60816
rect 129772 60872 131415 60874
rect 129772 60816 131354 60872
rect 131410 60816 131415 60872
rect 129772 60814 131415 60816
rect 223796 60872 225991 60874
rect 223796 60816 225930 60872
rect 225986 60816 225991 60872
rect 223796 60814 225991 60816
rect 79093 60811 79159 60814
rect 131349 60811 131415 60814
rect 225925 60811 225991 60814
rect 80197 60738 80263 60741
rect 76780 60736 80263 60738
rect 76780 60680 80202 60736
rect 80258 60680 80263 60736
rect 76780 60678 80263 60680
rect 80197 60675 80263 60678
rect 86913 60602 86979 60605
rect 89998 60602 90058 60776
rect 174037 60738 174103 60741
rect 170804 60736 174103 60738
rect 170804 60680 174042 60736
rect 174098 60680 174103 60736
rect 170804 60678 174103 60680
rect 174037 60675 174103 60678
rect 86913 60600 90058 60602
rect 86913 60544 86918 60600
rect 86974 60544 90058 60600
rect 86913 60542 90058 60544
rect 139629 60602 139695 60605
rect 182133 60602 182199 60605
rect 184022 60602 184082 60776
rect 139629 60600 143020 60602
rect 139629 60544 139634 60600
rect 139690 60544 143020 60600
rect 139629 60542 143020 60544
rect 182133 60600 184082 60602
rect 182133 60544 182138 60600
rect 182194 60544 184082 60600
rect 182133 60542 184082 60544
rect 86913 60539 86979 60542
rect 139629 60539 139695 60542
rect 182133 60539 182199 60542
rect 226385 60466 226451 60469
rect 223796 60464 226451 60466
rect 223796 60408 226390 60464
rect 226446 60408 226451 60464
rect 223796 60406 226451 60408
rect 226385 60403 226451 60406
rect 80105 60194 80171 60197
rect 76780 60192 80171 60194
rect 76780 60136 80110 60192
rect 80166 60136 80171 60192
rect 76780 60134 80171 60136
rect 80105 60131 80171 60134
rect 87005 60194 87071 60197
rect 89998 60194 90058 60368
rect 87005 60192 90058 60194
rect 87005 60136 87010 60192
rect 87066 60136 90058 60192
rect 87005 60134 90058 60136
rect 129742 60194 129802 60368
rect 131349 60194 131415 60197
rect 173669 60194 173735 60197
rect 129742 60192 131415 60194
rect 129742 60136 131354 60192
rect 131410 60136 131415 60192
rect 129742 60134 131415 60136
rect 170804 60192 173735 60194
rect 170804 60136 173674 60192
rect 173730 60136 173735 60192
rect 170804 60134 173735 60136
rect 87005 60131 87071 60134
rect 131349 60131 131415 60134
rect 173669 60131 173735 60134
rect 182225 60194 182291 60197
rect 184022 60194 184082 60368
rect 233561 60330 233627 60333
rect 233561 60328 237044 60330
rect 233561 60272 233566 60328
rect 233622 60272 237044 60328
rect 233561 60270 237044 60272
rect 233561 60267 233627 60270
rect 182225 60192 184082 60194
rect 182225 60136 182230 60192
rect 182286 60136 184082 60192
rect 182225 60134 184082 60136
rect 182225 60131 182291 60134
rect 86821 60058 86887 60061
rect 131809 60058 131875 60061
rect 86821 60056 90028 60058
rect 86821 60000 86826 60056
rect 86882 60000 90028 60056
rect 86821 59998 90028 60000
rect 129772 60056 131875 60058
rect 129772 60000 131814 60056
rect 131870 60000 131875 60056
rect 129772 59998 131875 60000
rect 86821 59995 86887 59998
rect 131809 59995 131875 59998
rect 182317 60058 182383 60061
rect 226293 60058 226359 60061
rect 182317 60056 184052 60058
rect 182317 60000 182322 60056
rect 182378 60000 184052 60056
rect 182317 59998 184052 60000
rect 223796 60056 226359 60058
rect 223796 60000 226298 60056
rect 226354 60000 226359 60056
rect 223796 59998 226359 60000
rect 182317 59995 182383 59998
rect 226293 59995 226359 59998
rect 139721 59922 139787 59925
rect 139721 59920 143020 59922
rect 139721 59864 139726 59920
rect 139782 59864 143020 59920
rect 139721 59862 143020 59864
rect 139721 59859 139787 59862
rect 233469 59786 233535 59789
rect 233469 59784 237044 59786
rect 233469 59728 233474 59784
rect 233530 59728 237044 59784
rect 233469 59726 237044 59728
rect 233469 59723 233535 59726
rect 80197 59650 80263 59653
rect 174037 59650 174103 59653
rect 76780 59648 80263 59650
rect 76780 59592 80202 59648
rect 80258 59592 80263 59648
rect 76780 59590 80263 59592
rect 170804 59648 174103 59650
rect 170804 59592 174042 59648
rect 174098 59592 174103 59648
rect 170804 59590 174103 59592
rect 80197 59587 80263 59590
rect 174037 59587 174103 59590
rect 180937 59650 181003 59653
rect 226201 59650 226267 59653
rect 180937 59648 184052 59650
rect 180937 59592 180942 59648
rect 180998 59592 184052 59648
rect 180937 59590 184052 59592
rect 223796 59648 226267 59650
rect 223796 59592 226206 59648
rect 226262 59592 226267 59648
rect 223796 59590 226267 59592
rect 180937 59587 181003 59590
rect 226201 59587 226267 59590
rect 87373 59378 87439 59381
rect 89998 59378 90058 59552
rect 87373 59376 90058 59378
rect 87373 59320 87378 59376
rect 87434 59320 90058 59376
rect 87373 59318 90058 59320
rect 129742 59378 129802 59552
rect 131533 59378 131599 59381
rect 129742 59376 131599 59378
rect 129742 59320 131538 59376
rect 131594 59320 131599 59376
rect 129742 59318 131599 59320
rect 87373 59315 87439 59318
rect 131533 59315 131599 59318
rect 139629 59242 139695 59245
rect 226385 59242 226451 59245
rect 139629 59240 143020 59242
rect 139629 59184 139634 59240
rect 139690 59184 143020 59240
rect 139629 59182 143020 59184
rect 223796 59240 226451 59242
rect 223796 59184 226390 59240
rect 226446 59184 226451 59240
rect 223796 59182 226451 59184
rect 139629 59179 139695 59182
rect 226385 59179 226451 59182
rect 80105 58970 80171 58973
rect 76780 58968 80171 58970
rect 76780 58912 80110 58968
rect 80166 58912 80171 58968
rect 76780 58910 80171 58912
rect 80105 58907 80171 58910
rect 87281 58970 87347 58973
rect 89998 58970 90058 59144
rect 87281 58968 90058 58970
rect 87281 58912 87286 58968
rect 87342 58912 90058 58968
rect 87281 58910 90058 58912
rect 129742 58970 129802 59144
rect 173669 59106 173735 59109
rect 170804 59104 173735 59106
rect 170804 59048 173674 59104
rect 173730 59048 173735 59104
rect 170804 59046 173735 59048
rect 173669 59043 173735 59046
rect 131441 58970 131507 58973
rect 129742 58968 131507 58970
rect 129742 58912 131446 58968
rect 131502 58912 131507 58968
rect 129742 58910 131507 58912
rect 87281 58907 87347 58910
rect 131441 58907 131507 58910
rect 182225 58970 182291 58973
rect 184022 58970 184082 59144
rect 233561 59106 233627 59109
rect 233561 59104 237044 59106
rect 233561 59048 233566 59104
rect 233622 59048 237044 59104
rect 233561 59046 237044 59048
rect 233561 59043 233627 59046
rect 182225 58968 184082 58970
rect 182225 58912 182230 58968
rect 182286 58912 184082 58968
rect 182225 58910 184082 58912
rect 182225 58907 182291 58910
rect 87189 58834 87255 58837
rect 131349 58834 131415 58837
rect 226293 58834 226359 58837
rect 87189 58832 90028 58834
rect 87189 58776 87194 58832
rect 87250 58776 90028 58832
rect 87189 58774 90028 58776
rect 129772 58832 131415 58834
rect 129772 58776 131354 58832
rect 131410 58776 131415 58832
rect 129772 58774 131415 58776
rect 223796 58832 226359 58834
rect 223796 58776 226298 58832
rect 226354 58776 226359 58832
rect 223796 58774 226359 58776
rect 87189 58771 87255 58774
rect 131349 58771 131415 58774
rect 226293 58771 226359 58774
rect 139721 58562 139787 58565
rect 173853 58562 173919 58565
rect 139721 58560 143020 58562
rect 139721 58504 139726 58560
rect 139782 58504 143020 58560
rect 139721 58502 143020 58504
rect 170804 58560 173919 58562
rect 170804 58504 173858 58560
rect 173914 58504 173919 58560
rect 170804 58502 173919 58504
rect 139721 58499 139787 58502
rect 173853 58499 173919 58502
rect 182041 58562 182107 58565
rect 184022 58562 184082 58736
rect 182041 58560 184082 58562
rect 182041 58504 182046 58560
rect 182102 58504 184082 58560
rect 182041 58502 184082 58504
rect 233745 58562 233811 58565
rect 233745 58560 237044 58562
rect 233745 58504 233750 58560
rect 233806 58504 237044 58560
rect 233745 58502 237044 58504
rect 182041 58499 182107 58502
rect 233745 58499 233811 58502
rect 80197 58426 80263 58429
rect 225741 58426 225807 58429
rect 76780 58424 80263 58426
rect 76780 58368 80202 58424
rect 80258 58368 80263 58424
rect 76780 58366 80263 58368
rect 223796 58424 225807 58426
rect 223796 58368 225746 58424
rect 225802 58368 225807 58424
rect 223796 58366 225807 58368
rect 80197 58363 80263 58366
rect 225741 58363 225807 58366
rect 87005 58154 87071 58157
rect 89998 58154 90058 58328
rect 87005 58152 90058 58154
rect 87005 58096 87010 58152
rect 87066 58096 90058 58152
rect 87005 58094 90058 58096
rect 129742 58154 129802 58328
rect 131533 58154 131599 58157
rect 129742 58152 131599 58154
rect 129742 58096 131538 58152
rect 131594 58096 131599 58152
rect 129742 58094 131599 58096
rect 87005 58091 87071 58094
rect 131533 58091 131599 58094
rect 182317 58154 182383 58157
rect 184022 58154 184082 58328
rect 182317 58152 184082 58154
rect 182317 58096 182322 58152
rect 182378 58096 184082 58152
rect 182317 58094 184082 58096
rect 182317 58091 182383 58094
rect 174037 58018 174103 58021
rect 225925 58018 225991 58021
rect 170804 58016 174103 58018
rect 170804 57960 174042 58016
rect 174098 57960 174103 58016
rect 170804 57958 174103 57960
rect 223796 58016 225991 58018
rect 223796 57960 225930 58016
rect 225986 57960 225991 58016
rect 223796 57958 225991 57960
rect 174037 57955 174103 57958
rect 225925 57955 225991 57958
rect 9896 57882 10376 57912
rect 13313 57882 13379 57885
rect 80105 57882 80171 57885
rect 9896 57880 13379 57882
rect 9896 57824 13318 57880
rect 13374 57824 13379 57880
rect 9896 57822 13379 57824
rect 76780 57880 80171 57882
rect 76780 57824 80110 57880
rect 80166 57824 80171 57880
rect 76780 57822 80171 57824
rect 9896 57792 10376 57822
rect 13313 57819 13379 57822
rect 80105 57819 80171 57822
rect 87097 57746 87163 57749
rect 89998 57746 90058 57920
rect 87097 57744 90058 57746
rect 87097 57688 87102 57744
rect 87158 57688 90058 57744
rect 87097 57686 90058 57688
rect 129742 57746 129802 57920
rect 139629 57882 139695 57885
rect 139629 57880 143020 57882
rect 139629 57824 139634 57880
rect 139690 57824 143020 57880
rect 139629 57822 143020 57824
rect 139629 57819 139695 57822
rect 131625 57746 131691 57749
rect 129742 57744 131691 57746
rect 129742 57688 131630 57744
rect 131686 57688 131691 57744
rect 129742 57686 131691 57688
rect 87097 57683 87163 57686
rect 131625 57683 131691 57686
rect 180293 57746 180359 57749
rect 181673 57746 181739 57749
rect 184022 57746 184082 57920
rect 233837 57882 233903 57885
rect 233837 57880 237044 57882
rect 233837 57824 233842 57880
rect 233898 57824 237044 57880
rect 233837 57822 237044 57824
rect 233837 57819 233903 57822
rect 180293 57744 181506 57746
rect 180293 57688 180298 57744
rect 180354 57688 181506 57744
rect 180293 57686 181506 57688
rect 180293 57683 180359 57686
rect 131441 57610 131507 57613
rect 129772 57608 131507 57610
rect 129772 57552 131446 57608
rect 131502 57552 131507 57608
rect 129772 57550 131507 57552
rect 131441 57547 131507 57550
rect 80197 57338 80263 57341
rect 76780 57336 80263 57338
rect 76780 57280 80202 57336
rect 80258 57280 80263 57336
rect 76780 57278 80263 57280
rect 80197 57275 80263 57278
rect 86729 57338 86795 57341
rect 89998 57338 90058 57512
rect 173761 57474 173827 57477
rect 170804 57472 173827 57474
rect 170804 57416 173766 57472
rect 173822 57416 173827 57472
rect 170804 57414 173827 57416
rect 181446 57474 181506 57686
rect 181673 57744 184082 57746
rect 181673 57688 181678 57744
rect 181734 57688 184082 57744
rect 181673 57686 184082 57688
rect 181673 57683 181739 57686
rect 225833 57610 225899 57613
rect 223796 57608 225899 57610
rect 223796 57552 225838 57608
rect 225894 57552 225899 57608
rect 223796 57550 225899 57552
rect 225833 57547 225899 57550
rect 183697 57474 183763 57477
rect 181446 57472 183763 57474
rect 181446 57416 183702 57472
rect 183758 57416 183763 57472
rect 181446 57414 183763 57416
rect 173761 57411 173827 57414
rect 183697 57411 183763 57414
rect 86729 57336 90058 57338
rect 86729 57280 86734 57336
rect 86790 57280 90058 57336
rect 86729 57278 90058 57280
rect 139721 57338 139787 57341
rect 181581 57338 181647 57341
rect 184022 57338 184082 57512
rect 139721 57336 143020 57338
rect 139721 57280 139726 57336
rect 139782 57280 143020 57336
rect 139721 57278 143020 57280
rect 181581 57336 184082 57338
rect 181581 57280 181586 57336
rect 181642 57280 184082 57336
rect 181581 57278 184082 57280
rect 233469 57338 233535 57341
rect 233469 57336 237044 57338
rect 233469 57280 233474 57336
rect 233530 57280 237044 57336
rect 233469 57278 237044 57280
rect 86729 57275 86795 57278
rect 139721 57275 139787 57278
rect 181581 57275 181647 57278
rect 233469 57275 233535 57278
rect 86545 57202 86611 57205
rect 131349 57202 131415 57205
rect 226477 57202 226543 57205
rect 86545 57200 90028 57202
rect 86545 57144 86550 57200
rect 86606 57144 90028 57200
rect 86545 57142 90028 57144
rect 129772 57200 131415 57202
rect 129772 57144 131354 57200
rect 131410 57144 131415 57200
rect 129772 57142 131415 57144
rect 223796 57200 226543 57202
rect 223796 57144 226482 57200
rect 226538 57144 226543 57200
rect 223796 57142 226543 57144
rect 86545 57139 86611 57142
rect 131349 57139 131415 57142
rect 226477 57139 226543 57142
rect 183697 57134 183763 57137
rect 183697 57132 184052 57134
rect 183697 57076 183702 57132
rect 183758 57076 184052 57132
rect 183697 57074 184052 57076
rect 183697 57071 183763 57074
rect 174037 57066 174103 57069
rect 170804 57064 174103 57066
rect 170804 57008 174042 57064
rect 174098 57008 174103 57064
rect 170804 57006 174103 57008
rect 174037 57003 174103 57006
rect 80197 56794 80263 56797
rect 225925 56794 225991 56797
rect 76780 56792 80263 56794
rect 76780 56736 80202 56792
rect 80258 56736 80263 56792
rect 76780 56734 80263 56736
rect 223796 56792 225991 56794
rect 223796 56736 225930 56792
rect 225986 56736 225991 56792
rect 223796 56734 225991 56736
rect 80197 56731 80263 56734
rect 225925 56731 225991 56734
rect 88201 56522 88267 56525
rect 89998 56522 90058 56696
rect 88201 56520 90058 56522
rect 88201 56464 88206 56520
rect 88262 56464 90058 56520
rect 88201 56462 90058 56464
rect 129742 56522 129802 56696
rect 139813 56658 139879 56661
rect 139813 56656 143020 56658
rect 139813 56600 139818 56656
rect 139874 56600 143020 56656
rect 139813 56598 143020 56600
rect 139813 56595 139879 56598
rect 131441 56522 131507 56525
rect 174037 56522 174103 56525
rect 129742 56520 131507 56522
rect 129742 56464 131446 56520
rect 131502 56464 131507 56520
rect 129742 56462 131507 56464
rect 170804 56520 174103 56522
rect 170804 56464 174042 56520
rect 174098 56464 174103 56520
rect 170804 56462 174103 56464
rect 88201 56459 88267 56462
rect 131441 56459 131507 56462
rect 174037 56459 174103 56462
rect 181305 56522 181371 56525
rect 184022 56522 184082 56696
rect 233561 56658 233627 56661
rect 233561 56656 237044 56658
rect 233561 56600 233566 56656
rect 233622 56600 237044 56656
rect 233561 56598 237044 56600
rect 233561 56595 233627 56598
rect 181305 56520 184082 56522
rect 181305 56464 181310 56520
rect 181366 56464 184082 56520
rect 181305 56462 184082 56464
rect 181305 56459 181371 56462
rect 226293 56386 226359 56389
rect 223796 56384 226359 56386
rect 223796 56328 226298 56384
rect 226354 56328 226359 56384
rect 223796 56326 226359 56328
rect 226293 56323 226359 56326
rect 80105 56114 80171 56117
rect 76780 56112 80171 56114
rect 76780 56056 80110 56112
rect 80166 56056 80171 56112
rect 76780 56054 80171 56056
rect 80105 56051 80171 56054
rect 88385 56114 88451 56117
rect 89998 56114 90058 56288
rect 88385 56112 90058 56114
rect 88385 56056 88390 56112
rect 88446 56056 90058 56112
rect 88385 56054 90058 56056
rect 129742 56114 129802 56288
rect 131533 56114 131599 56117
rect 129742 56112 131599 56114
rect 129742 56056 131538 56112
rect 131594 56056 131599 56112
rect 129742 56054 131599 56056
rect 88385 56051 88451 56054
rect 131533 56051 131599 56054
rect 181213 56114 181279 56117
rect 184022 56114 184082 56288
rect 181213 56112 184082 56114
rect 181213 56056 181218 56112
rect 181274 56056 184082 56112
rect 181213 56054 184082 56056
rect 233653 56114 233719 56117
rect 233653 56112 237044 56114
rect 233653 56056 233658 56112
rect 233714 56056 237044 56112
rect 233653 56054 237044 56056
rect 181213 56051 181279 56054
rect 233653 56051 233719 56054
rect 87925 55978 87991 55981
rect 131349 55978 131415 55981
rect 87925 55976 90028 55978
rect 87925 55920 87930 55976
rect 87986 55920 90028 55976
rect 87925 55918 90028 55920
rect 129772 55976 131415 55978
rect 129772 55920 131354 55976
rect 131410 55920 131415 55976
rect 129772 55918 131415 55920
rect 87925 55915 87991 55918
rect 131349 55915 131415 55918
rect 139629 55978 139695 55981
rect 172933 55978 172999 55981
rect 139629 55976 143020 55978
rect 139629 55920 139634 55976
rect 139690 55920 143020 55976
rect 139629 55918 143020 55920
rect 170804 55976 172999 55978
rect 170804 55920 172938 55976
rect 172994 55920 172999 55976
rect 170804 55918 172999 55920
rect 139629 55915 139695 55918
rect 172933 55915 172999 55918
rect 182317 55978 182383 55981
rect 226293 55978 226359 55981
rect 182317 55976 184052 55978
rect 182317 55920 182322 55976
rect 182378 55920 184052 55976
rect 182317 55918 184052 55920
rect 223796 55976 226359 55978
rect 223796 55920 226298 55976
rect 226354 55920 226359 55976
rect 223796 55918 226359 55920
rect 182317 55915 182383 55918
rect 226293 55915 226359 55918
rect 80013 55570 80079 55573
rect 225741 55570 225807 55573
rect 76780 55568 80079 55570
rect 76780 55512 80018 55568
rect 80074 55512 80079 55568
rect 76780 55510 80079 55512
rect 223796 55568 225807 55570
rect 223796 55512 225746 55568
rect 225802 55512 225807 55568
rect 223796 55510 225807 55512
rect 80013 55507 80079 55510
rect 225741 55507 225807 55510
rect 87281 55298 87347 55301
rect 89998 55298 90058 55472
rect 87281 55296 90058 55298
rect 87281 55240 87286 55296
rect 87342 55240 90058 55296
rect 87281 55238 90058 55240
rect 129742 55298 129802 55472
rect 173301 55434 173367 55437
rect 170804 55432 173367 55434
rect 170804 55376 173306 55432
rect 173362 55376 173367 55432
rect 170804 55374 173367 55376
rect 173301 55371 173367 55374
rect 131533 55298 131599 55301
rect 129742 55296 131599 55298
rect 129742 55240 131538 55296
rect 131594 55240 131599 55296
rect 129742 55238 131599 55240
rect 87281 55235 87347 55238
rect 131533 55235 131599 55238
rect 139721 55298 139787 55301
rect 181121 55298 181187 55301
rect 184022 55298 184082 55472
rect 233469 55434 233535 55437
rect 264749 55434 264815 55437
rect 233469 55432 237044 55434
rect 233469 55376 233474 55432
rect 233530 55376 237044 55432
rect 233469 55374 237044 55376
rect 264749 55432 264858 55434
rect 264749 55376 264754 55432
rect 264810 55376 264858 55432
rect 233469 55371 233535 55374
rect 264749 55371 264858 55376
rect 139721 55296 143020 55298
rect 139721 55240 139726 55296
rect 139782 55240 143020 55296
rect 139721 55238 143020 55240
rect 181121 55296 184082 55298
rect 181121 55240 181126 55296
rect 181182 55240 184082 55296
rect 181121 55238 184082 55240
rect 139721 55235 139787 55238
rect 181121 55235 181187 55238
rect 226385 55162 226451 55165
rect 223796 55160 226451 55162
rect 223796 55104 226390 55160
rect 226446 55104 226451 55160
rect 223796 55102 226451 55104
rect 226385 55099 226451 55102
rect 80197 55026 80263 55029
rect 76780 55024 80263 55026
rect 76780 54968 80202 55024
rect 80258 54968 80263 55024
rect 76780 54966 80263 54968
rect 80197 54963 80263 54966
rect 87189 54890 87255 54893
rect 89998 54890 90058 55064
rect 87189 54888 90058 54890
rect 87189 54832 87194 54888
rect 87250 54832 90058 54888
rect 87189 54830 90058 54832
rect 129742 54890 129802 55064
rect 131441 54890 131507 54893
rect 173761 54890 173827 54893
rect 129742 54888 131507 54890
rect 129742 54832 131446 54888
rect 131502 54832 131507 54888
rect 129742 54830 131507 54832
rect 170804 54888 173827 54890
rect 170804 54832 173766 54888
rect 173822 54832 173827 54888
rect 170804 54830 173827 54832
rect 87189 54827 87255 54830
rect 131441 54827 131507 54830
rect 173761 54827 173827 54830
rect 181673 54890 181739 54893
rect 184022 54890 184082 55064
rect 181673 54888 184082 54890
rect 181673 54832 181678 54888
rect 181734 54832 184082 54888
rect 181673 54830 184082 54832
rect 233561 54890 233627 54893
rect 233561 54888 237044 54890
rect 233561 54832 233566 54888
rect 233622 54832 237044 54888
rect 264798 54860 264858 55371
rect 233561 54830 237044 54832
rect 181673 54827 181739 54830
rect 233561 54827 233627 54830
rect 131349 54754 131415 54757
rect 226293 54754 226359 54757
rect 129772 54752 131415 54754
rect 129772 54696 131354 54752
rect 131410 54696 131415 54752
rect 129772 54694 131415 54696
rect 223796 54752 226359 54754
rect 223796 54696 226298 54752
rect 226354 54696 226359 54752
rect 223796 54694 226359 54696
rect 131349 54691 131415 54694
rect 226293 54691 226359 54694
rect 80105 54482 80171 54485
rect 76780 54480 80171 54482
rect 76780 54424 80110 54480
rect 80166 54424 80171 54480
rect 76780 54422 80171 54424
rect 80105 54419 80171 54422
rect 87281 54482 87347 54485
rect 89998 54482 90058 54656
rect 139905 54618 139971 54621
rect 139905 54616 143020 54618
rect 139905 54560 139910 54616
rect 139966 54560 143020 54616
rect 139905 54558 143020 54560
rect 139905 54555 139971 54558
rect 87281 54480 90058 54482
rect 87281 54424 87286 54480
rect 87342 54424 90058 54480
rect 87281 54422 90058 54424
rect 181581 54482 181647 54485
rect 184022 54482 184082 54656
rect 181581 54480 184082 54482
rect 181581 54424 181586 54480
rect 181642 54424 184082 54480
rect 181581 54422 184082 54424
rect 87281 54419 87347 54422
rect 181581 54419 181647 54422
rect 87097 54346 87163 54349
rect 131441 54346 131507 54349
rect 174037 54346 174103 54349
rect 87097 54344 90028 54346
rect 87097 54288 87102 54344
rect 87158 54288 90028 54344
rect 87097 54286 90028 54288
rect 129772 54344 131507 54346
rect 129772 54288 131446 54344
rect 131502 54288 131507 54344
rect 129772 54286 131507 54288
rect 170804 54344 174103 54346
rect 170804 54288 174042 54344
rect 174098 54288 174103 54344
rect 170804 54286 174103 54288
rect 87097 54283 87163 54286
rect 131441 54283 131507 54286
rect 174037 54283 174103 54286
rect 182317 54346 182383 54349
rect 226293 54346 226359 54349
rect 182317 54344 184052 54346
rect 182317 54288 182322 54344
rect 182378 54288 184052 54344
rect 182317 54286 184052 54288
rect 223796 54344 226359 54346
rect 223796 54288 226298 54344
rect 226354 54288 226359 54344
rect 223796 54286 226359 54288
rect 182317 54283 182383 54286
rect 226293 54283 226359 54286
rect 233469 54210 233535 54213
rect 233469 54208 237044 54210
rect 233469 54152 233474 54208
rect 233530 54152 237044 54208
rect 233469 54150 237044 54152
rect 233469 54147 233535 54150
rect 139721 54074 139787 54077
rect 225833 54074 225899 54077
rect 139721 54072 143020 54074
rect 139721 54016 139726 54072
rect 139782 54016 143020 54072
rect 139721 54014 143020 54016
rect 223796 54072 225899 54074
rect 223796 54016 225838 54072
rect 225894 54016 225899 54072
rect 223796 54014 225899 54016
rect 139721 54011 139787 54014
rect 225833 54011 225899 54014
rect 80197 53938 80263 53941
rect 76780 53936 80263 53938
rect 76780 53880 80202 53936
rect 80258 53880 80263 53936
rect 76780 53878 80263 53880
rect 80197 53875 80263 53878
rect 87189 53394 87255 53397
rect 89998 53394 90058 53976
rect 104342 53740 104348 53804
rect 104412 53802 104418 53804
rect 104577 53802 104643 53805
rect 104412 53800 104643 53802
rect 104412 53744 104582 53800
rect 104638 53744 104643 53800
rect 104412 53742 104643 53744
rect 104412 53740 104418 53742
rect 104577 53739 104643 53742
rect 129742 53530 129802 53976
rect 174037 53802 174103 53805
rect 170804 53800 174103 53802
rect 170804 53744 174042 53800
rect 174098 53744 174103 53800
rect 170804 53742 174103 53744
rect 174037 53739 174103 53742
rect 131349 53530 131415 53533
rect 129742 53528 131415 53530
rect 129742 53472 131354 53528
rect 131410 53472 131415 53528
rect 129742 53470 131415 53472
rect 131349 53467 131415 53470
rect 87189 53392 90058 53394
rect 87189 53336 87194 53392
rect 87250 53336 90058 53392
rect 87189 53334 90058 53336
rect 139997 53394 140063 53397
rect 139997 53392 143020 53394
rect 139997 53336 140002 53392
rect 140058 53336 143020 53392
rect 139997 53334 143020 53336
rect 87189 53331 87255 53334
rect 139997 53331 140063 53334
rect 80197 53258 80263 53261
rect 173485 53258 173551 53261
rect 76780 53256 80263 53258
rect 76780 53200 80202 53256
rect 80258 53200 80263 53256
rect 76780 53198 80263 53200
rect 170804 53256 173551 53258
rect 170804 53200 173490 53256
rect 173546 53200 173551 53256
rect 170804 53198 173551 53200
rect 80197 53195 80263 53198
rect 173485 53195 173551 53198
rect 180937 53122 181003 53125
rect 184022 53122 184082 53976
rect 233561 53666 233627 53669
rect 233561 53664 237044 53666
rect 233561 53608 233566 53664
rect 233622 53608 237044 53664
rect 233561 53606 237044 53608
rect 233561 53603 233627 53606
rect 180937 53120 184082 53122
rect 180937 53064 180942 53120
rect 180998 53064 184082 53120
rect 180937 53062 184082 53064
rect 180937 53059 181003 53062
rect 233469 52986 233535 52989
rect 233469 52984 237044 52986
rect 233469 52928 233474 52984
rect 233530 52928 237044 52984
rect 233469 52926 237044 52928
rect 233469 52923 233535 52926
rect 80197 52714 80263 52717
rect 76780 52712 80263 52714
rect 76780 52656 80202 52712
rect 80258 52656 80263 52712
rect 76780 52654 80263 52656
rect 80197 52651 80263 52654
rect 139537 52714 139603 52717
rect 173945 52714 174011 52717
rect 139537 52712 143020 52714
rect 139537 52656 139542 52712
rect 139598 52656 143020 52712
rect 139537 52654 143020 52656
rect 170804 52712 174011 52714
rect 170804 52656 173950 52712
rect 174006 52656 174011 52712
rect 170804 52654 174011 52656
rect 139537 52651 139603 52654
rect 173945 52651 174011 52654
rect 233653 52442 233719 52445
rect 233653 52440 237044 52442
rect 233653 52384 233658 52440
rect 233714 52384 237044 52440
rect 233653 52382 237044 52384
rect 233653 52379 233719 52382
rect 174037 52306 174103 52309
rect 170804 52304 174103 52306
rect 170804 52248 174042 52304
rect 174098 52248 174103 52304
rect 170804 52246 174103 52248
rect 174037 52243 174103 52246
rect 80105 52170 80171 52173
rect 76780 52168 80171 52170
rect 76780 52112 80110 52168
rect 80166 52112 80171 52168
rect 76780 52110 80171 52112
rect 80105 52107 80171 52110
rect 139445 52034 139511 52037
rect 139445 52032 143020 52034
rect 139445 51976 139450 52032
rect 139506 51976 143020 52032
rect 139445 51974 143020 51976
rect 139445 51971 139511 51974
rect 172841 51762 172907 51765
rect 170804 51760 172907 51762
rect 170804 51704 172846 51760
rect 172902 51704 172907 51760
rect 170804 51702 172907 51704
rect 172841 51699 172907 51702
rect 233469 51762 233535 51765
rect 233469 51760 237044 51762
rect 233469 51704 233474 51760
rect 233530 51704 237044 51760
rect 233469 51702 237044 51704
rect 233469 51699 233535 51702
rect 80197 51626 80263 51629
rect 76780 51624 80263 51626
rect 76780 51568 80202 51624
rect 80258 51568 80263 51624
rect 76780 51566 80263 51568
rect 80197 51563 80263 51566
rect 139629 51354 139695 51357
rect 139629 51352 143020 51354
rect 139629 51296 139634 51352
rect 139690 51296 143020 51352
rect 139629 51294 143020 51296
rect 139629 51291 139695 51294
rect 172933 51218 172999 51221
rect 170804 51216 172999 51218
rect 170804 51160 172938 51216
rect 172994 51160 172999 51216
rect 170804 51158 172999 51160
rect 172933 51155 172999 51158
rect 233469 51218 233535 51221
rect 233469 51216 237044 51218
rect 233469 51160 233474 51216
rect 233530 51160 237044 51216
rect 233469 51158 237044 51160
rect 233469 51155 233535 51158
rect 79737 51082 79803 51085
rect 76780 51080 79803 51082
rect 76780 51024 79742 51080
rect 79798 51024 79803 51080
rect 76780 51022 79803 51024
rect 79737 51019 79803 51022
rect 139905 50810 139971 50813
rect 139905 50808 143020 50810
rect 139905 50752 139910 50808
rect 139966 50752 143020 50808
rect 139905 50750 143020 50752
rect 139905 50747 139971 50750
rect 173945 50674 174011 50677
rect 170804 50672 174011 50674
rect 170804 50616 173950 50672
rect 174006 50616 174011 50672
rect 170804 50614 174011 50616
rect 173945 50611 174011 50614
rect 233653 50538 233719 50541
rect 233653 50536 237044 50538
rect 233653 50480 233658 50536
rect 233714 50480 237044 50536
rect 233653 50478 237044 50480
rect 233653 50475 233719 50478
rect 79461 50402 79527 50405
rect 76780 50400 79527 50402
rect 76780 50344 79466 50400
rect 79522 50344 79527 50400
rect 76780 50342 79527 50344
rect 79461 50339 79527 50342
rect 139629 50130 139695 50133
rect 173301 50130 173367 50133
rect 139629 50128 143020 50130
rect 139629 50072 139634 50128
rect 139690 50072 143020 50128
rect 139629 50070 143020 50072
rect 170804 50128 173367 50130
rect 170804 50072 173306 50128
rect 173362 50072 173367 50128
rect 170804 50070 173367 50072
rect 139629 50067 139695 50070
rect 173301 50067 173367 50070
rect 233653 49994 233719 49997
rect 233653 49992 237044 49994
rect 233653 49936 233658 49992
rect 233714 49936 237044 49992
rect 233653 49934 237044 49936
rect 233653 49931 233719 49934
rect 76750 49450 76810 49760
rect 172749 49586 172815 49589
rect 170804 49584 172815 49586
rect 170804 49528 172754 49584
rect 172810 49528 172815 49584
rect 170804 49526 172815 49528
rect 172749 49523 172815 49526
rect 80105 49450 80171 49453
rect 76750 49448 80171 49450
rect 76750 49392 80110 49448
rect 80166 49392 80171 49448
rect 76750 49390 80171 49392
rect 80105 49387 80171 49390
rect 139721 49450 139787 49453
rect 139721 49448 143020 49450
rect 139721 49392 139726 49448
rect 139782 49392 143020 49448
rect 139721 49390 143020 49392
rect 139721 49387 139787 49390
rect 80197 49314 80263 49317
rect 76780 49312 80263 49314
rect 76780 49256 80202 49312
rect 80258 49256 80263 49312
rect 76780 49254 80263 49256
rect 80197 49251 80263 49254
rect 233469 49314 233535 49317
rect 233469 49312 237044 49314
rect 233469 49256 233474 49312
rect 233530 49256 237044 49312
rect 233469 49254 237044 49256
rect 233469 49251 233535 49254
rect 173117 49042 173183 49045
rect 170804 49040 173183 49042
rect 170804 48984 173122 49040
rect 173178 48984 173183 49040
rect 170804 48982 173183 48984
rect 173117 48979 173183 48982
rect 80013 48770 80079 48773
rect 76780 48768 80079 48770
rect 76780 48712 80018 48768
rect 80074 48712 80079 48768
rect 76780 48710 80079 48712
rect 80013 48707 80079 48710
rect 139813 48770 139879 48773
rect 233561 48770 233627 48773
rect 139813 48768 143020 48770
rect 139813 48712 139818 48768
rect 139874 48712 143020 48768
rect 139813 48710 143020 48712
rect 233561 48768 237044 48770
rect 233561 48712 233566 48768
rect 233622 48712 237044 48768
rect 233561 48710 237044 48712
rect 139813 48707 139879 48710
rect 233561 48707 233627 48710
rect 173301 48498 173367 48501
rect 170804 48496 173367 48498
rect 170804 48440 173306 48496
rect 173362 48440 173367 48496
rect 170804 48438 173367 48440
rect 173301 48435 173367 48438
rect 139629 48226 139695 48229
rect 139629 48224 143020 48226
rect 139629 48168 139634 48224
rect 139690 48168 143020 48224
rect 139629 48166 143020 48168
rect 139629 48163 139695 48166
rect 76750 47546 76810 48128
rect 173393 48090 173459 48093
rect 170804 48088 173459 48090
rect 170804 48032 173398 48088
rect 173454 48032 173459 48088
rect 170804 48030 173459 48032
rect 173393 48027 173459 48030
rect 233469 47682 233535 47685
rect 237014 47682 237074 48128
rect 233469 47680 237074 47682
rect 233469 47624 233474 47680
rect 233530 47624 237074 47680
rect 233469 47622 237074 47624
rect 233469 47619 233535 47622
rect 79553 47546 79619 47549
rect 76750 47544 79619 47546
rect 76750 47488 79558 47544
rect 79614 47488 79619 47544
rect 76750 47486 79619 47488
rect 79553 47483 79619 47486
rect 236822 47484 236828 47548
rect 236892 47546 236898 47548
rect 241197 47546 241263 47549
rect 236892 47544 241263 47546
rect 236892 47488 241202 47544
rect 241258 47488 241263 47544
rect 236892 47486 241263 47488
rect 236892 47484 236898 47486
rect 241197 47483 241263 47486
rect 144270 45988 144276 46052
rect 144340 46050 144346 46052
rect 156557 46050 156623 46053
rect 144340 46048 156623 46050
rect 144340 45992 156562 46048
rect 156618 45992 156623 46048
rect 144340 45990 156623 45992
rect 144340 45988 144346 45990
rect 156557 45987 156623 45990
rect 237006 45852 237012 45916
rect 237076 45914 237082 45916
rect 250489 45914 250555 45917
rect 237076 45912 250555 45914
rect 237076 45856 250494 45912
rect 250550 45856 250555 45912
rect 237076 45854 250555 45856
rect 237076 45852 237082 45854
rect 250489 45851 250555 45854
rect 300169 45642 300235 45645
rect 303416 45642 303896 45672
rect 300169 45640 303896 45642
rect 300169 45584 300174 45640
rect 300230 45584 303896 45640
rect 300169 45582 303896 45584
rect 300169 45579 300235 45582
rect 303416 45552 303896 45582
rect 215529 34490 215595 34493
rect 218606 34490 218612 34492
rect 215529 34488 218612 34490
rect 215529 34432 215534 34488
rect 215590 34432 218612 34488
rect 215529 34430 218612 34432
rect 215529 34427 215595 34430
rect 218606 34428 218612 34430
rect 218676 34428 218682 34492
rect 129509 27554 129575 27557
rect 129509 27552 129618 27554
rect 129509 27496 129514 27552
rect 129570 27496 129618 27552
rect 129509 27491 129618 27496
rect 182174 27492 182180 27556
rect 182244 27554 182250 27556
rect 223533 27554 223599 27557
rect 182244 27494 184082 27554
rect 182244 27492 182250 27494
rect 129558 26916 129618 27491
rect 184022 26916 184082 27494
rect 223533 27552 223642 27554
rect 223533 27496 223538 27552
rect 223594 27496 223642 27552
rect 223533 27491 223642 27496
rect 223582 26912 223642 27491
rect 88477 26874 88543 26877
rect 89998 26874 90058 26912
rect 88477 26872 90058 26874
rect 88477 26816 88482 26872
rect 88538 26816 90058 26872
rect 88477 26814 90058 26816
rect 88477 26811 88543 26814
rect 9896 25242 10376 25272
rect 13313 25242 13379 25245
rect 9896 25240 13379 25242
rect 9896 25184 13318 25240
rect 13374 25184 13379 25240
rect 9896 25182 13379 25184
rect 9896 25152 10376 25182
rect 13313 25179 13379 25182
rect 299801 21162 299867 21165
rect 303416 21162 303896 21192
rect 299801 21160 303896 21162
rect 299801 21104 299806 21160
rect 299862 21104 303896 21160
rect 299801 21102 303896 21104
rect 299801 21099 299867 21102
rect 303416 21072 303896 21102
rect 211941 12322 212007 12325
rect 218606 12322 218612 12324
rect 211941 12320 218612 12322
rect 211941 12264 211946 12320
rect 212002 12264 218612 12320
rect 211941 12262 218612 12264
rect 211941 12259 212007 12262
rect 218606 12260 218612 12262
rect 218676 12260 218682 12324
rect 101725 12186 101791 12189
rect 131390 12186 131396 12188
rect 101725 12184 131396 12186
rect 101725 12128 101730 12184
rect 101786 12128 131396 12184
rect 101725 12126 131396 12128
rect 101725 12123 101791 12126
rect 131390 12124 131396 12126
rect 131460 12124 131466 12188
<< via3 >>
rect 131396 288204 131460 288268
rect 223580 288204 223644 288268
rect 90180 287796 90244 287860
rect 129556 287796 129620 287860
rect 184204 287796 184268 287860
rect 52460 265492 52524 265556
rect 52276 263724 52340 263788
rect 142252 263724 142316 263788
rect 226340 257604 226404 257668
rect 265164 256788 265228 256852
rect 142252 240468 142316 240532
rect 69756 224148 69820 224212
rect 241612 221564 241676 221628
rect 38108 218708 38172 218772
rect 265164 216592 265228 216596
rect 265164 216536 265214 216592
rect 265214 216536 265228 216592
rect 265164 216532 265228 216536
rect 293684 216532 293748 216596
rect 52276 216124 52340 216188
rect 81716 215172 81780 215236
rect 164884 212588 164948 212652
rect 135260 211772 135324 211836
rect 52460 202932 52524 202996
rect 20076 202252 20140 202316
rect 228916 202252 228980 202316
rect 242900 202252 242964 202316
rect 258908 202252 258972 202316
rect 278044 202252 278108 202316
rect 293684 202252 293748 202316
rect 35900 202116 35964 202180
rect 241612 181172 241676 181236
rect 85028 174644 85092 174708
rect 133236 174644 133300 174708
rect 128452 174508 128516 174572
rect 48228 144044 48292 144108
rect 109500 143968 109564 143972
rect 109500 143912 109550 143968
rect 109550 143912 109564 143968
rect 109500 143908 109564 143912
rect 128452 139828 128516 139892
rect 264980 138604 265044 138668
rect 20812 131532 20876 131596
rect 69756 130308 69820 130372
rect 288716 130308 288780 130372
rect 58164 130172 58228 130236
rect 61476 130172 61540 130236
rect 135444 130172 135508 130236
rect 138756 130172 138820 130236
rect 244004 130172 244068 130236
rect 245108 130172 245172 130236
rect 48596 129492 48660 129556
rect 57796 129492 57860 129556
rect 251364 129492 251428 129556
rect 269212 129492 269276 129556
rect 241612 127452 241676 127516
rect 48228 123236 48292 123300
rect 293684 122012 293748 122076
rect 81716 121332 81780 121396
rect 261116 120712 261180 120716
rect 261116 120656 261130 120712
rect 261130 120656 261180 120712
rect 261116 120652 261180 120656
rect 264980 120652 265044 120716
rect 229652 120244 229716 120308
rect 20076 108412 20140 108476
rect 35900 108276 35964 108340
rect 241612 87332 241676 87396
rect 85028 84068 85092 84132
rect 133236 83660 133300 83724
rect 182180 83720 182244 83724
rect 182180 83664 182194 83720
rect 182194 83664 182244 83720
rect 182180 83660 182244 83664
rect 237012 81348 237076 81412
rect 144276 81212 144340 81276
rect 236828 81212 236892 81276
rect 103980 77812 104044 77876
rect 104348 53740 104412 53804
rect 236828 47484 236892 47548
rect 144276 45988 144340 46052
rect 237012 45852 237076 45916
rect 218612 34428 218676 34492
rect 182180 27492 182244 27556
rect 218612 12260 218676 12324
rect 131396 12124 131460 12188
<< metal4 >>
rect 0 311286 4000 311408
rect 0 311050 122 311286
rect 358 311050 442 311286
rect 678 311050 762 311286
rect 998 311050 1082 311286
rect 1318 311050 1402 311286
rect 1638 311050 1722 311286
rect 1958 311050 2042 311286
rect 2278 311050 2362 311286
rect 2598 311050 2682 311286
rect 2918 311050 3002 311286
rect 3238 311050 3322 311286
rect 3558 311050 3642 311286
rect 3878 311050 4000 311286
rect 0 310966 4000 311050
rect 0 310730 122 310966
rect 358 310730 442 310966
rect 678 310730 762 310966
rect 998 310730 1082 310966
rect 1318 310730 1402 310966
rect 1638 310730 1722 310966
rect 1958 310730 2042 310966
rect 2278 310730 2362 310966
rect 2598 310730 2682 310966
rect 2918 310730 3002 310966
rect 3238 310730 3322 310966
rect 3558 310730 3642 310966
rect 3878 310730 4000 310966
rect 0 310646 4000 310730
rect 0 310410 122 310646
rect 358 310410 442 310646
rect 678 310410 762 310646
rect 998 310410 1082 310646
rect 1318 310410 1402 310646
rect 1638 310410 1722 310646
rect 1958 310410 2042 310646
rect 2278 310410 2362 310646
rect 2598 310410 2682 310646
rect 2918 310410 3002 310646
rect 3238 310410 3322 310646
rect 3558 310410 3642 310646
rect 3878 310410 4000 310646
rect 0 310326 4000 310410
rect 0 310090 122 310326
rect 358 310090 442 310326
rect 678 310090 762 310326
rect 998 310090 1082 310326
rect 1318 310090 1402 310326
rect 1638 310090 1722 310326
rect 1958 310090 2042 310326
rect 2278 310090 2362 310326
rect 2598 310090 2682 310326
rect 2918 310090 3002 310326
rect 3238 310090 3322 310326
rect 3558 310090 3642 310326
rect 3878 310090 4000 310326
rect 0 310006 4000 310090
rect 0 309770 122 310006
rect 358 309770 442 310006
rect 678 309770 762 310006
rect 998 309770 1082 310006
rect 1318 309770 1402 310006
rect 1638 309770 1722 310006
rect 1958 309770 2042 310006
rect 2278 309770 2362 310006
rect 2598 309770 2682 310006
rect 2918 309770 3002 310006
rect 3238 309770 3322 310006
rect 3558 309770 3642 310006
rect 3878 309770 4000 310006
rect 0 309686 4000 309770
rect 0 309450 122 309686
rect 358 309450 442 309686
rect 678 309450 762 309686
rect 998 309450 1082 309686
rect 1318 309450 1402 309686
rect 1638 309450 1722 309686
rect 1958 309450 2042 309686
rect 2278 309450 2362 309686
rect 2598 309450 2682 309686
rect 2918 309450 3002 309686
rect 3238 309450 3322 309686
rect 3558 309450 3642 309686
rect 3878 309450 4000 309686
rect 0 309366 4000 309450
rect 0 309130 122 309366
rect 358 309130 442 309366
rect 678 309130 762 309366
rect 998 309130 1082 309366
rect 1318 309130 1402 309366
rect 1638 309130 1722 309366
rect 1958 309130 2042 309366
rect 2278 309130 2362 309366
rect 2598 309130 2682 309366
rect 2918 309130 3002 309366
rect 3238 309130 3322 309366
rect 3558 309130 3642 309366
rect 3878 309130 4000 309366
rect 0 309046 4000 309130
rect 0 308810 122 309046
rect 358 308810 442 309046
rect 678 308810 762 309046
rect 998 308810 1082 309046
rect 1318 308810 1402 309046
rect 1638 308810 1722 309046
rect 1958 308810 2042 309046
rect 2278 308810 2362 309046
rect 2598 308810 2682 309046
rect 2918 308810 3002 309046
rect 3238 308810 3322 309046
rect 3558 308810 3642 309046
rect 3878 308810 4000 309046
rect 0 308726 4000 308810
rect 0 308490 122 308726
rect 358 308490 442 308726
rect 678 308490 762 308726
rect 998 308490 1082 308726
rect 1318 308490 1402 308726
rect 1638 308490 1722 308726
rect 1958 308490 2042 308726
rect 2278 308490 2362 308726
rect 2598 308490 2682 308726
rect 2918 308490 3002 308726
rect 3238 308490 3322 308726
rect 3558 308490 3642 308726
rect 3878 308490 4000 308726
rect 0 308406 4000 308490
rect 0 308170 122 308406
rect 358 308170 442 308406
rect 678 308170 762 308406
rect 998 308170 1082 308406
rect 1318 308170 1402 308406
rect 1638 308170 1722 308406
rect 1958 308170 2042 308406
rect 2278 308170 2362 308406
rect 2598 308170 2682 308406
rect 2918 308170 3002 308406
rect 3238 308170 3322 308406
rect 3558 308170 3642 308406
rect 3878 308170 4000 308406
rect 0 308086 4000 308170
rect 0 307850 122 308086
rect 358 307850 442 308086
rect 678 307850 762 308086
rect 998 307850 1082 308086
rect 1318 307850 1402 308086
rect 1638 307850 1722 308086
rect 1958 307850 2042 308086
rect 2278 307850 2362 308086
rect 2598 307850 2682 308086
rect 2918 307850 3002 308086
rect 3238 307850 3322 308086
rect 3558 307850 3642 308086
rect 3878 307850 4000 308086
rect 0 307766 4000 307850
rect 0 307530 122 307766
rect 358 307530 442 307766
rect 678 307530 762 307766
rect 998 307530 1082 307766
rect 1318 307530 1402 307766
rect 1638 307530 1722 307766
rect 1958 307530 2042 307766
rect 2278 307530 2362 307766
rect 2598 307530 2682 307766
rect 2918 307530 3002 307766
rect 3238 307530 3322 307766
rect 3558 307530 3642 307766
rect 3878 307530 4000 307766
rect 0 284524 4000 307530
rect 309732 311286 313732 311408
rect 309732 311050 309854 311286
rect 310090 311050 310174 311286
rect 310410 311050 310494 311286
rect 310730 311050 310814 311286
rect 311050 311050 311134 311286
rect 311370 311050 311454 311286
rect 311690 311050 311774 311286
rect 312010 311050 312094 311286
rect 312330 311050 312414 311286
rect 312650 311050 312734 311286
rect 312970 311050 313054 311286
rect 313290 311050 313374 311286
rect 313610 311050 313732 311286
rect 309732 310966 313732 311050
rect 309732 310730 309854 310966
rect 310090 310730 310174 310966
rect 310410 310730 310494 310966
rect 310730 310730 310814 310966
rect 311050 310730 311134 310966
rect 311370 310730 311454 310966
rect 311690 310730 311774 310966
rect 312010 310730 312094 310966
rect 312330 310730 312414 310966
rect 312650 310730 312734 310966
rect 312970 310730 313054 310966
rect 313290 310730 313374 310966
rect 313610 310730 313732 310966
rect 309732 310646 313732 310730
rect 309732 310410 309854 310646
rect 310090 310410 310174 310646
rect 310410 310410 310494 310646
rect 310730 310410 310814 310646
rect 311050 310410 311134 310646
rect 311370 310410 311454 310646
rect 311690 310410 311774 310646
rect 312010 310410 312094 310646
rect 312330 310410 312414 310646
rect 312650 310410 312734 310646
rect 312970 310410 313054 310646
rect 313290 310410 313374 310646
rect 313610 310410 313732 310646
rect 309732 310326 313732 310410
rect 309732 310090 309854 310326
rect 310090 310090 310174 310326
rect 310410 310090 310494 310326
rect 310730 310090 310814 310326
rect 311050 310090 311134 310326
rect 311370 310090 311454 310326
rect 311690 310090 311774 310326
rect 312010 310090 312094 310326
rect 312330 310090 312414 310326
rect 312650 310090 312734 310326
rect 312970 310090 313054 310326
rect 313290 310090 313374 310326
rect 313610 310090 313732 310326
rect 309732 310006 313732 310090
rect 309732 309770 309854 310006
rect 310090 309770 310174 310006
rect 310410 309770 310494 310006
rect 310730 309770 310814 310006
rect 311050 309770 311134 310006
rect 311370 309770 311454 310006
rect 311690 309770 311774 310006
rect 312010 309770 312094 310006
rect 312330 309770 312414 310006
rect 312650 309770 312734 310006
rect 312970 309770 313054 310006
rect 313290 309770 313374 310006
rect 313610 309770 313732 310006
rect 309732 309686 313732 309770
rect 309732 309450 309854 309686
rect 310090 309450 310174 309686
rect 310410 309450 310494 309686
rect 310730 309450 310814 309686
rect 311050 309450 311134 309686
rect 311370 309450 311454 309686
rect 311690 309450 311774 309686
rect 312010 309450 312094 309686
rect 312330 309450 312414 309686
rect 312650 309450 312734 309686
rect 312970 309450 313054 309686
rect 313290 309450 313374 309686
rect 313610 309450 313732 309686
rect 309732 309366 313732 309450
rect 309732 309130 309854 309366
rect 310090 309130 310174 309366
rect 310410 309130 310494 309366
rect 310730 309130 310814 309366
rect 311050 309130 311134 309366
rect 311370 309130 311454 309366
rect 311690 309130 311774 309366
rect 312010 309130 312094 309366
rect 312330 309130 312414 309366
rect 312650 309130 312734 309366
rect 312970 309130 313054 309366
rect 313290 309130 313374 309366
rect 313610 309130 313732 309366
rect 309732 309046 313732 309130
rect 309732 308810 309854 309046
rect 310090 308810 310174 309046
rect 310410 308810 310494 309046
rect 310730 308810 310814 309046
rect 311050 308810 311134 309046
rect 311370 308810 311454 309046
rect 311690 308810 311774 309046
rect 312010 308810 312094 309046
rect 312330 308810 312414 309046
rect 312650 308810 312734 309046
rect 312970 308810 313054 309046
rect 313290 308810 313374 309046
rect 313610 308810 313732 309046
rect 309732 308726 313732 308810
rect 309732 308490 309854 308726
rect 310090 308490 310174 308726
rect 310410 308490 310494 308726
rect 310730 308490 310814 308726
rect 311050 308490 311134 308726
rect 311370 308490 311454 308726
rect 311690 308490 311774 308726
rect 312010 308490 312094 308726
rect 312330 308490 312414 308726
rect 312650 308490 312734 308726
rect 312970 308490 313054 308726
rect 313290 308490 313374 308726
rect 313610 308490 313732 308726
rect 309732 308406 313732 308490
rect 309732 308170 309854 308406
rect 310090 308170 310174 308406
rect 310410 308170 310494 308406
rect 310730 308170 310814 308406
rect 311050 308170 311134 308406
rect 311370 308170 311454 308406
rect 311690 308170 311774 308406
rect 312010 308170 312094 308406
rect 312330 308170 312414 308406
rect 312650 308170 312734 308406
rect 312970 308170 313054 308406
rect 313290 308170 313374 308406
rect 313610 308170 313732 308406
rect 309732 308086 313732 308170
rect 309732 307850 309854 308086
rect 310090 307850 310174 308086
rect 310410 307850 310494 308086
rect 310730 307850 310814 308086
rect 311050 307850 311134 308086
rect 311370 307850 311454 308086
rect 311690 307850 311774 308086
rect 312010 307850 312094 308086
rect 312330 307850 312414 308086
rect 312650 307850 312734 308086
rect 312970 307850 313054 308086
rect 313290 307850 313374 308086
rect 313610 307850 313732 308086
rect 309732 307766 313732 307850
rect 309732 307530 309854 307766
rect 310090 307530 310174 307766
rect 310410 307530 310494 307766
rect 310730 307530 310814 307766
rect 311050 307530 311134 307766
rect 311370 307530 311454 307766
rect 311690 307530 311774 307766
rect 312010 307530 312094 307766
rect 312330 307530 312414 307766
rect 312650 307530 312734 307766
rect 312970 307530 313054 307766
rect 313290 307530 313374 307766
rect 313610 307530 313732 307766
rect 0 284288 122 284524
rect 358 284288 442 284524
rect 678 284288 762 284524
rect 998 284288 1082 284524
rect 1318 284288 1402 284524
rect 1638 284288 1722 284524
rect 1958 284288 2042 284524
rect 2278 284288 2362 284524
rect 2598 284288 2682 284524
rect 2918 284288 3002 284524
rect 3238 284288 3322 284524
rect 3558 284288 3642 284524
rect 3878 284288 4000 284524
rect 0 253888 4000 284288
rect 0 253652 122 253888
rect 358 253652 442 253888
rect 678 253652 762 253888
rect 998 253652 1082 253888
rect 1318 253652 1402 253888
rect 1638 253652 1722 253888
rect 1958 253652 2042 253888
rect 2278 253652 2362 253888
rect 2598 253652 2682 253888
rect 2918 253652 3002 253888
rect 3238 253652 3322 253888
rect 3558 253652 3642 253888
rect 3878 253652 4000 253888
rect 0 223252 4000 253652
rect 0 223016 122 223252
rect 358 223016 442 223252
rect 678 223016 762 223252
rect 998 223016 1082 223252
rect 1318 223016 1402 223252
rect 1638 223016 1722 223252
rect 1958 223016 2042 223252
rect 2278 223016 2362 223252
rect 2598 223016 2682 223252
rect 2918 223016 3002 223252
rect 3238 223016 3322 223252
rect 3558 223016 3642 223252
rect 3878 223016 4000 223252
rect 0 192616 4000 223016
rect 0 192380 122 192616
rect 358 192380 442 192616
rect 678 192380 762 192616
rect 998 192380 1082 192616
rect 1318 192380 1402 192616
rect 1638 192380 1722 192616
rect 1958 192380 2042 192616
rect 2278 192380 2362 192616
rect 2598 192380 2682 192616
rect 2918 192380 3002 192616
rect 3238 192380 3322 192616
rect 3558 192380 3642 192616
rect 3878 192380 4000 192616
rect 0 161980 4000 192380
rect 0 161744 122 161980
rect 358 161744 442 161980
rect 678 161744 762 161980
rect 998 161744 1082 161980
rect 1318 161744 1402 161980
rect 1638 161744 1722 161980
rect 1958 161744 2042 161980
rect 2278 161744 2362 161980
rect 2598 161744 2682 161980
rect 2918 161744 3002 161980
rect 3238 161744 3322 161980
rect 3558 161744 3642 161980
rect 3878 161744 4000 161980
rect 0 131344 4000 161744
rect 0 131108 122 131344
rect 358 131108 442 131344
rect 678 131108 762 131344
rect 998 131108 1082 131344
rect 1318 131108 1402 131344
rect 1638 131108 1722 131344
rect 1958 131108 2042 131344
rect 2278 131108 2362 131344
rect 2598 131108 2682 131344
rect 2918 131108 3002 131344
rect 3238 131108 3322 131344
rect 3558 131108 3642 131344
rect 3878 131108 4000 131344
rect 0 100708 4000 131108
rect 0 100472 122 100708
rect 358 100472 442 100708
rect 678 100472 762 100708
rect 998 100472 1082 100708
rect 1318 100472 1402 100708
rect 1638 100472 1722 100708
rect 1958 100472 2042 100708
rect 2278 100472 2362 100708
rect 2598 100472 2682 100708
rect 2918 100472 3002 100708
rect 3238 100472 3322 100708
rect 3558 100472 3642 100708
rect 3878 100472 4000 100708
rect 0 70072 4000 100472
rect 0 69836 122 70072
rect 358 69836 442 70072
rect 678 69836 762 70072
rect 998 69836 1082 70072
rect 1318 69836 1402 70072
rect 1638 69836 1722 70072
rect 1958 69836 2042 70072
rect 2278 69836 2362 70072
rect 2598 69836 2682 70072
rect 2918 69836 3002 70072
rect 3238 69836 3322 70072
rect 3558 69836 3642 70072
rect 3878 69836 4000 70072
rect 0 39436 4000 69836
rect 0 39200 122 39436
rect 358 39200 442 39436
rect 678 39200 762 39436
rect 998 39200 1082 39436
rect 1318 39200 1402 39436
rect 1638 39200 1722 39436
rect 1958 39200 2042 39436
rect 2278 39200 2362 39436
rect 2598 39200 2682 39436
rect 2918 39200 3002 39436
rect 3238 39200 3322 39436
rect 3558 39200 3642 39436
rect 3878 39200 4000 39436
rect 0 3878 4000 39200
rect 5000 306286 9000 306408
rect 5000 306050 5122 306286
rect 5358 306050 5442 306286
rect 5678 306050 5762 306286
rect 5998 306050 6082 306286
rect 6318 306050 6402 306286
rect 6638 306050 6722 306286
rect 6958 306050 7042 306286
rect 7278 306050 7362 306286
rect 7598 306050 7682 306286
rect 7918 306050 8002 306286
rect 8238 306050 8322 306286
rect 8558 306050 8642 306286
rect 8878 306050 9000 306286
rect 5000 305966 9000 306050
rect 5000 305730 5122 305966
rect 5358 305730 5442 305966
rect 5678 305730 5762 305966
rect 5998 305730 6082 305966
rect 6318 305730 6402 305966
rect 6638 305730 6722 305966
rect 6958 305730 7042 305966
rect 7278 305730 7362 305966
rect 7598 305730 7682 305966
rect 7918 305730 8002 305966
rect 8238 305730 8322 305966
rect 8558 305730 8642 305966
rect 8878 305730 9000 305966
rect 5000 305646 9000 305730
rect 5000 305410 5122 305646
rect 5358 305410 5442 305646
rect 5678 305410 5762 305646
rect 5998 305410 6082 305646
rect 6318 305410 6402 305646
rect 6638 305410 6722 305646
rect 6958 305410 7042 305646
rect 7278 305410 7362 305646
rect 7598 305410 7682 305646
rect 7918 305410 8002 305646
rect 8238 305410 8322 305646
rect 8558 305410 8642 305646
rect 8878 305410 9000 305646
rect 5000 305326 9000 305410
rect 5000 305090 5122 305326
rect 5358 305090 5442 305326
rect 5678 305090 5762 305326
rect 5998 305090 6082 305326
rect 6318 305090 6402 305326
rect 6638 305090 6722 305326
rect 6958 305090 7042 305326
rect 7278 305090 7362 305326
rect 7598 305090 7682 305326
rect 7918 305090 8002 305326
rect 8238 305090 8322 305326
rect 8558 305090 8642 305326
rect 8878 305090 9000 305326
rect 5000 305006 9000 305090
rect 5000 304770 5122 305006
rect 5358 304770 5442 305006
rect 5678 304770 5762 305006
rect 5998 304770 6082 305006
rect 6318 304770 6402 305006
rect 6638 304770 6722 305006
rect 6958 304770 7042 305006
rect 7278 304770 7362 305006
rect 7598 304770 7682 305006
rect 7918 304770 8002 305006
rect 8238 304770 8322 305006
rect 8558 304770 8642 305006
rect 8878 304770 9000 305006
rect 5000 304686 9000 304770
rect 5000 304450 5122 304686
rect 5358 304450 5442 304686
rect 5678 304450 5762 304686
rect 5998 304450 6082 304686
rect 6318 304450 6402 304686
rect 6638 304450 6722 304686
rect 6958 304450 7042 304686
rect 7278 304450 7362 304686
rect 7598 304450 7682 304686
rect 7918 304450 8002 304686
rect 8238 304450 8322 304686
rect 8558 304450 8642 304686
rect 8878 304450 9000 304686
rect 5000 304366 9000 304450
rect 5000 304130 5122 304366
rect 5358 304130 5442 304366
rect 5678 304130 5762 304366
rect 5998 304130 6082 304366
rect 6318 304130 6402 304366
rect 6638 304130 6722 304366
rect 6958 304130 7042 304366
rect 7278 304130 7362 304366
rect 7598 304130 7682 304366
rect 7918 304130 8002 304366
rect 8238 304130 8322 304366
rect 8558 304130 8642 304366
rect 8878 304130 9000 304366
rect 5000 304046 9000 304130
rect 5000 303810 5122 304046
rect 5358 303810 5442 304046
rect 5678 303810 5762 304046
rect 5998 303810 6082 304046
rect 6318 303810 6402 304046
rect 6638 303810 6722 304046
rect 6958 303810 7042 304046
rect 7278 303810 7362 304046
rect 7598 303810 7682 304046
rect 7918 303810 8002 304046
rect 8238 303810 8322 304046
rect 8558 303810 8642 304046
rect 8878 303810 9000 304046
rect 5000 303726 9000 303810
rect 5000 303490 5122 303726
rect 5358 303490 5442 303726
rect 5678 303490 5762 303726
rect 5998 303490 6082 303726
rect 6318 303490 6402 303726
rect 6638 303490 6722 303726
rect 6958 303490 7042 303726
rect 7278 303490 7362 303726
rect 7598 303490 7682 303726
rect 7918 303490 8002 303726
rect 8238 303490 8322 303726
rect 8558 303490 8642 303726
rect 8878 303490 9000 303726
rect 5000 303406 9000 303490
rect 5000 303170 5122 303406
rect 5358 303170 5442 303406
rect 5678 303170 5762 303406
rect 5998 303170 6082 303406
rect 6318 303170 6402 303406
rect 6638 303170 6722 303406
rect 6958 303170 7042 303406
rect 7278 303170 7362 303406
rect 7598 303170 7682 303406
rect 7918 303170 8002 303406
rect 8238 303170 8322 303406
rect 8558 303170 8642 303406
rect 8878 303170 9000 303406
rect 5000 303086 9000 303170
rect 5000 302850 5122 303086
rect 5358 302850 5442 303086
rect 5678 302850 5762 303086
rect 5998 302850 6082 303086
rect 6318 302850 6402 303086
rect 6638 302850 6722 303086
rect 6958 302850 7042 303086
rect 7278 302850 7362 303086
rect 7598 302850 7682 303086
rect 7918 302850 8002 303086
rect 8238 302850 8322 303086
rect 8558 302850 8642 303086
rect 8878 302850 9000 303086
rect 5000 302766 9000 302850
rect 5000 302530 5122 302766
rect 5358 302530 5442 302766
rect 5678 302530 5762 302766
rect 5998 302530 6082 302766
rect 6318 302530 6402 302766
rect 6638 302530 6722 302766
rect 6958 302530 7042 302766
rect 7278 302530 7362 302766
rect 7598 302530 7682 302766
rect 7918 302530 8002 302766
rect 8238 302530 8322 302766
rect 8558 302530 8642 302766
rect 8878 302530 9000 302766
rect 5000 299842 9000 302530
rect 5000 299606 5122 299842
rect 5358 299606 5442 299842
rect 5678 299606 5762 299842
rect 5998 299606 6082 299842
rect 6318 299606 6402 299842
rect 6638 299606 6722 299842
rect 6958 299606 7042 299842
rect 7278 299606 7362 299842
rect 7598 299606 7682 299842
rect 7918 299606 8002 299842
rect 8238 299606 8322 299842
rect 8558 299606 8642 299842
rect 8878 299606 9000 299842
rect 5000 269206 9000 299606
rect 304732 306286 308732 306408
rect 304732 306050 304854 306286
rect 305090 306050 305174 306286
rect 305410 306050 305494 306286
rect 305730 306050 305814 306286
rect 306050 306050 306134 306286
rect 306370 306050 306454 306286
rect 306690 306050 306774 306286
rect 307010 306050 307094 306286
rect 307330 306050 307414 306286
rect 307650 306050 307734 306286
rect 307970 306050 308054 306286
rect 308290 306050 308374 306286
rect 308610 306050 308732 306286
rect 304732 305966 308732 306050
rect 304732 305730 304854 305966
rect 305090 305730 305174 305966
rect 305410 305730 305494 305966
rect 305730 305730 305814 305966
rect 306050 305730 306134 305966
rect 306370 305730 306454 305966
rect 306690 305730 306774 305966
rect 307010 305730 307094 305966
rect 307330 305730 307414 305966
rect 307650 305730 307734 305966
rect 307970 305730 308054 305966
rect 308290 305730 308374 305966
rect 308610 305730 308732 305966
rect 304732 305646 308732 305730
rect 304732 305410 304854 305646
rect 305090 305410 305174 305646
rect 305410 305410 305494 305646
rect 305730 305410 305814 305646
rect 306050 305410 306134 305646
rect 306370 305410 306454 305646
rect 306690 305410 306774 305646
rect 307010 305410 307094 305646
rect 307330 305410 307414 305646
rect 307650 305410 307734 305646
rect 307970 305410 308054 305646
rect 308290 305410 308374 305646
rect 308610 305410 308732 305646
rect 304732 305326 308732 305410
rect 304732 305090 304854 305326
rect 305090 305090 305174 305326
rect 305410 305090 305494 305326
rect 305730 305090 305814 305326
rect 306050 305090 306134 305326
rect 306370 305090 306454 305326
rect 306690 305090 306774 305326
rect 307010 305090 307094 305326
rect 307330 305090 307414 305326
rect 307650 305090 307734 305326
rect 307970 305090 308054 305326
rect 308290 305090 308374 305326
rect 308610 305090 308732 305326
rect 304732 305006 308732 305090
rect 304732 304770 304854 305006
rect 305090 304770 305174 305006
rect 305410 304770 305494 305006
rect 305730 304770 305814 305006
rect 306050 304770 306134 305006
rect 306370 304770 306454 305006
rect 306690 304770 306774 305006
rect 307010 304770 307094 305006
rect 307330 304770 307414 305006
rect 307650 304770 307734 305006
rect 307970 304770 308054 305006
rect 308290 304770 308374 305006
rect 308610 304770 308732 305006
rect 304732 304686 308732 304770
rect 304732 304450 304854 304686
rect 305090 304450 305174 304686
rect 305410 304450 305494 304686
rect 305730 304450 305814 304686
rect 306050 304450 306134 304686
rect 306370 304450 306454 304686
rect 306690 304450 306774 304686
rect 307010 304450 307094 304686
rect 307330 304450 307414 304686
rect 307650 304450 307734 304686
rect 307970 304450 308054 304686
rect 308290 304450 308374 304686
rect 308610 304450 308732 304686
rect 304732 304366 308732 304450
rect 304732 304130 304854 304366
rect 305090 304130 305174 304366
rect 305410 304130 305494 304366
rect 305730 304130 305814 304366
rect 306050 304130 306134 304366
rect 306370 304130 306454 304366
rect 306690 304130 306774 304366
rect 307010 304130 307094 304366
rect 307330 304130 307414 304366
rect 307650 304130 307734 304366
rect 307970 304130 308054 304366
rect 308290 304130 308374 304366
rect 308610 304130 308732 304366
rect 304732 304046 308732 304130
rect 304732 303810 304854 304046
rect 305090 303810 305174 304046
rect 305410 303810 305494 304046
rect 305730 303810 305814 304046
rect 306050 303810 306134 304046
rect 306370 303810 306454 304046
rect 306690 303810 306774 304046
rect 307010 303810 307094 304046
rect 307330 303810 307414 304046
rect 307650 303810 307734 304046
rect 307970 303810 308054 304046
rect 308290 303810 308374 304046
rect 308610 303810 308732 304046
rect 304732 303726 308732 303810
rect 304732 303490 304854 303726
rect 305090 303490 305174 303726
rect 305410 303490 305494 303726
rect 305730 303490 305814 303726
rect 306050 303490 306134 303726
rect 306370 303490 306454 303726
rect 306690 303490 306774 303726
rect 307010 303490 307094 303726
rect 307330 303490 307414 303726
rect 307650 303490 307734 303726
rect 307970 303490 308054 303726
rect 308290 303490 308374 303726
rect 308610 303490 308732 303726
rect 304732 303406 308732 303490
rect 304732 303170 304854 303406
rect 305090 303170 305174 303406
rect 305410 303170 305494 303406
rect 305730 303170 305814 303406
rect 306050 303170 306134 303406
rect 306370 303170 306454 303406
rect 306690 303170 306774 303406
rect 307010 303170 307094 303406
rect 307330 303170 307414 303406
rect 307650 303170 307734 303406
rect 307970 303170 308054 303406
rect 308290 303170 308374 303406
rect 308610 303170 308732 303406
rect 304732 303086 308732 303170
rect 304732 302850 304854 303086
rect 305090 302850 305174 303086
rect 305410 302850 305494 303086
rect 305730 302850 305814 303086
rect 306050 302850 306134 303086
rect 306370 302850 306454 303086
rect 306690 302850 306774 303086
rect 307010 302850 307094 303086
rect 307330 302850 307414 303086
rect 307650 302850 307734 303086
rect 307970 302850 308054 303086
rect 308290 302850 308374 303086
rect 308610 302850 308732 303086
rect 304732 302766 308732 302850
rect 304732 302530 304854 302766
rect 305090 302530 305174 302766
rect 305410 302530 305494 302766
rect 305730 302530 305814 302766
rect 306050 302530 306134 302766
rect 306370 302530 306454 302766
rect 306690 302530 306774 302766
rect 307010 302530 307094 302766
rect 307330 302530 307414 302766
rect 307650 302530 307734 302766
rect 307970 302530 308054 302766
rect 308290 302530 308374 302766
rect 308610 302530 308732 302766
rect 304732 299842 308732 302530
rect 304732 299606 304854 299842
rect 305090 299606 305174 299842
rect 305410 299606 305494 299842
rect 305730 299606 305814 299842
rect 306050 299606 306134 299842
rect 306370 299606 306454 299842
rect 306690 299606 306774 299842
rect 307010 299606 307094 299842
rect 307330 299606 307414 299842
rect 307650 299606 307734 299842
rect 307970 299606 308054 299842
rect 308290 299606 308374 299842
rect 308610 299606 308732 299842
rect 131395 288268 131461 288269
rect 131395 288204 131396 288268
rect 131460 288204 131461 288268
rect 131395 288203 131461 288204
rect 223579 288268 223645 288269
rect 223579 288204 223580 288268
rect 223644 288204 223645 288268
rect 223579 288203 223645 288204
rect 90179 287796 90180 287846
rect 90244 287796 90245 287846
rect 90179 287795 90245 287796
rect 129555 287796 129556 287846
rect 129620 287796 129621 287846
rect 129555 287795 129621 287796
rect 5000 268970 5122 269206
rect 5358 268970 5442 269206
rect 5678 268970 5762 269206
rect 5998 268970 6082 269206
rect 6318 268970 6402 269206
rect 6638 268970 6722 269206
rect 6958 268970 7042 269206
rect 7278 268970 7362 269206
rect 7598 268970 7682 269206
rect 7918 268970 8002 269206
rect 8238 268970 8322 269206
rect 8558 268970 8642 269206
rect 8878 268970 9000 269206
rect 5000 238570 9000 268970
rect 52459 265556 52525 265557
rect 52459 265492 52460 265556
rect 52524 265492 52525 265556
rect 52459 265491 52525 265492
rect 52275 263788 52341 263789
rect 52275 263724 52276 263788
rect 52340 263724 52341 263788
rect 52275 263723 52341 263724
rect 5000 238334 5122 238570
rect 5358 238334 5442 238570
rect 5678 238334 5762 238570
rect 5998 238334 6082 238570
rect 6318 238334 6402 238570
rect 6638 238334 6722 238570
rect 6958 238334 7042 238570
rect 7278 238334 7362 238570
rect 7598 238334 7682 238570
rect 7918 238334 8002 238570
rect 8238 238334 8322 238570
rect 8558 238334 8642 238570
rect 8878 238334 9000 238570
rect 5000 207934 9000 238334
rect 38107 218772 38173 218773
rect 38107 218708 38108 218772
rect 38172 218708 38173 218772
rect 38107 218707 38173 218708
rect 5000 207698 5122 207934
rect 5358 207698 5442 207934
rect 5678 207698 5762 207934
rect 5998 207698 6082 207934
rect 6318 207698 6402 207934
rect 6638 207698 6722 207934
rect 6958 207698 7042 207934
rect 7278 207698 7362 207934
rect 7598 207698 7682 207934
rect 7918 207698 8002 207934
rect 8238 207698 8322 207934
rect 8558 207698 8642 207934
rect 8878 207698 9000 207934
rect 5000 177298 9000 207698
rect 38110 203082 38170 218707
rect 52278 216189 52338 263723
rect 52275 216188 52341 216189
rect 52275 216124 52276 216188
rect 52340 216124 52341 216188
rect 52275 216123 52341 216124
rect 52462 202997 52522 265491
rect 69755 224212 69821 224213
rect 69755 224148 69756 224212
rect 69820 224148 69821 224212
rect 69755 224147 69821 224148
rect 69758 215322 69818 224147
rect 52459 202996 52525 202997
rect 52459 202932 52460 202996
rect 52524 202932 52525 202996
rect 52459 202931 52525 202932
rect 35899 202116 35900 202166
rect 35964 202116 35965 202166
rect 35899 202115 35965 202116
rect 5000 177062 5122 177298
rect 5358 177062 5442 177298
rect 5678 177062 5762 177298
rect 5998 177062 6082 177298
rect 6318 177062 6402 177298
rect 6638 177062 6722 177298
rect 6958 177062 7042 177298
rect 7278 177062 7362 177298
rect 7598 177062 7682 177298
rect 7918 177062 8002 177298
rect 8238 177062 8322 177298
rect 8558 177062 8642 177298
rect 8878 177062 9000 177298
rect 5000 146662 9000 177062
rect 85027 174708 85093 174709
rect 85027 174644 85028 174708
rect 85092 174644 85093 174708
rect 85027 174643 85093 174644
rect 5000 146426 5122 146662
rect 5358 146426 5442 146662
rect 5678 146426 5762 146662
rect 5998 146426 6082 146662
rect 6318 146426 6402 146662
rect 6638 146426 6722 146662
rect 6958 146426 7042 146662
rect 7278 146426 7362 146662
rect 7598 146426 7682 146662
rect 7918 146426 8002 146662
rect 8238 146426 8322 146662
rect 8558 146426 8642 146662
rect 8878 146426 9000 146662
rect 5000 116026 9000 146426
rect 48227 144108 48293 144109
rect 48227 144044 48228 144108
rect 48292 144044 48293 144108
rect 48227 144043 48293 144044
rect 48230 142562 48290 144043
rect 20811 131596 20877 131597
rect 20811 131532 20812 131596
rect 20876 131532 20877 131596
rect 20811 131531 20877 131532
rect 20814 130322 20874 131531
rect 48230 123301 48290 142326
rect 69755 130372 69821 130373
rect 69755 130308 69756 130372
rect 69820 130308 69821 130372
rect 69755 130307 69821 130308
rect 61475 130236 61541 130237
rect 61475 130172 61476 130236
rect 61540 130172 61541 130236
rect 61475 130171 61541 130172
rect 48598 129557 48658 130086
rect 61478 129642 61538 130171
rect 48595 129556 48661 129557
rect 48595 129492 48596 129556
rect 48660 129492 48661 129556
rect 48595 129491 48661 129492
rect 48227 123300 48293 123301
rect 48227 123236 48228 123300
rect 48292 123236 48293 123300
rect 48227 123235 48293 123236
rect 69758 121482 69818 130307
rect 5000 115790 5122 116026
rect 5358 115790 5442 116026
rect 5678 115790 5762 116026
rect 5998 115790 6082 116026
rect 6318 115790 6402 116026
rect 6638 115790 6722 116026
rect 6958 115790 7042 116026
rect 7278 115790 7362 116026
rect 7598 115790 7682 116026
rect 7918 115790 8002 116026
rect 8238 115790 8322 116026
rect 8558 115790 8642 116026
rect 8878 115790 9000 116026
rect 5000 85390 9000 115790
rect 35899 108276 35900 108326
rect 35964 108276 35965 108326
rect 35899 108275 35965 108276
rect 5000 85154 5122 85390
rect 5358 85154 5442 85390
rect 5678 85154 5762 85390
rect 5998 85154 6082 85390
rect 6318 85154 6402 85390
rect 6638 85154 6722 85390
rect 6958 85154 7042 85390
rect 7278 85154 7362 85390
rect 7598 85154 7682 85390
rect 7918 85154 8002 85390
rect 8238 85154 8322 85390
rect 8558 85154 8642 85390
rect 8878 85154 9000 85390
rect 5000 54754 9000 85154
rect 85030 84133 85090 174643
rect 128451 174572 128517 174573
rect 128451 174508 128452 174572
rect 128516 174508 128517 174572
rect 128451 174507 128517 174508
rect 109499 143972 109565 143973
rect 109499 143908 109500 143972
rect 109564 143908 109565 143972
rect 109499 143907 109565 143908
rect 109502 142562 109562 143907
rect 128454 139893 128514 174507
rect 128451 139892 128517 139893
rect 128451 139828 128452 139892
rect 128516 139828 128517 139892
rect 128451 139827 128517 139828
rect 85027 84132 85093 84133
rect 85027 84068 85028 84132
rect 85092 84068 85093 84132
rect 85027 84067 85093 84068
rect 103979 77876 104045 77877
rect 103979 77812 103980 77876
rect 104044 77812 104045 77876
rect 103979 77811 104045 77812
rect 103982 68354 104042 77811
rect 103982 68294 104410 68354
rect 5000 54518 5122 54754
rect 5358 54518 5442 54754
rect 5678 54518 5762 54754
rect 5998 54518 6082 54754
rect 6318 54518 6402 54754
rect 6638 54518 6722 54754
rect 6958 54518 7042 54754
rect 7278 54518 7362 54754
rect 7598 54518 7682 54754
rect 7918 54518 8002 54754
rect 8238 54518 8322 54754
rect 8558 54518 8642 54754
rect 8878 54518 9000 54754
rect 5000 24118 9000 54518
rect 104350 53805 104410 68294
rect 104347 53804 104413 53805
rect 104347 53740 104348 53804
rect 104412 53740 104413 53804
rect 104347 53739 104413 53740
rect 5000 23882 5122 24118
rect 5358 23882 5442 24118
rect 5678 23882 5762 24118
rect 5998 23882 6082 24118
rect 6318 23882 6402 24118
rect 6638 23882 6722 24118
rect 6958 23882 7042 24118
rect 7278 23882 7362 24118
rect 7598 23882 7682 24118
rect 7918 23882 8002 24118
rect 8238 23882 8322 24118
rect 8558 23882 8642 24118
rect 8878 23882 9000 24118
rect 5000 8878 9000 23882
rect 131398 12189 131458 288203
rect 223582 288082 223642 288203
rect 184203 287796 184204 287846
rect 184268 287796 184269 287846
rect 184203 287795 184269 287796
rect 304732 269206 308732 299606
rect 304732 268970 304854 269206
rect 305090 268970 305174 269206
rect 305410 268970 305494 269206
rect 305730 268970 305814 269206
rect 306050 268970 306134 269206
rect 306370 268970 306454 269206
rect 306690 268970 306774 269206
rect 307010 268970 307094 269206
rect 307330 268970 307414 269206
rect 307650 268970 307734 269206
rect 307970 268970 308054 269206
rect 308290 268970 308374 269206
rect 308610 268970 308732 269206
rect 142251 263788 142317 263789
rect 142251 263724 142252 263788
rect 142316 263724 142317 263788
rect 142251 263723 142317 263724
rect 142254 240533 142314 263723
rect 226339 257668 226405 257669
rect 226339 257604 226340 257668
rect 226404 257604 226405 257668
rect 226339 257603 226405 257604
rect 226342 256122 226402 257603
rect 265163 256852 265229 256853
rect 265163 256788 265164 256852
rect 265228 256788 265229 256852
rect 265163 256787 265229 256788
rect 265166 256122 265226 256787
rect 142251 240532 142317 240533
rect 142251 240468 142252 240532
rect 142316 240468 142317 240532
rect 142251 240467 142317 240468
rect 241611 221628 241677 221629
rect 241611 221564 241612 221628
rect 241676 221564 241677 221628
rect 241611 221563 241677 221564
rect 164883 212652 164949 212653
rect 164883 212588 164884 212652
rect 164948 212588 164949 212652
rect 164883 212587 164949 212588
rect 164886 211922 164946 212587
rect 228918 202317 228978 202846
rect 228915 202316 228981 202317
rect 228915 202252 228916 202316
rect 228980 202252 228981 202316
rect 228915 202251 228981 202252
rect 241614 181237 241674 221563
rect 265166 216682 265226 255886
rect 304732 238570 308732 268970
rect 304732 238334 304854 238570
rect 305090 238334 305174 238570
rect 305410 238334 305494 238570
rect 305730 238334 305814 238570
rect 306050 238334 306134 238570
rect 306370 238334 306454 238570
rect 306690 238334 306774 238570
rect 307010 238334 307094 238570
rect 307330 238334 307414 238570
rect 307650 238334 307734 238570
rect 307970 238334 308054 238570
rect 308290 238334 308374 238570
rect 308610 238334 308732 238570
rect 265166 216404 265226 216446
rect 304732 207934 308732 238334
rect 304732 207698 304854 207934
rect 305090 207698 305174 207934
rect 305410 207698 305494 207934
rect 305730 207698 305814 207934
rect 306050 207698 306134 207934
rect 306370 207698 306454 207934
rect 306690 207698 306774 207934
rect 307010 207698 307094 207934
rect 307330 207698 307414 207934
rect 307650 207698 307734 207934
rect 307970 207698 308054 207934
rect 308290 207698 308374 207934
rect 308610 207698 308732 207934
rect 258907 202316 258973 202317
rect 258907 202314 258908 202316
rect 258690 202254 258908 202314
rect 258907 202252 258908 202254
rect 258972 202252 258973 202316
rect 258907 202251 258973 202252
rect 241611 181236 241677 181237
rect 241611 181172 241612 181236
rect 241676 181172 241677 181236
rect 241611 181171 241677 181172
rect 304732 177298 308732 207698
rect 304732 177062 304854 177298
rect 305090 177062 305174 177298
rect 305410 177062 305494 177298
rect 305730 177062 305814 177298
rect 306050 177062 306134 177298
rect 306370 177062 306454 177298
rect 306690 177062 306774 177298
rect 307010 177062 307094 177298
rect 307330 177062 307414 177298
rect 307650 177062 307734 177298
rect 307970 177062 308054 177298
rect 308290 177062 308374 177298
rect 308610 177062 308732 177298
rect 133235 174708 133301 174709
rect 133235 174644 133236 174708
rect 133300 174644 133301 174708
rect 133235 174643 133301 174644
rect 133238 83725 133298 174643
rect 304732 146662 308732 177062
rect 304732 146426 304854 146662
rect 305090 146426 305174 146662
rect 305410 146426 305494 146662
rect 305730 146426 305814 146662
rect 306050 146426 306134 146662
rect 306370 146426 306454 146662
rect 306690 146426 306774 146662
rect 307010 146426 307094 146662
rect 307330 146426 307414 146662
rect 307650 146426 307734 146662
rect 307970 146426 308054 146662
rect 308290 146426 308374 146662
rect 308610 146426 308732 146662
rect 264979 138668 265045 138669
rect 264979 138604 264980 138668
rect 265044 138604 265045 138668
rect 264979 138603 265045 138604
rect 138755 130236 138821 130237
rect 138755 130172 138756 130236
rect 138820 130172 138821 130236
rect 138755 130171 138821 130172
rect 138758 129642 138818 130171
rect 245107 130236 245173 130237
rect 245107 130172 245108 130236
rect 245172 130172 245173 130236
rect 245107 130171 245173 130172
rect 245110 129642 245170 130171
rect 241611 127516 241677 127517
rect 241611 127452 241612 127516
rect 241676 127452 241677 127516
rect 241611 127451 241677 127452
rect 229654 120309 229714 120566
rect 229651 120308 229717 120309
rect 229651 120244 229652 120308
rect 229716 120244 229717 120308
rect 229651 120243 229717 120244
rect 241614 87397 241674 127451
rect 264982 122162 265042 138603
rect 288715 130372 288781 130373
rect 288715 130322 288716 130372
rect 288780 130322 288781 130372
rect 269214 129557 269274 130086
rect 269211 129556 269277 129557
rect 269211 129492 269212 129556
rect 269276 129492 269277 129556
rect 269211 129491 269277 129492
rect 264982 120717 265042 121926
rect 264979 120716 265045 120717
rect 264979 120652 264980 120716
rect 265044 120652 265045 120716
rect 264979 120651 265045 120652
rect 304732 116026 308732 146426
rect 304732 115790 304854 116026
rect 305090 115790 305174 116026
rect 305410 115790 305494 116026
rect 305730 115790 305814 116026
rect 306050 115790 306134 116026
rect 306370 115790 306454 116026
rect 306690 115790 306774 116026
rect 307010 115790 307094 116026
rect 307330 115790 307414 116026
rect 307650 115790 307734 116026
rect 307970 115790 308054 116026
rect 308290 115790 308374 116026
rect 308610 115790 308732 116026
rect 241611 87396 241677 87397
rect 241611 87332 241612 87396
rect 241676 87332 241677 87396
rect 241611 87331 241677 87332
rect 304732 85390 308732 115790
rect 304732 85154 304854 85390
rect 305090 85154 305174 85390
rect 305410 85154 305494 85390
rect 305730 85154 305814 85390
rect 306050 85154 306134 85390
rect 306370 85154 306454 85390
rect 306690 85154 306774 85390
rect 307010 85154 307094 85390
rect 307330 85154 307414 85390
rect 307650 85154 307734 85390
rect 307970 85154 308054 85390
rect 308290 85154 308374 85390
rect 308610 85154 308732 85390
rect 133235 83724 133301 83725
rect 133235 83660 133236 83724
rect 133300 83660 133301 83724
rect 133235 83659 133301 83660
rect 182179 83724 182245 83725
rect 182179 83660 182180 83724
rect 182244 83660 182245 83724
rect 182179 83659 182245 83660
rect 144275 81276 144341 81277
rect 144275 81212 144276 81276
rect 144340 81212 144341 81276
rect 144275 81211 144341 81212
rect 144278 46053 144338 81211
rect 144275 46052 144341 46053
rect 144275 45988 144276 46052
rect 144340 45988 144341 46052
rect 144275 45987 144341 45988
rect 182182 27557 182242 83659
rect 237011 81412 237077 81413
rect 237011 81348 237012 81412
rect 237076 81348 237077 81412
rect 237011 81347 237077 81348
rect 236827 81276 236893 81277
rect 236827 81212 236828 81276
rect 236892 81212 236893 81276
rect 236827 81211 236893 81212
rect 236830 47549 236890 81211
rect 236827 47548 236893 47549
rect 236827 47484 236828 47548
rect 236892 47484 236893 47548
rect 236827 47483 236893 47484
rect 237014 45917 237074 81347
rect 304732 54754 308732 85154
rect 304732 54518 304854 54754
rect 305090 54518 305174 54754
rect 305410 54518 305494 54754
rect 305730 54518 305814 54754
rect 306050 54518 306134 54754
rect 306370 54518 306454 54754
rect 306690 54518 306774 54754
rect 307010 54518 307094 54754
rect 307330 54518 307414 54754
rect 307650 54518 307734 54754
rect 307970 54518 308054 54754
rect 308290 54518 308374 54754
rect 308610 54518 308732 54754
rect 237011 45916 237077 45917
rect 237011 45852 237012 45916
rect 237076 45852 237077 45916
rect 237011 45851 237077 45852
rect 218611 34492 218677 34493
rect 218611 34428 218612 34492
rect 218676 34428 218677 34492
rect 218611 34427 218677 34428
rect 182179 27556 182245 27557
rect 182179 27492 182180 27556
rect 182244 27492 182245 27556
rect 182179 27491 182245 27492
rect 218614 12325 218674 34427
rect 304732 24118 308732 54518
rect 304732 23882 304854 24118
rect 305090 23882 305174 24118
rect 305410 23882 305494 24118
rect 305730 23882 305814 24118
rect 306050 23882 306134 24118
rect 306370 23882 306454 24118
rect 306690 23882 306774 24118
rect 307010 23882 307094 24118
rect 307330 23882 307414 24118
rect 307650 23882 307734 24118
rect 307970 23882 308054 24118
rect 308290 23882 308374 24118
rect 308610 23882 308732 24118
rect 218611 12324 218677 12325
rect 218611 12260 218612 12324
rect 218676 12260 218677 12324
rect 218611 12259 218677 12260
rect 131395 12188 131461 12189
rect 131395 12124 131396 12188
rect 131460 12124 131461 12188
rect 131395 12123 131461 12124
rect 5000 8642 5122 8878
rect 5358 8642 5442 8878
rect 5678 8642 5762 8878
rect 5998 8642 6082 8878
rect 6318 8642 6402 8878
rect 6638 8642 6722 8878
rect 6958 8642 7042 8878
rect 7278 8642 7362 8878
rect 7598 8642 7682 8878
rect 7918 8642 8002 8878
rect 8238 8642 8322 8878
rect 8558 8642 8642 8878
rect 8878 8642 9000 8878
rect 5000 8558 9000 8642
rect 5000 8322 5122 8558
rect 5358 8322 5442 8558
rect 5678 8322 5762 8558
rect 5998 8322 6082 8558
rect 6318 8322 6402 8558
rect 6638 8322 6722 8558
rect 6958 8322 7042 8558
rect 7278 8322 7362 8558
rect 7598 8322 7682 8558
rect 7918 8322 8002 8558
rect 8238 8322 8322 8558
rect 8558 8322 8642 8558
rect 8878 8322 9000 8558
rect 5000 8238 9000 8322
rect 5000 8002 5122 8238
rect 5358 8002 5442 8238
rect 5678 8002 5762 8238
rect 5998 8002 6082 8238
rect 6318 8002 6402 8238
rect 6638 8002 6722 8238
rect 6958 8002 7042 8238
rect 7278 8002 7362 8238
rect 7598 8002 7682 8238
rect 7918 8002 8002 8238
rect 8238 8002 8322 8238
rect 8558 8002 8642 8238
rect 8878 8002 9000 8238
rect 5000 7918 9000 8002
rect 5000 7682 5122 7918
rect 5358 7682 5442 7918
rect 5678 7682 5762 7918
rect 5998 7682 6082 7918
rect 6318 7682 6402 7918
rect 6638 7682 6722 7918
rect 6958 7682 7042 7918
rect 7278 7682 7362 7918
rect 7598 7682 7682 7918
rect 7918 7682 8002 7918
rect 8238 7682 8322 7918
rect 8558 7682 8642 7918
rect 8878 7682 9000 7918
rect 5000 7598 9000 7682
rect 5000 7362 5122 7598
rect 5358 7362 5442 7598
rect 5678 7362 5762 7598
rect 5998 7362 6082 7598
rect 6318 7362 6402 7598
rect 6638 7362 6722 7598
rect 6958 7362 7042 7598
rect 7278 7362 7362 7598
rect 7598 7362 7682 7598
rect 7918 7362 8002 7598
rect 8238 7362 8322 7598
rect 8558 7362 8642 7598
rect 8878 7362 9000 7598
rect 5000 7278 9000 7362
rect 5000 7042 5122 7278
rect 5358 7042 5442 7278
rect 5678 7042 5762 7278
rect 5998 7042 6082 7278
rect 6318 7042 6402 7278
rect 6638 7042 6722 7278
rect 6958 7042 7042 7278
rect 7278 7042 7362 7278
rect 7598 7042 7682 7278
rect 7918 7042 8002 7278
rect 8238 7042 8322 7278
rect 8558 7042 8642 7278
rect 8878 7042 9000 7278
rect 5000 6958 9000 7042
rect 5000 6722 5122 6958
rect 5358 6722 5442 6958
rect 5678 6722 5762 6958
rect 5998 6722 6082 6958
rect 6318 6722 6402 6958
rect 6638 6722 6722 6958
rect 6958 6722 7042 6958
rect 7278 6722 7362 6958
rect 7598 6722 7682 6958
rect 7918 6722 8002 6958
rect 8238 6722 8322 6958
rect 8558 6722 8642 6958
rect 8878 6722 9000 6958
rect 5000 6638 9000 6722
rect 5000 6402 5122 6638
rect 5358 6402 5442 6638
rect 5678 6402 5762 6638
rect 5998 6402 6082 6638
rect 6318 6402 6402 6638
rect 6638 6402 6722 6638
rect 6958 6402 7042 6638
rect 7278 6402 7362 6638
rect 7598 6402 7682 6638
rect 7918 6402 8002 6638
rect 8238 6402 8322 6638
rect 8558 6402 8642 6638
rect 8878 6402 9000 6638
rect 5000 6318 9000 6402
rect 5000 6082 5122 6318
rect 5358 6082 5442 6318
rect 5678 6082 5762 6318
rect 5998 6082 6082 6318
rect 6318 6082 6402 6318
rect 6638 6082 6722 6318
rect 6958 6082 7042 6318
rect 7278 6082 7362 6318
rect 7598 6082 7682 6318
rect 7918 6082 8002 6318
rect 8238 6082 8322 6318
rect 8558 6082 8642 6318
rect 8878 6082 9000 6318
rect 5000 5998 9000 6082
rect 5000 5762 5122 5998
rect 5358 5762 5442 5998
rect 5678 5762 5762 5998
rect 5998 5762 6082 5998
rect 6318 5762 6402 5998
rect 6638 5762 6722 5998
rect 6958 5762 7042 5998
rect 7278 5762 7362 5998
rect 7598 5762 7682 5998
rect 7918 5762 8002 5998
rect 8238 5762 8322 5998
rect 8558 5762 8642 5998
rect 8878 5762 9000 5998
rect 5000 5678 9000 5762
rect 5000 5442 5122 5678
rect 5358 5442 5442 5678
rect 5678 5442 5762 5678
rect 5998 5442 6082 5678
rect 6318 5442 6402 5678
rect 6638 5442 6722 5678
rect 6958 5442 7042 5678
rect 7278 5442 7362 5678
rect 7598 5442 7682 5678
rect 7918 5442 8002 5678
rect 8238 5442 8322 5678
rect 8558 5442 8642 5678
rect 8878 5442 9000 5678
rect 5000 5358 9000 5442
rect 5000 5122 5122 5358
rect 5358 5122 5442 5358
rect 5678 5122 5762 5358
rect 5998 5122 6082 5358
rect 6318 5122 6402 5358
rect 6638 5122 6722 5358
rect 6958 5122 7042 5358
rect 7278 5122 7362 5358
rect 7598 5122 7682 5358
rect 7918 5122 8002 5358
rect 8238 5122 8322 5358
rect 8558 5122 8642 5358
rect 8878 5122 9000 5358
rect 5000 5000 9000 5122
rect 304732 8878 308732 23882
rect 304732 8642 304854 8878
rect 305090 8642 305174 8878
rect 305410 8642 305494 8878
rect 305730 8642 305814 8878
rect 306050 8642 306134 8878
rect 306370 8642 306454 8878
rect 306690 8642 306774 8878
rect 307010 8642 307094 8878
rect 307330 8642 307414 8878
rect 307650 8642 307734 8878
rect 307970 8642 308054 8878
rect 308290 8642 308374 8878
rect 308610 8642 308732 8878
rect 304732 8558 308732 8642
rect 304732 8322 304854 8558
rect 305090 8322 305174 8558
rect 305410 8322 305494 8558
rect 305730 8322 305814 8558
rect 306050 8322 306134 8558
rect 306370 8322 306454 8558
rect 306690 8322 306774 8558
rect 307010 8322 307094 8558
rect 307330 8322 307414 8558
rect 307650 8322 307734 8558
rect 307970 8322 308054 8558
rect 308290 8322 308374 8558
rect 308610 8322 308732 8558
rect 304732 8238 308732 8322
rect 304732 8002 304854 8238
rect 305090 8002 305174 8238
rect 305410 8002 305494 8238
rect 305730 8002 305814 8238
rect 306050 8002 306134 8238
rect 306370 8002 306454 8238
rect 306690 8002 306774 8238
rect 307010 8002 307094 8238
rect 307330 8002 307414 8238
rect 307650 8002 307734 8238
rect 307970 8002 308054 8238
rect 308290 8002 308374 8238
rect 308610 8002 308732 8238
rect 304732 7918 308732 8002
rect 304732 7682 304854 7918
rect 305090 7682 305174 7918
rect 305410 7682 305494 7918
rect 305730 7682 305814 7918
rect 306050 7682 306134 7918
rect 306370 7682 306454 7918
rect 306690 7682 306774 7918
rect 307010 7682 307094 7918
rect 307330 7682 307414 7918
rect 307650 7682 307734 7918
rect 307970 7682 308054 7918
rect 308290 7682 308374 7918
rect 308610 7682 308732 7918
rect 304732 7598 308732 7682
rect 304732 7362 304854 7598
rect 305090 7362 305174 7598
rect 305410 7362 305494 7598
rect 305730 7362 305814 7598
rect 306050 7362 306134 7598
rect 306370 7362 306454 7598
rect 306690 7362 306774 7598
rect 307010 7362 307094 7598
rect 307330 7362 307414 7598
rect 307650 7362 307734 7598
rect 307970 7362 308054 7598
rect 308290 7362 308374 7598
rect 308610 7362 308732 7598
rect 304732 7278 308732 7362
rect 304732 7042 304854 7278
rect 305090 7042 305174 7278
rect 305410 7042 305494 7278
rect 305730 7042 305814 7278
rect 306050 7042 306134 7278
rect 306370 7042 306454 7278
rect 306690 7042 306774 7278
rect 307010 7042 307094 7278
rect 307330 7042 307414 7278
rect 307650 7042 307734 7278
rect 307970 7042 308054 7278
rect 308290 7042 308374 7278
rect 308610 7042 308732 7278
rect 304732 6958 308732 7042
rect 304732 6722 304854 6958
rect 305090 6722 305174 6958
rect 305410 6722 305494 6958
rect 305730 6722 305814 6958
rect 306050 6722 306134 6958
rect 306370 6722 306454 6958
rect 306690 6722 306774 6958
rect 307010 6722 307094 6958
rect 307330 6722 307414 6958
rect 307650 6722 307734 6958
rect 307970 6722 308054 6958
rect 308290 6722 308374 6958
rect 308610 6722 308732 6958
rect 304732 6638 308732 6722
rect 304732 6402 304854 6638
rect 305090 6402 305174 6638
rect 305410 6402 305494 6638
rect 305730 6402 305814 6638
rect 306050 6402 306134 6638
rect 306370 6402 306454 6638
rect 306690 6402 306774 6638
rect 307010 6402 307094 6638
rect 307330 6402 307414 6638
rect 307650 6402 307734 6638
rect 307970 6402 308054 6638
rect 308290 6402 308374 6638
rect 308610 6402 308732 6638
rect 304732 6318 308732 6402
rect 304732 6082 304854 6318
rect 305090 6082 305174 6318
rect 305410 6082 305494 6318
rect 305730 6082 305814 6318
rect 306050 6082 306134 6318
rect 306370 6082 306454 6318
rect 306690 6082 306774 6318
rect 307010 6082 307094 6318
rect 307330 6082 307414 6318
rect 307650 6082 307734 6318
rect 307970 6082 308054 6318
rect 308290 6082 308374 6318
rect 308610 6082 308732 6318
rect 304732 5998 308732 6082
rect 304732 5762 304854 5998
rect 305090 5762 305174 5998
rect 305410 5762 305494 5998
rect 305730 5762 305814 5998
rect 306050 5762 306134 5998
rect 306370 5762 306454 5998
rect 306690 5762 306774 5998
rect 307010 5762 307094 5998
rect 307330 5762 307414 5998
rect 307650 5762 307734 5998
rect 307970 5762 308054 5998
rect 308290 5762 308374 5998
rect 308610 5762 308732 5998
rect 304732 5678 308732 5762
rect 304732 5442 304854 5678
rect 305090 5442 305174 5678
rect 305410 5442 305494 5678
rect 305730 5442 305814 5678
rect 306050 5442 306134 5678
rect 306370 5442 306454 5678
rect 306690 5442 306774 5678
rect 307010 5442 307094 5678
rect 307330 5442 307414 5678
rect 307650 5442 307734 5678
rect 307970 5442 308054 5678
rect 308290 5442 308374 5678
rect 308610 5442 308732 5678
rect 304732 5358 308732 5442
rect 304732 5122 304854 5358
rect 305090 5122 305174 5358
rect 305410 5122 305494 5358
rect 305730 5122 305814 5358
rect 306050 5122 306134 5358
rect 306370 5122 306454 5358
rect 306690 5122 306774 5358
rect 307010 5122 307094 5358
rect 307330 5122 307414 5358
rect 307650 5122 307734 5358
rect 307970 5122 308054 5358
rect 308290 5122 308374 5358
rect 308610 5122 308732 5358
rect 304732 5000 308732 5122
rect 309732 284524 313732 307530
rect 309732 284288 309854 284524
rect 310090 284288 310174 284524
rect 310410 284288 310494 284524
rect 310730 284288 310814 284524
rect 311050 284288 311134 284524
rect 311370 284288 311454 284524
rect 311690 284288 311774 284524
rect 312010 284288 312094 284524
rect 312330 284288 312414 284524
rect 312650 284288 312734 284524
rect 312970 284288 313054 284524
rect 313290 284288 313374 284524
rect 313610 284288 313732 284524
rect 309732 253888 313732 284288
rect 309732 253652 309854 253888
rect 310090 253652 310174 253888
rect 310410 253652 310494 253888
rect 310730 253652 310814 253888
rect 311050 253652 311134 253888
rect 311370 253652 311454 253888
rect 311690 253652 311774 253888
rect 312010 253652 312094 253888
rect 312330 253652 312414 253888
rect 312650 253652 312734 253888
rect 312970 253652 313054 253888
rect 313290 253652 313374 253888
rect 313610 253652 313732 253888
rect 309732 223252 313732 253652
rect 309732 223016 309854 223252
rect 310090 223016 310174 223252
rect 310410 223016 310494 223252
rect 310730 223016 310814 223252
rect 311050 223016 311134 223252
rect 311370 223016 311454 223252
rect 311690 223016 311774 223252
rect 312010 223016 312094 223252
rect 312330 223016 312414 223252
rect 312650 223016 312734 223252
rect 312970 223016 313054 223252
rect 313290 223016 313374 223252
rect 313610 223016 313732 223252
rect 309732 192616 313732 223016
rect 309732 192380 309854 192616
rect 310090 192380 310174 192616
rect 310410 192380 310494 192616
rect 310730 192380 310814 192616
rect 311050 192380 311134 192616
rect 311370 192380 311454 192616
rect 311690 192380 311774 192616
rect 312010 192380 312094 192616
rect 312330 192380 312414 192616
rect 312650 192380 312734 192616
rect 312970 192380 313054 192616
rect 313290 192380 313374 192616
rect 313610 192380 313732 192616
rect 309732 161980 313732 192380
rect 309732 161744 309854 161980
rect 310090 161744 310174 161980
rect 310410 161744 310494 161980
rect 310730 161744 310814 161980
rect 311050 161744 311134 161980
rect 311370 161744 311454 161980
rect 311690 161744 311774 161980
rect 312010 161744 312094 161980
rect 312330 161744 312414 161980
rect 312650 161744 312734 161980
rect 312970 161744 313054 161980
rect 313290 161744 313374 161980
rect 313610 161744 313732 161980
rect 309732 131344 313732 161744
rect 309732 131108 309854 131344
rect 310090 131108 310174 131344
rect 310410 131108 310494 131344
rect 310730 131108 310814 131344
rect 311050 131108 311134 131344
rect 311370 131108 311454 131344
rect 311690 131108 311774 131344
rect 312010 131108 312094 131344
rect 312330 131108 312414 131344
rect 312650 131108 312734 131344
rect 312970 131108 313054 131344
rect 313290 131108 313374 131344
rect 313610 131108 313732 131344
rect 309732 100708 313732 131108
rect 309732 100472 309854 100708
rect 310090 100472 310174 100708
rect 310410 100472 310494 100708
rect 310730 100472 310814 100708
rect 311050 100472 311134 100708
rect 311370 100472 311454 100708
rect 311690 100472 311774 100708
rect 312010 100472 312094 100708
rect 312330 100472 312414 100708
rect 312650 100472 312734 100708
rect 312970 100472 313054 100708
rect 313290 100472 313374 100708
rect 313610 100472 313732 100708
rect 309732 70072 313732 100472
rect 309732 69836 309854 70072
rect 310090 69836 310174 70072
rect 310410 69836 310494 70072
rect 310730 69836 310814 70072
rect 311050 69836 311134 70072
rect 311370 69836 311454 70072
rect 311690 69836 311774 70072
rect 312010 69836 312094 70072
rect 312330 69836 312414 70072
rect 312650 69836 312734 70072
rect 312970 69836 313054 70072
rect 313290 69836 313374 70072
rect 313610 69836 313732 70072
rect 309732 39436 313732 69836
rect 309732 39200 309854 39436
rect 310090 39200 310174 39436
rect 310410 39200 310494 39436
rect 310730 39200 310814 39436
rect 311050 39200 311134 39436
rect 311370 39200 311454 39436
rect 311690 39200 311774 39436
rect 312010 39200 312094 39436
rect 312330 39200 312414 39436
rect 312650 39200 312734 39436
rect 312970 39200 313054 39436
rect 313290 39200 313374 39436
rect 313610 39200 313732 39436
rect 0 3642 122 3878
rect 358 3642 442 3878
rect 678 3642 762 3878
rect 998 3642 1082 3878
rect 1318 3642 1402 3878
rect 1638 3642 1722 3878
rect 1958 3642 2042 3878
rect 2278 3642 2362 3878
rect 2598 3642 2682 3878
rect 2918 3642 3002 3878
rect 3238 3642 3322 3878
rect 3558 3642 3642 3878
rect 3878 3642 4000 3878
rect 0 3558 4000 3642
rect 0 3322 122 3558
rect 358 3322 442 3558
rect 678 3322 762 3558
rect 998 3322 1082 3558
rect 1318 3322 1402 3558
rect 1638 3322 1722 3558
rect 1958 3322 2042 3558
rect 2278 3322 2362 3558
rect 2598 3322 2682 3558
rect 2918 3322 3002 3558
rect 3238 3322 3322 3558
rect 3558 3322 3642 3558
rect 3878 3322 4000 3558
rect 0 3238 4000 3322
rect 0 3002 122 3238
rect 358 3002 442 3238
rect 678 3002 762 3238
rect 998 3002 1082 3238
rect 1318 3002 1402 3238
rect 1638 3002 1722 3238
rect 1958 3002 2042 3238
rect 2278 3002 2362 3238
rect 2598 3002 2682 3238
rect 2918 3002 3002 3238
rect 3238 3002 3322 3238
rect 3558 3002 3642 3238
rect 3878 3002 4000 3238
rect 0 2918 4000 3002
rect 0 2682 122 2918
rect 358 2682 442 2918
rect 678 2682 762 2918
rect 998 2682 1082 2918
rect 1318 2682 1402 2918
rect 1638 2682 1722 2918
rect 1958 2682 2042 2918
rect 2278 2682 2362 2918
rect 2598 2682 2682 2918
rect 2918 2682 3002 2918
rect 3238 2682 3322 2918
rect 3558 2682 3642 2918
rect 3878 2682 4000 2918
rect 0 2598 4000 2682
rect 0 2362 122 2598
rect 358 2362 442 2598
rect 678 2362 762 2598
rect 998 2362 1082 2598
rect 1318 2362 1402 2598
rect 1638 2362 1722 2598
rect 1958 2362 2042 2598
rect 2278 2362 2362 2598
rect 2598 2362 2682 2598
rect 2918 2362 3002 2598
rect 3238 2362 3322 2598
rect 3558 2362 3642 2598
rect 3878 2362 4000 2598
rect 0 2278 4000 2362
rect 0 2042 122 2278
rect 358 2042 442 2278
rect 678 2042 762 2278
rect 998 2042 1082 2278
rect 1318 2042 1402 2278
rect 1638 2042 1722 2278
rect 1958 2042 2042 2278
rect 2278 2042 2362 2278
rect 2598 2042 2682 2278
rect 2918 2042 3002 2278
rect 3238 2042 3322 2278
rect 3558 2042 3642 2278
rect 3878 2042 4000 2278
rect 0 1958 4000 2042
rect 0 1722 122 1958
rect 358 1722 442 1958
rect 678 1722 762 1958
rect 998 1722 1082 1958
rect 1318 1722 1402 1958
rect 1638 1722 1722 1958
rect 1958 1722 2042 1958
rect 2278 1722 2362 1958
rect 2598 1722 2682 1958
rect 2918 1722 3002 1958
rect 3238 1722 3322 1958
rect 3558 1722 3642 1958
rect 3878 1722 4000 1958
rect 0 1638 4000 1722
rect 0 1402 122 1638
rect 358 1402 442 1638
rect 678 1402 762 1638
rect 998 1402 1082 1638
rect 1318 1402 1402 1638
rect 1638 1402 1722 1638
rect 1958 1402 2042 1638
rect 2278 1402 2362 1638
rect 2598 1402 2682 1638
rect 2918 1402 3002 1638
rect 3238 1402 3322 1638
rect 3558 1402 3642 1638
rect 3878 1402 4000 1638
rect 0 1318 4000 1402
rect 0 1082 122 1318
rect 358 1082 442 1318
rect 678 1082 762 1318
rect 998 1082 1082 1318
rect 1318 1082 1402 1318
rect 1638 1082 1722 1318
rect 1958 1082 2042 1318
rect 2278 1082 2362 1318
rect 2598 1082 2682 1318
rect 2918 1082 3002 1318
rect 3238 1082 3322 1318
rect 3558 1082 3642 1318
rect 3878 1082 4000 1318
rect 0 998 4000 1082
rect 0 762 122 998
rect 358 762 442 998
rect 678 762 762 998
rect 998 762 1082 998
rect 1318 762 1402 998
rect 1638 762 1722 998
rect 1958 762 2042 998
rect 2278 762 2362 998
rect 2598 762 2682 998
rect 2918 762 3002 998
rect 3238 762 3322 998
rect 3558 762 3642 998
rect 3878 762 4000 998
rect 0 678 4000 762
rect 0 442 122 678
rect 358 442 442 678
rect 678 442 762 678
rect 998 442 1082 678
rect 1318 442 1402 678
rect 1638 442 1722 678
rect 1958 442 2042 678
rect 2278 442 2362 678
rect 2598 442 2682 678
rect 2918 442 3002 678
rect 3238 442 3322 678
rect 3558 442 3642 678
rect 3878 442 4000 678
rect 0 358 4000 442
rect 0 122 122 358
rect 358 122 442 358
rect 678 122 762 358
rect 998 122 1082 358
rect 1318 122 1402 358
rect 1638 122 1722 358
rect 1958 122 2042 358
rect 2278 122 2362 358
rect 2598 122 2682 358
rect 2918 122 3002 358
rect 3238 122 3322 358
rect 3558 122 3642 358
rect 3878 122 4000 358
rect 0 0 4000 122
rect 309732 3878 313732 39200
rect 309732 3642 309854 3878
rect 310090 3642 310174 3878
rect 310410 3642 310494 3878
rect 310730 3642 310814 3878
rect 311050 3642 311134 3878
rect 311370 3642 311454 3878
rect 311690 3642 311774 3878
rect 312010 3642 312094 3878
rect 312330 3642 312414 3878
rect 312650 3642 312734 3878
rect 312970 3642 313054 3878
rect 313290 3642 313374 3878
rect 313610 3642 313732 3878
rect 309732 3558 313732 3642
rect 309732 3322 309854 3558
rect 310090 3322 310174 3558
rect 310410 3322 310494 3558
rect 310730 3322 310814 3558
rect 311050 3322 311134 3558
rect 311370 3322 311454 3558
rect 311690 3322 311774 3558
rect 312010 3322 312094 3558
rect 312330 3322 312414 3558
rect 312650 3322 312734 3558
rect 312970 3322 313054 3558
rect 313290 3322 313374 3558
rect 313610 3322 313732 3558
rect 309732 3238 313732 3322
rect 309732 3002 309854 3238
rect 310090 3002 310174 3238
rect 310410 3002 310494 3238
rect 310730 3002 310814 3238
rect 311050 3002 311134 3238
rect 311370 3002 311454 3238
rect 311690 3002 311774 3238
rect 312010 3002 312094 3238
rect 312330 3002 312414 3238
rect 312650 3002 312734 3238
rect 312970 3002 313054 3238
rect 313290 3002 313374 3238
rect 313610 3002 313732 3238
rect 309732 2918 313732 3002
rect 309732 2682 309854 2918
rect 310090 2682 310174 2918
rect 310410 2682 310494 2918
rect 310730 2682 310814 2918
rect 311050 2682 311134 2918
rect 311370 2682 311454 2918
rect 311690 2682 311774 2918
rect 312010 2682 312094 2918
rect 312330 2682 312414 2918
rect 312650 2682 312734 2918
rect 312970 2682 313054 2918
rect 313290 2682 313374 2918
rect 313610 2682 313732 2918
rect 309732 2598 313732 2682
rect 309732 2362 309854 2598
rect 310090 2362 310174 2598
rect 310410 2362 310494 2598
rect 310730 2362 310814 2598
rect 311050 2362 311134 2598
rect 311370 2362 311454 2598
rect 311690 2362 311774 2598
rect 312010 2362 312094 2598
rect 312330 2362 312414 2598
rect 312650 2362 312734 2598
rect 312970 2362 313054 2598
rect 313290 2362 313374 2598
rect 313610 2362 313732 2598
rect 309732 2278 313732 2362
rect 309732 2042 309854 2278
rect 310090 2042 310174 2278
rect 310410 2042 310494 2278
rect 310730 2042 310814 2278
rect 311050 2042 311134 2278
rect 311370 2042 311454 2278
rect 311690 2042 311774 2278
rect 312010 2042 312094 2278
rect 312330 2042 312414 2278
rect 312650 2042 312734 2278
rect 312970 2042 313054 2278
rect 313290 2042 313374 2278
rect 313610 2042 313732 2278
rect 309732 1958 313732 2042
rect 309732 1722 309854 1958
rect 310090 1722 310174 1958
rect 310410 1722 310494 1958
rect 310730 1722 310814 1958
rect 311050 1722 311134 1958
rect 311370 1722 311454 1958
rect 311690 1722 311774 1958
rect 312010 1722 312094 1958
rect 312330 1722 312414 1958
rect 312650 1722 312734 1958
rect 312970 1722 313054 1958
rect 313290 1722 313374 1958
rect 313610 1722 313732 1958
rect 309732 1638 313732 1722
rect 309732 1402 309854 1638
rect 310090 1402 310174 1638
rect 310410 1402 310494 1638
rect 310730 1402 310814 1638
rect 311050 1402 311134 1638
rect 311370 1402 311454 1638
rect 311690 1402 311774 1638
rect 312010 1402 312094 1638
rect 312330 1402 312414 1638
rect 312650 1402 312734 1638
rect 312970 1402 313054 1638
rect 313290 1402 313374 1638
rect 313610 1402 313732 1638
rect 309732 1318 313732 1402
rect 309732 1082 309854 1318
rect 310090 1082 310174 1318
rect 310410 1082 310494 1318
rect 310730 1082 310814 1318
rect 311050 1082 311134 1318
rect 311370 1082 311454 1318
rect 311690 1082 311774 1318
rect 312010 1082 312094 1318
rect 312330 1082 312414 1318
rect 312650 1082 312734 1318
rect 312970 1082 313054 1318
rect 313290 1082 313374 1318
rect 313610 1082 313732 1318
rect 309732 998 313732 1082
rect 309732 762 309854 998
rect 310090 762 310174 998
rect 310410 762 310494 998
rect 310730 762 310814 998
rect 311050 762 311134 998
rect 311370 762 311454 998
rect 311690 762 311774 998
rect 312010 762 312094 998
rect 312330 762 312414 998
rect 312650 762 312734 998
rect 312970 762 313054 998
rect 313290 762 313374 998
rect 313610 762 313732 998
rect 309732 678 313732 762
rect 309732 442 309854 678
rect 310090 442 310174 678
rect 310410 442 310494 678
rect 310730 442 310814 678
rect 311050 442 311134 678
rect 311370 442 311454 678
rect 311690 442 311774 678
rect 312010 442 312094 678
rect 312330 442 312414 678
rect 312650 442 312734 678
rect 312970 442 313054 678
rect 313290 442 313374 678
rect 313610 442 313732 678
rect 309732 358 313732 442
rect 309732 122 309854 358
rect 310090 122 310174 358
rect 310410 122 310494 358
rect 310730 122 310814 358
rect 311050 122 311134 358
rect 311370 122 311454 358
rect 311690 122 311774 358
rect 312010 122 312094 358
rect 312330 122 312414 358
rect 312650 122 312734 358
rect 312970 122 313054 358
rect 313290 122 313374 358
rect 313610 122 313732 358
rect 309732 0 313732 122
<< via4 >>
rect 122 311050 358 311286
rect 442 311050 678 311286
rect 762 311050 998 311286
rect 1082 311050 1318 311286
rect 1402 311050 1638 311286
rect 1722 311050 1958 311286
rect 2042 311050 2278 311286
rect 2362 311050 2598 311286
rect 2682 311050 2918 311286
rect 3002 311050 3238 311286
rect 3322 311050 3558 311286
rect 3642 311050 3878 311286
rect 122 310730 358 310966
rect 442 310730 678 310966
rect 762 310730 998 310966
rect 1082 310730 1318 310966
rect 1402 310730 1638 310966
rect 1722 310730 1958 310966
rect 2042 310730 2278 310966
rect 2362 310730 2598 310966
rect 2682 310730 2918 310966
rect 3002 310730 3238 310966
rect 3322 310730 3558 310966
rect 3642 310730 3878 310966
rect 122 310410 358 310646
rect 442 310410 678 310646
rect 762 310410 998 310646
rect 1082 310410 1318 310646
rect 1402 310410 1638 310646
rect 1722 310410 1958 310646
rect 2042 310410 2278 310646
rect 2362 310410 2598 310646
rect 2682 310410 2918 310646
rect 3002 310410 3238 310646
rect 3322 310410 3558 310646
rect 3642 310410 3878 310646
rect 122 310090 358 310326
rect 442 310090 678 310326
rect 762 310090 998 310326
rect 1082 310090 1318 310326
rect 1402 310090 1638 310326
rect 1722 310090 1958 310326
rect 2042 310090 2278 310326
rect 2362 310090 2598 310326
rect 2682 310090 2918 310326
rect 3002 310090 3238 310326
rect 3322 310090 3558 310326
rect 3642 310090 3878 310326
rect 122 309770 358 310006
rect 442 309770 678 310006
rect 762 309770 998 310006
rect 1082 309770 1318 310006
rect 1402 309770 1638 310006
rect 1722 309770 1958 310006
rect 2042 309770 2278 310006
rect 2362 309770 2598 310006
rect 2682 309770 2918 310006
rect 3002 309770 3238 310006
rect 3322 309770 3558 310006
rect 3642 309770 3878 310006
rect 122 309450 358 309686
rect 442 309450 678 309686
rect 762 309450 998 309686
rect 1082 309450 1318 309686
rect 1402 309450 1638 309686
rect 1722 309450 1958 309686
rect 2042 309450 2278 309686
rect 2362 309450 2598 309686
rect 2682 309450 2918 309686
rect 3002 309450 3238 309686
rect 3322 309450 3558 309686
rect 3642 309450 3878 309686
rect 122 309130 358 309366
rect 442 309130 678 309366
rect 762 309130 998 309366
rect 1082 309130 1318 309366
rect 1402 309130 1638 309366
rect 1722 309130 1958 309366
rect 2042 309130 2278 309366
rect 2362 309130 2598 309366
rect 2682 309130 2918 309366
rect 3002 309130 3238 309366
rect 3322 309130 3558 309366
rect 3642 309130 3878 309366
rect 122 308810 358 309046
rect 442 308810 678 309046
rect 762 308810 998 309046
rect 1082 308810 1318 309046
rect 1402 308810 1638 309046
rect 1722 308810 1958 309046
rect 2042 308810 2278 309046
rect 2362 308810 2598 309046
rect 2682 308810 2918 309046
rect 3002 308810 3238 309046
rect 3322 308810 3558 309046
rect 3642 308810 3878 309046
rect 122 308490 358 308726
rect 442 308490 678 308726
rect 762 308490 998 308726
rect 1082 308490 1318 308726
rect 1402 308490 1638 308726
rect 1722 308490 1958 308726
rect 2042 308490 2278 308726
rect 2362 308490 2598 308726
rect 2682 308490 2918 308726
rect 3002 308490 3238 308726
rect 3322 308490 3558 308726
rect 3642 308490 3878 308726
rect 122 308170 358 308406
rect 442 308170 678 308406
rect 762 308170 998 308406
rect 1082 308170 1318 308406
rect 1402 308170 1638 308406
rect 1722 308170 1958 308406
rect 2042 308170 2278 308406
rect 2362 308170 2598 308406
rect 2682 308170 2918 308406
rect 3002 308170 3238 308406
rect 3322 308170 3558 308406
rect 3642 308170 3878 308406
rect 122 307850 358 308086
rect 442 307850 678 308086
rect 762 307850 998 308086
rect 1082 307850 1318 308086
rect 1402 307850 1638 308086
rect 1722 307850 1958 308086
rect 2042 307850 2278 308086
rect 2362 307850 2598 308086
rect 2682 307850 2918 308086
rect 3002 307850 3238 308086
rect 3322 307850 3558 308086
rect 3642 307850 3878 308086
rect 122 307530 358 307766
rect 442 307530 678 307766
rect 762 307530 998 307766
rect 1082 307530 1318 307766
rect 1402 307530 1638 307766
rect 1722 307530 1958 307766
rect 2042 307530 2278 307766
rect 2362 307530 2598 307766
rect 2682 307530 2918 307766
rect 3002 307530 3238 307766
rect 3322 307530 3558 307766
rect 3642 307530 3878 307766
rect 309854 311050 310090 311286
rect 310174 311050 310410 311286
rect 310494 311050 310730 311286
rect 310814 311050 311050 311286
rect 311134 311050 311370 311286
rect 311454 311050 311690 311286
rect 311774 311050 312010 311286
rect 312094 311050 312330 311286
rect 312414 311050 312650 311286
rect 312734 311050 312970 311286
rect 313054 311050 313290 311286
rect 313374 311050 313610 311286
rect 309854 310730 310090 310966
rect 310174 310730 310410 310966
rect 310494 310730 310730 310966
rect 310814 310730 311050 310966
rect 311134 310730 311370 310966
rect 311454 310730 311690 310966
rect 311774 310730 312010 310966
rect 312094 310730 312330 310966
rect 312414 310730 312650 310966
rect 312734 310730 312970 310966
rect 313054 310730 313290 310966
rect 313374 310730 313610 310966
rect 309854 310410 310090 310646
rect 310174 310410 310410 310646
rect 310494 310410 310730 310646
rect 310814 310410 311050 310646
rect 311134 310410 311370 310646
rect 311454 310410 311690 310646
rect 311774 310410 312010 310646
rect 312094 310410 312330 310646
rect 312414 310410 312650 310646
rect 312734 310410 312970 310646
rect 313054 310410 313290 310646
rect 313374 310410 313610 310646
rect 309854 310090 310090 310326
rect 310174 310090 310410 310326
rect 310494 310090 310730 310326
rect 310814 310090 311050 310326
rect 311134 310090 311370 310326
rect 311454 310090 311690 310326
rect 311774 310090 312010 310326
rect 312094 310090 312330 310326
rect 312414 310090 312650 310326
rect 312734 310090 312970 310326
rect 313054 310090 313290 310326
rect 313374 310090 313610 310326
rect 309854 309770 310090 310006
rect 310174 309770 310410 310006
rect 310494 309770 310730 310006
rect 310814 309770 311050 310006
rect 311134 309770 311370 310006
rect 311454 309770 311690 310006
rect 311774 309770 312010 310006
rect 312094 309770 312330 310006
rect 312414 309770 312650 310006
rect 312734 309770 312970 310006
rect 313054 309770 313290 310006
rect 313374 309770 313610 310006
rect 309854 309450 310090 309686
rect 310174 309450 310410 309686
rect 310494 309450 310730 309686
rect 310814 309450 311050 309686
rect 311134 309450 311370 309686
rect 311454 309450 311690 309686
rect 311774 309450 312010 309686
rect 312094 309450 312330 309686
rect 312414 309450 312650 309686
rect 312734 309450 312970 309686
rect 313054 309450 313290 309686
rect 313374 309450 313610 309686
rect 309854 309130 310090 309366
rect 310174 309130 310410 309366
rect 310494 309130 310730 309366
rect 310814 309130 311050 309366
rect 311134 309130 311370 309366
rect 311454 309130 311690 309366
rect 311774 309130 312010 309366
rect 312094 309130 312330 309366
rect 312414 309130 312650 309366
rect 312734 309130 312970 309366
rect 313054 309130 313290 309366
rect 313374 309130 313610 309366
rect 309854 308810 310090 309046
rect 310174 308810 310410 309046
rect 310494 308810 310730 309046
rect 310814 308810 311050 309046
rect 311134 308810 311370 309046
rect 311454 308810 311690 309046
rect 311774 308810 312010 309046
rect 312094 308810 312330 309046
rect 312414 308810 312650 309046
rect 312734 308810 312970 309046
rect 313054 308810 313290 309046
rect 313374 308810 313610 309046
rect 309854 308490 310090 308726
rect 310174 308490 310410 308726
rect 310494 308490 310730 308726
rect 310814 308490 311050 308726
rect 311134 308490 311370 308726
rect 311454 308490 311690 308726
rect 311774 308490 312010 308726
rect 312094 308490 312330 308726
rect 312414 308490 312650 308726
rect 312734 308490 312970 308726
rect 313054 308490 313290 308726
rect 313374 308490 313610 308726
rect 309854 308170 310090 308406
rect 310174 308170 310410 308406
rect 310494 308170 310730 308406
rect 310814 308170 311050 308406
rect 311134 308170 311370 308406
rect 311454 308170 311690 308406
rect 311774 308170 312010 308406
rect 312094 308170 312330 308406
rect 312414 308170 312650 308406
rect 312734 308170 312970 308406
rect 313054 308170 313290 308406
rect 313374 308170 313610 308406
rect 309854 307850 310090 308086
rect 310174 307850 310410 308086
rect 310494 307850 310730 308086
rect 310814 307850 311050 308086
rect 311134 307850 311370 308086
rect 311454 307850 311690 308086
rect 311774 307850 312010 308086
rect 312094 307850 312330 308086
rect 312414 307850 312650 308086
rect 312734 307850 312970 308086
rect 313054 307850 313290 308086
rect 313374 307850 313610 308086
rect 309854 307530 310090 307766
rect 310174 307530 310410 307766
rect 310494 307530 310730 307766
rect 310814 307530 311050 307766
rect 311134 307530 311370 307766
rect 311454 307530 311690 307766
rect 311774 307530 312010 307766
rect 312094 307530 312330 307766
rect 312414 307530 312650 307766
rect 312734 307530 312970 307766
rect 313054 307530 313290 307766
rect 313374 307530 313610 307766
rect 122 284288 358 284524
rect 442 284288 678 284524
rect 762 284288 998 284524
rect 1082 284288 1318 284524
rect 1402 284288 1638 284524
rect 1722 284288 1958 284524
rect 2042 284288 2278 284524
rect 2362 284288 2598 284524
rect 2682 284288 2918 284524
rect 3002 284288 3238 284524
rect 3322 284288 3558 284524
rect 3642 284288 3878 284524
rect 122 253652 358 253888
rect 442 253652 678 253888
rect 762 253652 998 253888
rect 1082 253652 1318 253888
rect 1402 253652 1638 253888
rect 1722 253652 1958 253888
rect 2042 253652 2278 253888
rect 2362 253652 2598 253888
rect 2682 253652 2918 253888
rect 3002 253652 3238 253888
rect 3322 253652 3558 253888
rect 3642 253652 3878 253888
rect 122 223016 358 223252
rect 442 223016 678 223252
rect 762 223016 998 223252
rect 1082 223016 1318 223252
rect 1402 223016 1638 223252
rect 1722 223016 1958 223252
rect 2042 223016 2278 223252
rect 2362 223016 2598 223252
rect 2682 223016 2918 223252
rect 3002 223016 3238 223252
rect 3322 223016 3558 223252
rect 3642 223016 3878 223252
rect 122 192380 358 192616
rect 442 192380 678 192616
rect 762 192380 998 192616
rect 1082 192380 1318 192616
rect 1402 192380 1638 192616
rect 1722 192380 1958 192616
rect 2042 192380 2278 192616
rect 2362 192380 2598 192616
rect 2682 192380 2918 192616
rect 3002 192380 3238 192616
rect 3322 192380 3558 192616
rect 3642 192380 3878 192616
rect 122 161744 358 161980
rect 442 161744 678 161980
rect 762 161744 998 161980
rect 1082 161744 1318 161980
rect 1402 161744 1638 161980
rect 1722 161744 1958 161980
rect 2042 161744 2278 161980
rect 2362 161744 2598 161980
rect 2682 161744 2918 161980
rect 3002 161744 3238 161980
rect 3322 161744 3558 161980
rect 3642 161744 3878 161980
rect 122 131108 358 131344
rect 442 131108 678 131344
rect 762 131108 998 131344
rect 1082 131108 1318 131344
rect 1402 131108 1638 131344
rect 1722 131108 1958 131344
rect 2042 131108 2278 131344
rect 2362 131108 2598 131344
rect 2682 131108 2918 131344
rect 3002 131108 3238 131344
rect 3322 131108 3558 131344
rect 3642 131108 3878 131344
rect 122 100472 358 100708
rect 442 100472 678 100708
rect 762 100472 998 100708
rect 1082 100472 1318 100708
rect 1402 100472 1638 100708
rect 1722 100472 1958 100708
rect 2042 100472 2278 100708
rect 2362 100472 2598 100708
rect 2682 100472 2918 100708
rect 3002 100472 3238 100708
rect 3322 100472 3558 100708
rect 3642 100472 3878 100708
rect 122 69836 358 70072
rect 442 69836 678 70072
rect 762 69836 998 70072
rect 1082 69836 1318 70072
rect 1402 69836 1638 70072
rect 1722 69836 1958 70072
rect 2042 69836 2278 70072
rect 2362 69836 2598 70072
rect 2682 69836 2918 70072
rect 3002 69836 3238 70072
rect 3322 69836 3558 70072
rect 3642 69836 3878 70072
rect 122 39200 358 39436
rect 442 39200 678 39436
rect 762 39200 998 39436
rect 1082 39200 1318 39436
rect 1402 39200 1638 39436
rect 1722 39200 1958 39436
rect 2042 39200 2278 39436
rect 2362 39200 2598 39436
rect 2682 39200 2918 39436
rect 3002 39200 3238 39436
rect 3322 39200 3558 39436
rect 3642 39200 3878 39436
rect 5122 306050 5358 306286
rect 5442 306050 5678 306286
rect 5762 306050 5998 306286
rect 6082 306050 6318 306286
rect 6402 306050 6638 306286
rect 6722 306050 6958 306286
rect 7042 306050 7278 306286
rect 7362 306050 7598 306286
rect 7682 306050 7918 306286
rect 8002 306050 8238 306286
rect 8322 306050 8558 306286
rect 8642 306050 8878 306286
rect 5122 305730 5358 305966
rect 5442 305730 5678 305966
rect 5762 305730 5998 305966
rect 6082 305730 6318 305966
rect 6402 305730 6638 305966
rect 6722 305730 6958 305966
rect 7042 305730 7278 305966
rect 7362 305730 7598 305966
rect 7682 305730 7918 305966
rect 8002 305730 8238 305966
rect 8322 305730 8558 305966
rect 8642 305730 8878 305966
rect 5122 305410 5358 305646
rect 5442 305410 5678 305646
rect 5762 305410 5998 305646
rect 6082 305410 6318 305646
rect 6402 305410 6638 305646
rect 6722 305410 6958 305646
rect 7042 305410 7278 305646
rect 7362 305410 7598 305646
rect 7682 305410 7918 305646
rect 8002 305410 8238 305646
rect 8322 305410 8558 305646
rect 8642 305410 8878 305646
rect 5122 305090 5358 305326
rect 5442 305090 5678 305326
rect 5762 305090 5998 305326
rect 6082 305090 6318 305326
rect 6402 305090 6638 305326
rect 6722 305090 6958 305326
rect 7042 305090 7278 305326
rect 7362 305090 7598 305326
rect 7682 305090 7918 305326
rect 8002 305090 8238 305326
rect 8322 305090 8558 305326
rect 8642 305090 8878 305326
rect 5122 304770 5358 305006
rect 5442 304770 5678 305006
rect 5762 304770 5998 305006
rect 6082 304770 6318 305006
rect 6402 304770 6638 305006
rect 6722 304770 6958 305006
rect 7042 304770 7278 305006
rect 7362 304770 7598 305006
rect 7682 304770 7918 305006
rect 8002 304770 8238 305006
rect 8322 304770 8558 305006
rect 8642 304770 8878 305006
rect 5122 304450 5358 304686
rect 5442 304450 5678 304686
rect 5762 304450 5998 304686
rect 6082 304450 6318 304686
rect 6402 304450 6638 304686
rect 6722 304450 6958 304686
rect 7042 304450 7278 304686
rect 7362 304450 7598 304686
rect 7682 304450 7918 304686
rect 8002 304450 8238 304686
rect 8322 304450 8558 304686
rect 8642 304450 8878 304686
rect 5122 304130 5358 304366
rect 5442 304130 5678 304366
rect 5762 304130 5998 304366
rect 6082 304130 6318 304366
rect 6402 304130 6638 304366
rect 6722 304130 6958 304366
rect 7042 304130 7278 304366
rect 7362 304130 7598 304366
rect 7682 304130 7918 304366
rect 8002 304130 8238 304366
rect 8322 304130 8558 304366
rect 8642 304130 8878 304366
rect 5122 303810 5358 304046
rect 5442 303810 5678 304046
rect 5762 303810 5998 304046
rect 6082 303810 6318 304046
rect 6402 303810 6638 304046
rect 6722 303810 6958 304046
rect 7042 303810 7278 304046
rect 7362 303810 7598 304046
rect 7682 303810 7918 304046
rect 8002 303810 8238 304046
rect 8322 303810 8558 304046
rect 8642 303810 8878 304046
rect 5122 303490 5358 303726
rect 5442 303490 5678 303726
rect 5762 303490 5998 303726
rect 6082 303490 6318 303726
rect 6402 303490 6638 303726
rect 6722 303490 6958 303726
rect 7042 303490 7278 303726
rect 7362 303490 7598 303726
rect 7682 303490 7918 303726
rect 8002 303490 8238 303726
rect 8322 303490 8558 303726
rect 8642 303490 8878 303726
rect 5122 303170 5358 303406
rect 5442 303170 5678 303406
rect 5762 303170 5998 303406
rect 6082 303170 6318 303406
rect 6402 303170 6638 303406
rect 6722 303170 6958 303406
rect 7042 303170 7278 303406
rect 7362 303170 7598 303406
rect 7682 303170 7918 303406
rect 8002 303170 8238 303406
rect 8322 303170 8558 303406
rect 8642 303170 8878 303406
rect 5122 302850 5358 303086
rect 5442 302850 5678 303086
rect 5762 302850 5998 303086
rect 6082 302850 6318 303086
rect 6402 302850 6638 303086
rect 6722 302850 6958 303086
rect 7042 302850 7278 303086
rect 7362 302850 7598 303086
rect 7682 302850 7918 303086
rect 8002 302850 8238 303086
rect 8322 302850 8558 303086
rect 8642 302850 8878 303086
rect 5122 302530 5358 302766
rect 5442 302530 5678 302766
rect 5762 302530 5998 302766
rect 6082 302530 6318 302766
rect 6402 302530 6638 302766
rect 6722 302530 6958 302766
rect 7042 302530 7278 302766
rect 7362 302530 7598 302766
rect 7682 302530 7918 302766
rect 8002 302530 8238 302766
rect 8322 302530 8558 302766
rect 8642 302530 8878 302766
rect 5122 299606 5358 299842
rect 5442 299606 5678 299842
rect 5762 299606 5998 299842
rect 6082 299606 6318 299842
rect 6402 299606 6638 299842
rect 6722 299606 6958 299842
rect 7042 299606 7278 299842
rect 7362 299606 7598 299842
rect 7682 299606 7918 299842
rect 8002 299606 8238 299842
rect 8322 299606 8558 299842
rect 8642 299606 8878 299842
rect 304854 306050 305090 306286
rect 305174 306050 305410 306286
rect 305494 306050 305730 306286
rect 305814 306050 306050 306286
rect 306134 306050 306370 306286
rect 306454 306050 306690 306286
rect 306774 306050 307010 306286
rect 307094 306050 307330 306286
rect 307414 306050 307650 306286
rect 307734 306050 307970 306286
rect 308054 306050 308290 306286
rect 308374 306050 308610 306286
rect 304854 305730 305090 305966
rect 305174 305730 305410 305966
rect 305494 305730 305730 305966
rect 305814 305730 306050 305966
rect 306134 305730 306370 305966
rect 306454 305730 306690 305966
rect 306774 305730 307010 305966
rect 307094 305730 307330 305966
rect 307414 305730 307650 305966
rect 307734 305730 307970 305966
rect 308054 305730 308290 305966
rect 308374 305730 308610 305966
rect 304854 305410 305090 305646
rect 305174 305410 305410 305646
rect 305494 305410 305730 305646
rect 305814 305410 306050 305646
rect 306134 305410 306370 305646
rect 306454 305410 306690 305646
rect 306774 305410 307010 305646
rect 307094 305410 307330 305646
rect 307414 305410 307650 305646
rect 307734 305410 307970 305646
rect 308054 305410 308290 305646
rect 308374 305410 308610 305646
rect 304854 305090 305090 305326
rect 305174 305090 305410 305326
rect 305494 305090 305730 305326
rect 305814 305090 306050 305326
rect 306134 305090 306370 305326
rect 306454 305090 306690 305326
rect 306774 305090 307010 305326
rect 307094 305090 307330 305326
rect 307414 305090 307650 305326
rect 307734 305090 307970 305326
rect 308054 305090 308290 305326
rect 308374 305090 308610 305326
rect 304854 304770 305090 305006
rect 305174 304770 305410 305006
rect 305494 304770 305730 305006
rect 305814 304770 306050 305006
rect 306134 304770 306370 305006
rect 306454 304770 306690 305006
rect 306774 304770 307010 305006
rect 307094 304770 307330 305006
rect 307414 304770 307650 305006
rect 307734 304770 307970 305006
rect 308054 304770 308290 305006
rect 308374 304770 308610 305006
rect 304854 304450 305090 304686
rect 305174 304450 305410 304686
rect 305494 304450 305730 304686
rect 305814 304450 306050 304686
rect 306134 304450 306370 304686
rect 306454 304450 306690 304686
rect 306774 304450 307010 304686
rect 307094 304450 307330 304686
rect 307414 304450 307650 304686
rect 307734 304450 307970 304686
rect 308054 304450 308290 304686
rect 308374 304450 308610 304686
rect 304854 304130 305090 304366
rect 305174 304130 305410 304366
rect 305494 304130 305730 304366
rect 305814 304130 306050 304366
rect 306134 304130 306370 304366
rect 306454 304130 306690 304366
rect 306774 304130 307010 304366
rect 307094 304130 307330 304366
rect 307414 304130 307650 304366
rect 307734 304130 307970 304366
rect 308054 304130 308290 304366
rect 308374 304130 308610 304366
rect 304854 303810 305090 304046
rect 305174 303810 305410 304046
rect 305494 303810 305730 304046
rect 305814 303810 306050 304046
rect 306134 303810 306370 304046
rect 306454 303810 306690 304046
rect 306774 303810 307010 304046
rect 307094 303810 307330 304046
rect 307414 303810 307650 304046
rect 307734 303810 307970 304046
rect 308054 303810 308290 304046
rect 308374 303810 308610 304046
rect 304854 303490 305090 303726
rect 305174 303490 305410 303726
rect 305494 303490 305730 303726
rect 305814 303490 306050 303726
rect 306134 303490 306370 303726
rect 306454 303490 306690 303726
rect 306774 303490 307010 303726
rect 307094 303490 307330 303726
rect 307414 303490 307650 303726
rect 307734 303490 307970 303726
rect 308054 303490 308290 303726
rect 308374 303490 308610 303726
rect 304854 303170 305090 303406
rect 305174 303170 305410 303406
rect 305494 303170 305730 303406
rect 305814 303170 306050 303406
rect 306134 303170 306370 303406
rect 306454 303170 306690 303406
rect 306774 303170 307010 303406
rect 307094 303170 307330 303406
rect 307414 303170 307650 303406
rect 307734 303170 307970 303406
rect 308054 303170 308290 303406
rect 308374 303170 308610 303406
rect 304854 302850 305090 303086
rect 305174 302850 305410 303086
rect 305494 302850 305730 303086
rect 305814 302850 306050 303086
rect 306134 302850 306370 303086
rect 306454 302850 306690 303086
rect 306774 302850 307010 303086
rect 307094 302850 307330 303086
rect 307414 302850 307650 303086
rect 307734 302850 307970 303086
rect 308054 302850 308290 303086
rect 308374 302850 308610 303086
rect 304854 302530 305090 302766
rect 305174 302530 305410 302766
rect 305494 302530 305730 302766
rect 305814 302530 306050 302766
rect 306134 302530 306370 302766
rect 306454 302530 306690 302766
rect 306774 302530 307010 302766
rect 307094 302530 307330 302766
rect 307414 302530 307650 302766
rect 307734 302530 307970 302766
rect 308054 302530 308290 302766
rect 308374 302530 308610 302766
rect 304854 299606 305090 299842
rect 305174 299606 305410 299842
rect 305494 299606 305730 299842
rect 305814 299606 306050 299842
rect 306134 299606 306370 299842
rect 306454 299606 306690 299842
rect 306774 299606 307010 299842
rect 307094 299606 307330 299842
rect 307414 299606 307650 299842
rect 307734 299606 307970 299842
rect 308054 299606 308290 299842
rect 308374 299606 308610 299842
rect 90094 287860 90330 288082
rect 90094 287846 90180 287860
rect 90180 287846 90244 287860
rect 90244 287846 90330 287860
rect 129470 287860 129706 288082
rect 129470 287846 129556 287860
rect 129556 287846 129620 287860
rect 129620 287846 129706 287860
rect 5122 268970 5358 269206
rect 5442 268970 5678 269206
rect 5762 268970 5998 269206
rect 6082 268970 6318 269206
rect 6402 268970 6638 269206
rect 6722 268970 6958 269206
rect 7042 268970 7278 269206
rect 7362 268970 7598 269206
rect 7682 268970 7918 269206
rect 8002 268970 8238 269206
rect 8322 268970 8558 269206
rect 8642 268970 8878 269206
rect 5122 238334 5358 238570
rect 5442 238334 5678 238570
rect 5762 238334 5998 238570
rect 6082 238334 6318 238570
rect 6402 238334 6638 238570
rect 6722 238334 6958 238570
rect 7042 238334 7278 238570
rect 7362 238334 7598 238570
rect 7682 238334 7918 238570
rect 8002 238334 8238 238570
rect 8322 238334 8558 238570
rect 8642 238334 8878 238570
rect 5122 207698 5358 207934
rect 5442 207698 5678 207934
rect 5762 207698 5998 207934
rect 6082 207698 6318 207934
rect 6402 207698 6638 207934
rect 6722 207698 6958 207934
rect 7042 207698 7278 207934
rect 7362 207698 7598 207934
rect 7682 207698 7918 207934
rect 8002 207698 8238 207934
rect 8322 207698 8558 207934
rect 8642 207698 8878 207934
rect 38022 202846 38258 203082
rect 69670 215086 69906 215322
rect 81630 215236 81866 215322
rect 81630 215172 81716 215236
rect 81716 215172 81780 215236
rect 81780 215172 81866 215236
rect 81630 215086 81866 215172
rect 19990 202316 20226 202402
rect 19990 202252 20076 202316
rect 20076 202252 20140 202316
rect 20140 202252 20226 202316
rect 19990 202166 20226 202252
rect 35814 202180 36050 202402
rect 35814 202166 35900 202180
rect 35900 202166 35964 202180
rect 35964 202166 36050 202180
rect 5122 177062 5358 177298
rect 5442 177062 5678 177298
rect 5762 177062 5998 177298
rect 6082 177062 6318 177298
rect 6402 177062 6638 177298
rect 6722 177062 6958 177298
rect 7042 177062 7278 177298
rect 7362 177062 7598 177298
rect 7682 177062 7918 177298
rect 8002 177062 8238 177298
rect 8322 177062 8558 177298
rect 8642 177062 8878 177298
rect 5122 146426 5358 146662
rect 5442 146426 5678 146662
rect 5762 146426 5998 146662
rect 6082 146426 6318 146662
rect 6402 146426 6638 146662
rect 6722 146426 6958 146662
rect 7042 146426 7278 146662
rect 7362 146426 7598 146662
rect 7682 146426 7918 146662
rect 8002 146426 8238 146662
rect 8322 146426 8558 146662
rect 8642 146426 8878 146662
rect 48142 142326 48378 142562
rect 20726 130086 20962 130322
rect 48510 130086 48746 130322
rect 58078 130236 58314 130322
rect 58078 130172 58164 130236
rect 58164 130172 58228 130236
rect 58228 130172 58314 130236
rect 58078 130086 58314 130172
rect 57710 129556 57946 129642
rect 57710 129492 57796 129556
rect 57796 129492 57860 129556
rect 57860 129492 57946 129556
rect 57710 129406 57946 129492
rect 61390 129406 61626 129642
rect 69670 121246 69906 121482
rect 81630 121396 81866 121482
rect 81630 121332 81716 121396
rect 81716 121332 81780 121396
rect 81780 121332 81866 121396
rect 81630 121246 81866 121332
rect 5122 115790 5358 116026
rect 5442 115790 5678 116026
rect 5762 115790 5998 116026
rect 6082 115790 6318 116026
rect 6402 115790 6638 116026
rect 6722 115790 6958 116026
rect 7042 115790 7278 116026
rect 7362 115790 7598 116026
rect 7682 115790 7918 116026
rect 8002 115790 8238 116026
rect 8322 115790 8558 116026
rect 8642 115790 8878 116026
rect 19990 108476 20226 108562
rect 19990 108412 20076 108476
rect 20076 108412 20140 108476
rect 20140 108412 20226 108476
rect 19990 108326 20226 108412
rect 35814 108340 36050 108562
rect 35814 108326 35900 108340
rect 35900 108326 35964 108340
rect 35964 108326 36050 108340
rect 5122 85154 5358 85390
rect 5442 85154 5678 85390
rect 5762 85154 5998 85390
rect 6082 85154 6318 85390
rect 6402 85154 6638 85390
rect 6722 85154 6958 85390
rect 7042 85154 7278 85390
rect 7362 85154 7598 85390
rect 7682 85154 7918 85390
rect 8002 85154 8238 85390
rect 8322 85154 8558 85390
rect 8642 85154 8878 85390
rect 109414 142326 109650 142562
rect 5122 54518 5358 54754
rect 5442 54518 5678 54754
rect 5762 54518 5998 54754
rect 6082 54518 6318 54754
rect 6402 54518 6638 54754
rect 6722 54518 6958 54754
rect 7042 54518 7278 54754
rect 7362 54518 7598 54754
rect 7682 54518 7918 54754
rect 8002 54518 8238 54754
rect 8322 54518 8558 54754
rect 8642 54518 8878 54754
rect 5122 23882 5358 24118
rect 5442 23882 5678 24118
rect 5762 23882 5998 24118
rect 6082 23882 6318 24118
rect 6402 23882 6638 24118
rect 6722 23882 6958 24118
rect 7042 23882 7278 24118
rect 7362 23882 7598 24118
rect 7682 23882 7918 24118
rect 8002 23882 8238 24118
rect 8322 23882 8558 24118
rect 8642 23882 8878 24118
rect 184118 287860 184354 288082
rect 184118 287846 184204 287860
rect 184204 287846 184268 287860
rect 184268 287846 184354 287860
rect 223494 287846 223730 288082
rect 304854 268970 305090 269206
rect 305174 268970 305410 269206
rect 305494 268970 305730 269206
rect 305814 268970 306050 269206
rect 306134 268970 306370 269206
rect 306454 268970 306690 269206
rect 306774 268970 307010 269206
rect 307094 268970 307330 269206
rect 307414 268970 307650 269206
rect 307734 268970 307970 269206
rect 308054 268970 308290 269206
rect 308374 268970 308610 269206
rect 226254 255886 226490 256122
rect 265078 255886 265314 256122
rect 135174 211836 135410 211922
rect 135174 211772 135260 211836
rect 135260 211772 135324 211836
rect 135324 211772 135410 211836
rect 135174 211686 135410 211772
rect 164798 211686 165034 211922
rect 228830 202846 229066 203082
rect 304854 238334 305090 238570
rect 305174 238334 305410 238570
rect 305494 238334 305730 238570
rect 305814 238334 306050 238570
rect 306134 238334 306370 238570
rect 306454 238334 306690 238570
rect 306774 238334 307010 238570
rect 307094 238334 307330 238570
rect 307414 238334 307650 238570
rect 307734 238334 307970 238570
rect 308054 238334 308290 238570
rect 308374 238334 308610 238570
rect 265078 216596 265314 216682
rect 265078 216532 265164 216596
rect 265164 216532 265228 216596
rect 265228 216532 265314 216596
rect 265078 216446 265314 216532
rect 293598 216596 293834 216682
rect 293598 216532 293684 216596
rect 293684 216532 293748 216596
rect 293748 216532 293834 216596
rect 293598 216446 293834 216532
rect 304854 207698 305090 207934
rect 305174 207698 305410 207934
rect 305494 207698 305730 207934
rect 305814 207698 306050 207934
rect 306134 207698 306370 207934
rect 306454 207698 306690 207934
rect 306774 207698 307010 207934
rect 307094 207698 307330 207934
rect 307414 207698 307650 207934
rect 307734 207698 307970 207934
rect 308054 207698 308290 207934
rect 308374 207698 308610 207934
rect 242814 202316 243050 202402
rect 242814 202252 242900 202316
rect 242900 202252 242964 202316
rect 242964 202252 243050 202316
rect 242814 202166 243050 202252
rect 258454 202166 258690 202402
rect 277958 202316 278194 202402
rect 277958 202252 278044 202316
rect 278044 202252 278108 202316
rect 278108 202252 278194 202316
rect 277958 202166 278194 202252
rect 293598 202316 293834 202402
rect 293598 202252 293684 202316
rect 293684 202252 293748 202316
rect 293748 202252 293834 202316
rect 293598 202166 293834 202252
rect 304854 177062 305090 177298
rect 305174 177062 305410 177298
rect 305494 177062 305730 177298
rect 305814 177062 306050 177298
rect 306134 177062 306370 177298
rect 306454 177062 306690 177298
rect 306774 177062 307010 177298
rect 307094 177062 307330 177298
rect 307414 177062 307650 177298
rect 307734 177062 307970 177298
rect 308054 177062 308290 177298
rect 308374 177062 308610 177298
rect 304854 146426 305090 146662
rect 305174 146426 305410 146662
rect 305494 146426 305730 146662
rect 305814 146426 306050 146662
rect 306134 146426 306370 146662
rect 306454 146426 306690 146662
rect 306774 146426 307010 146662
rect 307094 146426 307330 146662
rect 307414 146426 307650 146662
rect 307734 146426 307970 146662
rect 308054 146426 308290 146662
rect 308374 146426 308610 146662
rect 135358 130236 135594 130322
rect 135358 130172 135444 130236
rect 135444 130172 135508 130236
rect 135508 130172 135594 130236
rect 135358 130086 135594 130172
rect 243918 130236 244154 130322
rect 243918 130172 244004 130236
rect 244004 130172 244068 130236
rect 244068 130172 244154 130236
rect 243918 130086 244154 130172
rect 138670 129406 138906 129642
rect 245022 129406 245258 129642
rect 251278 129556 251514 129642
rect 251278 129492 251364 129556
rect 251364 129492 251428 129556
rect 251428 129492 251514 129556
rect 251278 129406 251514 129492
rect 229566 120566 229802 120802
rect 269126 130086 269362 130322
rect 288630 130308 288716 130322
rect 288716 130308 288780 130322
rect 288780 130308 288866 130322
rect 288630 130086 288866 130308
rect 264894 121926 265130 122162
rect 293598 122076 293834 122162
rect 293598 122012 293684 122076
rect 293684 122012 293748 122076
rect 293748 122012 293834 122076
rect 293598 121926 293834 122012
rect 261030 120716 261266 120802
rect 261030 120652 261116 120716
rect 261116 120652 261180 120716
rect 261180 120652 261266 120716
rect 261030 120566 261266 120652
rect 304854 115790 305090 116026
rect 305174 115790 305410 116026
rect 305494 115790 305730 116026
rect 305814 115790 306050 116026
rect 306134 115790 306370 116026
rect 306454 115790 306690 116026
rect 306774 115790 307010 116026
rect 307094 115790 307330 116026
rect 307414 115790 307650 116026
rect 307734 115790 307970 116026
rect 308054 115790 308290 116026
rect 308374 115790 308610 116026
rect 304854 85154 305090 85390
rect 305174 85154 305410 85390
rect 305494 85154 305730 85390
rect 305814 85154 306050 85390
rect 306134 85154 306370 85390
rect 306454 85154 306690 85390
rect 306774 85154 307010 85390
rect 307094 85154 307330 85390
rect 307414 85154 307650 85390
rect 307734 85154 307970 85390
rect 308054 85154 308290 85390
rect 308374 85154 308610 85390
rect 304854 54518 305090 54754
rect 305174 54518 305410 54754
rect 305494 54518 305730 54754
rect 305814 54518 306050 54754
rect 306134 54518 306370 54754
rect 306454 54518 306690 54754
rect 306774 54518 307010 54754
rect 307094 54518 307330 54754
rect 307414 54518 307650 54754
rect 307734 54518 307970 54754
rect 308054 54518 308290 54754
rect 308374 54518 308610 54754
rect 304854 23882 305090 24118
rect 305174 23882 305410 24118
rect 305494 23882 305730 24118
rect 305814 23882 306050 24118
rect 306134 23882 306370 24118
rect 306454 23882 306690 24118
rect 306774 23882 307010 24118
rect 307094 23882 307330 24118
rect 307414 23882 307650 24118
rect 307734 23882 307970 24118
rect 308054 23882 308290 24118
rect 308374 23882 308610 24118
rect 5122 8642 5358 8878
rect 5442 8642 5678 8878
rect 5762 8642 5998 8878
rect 6082 8642 6318 8878
rect 6402 8642 6638 8878
rect 6722 8642 6958 8878
rect 7042 8642 7278 8878
rect 7362 8642 7598 8878
rect 7682 8642 7918 8878
rect 8002 8642 8238 8878
rect 8322 8642 8558 8878
rect 8642 8642 8878 8878
rect 5122 8322 5358 8558
rect 5442 8322 5678 8558
rect 5762 8322 5998 8558
rect 6082 8322 6318 8558
rect 6402 8322 6638 8558
rect 6722 8322 6958 8558
rect 7042 8322 7278 8558
rect 7362 8322 7598 8558
rect 7682 8322 7918 8558
rect 8002 8322 8238 8558
rect 8322 8322 8558 8558
rect 8642 8322 8878 8558
rect 5122 8002 5358 8238
rect 5442 8002 5678 8238
rect 5762 8002 5998 8238
rect 6082 8002 6318 8238
rect 6402 8002 6638 8238
rect 6722 8002 6958 8238
rect 7042 8002 7278 8238
rect 7362 8002 7598 8238
rect 7682 8002 7918 8238
rect 8002 8002 8238 8238
rect 8322 8002 8558 8238
rect 8642 8002 8878 8238
rect 5122 7682 5358 7918
rect 5442 7682 5678 7918
rect 5762 7682 5998 7918
rect 6082 7682 6318 7918
rect 6402 7682 6638 7918
rect 6722 7682 6958 7918
rect 7042 7682 7278 7918
rect 7362 7682 7598 7918
rect 7682 7682 7918 7918
rect 8002 7682 8238 7918
rect 8322 7682 8558 7918
rect 8642 7682 8878 7918
rect 5122 7362 5358 7598
rect 5442 7362 5678 7598
rect 5762 7362 5998 7598
rect 6082 7362 6318 7598
rect 6402 7362 6638 7598
rect 6722 7362 6958 7598
rect 7042 7362 7278 7598
rect 7362 7362 7598 7598
rect 7682 7362 7918 7598
rect 8002 7362 8238 7598
rect 8322 7362 8558 7598
rect 8642 7362 8878 7598
rect 5122 7042 5358 7278
rect 5442 7042 5678 7278
rect 5762 7042 5998 7278
rect 6082 7042 6318 7278
rect 6402 7042 6638 7278
rect 6722 7042 6958 7278
rect 7042 7042 7278 7278
rect 7362 7042 7598 7278
rect 7682 7042 7918 7278
rect 8002 7042 8238 7278
rect 8322 7042 8558 7278
rect 8642 7042 8878 7278
rect 5122 6722 5358 6958
rect 5442 6722 5678 6958
rect 5762 6722 5998 6958
rect 6082 6722 6318 6958
rect 6402 6722 6638 6958
rect 6722 6722 6958 6958
rect 7042 6722 7278 6958
rect 7362 6722 7598 6958
rect 7682 6722 7918 6958
rect 8002 6722 8238 6958
rect 8322 6722 8558 6958
rect 8642 6722 8878 6958
rect 5122 6402 5358 6638
rect 5442 6402 5678 6638
rect 5762 6402 5998 6638
rect 6082 6402 6318 6638
rect 6402 6402 6638 6638
rect 6722 6402 6958 6638
rect 7042 6402 7278 6638
rect 7362 6402 7598 6638
rect 7682 6402 7918 6638
rect 8002 6402 8238 6638
rect 8322 6402 8558 6638
rect 8642 6402 8878 6638
rect 5122 6082 5358 6318
rect 5442 6082 5678 6318
rect 5762 6082 5998 6318
rect 6082 6082 6318 6318
rect 6402 6082 6638 6318
rect 6722 6082 6958 6318
rect 7042 6082 7278 6318
rect 7362 6082 7598 6318
rect 7682 6082 7918 6318
rect 8002 6082 8238 6318
rect 8322 6082 8558 6318
rect 8642 6082 8878 6318
rect 5122 5762 5358 5998
rect 5442 5762 5678 5998
rect 5762 5762 5998 5998
rect 6082 5762 6318 5998
rect 6402 5762 6638 5998
rect 6722 5762 6958 5998
rect 7042 5762 7278 5998
rect 7362 5762 7598 5998
rect 7682 5762 7918 5998
rect 8002 5762 8238 5998
rect 8322 5762 8558 5998
rect 8642 5762 8878 5998
rect 5122 5442 5358 5678
rect 5442 5442 5678 5678
rect 5762 5442 5998 5678
rect 6082 5442 6318 5678
rect 6402 5442 6638 5678
rect 6722 5442 6958 5678
rect 7042 5442 7278 5678
rect 7362 5442 7598 5678
rect 7682 5442 7918 5678
rect 8002 5442 8238 5678
rect 8322 5442 8558 5678
rect 8642 5442 8878 5678
rect 5122 5122 5358 5358
rect 5442 5122 5678 5358
rect 5762 5122 5998 5358
rect 6082 5122 6318 5358
rect 6402 5122 6638 5358
rect 6722 5122 6958 5358
rect 7042 5122 7278 5358
rect 7362 5122 7598 5358
rect 7682 5122 7918 5358
rect 8002 5122 8238 5358
rect 8322 5122 8558 5358
rect 8642 5122 8878 5358
rect 304854 8642 305090 8878
rect 305174 8642 305410 8878
rect 305494 8642 305730 8878
rect 305814 8642 306050 8878
rect 306134 8642 306370 8878
rect 306454 8642 306690 8878
rect 306774 8642 307010 8878
rect 307094 8642 307330 8878
rect 307414 8642 307650 8878
rect 307734 8642 307970 8878
rect 308054 8642 308290 8878
rect 308374 8642 308610 8878
rect 304854 8322 305090 8558
rect 305174 8322 305410 8558
rect 305494 8322 305730 8558
rect 305814 8322 306050 8558
rect 306134 8322 306370 8558
rect 306454 8322 306690 8558
rect 306774 8322 307010 8558
rect 307094 8322 307330 8558
rect 307414 8322 307650 8558
rect 307734 8322 307970 8558
rect 308054 8322 308290 8558
rect 308374 8322 308610 8558
rect 304854 8002 305090 8238
rect 305174 8002 305410 8238
rect 305494 8002 305730 8238
rect 305814 8002 306050 8238
rect 306134 8002 306370 8238
rect 306454 8002 306690 8238
rect 306774 8002 307010 8238
rect 307094 8002 307330 8238
rect 307414 8002 307650 8238
rect 307734 8002 307970 8238
rect 308054 8002 308290 8238
rect 308374 8002 308610 8238
rect 304854 7682 305090 7918
rect 305174 7682 305410 7918
rect 305494 7682 305730 7918
rect 305814 7682 306050 7918
rect 306134 7682 306370 7918
rect 306454 7682 306690 7918
rect 306774 7682 307010 7918
rect 307094 7682 307330 7918
rect 307414 7682 307650 7918
rect 307734 7682 307970 7918
rect 308054 7682 308290 7918
rect 308374 7682 308610 7918
rect 304854 7362 305090 7598
rect 305174 7362 305410 7598
rect 305494 7362 305730 7598
rect 305814 7362 306050 7598
rect 306134 7362 306370 7598
rect 306454 7362 306690 7598
rect 306774 7362 307010 7598
rect 307094 7362 307330 7598
rect 307414 7362 307650 7598
rect 307734 7362 307970 7598
rect 308054 7362 308290 7598
rect 308374 7362 308610 7598
rect 304854 7042 305090 7278
rect 305174 7042 305410 7278
rect 305494 7042 305730 7278
rect 305814 7042 306050 7278
rect 306134 7042 306370 7278
rect 306454 7042 306690 7278
rect 306774 7042 307010 7278
rect 307094 7042 307330 7278
rect 307414 7042 307650 7278
rect 307734 7042 307970 7278
rect 308054 7042 308290 7278
rect 308374 7042 308610 7278
rect 304854 6722 305090 6958
rect 305174 6722 305410 6958
rect 305494 6722 305730 6958
rect 305814 6722 306050 6958
rect 306134 6722 306370 6958
rect 306454 6722 306690 6958
rect 306774 6722 307010 6958
rect 307094 6722 307330 6958
rect 307414 6722 307650 6958
rect 307734 6722 307970 6958
rect 308054 6722 308290 6958
rect 308374 6722 308610 6958
rect 304854 6402 305090 6638
rect 305174 6402 305410 6638
rect 305494 6402 305730 6638
rect 305814 6402 306050 6638
rect 306134 6402 306370 6638
rect 306454 6402 306690 6638
rect 306774 6402 307010 6638
rect 307094 6402 307330 6638
rect 307414 6402 307650 6638
rect 307734 6402 307970 6638
rect 308054 6402 308290 6638
rect 308374 6402 308610 6638
rect 304854 6082 305090 6318
rect 305174 6082 305410 6318
rect 305494 6082 305730 6318
rect 305814 6082 306050 6318
rect 306134 6082 306370 6318
rect 306454 6082 306690 6318
rect 306774 6082 307010 6318
rect 307094 6082 307330 6318
rect 307414 6082 307650 6318
rect 307734 6082 307970 6318
rect 308054 6082 308290 6318
rect 308374 6082 308610 6318
rect 304854 5762 305090 5998
rect 305174 5762 305410 5998
rect 305494 5762 305730 5998
rect 305814 5762 306050 5998
rect 306134 5762 306370 5998
rect 306454 5762 306690 5998
rect 306774 5762 307010 5998
rect 307094 5762 307330 5998
rect 307414 5762 307650 5998
rect 307734 5762 307970 5998
rect 308054 5762 308290 5998
rect 308374 5762 308610 5998
rect 304854 5442 305090 5678
rect 305174 5442 305410 5678
rect 305494 5442 305730 5678
rect 305814 5442 306050 5678
rect 306134 5442 306370 5678
rect 306454 5442 306690 5678
rect 306774 5442 307010 5678
rect 307094 5442 307330 5678
rect 307414 5442 307650 5678
rect 307734 5442 307970 5678
rect 308054 5442 308290 5678
rect 308374 5442 308610 5678
rect 304854 5122 305090 5358
rect 305174 5122 305410 5358
rect 305494 5122 305730 5358
rect 305814 5122 306050 5358
rect 306134 5122 306370 5358
rect 306454 5122 306690 5358
rect 306774 5122 307010 5358
rect 307094 5122 307330 5358
rect 307414 5122 307650 5358
rect 307734 5122 307970 5358
rect 308054 5122 308290 5358
rect 308374 5122 308610 5358
rect 309854 284288 310090 284524
rect 310174 284288 310410 284524
rect 310494 284288 310730 284524
rect 310814 284288 311050 284524
rect 311134 284288 311370 284524
rect 311454 284288 311690 284524
rect 311774 284288 312010 284524
rect 312094 284288 312330 284524
rect 312414 284288 312650 284524
rect 312734 284288 312970 284524
rect 313054 284288 313290 284524
rect 313374 284288 313610 284524
rect 309854 253652 310090 253888
rect 310174 253652 310410 253888
rect 310494 253652 310730 253888
rect 310814 253652 311050 253888
rect 311134 253652 311370 253888
rect 311454 253652 311690 253888
rect 311774 253652 312010 253888
rect 312094 253652 312330 253888
rect 312414 253652 312650 253888
rect 312734 253652 312970 253888
rect 313054 253652 313290 253888
rect 313374 253652 313610 253888
rect 309854 223016 310090 223252
rect 310174 223016 310410 223252
rect 310494 223016 310730 223252
rect 310814 223016 311050 223252
rect 311134 223016 311370 223252
rect 311454 223016 311690 223252
rect 311774 223016 312010 223252
rect 312094 223016 312330 223252
rect 312414 223016 312650 223252
rect 312734 223016 312970 223252
rect 313054 223016 313290 223252
rect 313374 223016 313610 223252
rect 309854 192380 310090 192616
rect 310174 192380 310410 192616
rect 310494 192380 310730 192616
rect 310814 192380 311050 192616
rect 311134 192380 311370 192616
rect 311454 192380 311690 192616
rect 311774 192380 312010 192616
rect 312094 192380 312330 192616
rect 312414 192380 312650 192616
rect 312734 192380 312970 192616
rect 313054 192380 313290 192616
rect 313374 192380 313610 192616
rect 309854 161744 310090 161980
rect 310174 161744 310410 161980
rect 310494 161744 310730 161980
rect 310814 161744 311050 161980
rect 311134 161744 311370 161980
rect 311454 161744 311690 161980
rect 311774 161744 312010 161980
rect 312094 161744 312330 161980
rect 312414 161744 312650 161980
rect 312734 161744 312970 161980
rect 313054 161744 313290 161980
rect 313374 161744 313610 161980
rect 309854 131108 310090 131344
rect 310174 131108 310410 131344
rect 310494 131108 310730 131344
rect 310814 131108 311050 131344
rect 311134 131108 311370 131344
rect 311454 131108 311690 131344
rect 311774 131108 312010 131344
rect 312094 131108 312330 131344
rect 312414 131108 312650 131344
rect 312734 131108 312970 131344
rect 313054 131108 313290 131344
rect 313374 131108 313610 131344
rect 309854 100472 310090 100708
rect 310174 100472 310410 100708
rect 310494 100472 310730 100708
rect 310814 100472 311050 100708
rect 311134 100472 311370 100708
rect 311454 100472 311690 100708
rect 311774 100472 312010 100708
rect 312094 100472 312330 100708
rect 312414 100472 312650 100708
rect 312734 100472 312970 100708
rect 313054 100472 313290 100708
rect 313374 100472 313610 100708
rect 309854 69836 310090 70072
rect 310174 69836 310410 70072
rect 310494 69836 310730 70072
rect 310814 69836 311050 70072
rect 311134 69836 311370 70072
rect 311454 69836 311690 70072
rect 311774 69836 312010 70072
rect 312094 69836 312330 70072
rect 312414 69836 312650 70072
rect 312734 69836 312970 70072
rect 313054 69836 313290 70072
rect 313374 69836 313610 70072
rect 309854 39200 310090 39436
rect 310174 39200 310410 39436
rect 310494 39200 310730 39436
rect 310814 39200 311050 39436
rect 311134 39200 311370 39436
rect 311454 39200 311690 39436
rect 311774 39200 312010 39436
rect 312094 39200 312330 39436
rect 312414 39200 312650 39436
rect 312734 39200 312970 39436
rect 313054 39200 313290 39436
rect 313374 39200 313610 39436
rect 122 3642 358 3878
rect 442 3642 678 3878
rect 762 3642 998 3878
rect 1082 3642 1318 3878
rect 1402 3642 1638 3878
rect 1722 3642 1958 3878
rect 2042 3642 2278 3878
rect 2362 3642 2598 3878
rect 2682 3642 2918 3878
rect 3002 3642 3238 3878
rect 3322 3642 3558 3878
rect 3642 3642 3878 3878
rect 122 3322 358 3558
rect 442 3322 678 3558
rect 762 3322 998 3558
rect 1082 3322 1318 3558
rect 1402 3322 1638 3558
rect 1722 3322 1958 3558
rect 2042 3322 2278 3558
rect 2362 3322 2598 3558
rect 2682 3322 2918 3558
rect 3002 3322 3238 3558
rect 3322 3322 3558 3558
rect 3642 3322 3878 3558
rect 122 3002 358 3238
rect 442 3002 678 3238
rect 762 3002 998 3238
rect 1082 3002 1318 3238
rect 1402 3002 1638 3238
rect 1722 3002 1958 3238
rect 2042 3002 2278 3238
rect 2362 3002 2598 3238
rect 2682 3002 2918 3238
rect 3002 3002 3238 3238
rect 3322 3002 3558 3238
rect 3642 3002 3878 3238
rect 122 2682 358 2918
rect 442 2682 678 2918
rect 762 2682 998 2918
rect 1082 2682 1318 2918
rect 1402 2682 1638 2918
rect 1722 2682 1958 2918
rect 2042 2682 2278 2918
rect 2362 2682 2598 2918
rect 2682 2682 2918 2918
rect 3002 2682 3238 2918
rect 3322 2682 3558 2918
rect 3642 2682 3878 2918
rect 122 2362 358 2598
rect 442 2362 678 2598
rect 762 2362 998 2598
rect 1082 2362 1318 2598
rect 1402 2362 1638 2598
rect 1722 2362 1958 2598
rect 2042 2362 2278 2598
rect 2362 2362 2598 2598
rect 2682 2362 2918 2598
rect 3002 2362 3238 2598
rect 3322 2362 3558 2598
rect 3642 2362 3878 2598
rect 122 2042 358 2278
rect 442 2042 678 2278
rect 762 2042 998 2278
rect 1082 2042 1318 2278
rect 1402 2042 1638 2278
rect 1722 2042 1958 2278
rect 2042 2042 2278 2278
rect 2362 2042 2598 2278
rect 2682 2042 2918 2278
rect 3002 2042 3238 2278
rect 3322 2042 3558 2278
rect 3642 2042 3878 2278
rect 122 1722 358 1958
rect 442 1722 678 1958
rect 762 1722 998 1958
rect 1082 1722 1318 1958
rect 1402 1722 1638 1958
rect 1722 1722 1958 1958
rect 2042 1722 2278 1958
rect 2362 1722 2598 1958
rect 2682 1722 2918 1958
rect 3002 1722 3238 1958
rect 3322 1722 3558 1958
rect 3642 1722 3878 1958
rect 122 1402 358 1638
rect 442 1402 678 1638
rect 762 1402 998 1638
rect 1082 1402 1318 1638
rect 1402 1402 1638 1638
rect 1722 1402 1958 1638
rect 2042 1402 2278 1638
rect 2362 1402 2598 1638
rect 2682 1402 2918 1638
rect 3002 1402 3238 1638
rect 3322 1402 3558 1638
rect 3642 1402 3878 1638
rect 122 1082 358 1318
rect 442 1082 678 1318
rect 762 1082 998 1318
rect 1082 1082 1318 1318
rect 1402 1082 1638 1318
rect 1722 1082 1958 1318
rect 2042 1082 2278 1318
rect 2362 1082 2598 1318
rect 2682 1082 2918 1318
rect 3002 1082 3238 1318
rect 3322 1082 3558 1318
rect 3642 1082 3878 1318
rect 122 762 358 998
rect 442 762 678 998
rect 762 762 998 998
rect 1082 762 1318 998
rect 1402 762 1638 998
rect 1722 762 1958 998
rect 2042 762 2278 998
rect 2362 762 2598 998
rect 2682 762 2918 998
rect 3002 762 3238 998
rect 3322 762 3558 998
rect 3642 762 3878 998
rect 122 442 358 678
rect 442 442 678 678
rect 762 442 998 678
rect 1082 442 1318 678
rect 1402 442 1638 678
rect 1722 442 1958 678
rect 2042 442 2278 678
rect 2362 442 2598 678
rect 2682 442 2918 678
rect 3002 442 3238 678
rect 3322 442 3558 678
rect 3642 442 3878 678
rect 122 122 358 358
rect 442 122 678 358
rect 762 122 998 358
rect 1082 122 1318 358
rect 1402 122 1638 358
rect 1722 122 1958 358
rect 2042 122 2278 358
rect 2362 122 2598 358
rect 2682 122 2918 358
rect 3002 122 3238 358
rect 3322 122 3558 358
rect 3642 122 3878 358
rect 309854 3642 310090 3878
rect 310174 3642 310410 3878
rect 310494 3642 310730 3878
rect 310814 3642 311050 3878
rect 311134 3642 311370 3878
rect 311454 3642 311690 3878
rect 311774 3642 312010 3878
rect 312094 3642 312330 3878
rect 312414 3642 312650 3878
rect 312734 3642 312970 3878
rect 313054 3642 313290 3878
rect 313374 3642 313610 3878
rect 309854 3322 310090 3558
rect 310174 3322 310410 3558
rect 310494 3322 310730 3558
rect 310814 3322 311050 3558
rect 311134 3322 311370 3558
rect 311454 3322 311690 3558
rect 311774 3322 312010 3558
rect 312094 3322 312330 3558
rect 312414 3322 312650 3558
rect 312734 3322 312970 3558
rect 313054 3322 313290 3558
rect 313374 3322 313610 3558
rect 309854 3002 310090 3238
rect 310174 3002 310410 3238
rect 310494 3002 310730 3238
rect 310814 3002 311050 3238
rect 311134 3002 311370 3238
rect 311454 3002 311690 3238
rect 311774 3002 312010 3238
rect 312094 3002 312330 3238
rect 312414 3002 312650 3238
rect 312734 3002 312970 3238
rect 313054 3002 313290 3238
rect 313374 3002 313610 3238
rect 309854 2682 310090 2918
rect 310174 2682 310410 2918
rect 310494 2682 310730 2918
rect 310814 2682 311050 2918
rect 311134 2682 311370 2918
rect 311454 2682 311690 2918
rect 311774 2682 312010 2918
rect 312094 2682 312330 2918
rect 312414 2682 312650 2918
rect 312734 2682 312970 2918
rect 313054 2682 313290 2918
rect 313374 2682 313610 2918
rect 309854 2362 310090 2598
rect 310174 2362 310410 2598
rect 310494 2362 310730 2598
rect 310814 2362 311050 2598
rect 311134 2362 311370 2598
rect 311454 2362 311690 2598
rect 311774 2362 312010 2598
rect 312094 2362 312330 2598
rect 312414 2362 312650 2598
rect 312734 2362 312970 2598
rect 313054 2362 313290 2598
rect 313374 2362 313610 2598
rect 309854 2042 310090 2278
rect 310174 2042 310410 2278
rect 310494 2042 310730 2278
rect 310814 2042 311050 2278
rect 311134 2042 311370 2278
rect 311454 2042 311690 2278
rect 311774 2042 312010 2278
rect 312094 2042 312330 2278
rect 312414 2042 312650 2278
rect 312734 2042 312970 2278
rect 313054 2042 313290 2278
rect 313374 2042 313610 2278
rect 309854 1722 310090 1958
rect 310174 1722 310410 1958
rect 310494 1722 310730 1958
rect 310814 1722 311050 1958
rect 311134 1722 311370 1958
rect 311454 1722 311690 1958
rect 311774 1722 312010 1958
rect 312094 1722 312330 1958
rect 312414 1722 312650 1958
rect 312734 1722 312970 1958
rect 313054 1722 313290 1958
rect 313374 1722 313610 1958
rect 309854 1402 310090 1638
rect 310174 1402 310410 1638
rect 310494 1402 310730 1638
rect 310814 1402 311050 1638
rect 311134 1402 311370 1638
rect 311454 1402 311690 1638
rect 311774 1402 312010 1638
rect 312094 1402 312330 1638
rect 312414 1402 312650 1638
rect 312734 1402 312970 1638
rect 313054 1402 313290 1638
rect 313374 1402 313610 1638
rect 309854 1082 310090 1318
rect 310174 1082 310410 1318
rect 310494 1082 310730 1318
rect 310814 1082 311050 1318
rect 311134 1082 311370 1318
rect 311454 1082 311690 1318
rect 311774 1082 312010 1318
rect 312094 1082 312330 1318
rect 312414 1082 312650 1318
rect 312734 1082 312970 1318
rect 313054 1082 313290 1318
rect 313374 1082 313610 1318
rect 309854 762 310090 998
rect 310174 762 310410 998
rect 310494 762 310730 998
rect 310814 762 311050 998
rect 311134 762 311370 998
rect 311454 762 311690 998
rect 311774 762 312010 998
rect 312094 762 312330 998
rect 312414 762 312650 998
rect 312734 762 312970 998
rect 313054 762 313290 998
rect 313374 762 313610 998
rect 309854 442 310090 678
rect 310174 442 310410 678
rect 310494 442 310730 678
rect 310814 442 311050 678
rect 311134 442 311370 678
rect 311454 442 311690 678
rect 311774 442 312010 678
rect 312094 442 312330 678
rect 312414 442 312650 678
rect 312734 442 312970 678
rect 313054 442 313290 678
rect 313374 442 313610 678
rect 309854 122 310090 358
rect 310174 122 310410 358
rect 310494 122 310730 358
rect 310814 122 311050 358
rect 311134 122 311370 358
rect 311454 122 311690 358
rect 311774 122 312010 358
rect 312094 122 312330 358
rect 312414 122 312650 358
rect 312734 122 312970 358
rect 313054 122 313290 358
rect 313374 122 313610 358
<< metal5 >>
rect 0 311286 313732 311408
rect 0 311050 122 311286
rect 358 311050 442 311286
rect 678 311050 762 311286
rect 998 311050 1082 311286
rect 1318 311050 1402 311286
rect 1638 311050 1722 311286
rect 1958 311050 2042 311286
rect 2278 311050 2362 311286
rect 2598 311050 2682 311286
rect 2918 311050 3002 311286
rect 3238 311050 3322 311286
rect 3558 311050 3642 311286
rect 3878 311050 309854 311286
rect 310090 311050 310174 311286
rect 310410 311050 310494 311286
rect 310730 311050 310814 311286
rect 311050 311050 311134 311286
rect 311370 311050 311454 311286
rect 311690 311050 311774 311286
rect 312010 311050 312094 311286
rect 312330 311050 312414 311286
rect 312650 311050 312734 311286
rect 312970 311050 313054 311286
rect 313290 311050 313374 311286
rect 313610 311050 313732 311286
rect 0 310966 313732 311050
rect 0 310730 122 310966
rect 358 310730 442 310966
rect 678 310730 762 310966
rect 998 310730 1082 310966
rect 1318 310730 1402 310966
rect 1638 310730 1722 310966
rect 1958 310730 2042 310966
rect 2278 310730 2362 310966
rect 2598 310730 2682 310966
rect 2918 310730 3002 310966
rect 3238 310730 3322 310966
rect 3558 310730 3642 310966
rect 3878 310730 309854 310966
rect 310090 310730 310174 310966
rect 310410 310730 310494 310966
rect 310730 310730 310814 310966
rect 311050 310730 311134 310966
rect 311370 310730 311454 310966
rect 311690 310730 311774 310966
rect 312010 310730 312094 310966
rect 312330 310730 312414 310966
rect 312650 310730 312734 310966
rect 312970 310730 313054 310966
rect 313290 310730 313374 310966
rect 313610 310730 313732 310966
rect 0 310646 313732 310730
rect 0 310410 122 310646
rect 358 310410 442 310646
rect 678 310410 762 310646
rect 998 310410 1082 310646
rect 1318 310410 1402 310646
rect 1638 310410 1722 310646
rect 1958 310410 2042 310646
rect 2278 310410 2362 310646
rect 2598 310410 2682 310646
rect 2918 310410 3002 310646
rect 3238 310410 3322 310646
rect 3558 310410 3642 310646
rect 3878 310410 309854 310646
rect 310090 310410 310174 310646
rect 310410 310410 310494 310646
rect 310730 310410 310814 310646
rect 311050 310410 311134 310646
rect 311370 310410 311454 310646
rect 311690 310410 311774 310646
rect 312010 310410 312094 310646
rect 312330 310410 312414 310646
rect 312650 310410 312734 310646
rect 312970 310410 313054 310646
rect 313290 310410 313374 310646
rect 313610 310410 313732 310646
rect 0 310326 313732 310410
rect 0 310090 122 310326
rect 358 310090 442 310326
rect 678 310090 762 310326
rect 998 310090 1082 310326
rect 1318 310090 1402 310326
rect 1638 310090 1722 310326
rect 1958 310090 2042 310326
rect 2278 310090 2362 310326
rect 2598 310090 2682 310326
rect 2918 310090 3002 310326
rect 3238 310090 3322 310326
rect 3558 310090 3642 310326
rect 3878 310090 309854 310326
rect 310090 310090 310174 310326
rect 310410 310090 310494 310326
rect 310730 310090 310814 310326
rect 311050 310090 311134 310326
rect 311370 310090 311454 310326
rect 311690 310090 311774 310326
rect 312010 310090 312094 310326
rect 312330 310090 312414 310326
rect 312650 310090 312734 310326
rect 312970 310090 313054 310326
rect 313290 310090 313374 310326
rect 313610 310090 313732 310326
rect 0 310006 313732 310090
rect 0 309770 122 310006
rect 358 309770 442 310006
rect 678 309770 762 310006
rect 998 309770 1082 310006
rect 1318 309770 1402 310006
rect 1638 309770 1722 310006
rect 1958 309770 2042 310006
rect 2278 309770 2362 310006
rect 2598 309770 2682 310006
rect 2918 309770 3002 310006
rect 3238 309770 3322 310006
rect 3558 309770 3642 310006
rect 3878 309770 309854 310006
rect 310090 309770 310174 310006
rect 310410 309770 310494 310006
rect 310730 309770 310814 310006
rect 311050 309770 311134 310006
rect 311370 309770 311454 310006
rect 311690 309770 311774 310006
rect 312010 309770 312094 310006
rect 312330 309770 312414 310006
rect 312650 309770 312734 310006
rect 312970 309770 313054 310006
rect 313290 309770 313374 310006
rect 313610 309770 313732 310006
rect 0 309686 313732 309770
rect 0 309450 122 309686
rect 358 309450 442 309686
rect 678 309450 762 309686
rect 998 309450 1082 309686
rect 1318 309450 1402 309686
rect 1638 309450 1722 309686
rect 1958 309450 2042 309686
rect 2278 309450 2362 309686
rect 2598 309450 2682 309686
rect 2918 309450 3002 309686
rect 3238 309450 3322 309686
rect 3558 309450 3642 309686
rect 3878 309450 309854 309686
rect 310090 309450 310174 309686
rect 310410 309450 310494 309686
rect 310730 309450 310814 309686
rect 311050 309450 311134 309686
rect 311370 309450 311454 309686
rect 311690 309450 311774 309686
rect 312010 309450 312094 309686
rect 312330 309450 312414 309686
rect 312650 309450 312734 309686
rect 312970 309450 313054 309686
rect 313290 309450 313374 309686
rect 313610 309450 313732 309686
rect 0 309366 313732 309450
rect 0 309130 122 309366
rect 358 309130 442 309366
rect 678 309130 762 309366
rect 998 309130 1082 309366
rect 1318 309130 1402 309366
rect 1638 309130 1722 309366
rect 1958 309130 2042 309366
rect 2278 309130 2362 309366
rect 2598 309130 2682 309366
rect 2918 309130 3002 309366
rect 3238 309130 3322 309366
rect 3558 309130 3642 309366
rect 3878 309130 309854 309366
rect 310090 309130 310174 309366
rect 310410 309130 310494 309366
rect 310730 309130 310814 309366
rect 311050 309130 311134 309366
rect 311370 309130 311454 309366
rect 311690 309130 311774 309366
rect 312010 309130 312094 309366
rect 312330 309130 312414 309366
rect 312650 309130 312734 309366
rect 312970 309130 313054 309366
rect 313290 309130 313374 309366
rect 313610 309130 313732 309366
rect 0 309046 313732 309130
rect 0 308810 122 309046
rect 358 308810 442 309046
rect 678 308810 762 309046
rect 998 308810 1082 309046
rect 1318 308810 1402 309046
rect 1638 308810 1722 309046
rect 1958 308810 2042 309046
rect 2278 308810 2362 309046
rect 2598 308810 2682 309046
rect 2918 308810 3002 309046
rect 3238 308810 3322 309046
rect 3558 308810 3642 309046
rect 3878 308810 309854 309046
rect 310090 308810 310174 309046
rect 310410 308810 310494 309046
rect 310730 308810 310814 309046
rect 311050 308810 311134 309046
rect 311370 308810 311454 309046
rect 311690 308810 311774 309046
rect 312010 308810 312094 309046
rect 312330 308810 312414 309046
rect 312650 308810 312734 309046
rect 312970 308810 313054 309046
rect 313290 308810 313374 309046
rect 313610 308810 313732 309046
rect 0 308726 313732 308810
rect 0 308490 122 308726
rect 358 308490 442 308726
rect 678 308490 762 308726
rect 998 308490 1082 308726
rect 1318 308490 1402 308726
rect 1638 308490 1722 308726
rect 1958 308490 2042 308726
rect 2278 308490 2362 308726
rect 2598 308490 2682 308726
rect 2918 308490 3002 308726
rect 3238 308490 3322 308726
rect 3558 308490 3642 308726
rect 3878 308490 309854 308726
rect 310090 308490 310174 308726
rect 310410 308490 310494 308726
rect 310730 308490 310814 308726
rect 311050 308490 311134 308726
rect 311370 308490 311454 308726
rect 311690 308490 311774 308726
rect 312010 308490 312094 308726
rect 312330 308490 312414 308726
rect 312650 308490 312734 308726
rect 312970 308490 313054 308726
rect 313290 308490 313374 308726
rect 313610 308490 313732 308726
rect 0 308406 313732 308490
rect 0 308170 122 308406
rect 358 308170 442 308406
rect 678 308170 762 308406
rect 998 308170 1082 308406
rect 1318 308170 1402 308406
rect 1638 308170 1722 308406
rect 1958 308170 2042 308406
rect 2278 308170 2362 308406
rect 2598 308170 2682 308406
rect 2918 308170 3002 308406
rect 3238 308170 3322 308406
rect 3558 308170 3642 308406
rect 3878 308170 309854 308406
rect 310090 308170 310174 308406
rect 310410 308170 310494 308406
rect 310730 308170 310814 308406
rect 311050 308170 311134 308406
rect 311370 308170 311454 308406
rect 311690 308170 311774 308406
rect 312010 308170 312094 308406
rect 312330 308170 312414 308406
rect 312650 308170 312734 308406
rect 312970 308170 313054 308406
rect 313290 308170 313374 308406
rect 313610 308170 313732 308406
rect 0 308086 313732 308170
rect 0 307850 122 308086
rect 358 307850 442 308086
rect 678 307850 762 308086
rect 998 307850 1082 308086
rect 1318 307850 1402 308086
rect 1638 307850 1722 308086
rect 1958 307850 2042 308086
rect 2278 307850 2362 308086
rect 2598 307850 2682 308086
rect 2918 307850 3002 308086
rect 3238 307850 3322 308086
rect 3558 307850 3642 308086
rect 3878 307850 309854 308086
rect 310090 307850 310174 308086
rect 310410 307850 310494 308086
rect 310730 307850 310814 308086
rect 311050 307850 311134 308086
rect 311370 307850 311454 308086
rect 311690 307850 311774 308086
rect 312010 307850 312094 308086
rect 312330 307850 312414 308086
rect 312650 307850 312734 308086
rect 312970 307850 313054 308086
rect 313290 307850 313374 308086
rect 313610 307850 313732 308086
rect 0 307766 313732 307850
rect 0 307530 122 307766
rect 358 307530 442 307766
rect 678 307530 762 307766
rect 998 307530 1082 307766
rect 1318 307530 1402 307766
rect 1638 307530 1722 307766
rect 1958 307530 2042 307766
rect 2278 307530 2362 307766
rect 2598 307530 2682 307766
rect 2918 307530 3002 307766
rect 3238 307530 3322 307766
rect 3558 307530 3642 307766
rect 3878 307530 309854 307766
rect 310090 307530 310174 307766
rect 310410 307530 310494 307766
rect 310730 307530 310814 307766
rect 311050 307530 311134 307766
rect 311370 307530 311454 307766
rect 311690 307530 311774 307766
rect 312010 307530 312094 307766
rect 312330 307530 312414 307766
rect 312650 307530 312734 307766
rect 312970 307530 313054 307766
rect 313290 307530 313374 307766
rect 313610 307530 313732 307766
rect 0 307408 313732 307530
rect 5000 306286 308732 306408
rect 5000 306050 5122 306286
rect 5358 306050 5442 306286
rect 5678 306050 5762 306286
rect 5998 306050 6082 306286
rect 6318 306050 6402 306286
rect 6638 306050 6722 306286
rect 6958 306050 7042 306286
rect 7278 306050 7362 306286
rect 7598 306050 7682 306286
rect 7918 306050 8002 306286
rect 8238 306050 8322 306286
rect 8558 306050 8642 306286
rect 8878 306050 304854 306286
rect 305090 306050 305174 306286
rect 305410 306050 305494 306286
rect 305730 306050 305814 306286
rect 306050 306050 306134 306286
rect 306370 306050 306454 306286
rect 306690 306050 306774 306286
rect 307010 306050 307094 306286
rect 307330 306050 307414 306286
rect 307650 306050 307734 306286
rect 307970 306050 308054 306286
rect 308290 306050 308374 306286
rect 308610 306050 308732 306286
rect 5000 305966 308732 306050
rect 5000 305730 5122 305966
rect 5358 305730 5442 305966
rect 5678 305730 5762 305966
rect 5998 305730 6082 305966
rect 6318 305730 6402 305966
rect 6638 305730 6722 305966
rect 6958 305730 7042 305966
rect 7278 305730 7362 305966
rect 7598 305730 7682 305966
rect 7918 305730 8002 305966
rect 8238 305730 8322 305966
rect 8558 305730 8642 305966
rect 8878 305730 304854 305966
rect 305090 305730 305174 305966
rect 305410 305730 305494 305966
rect 305730 305730 305814 305966
rect 306050 305730 306134 305966
rect 306370 305730 306454 305966
rect 306690 305730 306774 305966
rect 307010 305730 307094 305966
rect 307330 305730 307414 305966
rect 307650 305730 307734 305966
rect 307970 305730 308054 305966
rect 308290 305730 308374 305966
rect 308610 305730 308732 305966
rect 5000 305646 308732 305730
rect 5000 305410 5122 305646
rect 5358 305410 5442 305646
rect 5678 305410 5762 305646
rect 5998 305410 6082 305646
rect 6318 305410 6402 305646
rect 6638 305410 6722 305646
rect 6958 305410 7042 305646
rect 7278 305410 7362 305646
rect 7598 305410 7682 305646
rect 7918 305410 8002 305646
rect 8238 305410 8322 305646
rect 8558 305410 8642 305646
rect 8878 305410 304854 305646
rect 305090 305410 305174 305646
rect 305410 305410 305494 305646
rect 305730 305410 305814 305646
rect 306050 305410 306134 305646
rect 306370 305410 306454 305646
rect 306690 305410 306774 305646
rect 307010 305410 307094 305646
rect 307330 305410 307414 305646
rect 307650 305410 307734 305646
rect 307970 305410 308054 305646
rect 308290 305410 308374 305646
rect 308610 305410 308732 305646
rect 5000 305326 308732 305410
rect 5000 305090 5122 305326
rect 5358 305090 5442 305326
rect 5678 305090 5762 305326
rect 5998 305090 6082 305326
rect 6318 305090 6402 305326
rect 6638 305090 6722 305326
rect 6958 305090 7042 305326
rect 7278 305090 7362 305326
rect 7598 305090 7682 305326
rect 7918 305090 8002 305326
rect 8238 305090 8322 305326
rect 8558 305090 8642 305326
rect 8878 305090 304854 305326
rect 305090 305090 305174 305326
rect 305410 305090 305494 305326
rect 305730 305090 305814 305326
rect 306050 305090 306134 305326
rect 306370 305090 306454 305326
rect 306690 305090 306774 305326
rect 307010 305090 307094 305326
rect 307330 305090 307414 305326
rect 307650 305090 307734 305326
rect 307970 305090 308054 305326
rect 308290 305090 308374 305326
rect 308610 305090 308732 305326
rect 5000 305006 308732 305090
rect 5000 304770 5122 305006
rect 5358 304770 5442 305006
rect 5678 304770 5762 305006
rect 5998 304770 6082 305006
rect 6318 304770 6402 305006
rect 6638 304770 6722 305006
rect 6958 304770 7042 305006
rect 7278 304770 7362 305006
rect 7598 304770 7682 305006
rect 7918 304770 8002 305006
rect 8238 304770 8322 305006
rect 8558 304770 8642 305006
rect 8878 304770 304854 305006
rect 305090 304770 305174 305006
rect 305410 304770 305494 305006
rect 305730 304770 305814 305006
rect 306050 304770 306134 305006
rect 306370 304770 306454 305006
rect 306690 304770 306774 305006
rect 307010 304770 307094 305006
rect 307330 304770 307414 305006
rect 307650 304770 307734 305006
rect 307970 304770 308054 305006
rect 308290 304770 308374 305006
rect 308610 304770 308732 305006
rect 5000 304686 308732 304770
rect 5000 304450 5122 304686
rect 5358 304450 5442 304686
rect 5678 304450 5762 304686
rect 5998 304450 6082 304686
rect 6318 304450 6402 304686
rect 6638 304450 6722 304686
rect 6958 304450 7042 304686
rect 7278 304450 7362 304686
rect 7598 304450 7682 304686
rect 7918 304450 8002 304686
rect 8238 304450 8322 304686
rect 8558 304450 8642 304686
rect 8878 304450 304854 304686
rect 305090 304450 305174 304686
rect 305410 304450 305494 304686
rect 305730 304450 305814 304686
rect 306050 304450 306134 304686
rect 306370 304450 306454 304686
rect 306690 304450 306774 304686
rect 307010 304450 307094 304686
rect 307330 304450 307414 304686
rect 307650 304450 307734 304686
rect 307970 304450 308054 304686
rect 308290 304450 308374 304686
rect 308610 304450 308732 304686
rect 5000 304366 308732 304450
rect 5000 304130 5122 304366
rect 5358 304130 5442 304366
rect 5678 304130 5762 304366
rect 5998 304130 6082 304366
rect 6318 304130 6402 304366
rect 6638 304130 6722 304366
rect 6958 304130 7042 304366
rect 7278 304130 7362 304366
rect 7598 304130 7682 304366
rect 7918 304130 8002 304366
rect 8238 304130 8322 304366
rect 8558 304130 8642 304366
rect 8878 304130 304854 304366
rect 305090 304130 305174 304366
rect 305410 304130 305494 304366
rect 305730 304130 305814 304366
rect 306050 304130 306134 304366
rect 306370 304130 306454 304366
rect 306690 304130 306774 304366
rect 307010 304130 307094 304366
rect 307330 304130 307414 304366
rect 307650 304130 307734 304366
rect 307970 304130 308054 304366
rect 308290 304130 308374 304366
rect 308610 304130 308732 304366
rect 5000 304046 308732 304130
rect 5000 303810 5122 304046
rect 5358 303810 5442 304046
rect 5678 303810 5762 304046
rect 5998 303810 6082 304046
rect 6318 303810 6402 304046
rect 6638 303810 6722 304046
rect 6958 303810 7042 304046
rect 7278 303810 7362 304046
rect 7598 303810 7682 304046
rect 7918 303810 8002 304046
rect 8238 303810 8322 304046
rect 8558 303810 8642 304046
rect 8878 303810 304854 304046
rect 305090 303810 305174 304046
rect 305410 303810 305494 304046
rect 305730 303810 305814 304046
rect 306050 303810 306134 304046
rect 306370 303810 306454 304046
rect 306690 303810 306774 304046
rect 307010 303810 307094 304046
rect 307330 303810 307414 304046
rect 307650 303810 307734 304046
rect 307970 303810 308054 304046
rect 308290 303810 308374 304046
rect 308610 303810 308732 304046
rect 5000 303726 308732 303810
rect 5000 303490 5122 303726
rect 5358 303490 5442 303726
rect 5678 303490 5762 303726
rect 5998 303490 6082 303726
rect 6318 303490 6402 303726
rect 6638 303490 6722 303726
rect 6958 303490 7042 303726
rect 7278 303490 7362 303726
rect 7598 303490 7682 303726
rect 7918 303490 8002 303726
rect 8238 303490 8322 303726
rect 8558 303490 8642 303726
rect 8878 303490 304854 303726
rect 305090 303490 305174 303726
rect 305410 303490 305494 303726
rect 305730 303490 305814 303726
rect 306050 303490 306134 303726
rect 306370 303490 306454 303726
rect 306690 303490 306774 303726
rect 307010 303490 307094 303726
rect 307330 303490 307414 303726
rect 307650 303490 307734 303726
rect 307970 303490 308054 303726
rect 308290 303490 308374 303726
rect 308610 303490 308732 303726
rect 5000 303406 308732 303490
rect 5000 303170 5122 303406
rect 5358 303170 5442 303406
rect 5678 303170 5762 303406
rect 5998 303170 6082 303406
rect 6318 303170 6402 303406
rect 6638 303170 6722 303406
rect 6958 303170 7042 303406
rect 7278 303170 7362 303406
rect 7598 303170 7682 303406
rect 7918 303170 8002 303406
rect 8238 303170 8322 303406
rect 8558 303170 8642 303406
rect 8878 303170 304854 303406
rect 305090 303170 305174 303406
rect 305410 303170 305494 303406
rect 305730 303170 305814 303406
rect 306050 303170 306134 303406
rect 306370 303170 306454 303406
rect 306690 303170 306774 303406
rect 307010 303170 307094 303406
rect 307330 303170 307414 303406
rect 307650 303170 307734 303406
rect 307970 303170 308054 303406
rect 308290 303170 308374 303406
rect 308610 303170 308732 303406
rect 5000 303086 308732 303170
rect 5000 302850 5122 303086
rect 5358 302850 5442 303086
rect 5678 302850 5762 303086
rect 5998 302850 6082 303086
rect 6318 302850 6402 303086
rect 6638 302850 6722 303086
rect 6958 302850 7042 303086
rect 7278 302850 7362 303086
rect 7598 302850 7682 303086
rect 7918 302850 8002 303086
rect 8238 302850 8322 303086
rect 8558 302850 8642 303086
rect 8878 302850 304854 303086
rect 305090 302850 305174 303086
rect 305410 302850 305494 303086
rect 305730 302850 305814 303086
rect 306050 302850 306134 303086
rect 306370 302850 306454 303086
rect 306690 302850 306774 303086
rect 307010 302850 307094 303086
rect 307330 302850 307414 303086
rect 307650 302850 307734 303086
rect 307970 302850 308054 303086
rect 308290 302850 308374 303086
rect 308610 302850 308732 303086
rect 5000 302766 308732 302850
rect 5000 302530 5122 302766
rect 5358 302530 5442 302766
rect 5678 302530 5762 302766
rect 5998 302530 6082 302766
rect 6318 302530 6402 302766
rect 6638 302530 6722 302766
rect 6958 302530 7042 302766
rect 7278 302530 7362 302766
rect 7598 302530 7682 302766
rect 7918 302530 8002 302766
rect 8238 302530 8322 302766
rect 8558 302530 8642 302766
rect 8878 302530 304854 302766
rect 305090 302530 305174 302766
rect 305410 302530 305494 302766
rect 305730 302530 305814 302766
rect 306050 302530 306134 302766
rect 306370 302530 306454 302766
rect 306690 302530 306774 302766
rect 307010 302530 307094 302766
rect 307330 302530 307414 302766
rect 307650 302530 307734 302766
rect 307970 302530 308054 302766
rect 308290 302530 308374 302766
rect 308610 302530 308732 302766
rect 5000 302408 308732 302530
rect 0 299842 313732 299884
rect 0 299606 5122 299842
rect 5358 299606 5442 299842
rect 5678 299606 5762 299842
rect 5998 299606 6082 299842
rect 6318 299606 6402 299842
rect 6638 299606 6722 299842
rect 6958 299606 7042 299842
rect 7278 299606 7362 299842
rect 7598 299606 7682 299842
rect 7918 299606 8002 299842
rect 8238 299606 8322 299842
rect 8558 299606 8642 299842
rect 8878 299606 304854 299842
rect 305090 299606 305174 299842
rect 305410 299606 305494 299842
rect 305730 299606 305814 299842
rect 306050 299606 306134 299842
rect 306370 299606 306454 299842
rect 306690 299606 306774 299842
rect 307010 299606 307094 299842
rect 307330 299606 307414 299842
rect 307650 299606 307734 299842
rect 307970 299606 308054 299842
rect 308290 299606 308374 299842
rect 308610 299606 313732 299842
rect 0 299564 313732 299606
rect 118572 288804 119076 289484
rect 109188 288484 119076 288804
rect 109188 288124 109508 288484
rect 90052 288082 109508 288124
rect 90052 287846 90094 288082
rect 90330 287846 109508 288082
rect 90052 287804 109508 287846
rect 118756 288124 119076 288484
rect 118756 288082 129748 288124
rect 118756 287846 129470 288082
rect 129706 287846 129748 288082
rect 118756 287804 129748 287846
rect 184076 288082 186788 288124
rect 184076 287846 184118 288082
rect 184354 287846 186788 288082
rect 184076 287804 186788 287846
rect 186468 287444 186788 287804
rect 196036 287804 206844 288124
rect 196036 287444 196356 287804
rect 186468 287124 196356 287444
rect 206524 287444 206844 287804
rect 215356 288082 223772 288124
rect 215356 287846 223494 288082
rect 223730 287846 223772 288082
rect 215356 287804 223772 287846
rect 215356 287444 215676 287804
rect 206524 287124 215676 287444
rect 195852 286444 196356 287124
rect 215172 286444 215676 287124
rect 0 284524 313732 284566
rect 0 284288 122 284524
rect 358 284288 442 284524
rect 678 284288 762 284524
rect 998 284288 1082 284524
rect 1318 284288 1402 284524
rect 1638 284288 1722 284524
rect 1958 284288 2042 284524
rect 2278 284288 2362 284524
rect 2598 284288 2682 284524
rect 2918 284288 3002 284524
rect 3238 284288 3322 284524
rect 3558 284288 3642 284524
rect 3878 284288 309854 284524
rect 310090 284288 310174 284524
rect 310410 284288 310494 284524
rect 310730 284288 310814 284524
rect 311050 284288 311134 284524
rect 311370 284288 311454 284524
rect 311690 284288 311774 284524
rect 312010 284288 312094 284524
rect 312330 284288 312414 284524
rect 312650 284288 312734 284524
rect 312970 284288 313054 284524
rect 313290 284288 313374 284524
rect 313610 284288 313732 284524
rect 0 284246 313732 284288
rect 0 269206 313732 269248
rect 0 268970 5122 269206
rect 5358 268970 5442 269206
rect 5678 268970 5762 269206
rect 5998 268970 6082 269206
rect 6318 268970 6402 269206
rect 6638 268970 6722 269206
rect 6958 268970 7042 269206
rect 7278 268970 7362 269206
rect 7598 268970 7682 269206
rect 7918 268970 8002 269206
rect 8238 268970 8322 269206
rect 8558 268970 8642 269206
rect 8878 268970 304854 269206
rect 305090 268970 305174 269206
rect 305410 268970 305494 269206
rect 305730 268970 305814 269206
rect 306050 268970 306134 269206
rect 306370 268970 306454 269206
rect 306690 268970 306774 269206
rect 307010 268970 307094 269206
rect 307330 268970 307414 269206
rect 307650 268970 307734 269206
rect 307970 268970 308054 269206
rect 308290 268970 308374 269206
rect 308610 268970 313732 269206
rect 0 268928 313732 268970
rect 226212 256122 265356 256164
rect 226212 255886 226254 256122
rect 226490 255886 265078 256122
rect 265314 255886 265356 256122
rect 226212 255844 265356 255886
rect 0 253888 313732 253930
rect 0 253652 122 253888
rect 358 253652 442 253888
rect 678 253652 762 253888
rect 998 253652 1082 253888
rect 1318 253652 1402 253888
rect 1638 253652 1722 253888
rect 1958 253652 2042 253888
rect 2278 253652 2362 253888
rect 2598 253652 2682 253888
rect 2918 253652 3002 253888
rect 3238 253652 3322 253888
rect 3558 253652 3642 253888
rect 3878 253652 309854 253888
rect 310090 253652 310174 253888
rect 310410 253652 310494 253888
rect 310730 253652 310814 253888
rect 311050 253652 311134 253888
rect 311370 253652 311454 253888
rect 311690 253652 311774 253888
rect 312010 253652 312094 253888
rect 312330 253652 312414 253888
rect 312650 253652 312734 253888
rect 312970 253652 313054 253888
rect 313290 253652 313374 253888
rect 313610 253652 313732 253888
rect 0 253610 313732 253652
rect 0 238570 313732 238612
rect 0 238334 5122 238570
rect 5358 238334 5442 238570
rect 5678 238334 5762 238570
rect 5998 238334 6082 238570
rect 6318 238334 6402 238570
rect 6638 238334 6722 238570
rect 6958 238334 7042 238570
rect 7278 238334 7362 238570
rect 7598 238334 7682 238570
rect 7918 238334 8002 238570
rect 8238 238334 8322 238570
rect 8558 238334 8642 238570
rect 8878 238334 304854 238570
rect 305090 238334 305174 238570
rect 305410 238334 305494 238570
rect 305730 238334 305814 238570
rect 306050 238334 306134 238570
rect 306370 238334 306454 238570
rect 306690 238334 306774 238570
rect 307010 238334 307094 238570
rect 307330 238334 307414 238570
rect 307650 238334 307734 238570
rect 307970 238334 308054 238570
rect 308290 238334 308374 238570
rect 308610 238334 313732 238570
rect 0 238292 313732 238334
rect 0 223252 313732 223294
rect 0 223016 122 223252
rect 358 223016 442 223252
rect 678 223016 762 223252
rect 998 223016 1082 223252
rect 1318 223016 1402 223252
rect 1638 223016 1722 223252
rect 1958 223016 2042 223252
rect 2278 223016 2362 223252
rect 2598 223016 2682 223252
rect 2918 223016 3002 223252
rect 3238 223016 3322 223252
rect 3558 223016 3642 223252
rect 3878 223016 309854 223252
rect 310090 223016 310174 223252
rect 310410 223016 310494 223252
rect 310730 223016 310814 223252
rect 311050 223016 311134 223252
rect 311370 223016 311454 223252
rect 311690 223016 311774 223252
rect 312010 223016 312094 223252
rect 312330 223016 312414 223252
rect 312650 223016 312734 223252
rect 312970 223016 313054 223252
rect 313290 223016 313374 223252
rect 313610 223016 313732 223252
rect 0 222974 313732 223016
rect 265036 216682 293876 216724
rect 265036 216446 265078 216682
rect 265314 216446 293598 216682
rect 293834 216446 293876 216682
rect 265036 216404 293876 216446
rect 69628 215322 81908 215364
rect 69628 215086 69670 215322
rect 69906 215086 81630 215322
rect 81866 215086 81908 215322
rect 69628 215044 81908 215086
rect 135132 211922 165076 211964
rect 135132 211686 135174 211922
rect 135410 211686 164798 211922
rect 165034 211686 165076 211922
rect 135132 211644 165076 211686
rect 0 207934 313732 207976
rect 0 207698 5122 207934
rect 5358 207698 5442 207934
rect 5678 207698 5762 207934
rect 5998 207698 6082 207934
rect 6318 207698 6402 207934
rect 6638 207698 6722 207934
rect 6958 207698 7042 207934
rect 7278 207698 7362 207934
rect 7598 207698 7682 207934
rect 7918 207698 8002 207934
rect 8238 207698 8322 207934
rect 8558 207698 8642 207934
rect 8878 207698 304854 207934
rect 305090 207698 305174 207934
rect 305410 207698 305494 207934
rect 305730 207698 305814 207934
rect 306050 207698 306134 207934
rect 306370 207698 306454 207934
rect 306690 207698 306774 207934
rect 307010 207698 307094 207934
rect 307330 207698 307414 207934
rect 307650 207698 307734 207934
rect 307970 207698 308054 207934
rect 308290 207698 308374 207934
rect 308610 207698 313732 207934
rect 0 207656 313732 207698
rect 37980 203082 229108 203124
rect 37980 202846 38022 203082
rect 38258 202846 228830 203082
rect 229066 202846 229108 203082
rect 37980 202804 229108 202846
rect 19948 202402 36092 202444
rect 19948 202166 19990 202402
rect 20226 202166 35814 202402
rect 36050 202166 36092 202402
rect 19948 202124 36092 202166
rect 242772 202402 258732 202444
rect 242772 202166 242814 202402
rect 243050 202166 258454 202402
rect 258690 202166 258732 202402
rect 242772 202124 258732 202166
rect 277916 202402 293876 202444
rect 277916 202166 277958 202402
rect 278194 202166 293598 202402
rect 293834 202166 293876 202402
rect 277916 202124 293876 202166
rect 0 192616 313732 192658
rect 0 192380 122 192616
rect 358 192380 442 192616
rect 678 192380 762 192616
rect 998 192380 1082 192616
rect 1318 192380 1402 192616
rect 1638 192380 1722 192616
rect 1958 192380 2042 192616
rect 2278 192380 2362 192616
rect 2598 192380 2682 192616
rect 2918 192380 3002 192616
rect 3238 192380 3322 192616
rect 3558 192380 3642 192616
rect 3878 192380 309854 192616
rect 310090 192380 310174 192616
rect 310410 192380 310494 192616
rect 310730 192380 310814 192616
rect 311050 192380 311134 192616
rect 311370 192380 311454 192616
rect 311690 192380 311774 192616
rect 312010 192380 312094 192616
rect 312330 192380 312414 192616
rect 312650 192380 312734 192616
rect 312970 192380 313054 192616
rect 313290 192380 313374 192616
rect 313610 192380 313732 192616
rect 0 192338 313732 192380
rect 0 177298 313732 177340
rect 0 177062 5122 177298
rect 5358 177062 5442 177298
rect 5678 177062 5762 177298
rect 5998 177062 6082 177298
rect 6318 177062 6402 177298
rect 6638 177062 6722 177298
rect 6958 177062 7042 177298
rect 7278 177062 7362 177298
rect 7598 177062 7682 177298
rect 7918 177062 8002 177298
rect 8238 177062 8322 177298
rect 8558 177062 8642 177298
rect 8878 177062 304854 177298
rect 305090 177062 305174 177298
rect 305410 177062 305494 177298
rect 305730 177062 305814 177298
rect 306050 177062 306134 177298
rect 306370 177062 306454 177298
rect 306690 177062 306774 177298
rect 307010 177062 307094 177298
rect 307330 177062 307414 177298
rect 307650 177062 307734 177298
rect 307970 177062 308054 177298
rect 308290 177062 308374 177298
rect 308610 177062 313732 177298
rect 0 177020 313732 177062
rect 0 161980 313732 162022
rect 0 161744 122 161980
rect 358 161744 442 161980
rect 678 161744 762 161980
rect 998 161744 1082 161980
rect 1318 161744 1402 161980
rect 1638 161744 1722 161980
rect 1958 161744 2042 161980
rect 2278 161744 2362 161980
rect 2598 161744 2682 161980
rect 2918 161744 3002 161980
rect 3238 161744 3322 161980
rect 3558 161744 3642 161980
rect 3878 161744 309854 161980
rect 310090 161744 310174 161980
rect 310410 161744 310494 161980
rect 310730 161744 310814 161980
rect 311050 161744 311134 161980
rect 311370 161744 311454 161980
rect 311690 161744 311774 161980
rect 312010 161744 312094 161980
rect 312330 161744 312414 161980
rect 312650 161744 312734 161980
rect 312970 161744 313054 161980
rect 313290 161744 313374 161980
rect 313610 161744 313732 161980
rect 0 161702 313732 161744
rect 0 146662 313732 146704
rect 0 146426 5122 146662
rect 5358 146426 5442 146662
rect 5678 146426 5762 146662
rect 5998 146426 6082 146662
rect 6318 146426 6402 146662
rect 6638 146426 6722 146662
rect 6958 146426 7042 146662
rect 7278 146426 7362 146662
rect 7598 146426 7682 146662
rect 7918 146426 8002 146662
rect 8238 146426 8322 146662
rect 8558 146426 8642 146662
rect 8878 146426 304854 146662
rect 305090 146426 305174 146662
rect 305410 146426 305494 146662
rect 305730 146426 305814 146662
rect 306050 146426 306134 146662
rect 306370 146426 306454 146662
rect 306690 146426 306774 146662
rect 307010 146426 307094 146662
rect 307330 146426 307414 146662
rect 307650 146426 307734 146662
rect 307970 146426 308054 146662
rect 308290 146426 308374 146662
rect 308610 146426 313732 146662
rect 0 146384 313732 146426
rect 48100 142562 109692 142604
rect 48100 142326 48142 142562
rect 48378 142326 109414 142562
rect 109650 142326 109692 142562
rect 48100 142284 109692 142326
rect 0 131344 313732 131386
rect 0 131108 122 131344
rect 358 131108 442 131344
rect 678 131108 762 131344
rect 998 131108 1082 131344
rect 1318 131108 1402 131344
rect 1638 131108 1722 131344
rect 1958 131108 2042 131344
rect 2278 131108 2362 131344
rect 2598 131108 2682 131344
rect 2918 131108 3002 131344
rect 3238 131108 3322 131344
rect 3558 131108 3642 131344
rect 3878 131108 309854 131344
rect 310090 131108 310174 131344
rect 310410 131108 310494 131344
rect 310730 131108 310814 131344
rect 311050 131108 311134 131344
rect 311370 131108 311454 131344
rect 311690 131108 311774 131344
rect 312010 131108 312094 131344
rect 312330 131108 312414 131344
rect 312650 131108 312734 131344
rect 312970 131108 313054 131344
rect 313290 131108 313374 131344
rect 313610 131108 313732 131344
rect 0 131066 313732 131108
rect 20684 130322 32228 130364
rect 20684 130086 20726 130322
rect 20962 130086 32228 130322
rect 20684 130044 32228 130086
rect 31908 129684 32228 130044
rect 41476 130322 48788 130364
rect 41476 130086 48510 130322
rect 48746 130086 48788 130322
rect 41476 130044 48788 130086
rect 57668 130322 58356 130364
rect 57668 130086 58078 130322
rect 58314 130086 58356 130322
rect 57668 130044 58356 130086
rect 93732 130044 103988 130364
rect 41476 129684 41796 130044
rect 31908 129364 41796 129684
rect 57668 129642 57988 130044
rect 57668 129406 57710 129642
rect 57946 129406 57988 129642
rect 57668 129364 57988 129406
rect 61348 129642 68292 129684
rect 61348 129406 61390 129642
rect 61626 129406 68292 129642
rect 61348 129364 68292 129406
rect 41292 128684 41796 129364
rect 67972 128324 68292 129364
rect 93732 129004 94052 130044
rect 77356 128684 80436 129004
rect 77356 128324 77676 128684
rect 67972 128004 77676 128324
rect 80116 128324 80436 128684
rect 84716 128684 94052 129004
rect 103668 129004 103988 130044
rect 113052 130044 116316 130364
rect 113052 129004 113372 130044
rect 115996 129684 116316 130044
rect 125748 130322 135636 130364
rect 125748 130086 135358 130322
rect 135594 130086 135636 130322
rect 125748 130044 135636 130086
rect 190332 130044 200588 130364
rect 125748 129684 126068 130044
rect 115996 129364 126068 129684
rect 138628 129642 167468 129684
rect 138628 129406 138670 129642
rect 138906 129406 167468 129642
rect 138628 129364 167468 129406
rect 103668 128684 113372 129004
rect 125564 128684 126068 129364
rect 84716 128324 85036 128684
rect 80116 128004 85036 128324
rect 167148 128324 167468 129364
rect 190332 129004 190652 130044
rect 173956 128684 177036 129004
rect 173956 128324 174276 128684
rect 167148 128004 174276 128324
rect 176716 128324 177036 128684
rect 181316 128684 190652 129004
rect 200268 129004 200588 130044
rect 209652 130044 219908 130364
rect 209652 129004 209972 130044
rect 200268 128684 209972 129004
rect 219588 129004 219908 130044
rect 234492 130322 244196 130364
rect 234492 130086 243918 130322
rect 244154 130086 244196 130322
rect 234492 130044 244196 130086
rect 269084 130322 270692 130364
rect 269084 130086 269126 130322
rect 269362 130086 270692 130322
rect 269084 130044 270692 130086
rect 234492 129684 234812 130044
rect 225108 129364 234812 129684
rect 244980 129642 251556 129684
rect 244980 129406 245022 129642
rect 245258 129406 251278 129642
rect 251514 129406 251556 129642
rect 244980 129364 251556 129406
rect 225108 129004 225428 129364
rect 219588 128684 225428 129004
rect 270372 129004 270692 130044
rect 286932 130322 288908 130364
rect 286932 130086 288630 130322
rect 288866 130086 288908 130322
rect 286932 130044 288908 130086
rect 286932 129004 287252 130044
rect 270372 128684 287252 129004
rect 181316 128324 181636 128684
rect 176716 128004 181636 128324
rect 264852 122162 293876 122204
rect 264852 121926 264894 122162
rect 265130 121926 293598 122162
rect 293834 121926 293876 122162
rect 264852 121884 293876 121926
rect 69628 121482 81908 121524
rect 69628 121246 69670 121482
rect 69906 121246 81630 121482
rect 81866 121246 81908 121482
rect 69628 121204 81908 121246
rect 229524 120802 261308 120844
rect 229524 120566 229566 120802
rect 229802 120566 261030 120802
rect 261266 120566 261308 120802
rect 229524 120524 261308 120566
rect 0 116026 313732 116068
rect 0 115790 5122 116026
rect 5358 115790 5442 116026
rect 5678 115790 5762 116026
rect 5998 115790 6082 116026
rect 6318 115790 6402 116026
rect 6638 115790 6722 116026
rect 6958 115790 7042 116026
rect 7278 115790 7362 116026
rect 7598 115790 7682 116026
rect 7918 115790 8002 116026
rect 8238 115790 8322 116026
rect 8558 115790 8642 116026
rect 8878 115790 304854 116026
rect 305090 115790 305174 116026
rect 305410 115790 305494 116026
rect 305730 115790 305814 116026
rect 306050 115790 306134 116026
rect 306370 115790 306454 116026
rect 306690 115790 306774 116026
rect 307010 115790 307094 116026
rect 307330 115790 307414 116026
rect 307650 115790 307734 116026
rect 307970 115790 308054 116026
rect 308290 115790 308374 116026
rect 308610 115790 313732 116026
rect 0 115748 313732 115790
rect 19948 108562 36092 108604
rect 19948 108326 19990 108562
rect 20226 108326 35814 108562
rect 36050 108326 36092 108562
rect 19948 108284 36092 108326
rect 0 100708 313732 100750
rect 0 100472 122 100708
rect 358 100472 442 100708
rect 678 100472 762 100708
rect 998 100472 1082 100708
rect 1318 100472 1402 100708
rect 1638 100472 1722 100708
rect 1958 100472 2042 100708
rect 2278 100472 2362 100708
rect 2598 100472 2682 100708
rect 2918 100472 3002 100708
rect 3238 100472 3322 100708
rect 3558 100472 3642 100708
rect 3878 100472 309854 100708
rect 310090 100472 310174 100708
rect 310410 100472 310494 100708
rect 310730 100472 310814 100708
rect 311050 100472 311134 100708
rect 311370 100472 311454 100708
rect 311690 100472 311774 100708
rect 312010 100472 312094 100708
rect 312330 100472 312414 100708
rect 312650 100472 312734 100708
rect 312970 100472 313054 100708
rect 313290 100472 313374 100708
rect 313610 100472 313732 100708
rect 0 100430 313732 100472
rect 0 85390 313732 85432
rect 0 85154 5122 85390
rect 5358 85154 5442 85390
rect 5678 85154 5762 85390
rect 5998 85154 6082 85390
rect 6318 85154 6402 85390
rect 6638 85154 6722 85390
rect 6958 85154 7042 85390
rect 7278 85154 7362 85390
rect 7598 85154 7682 85390
rect 7918 85154 8002 85390
rect 8238 85154 8322 85390
rect 8558 85154 8642 85390
rect 8878 85154 304854 85390
rect 305090 85154 305174 85390
rect 305410 85154 305494 85390
rect 305730 85154 305814 85390
rect 306050 85154 306134 85390
rect 306370 85154 306454 85390
rect 306690 85154 306774 85390
rect 307010 85154 307094 85390
rect 307330 85154 307414 85390
rect 307650 85154 307734 85390
rect 307970 85154 308054 85390
rect 308290 85154 308374 85390
rect 308610 85154 313732 85390
rect 0 85112 313732 85154
rect 0 70072 313732 70114
rect 0 69836 122 70072
rect 358 69836 442 70072
rect 678 69836 762 70072
rect 998 69836 1082 70072
rect 1318 69836 1402 70072
rect 1638 69836 1722 70072
rect 1958 69836 2042 70072
rect 2278 69836 2362 70072
rect 2598 69836 2682 70072
rect 2918 69836 3002 70072
rect 3238 69836 3322 70072
rect 3558 69836 3642 70072
rect 3878 69836 309854 70072
rect 310090 69836 310174 70072
rect 310410 69836 310494 70072
rect 310730 69836 310814 70072
rect 311050 69836 311134 70072
rect 311370 69836 311454 70072
rect 311690 69836 311774 70072
rect 312010 69836 312094 70072
rect 312330 69836 312414 70072
rect 312650 69836 312734 70072
rect 312970 69836 313054 70072
rect 313290 69836 313374 70072
rect 313610 69836 313732 70072
rect 0 69794 313732 69836
rect 0 54754 313732 54796
rect 0 54518 5122 54754
rect 5358 54518 5442 54754
rect 5678 54518 5762 54754
rect 5998 54518 6082 54754
rect 6318 54518 6402 54754
rect 6638 54518 6722 54754
rect 6958 54518 7042 54754
rect 7278 54518 7362 54754
rect 7598 54518 7682 54754
rect 7918 54518 8002 54754
rect 8238 54518 8322 54754
rect 8558 54518 8642 54754
rect 8878 54518 304854 54754
rect 305090 54518 305174 54754
rect 305410 54518 305494 54754
rect 305730 54518 305814 54754
rect 306050 54518 306134 54754
rect 306370 54518 306454 54754
rect 306690 54518 306774 54754
rect 307010 54518 307094 54754
rect 307330 54518 307414 54754
rect 307650 54518 307734 54754
rect 307970 54518 308054 54754
rect 308290 54518 308374 54754
rect 308610 54518 313732 54754
rect 0 54476 313732 54518
rect 0 39436 313732 39478
rect 0 39200 122 39436
rect 358 39200 442 39436
rect 678 39200 762 39436
rect 998 39200 1082 39436
rect 1318 39200 1402 39436
rect 1638 39200 1722 39436
rect 1958 39200 2042 39436
rect 2278 39200 2362 39436
rect 2598 39200 2682 39436
rect 2918 39200 3002 39436
rect 3238 39200 3322 39436
rect 3558 39200 3642 39436
rect 3878 39200 309854 39436
rect 310090 39200 310174 39436
rect 310410 39200 310494 39436
rect 310730 39200 310814 39436
rect 311050 39200 311134 39436
rect 311370 39200 311454 39436
rect 311690 39200 311774 39436
rect 312010 39200 312094 39436
rect 312330 39200 312414 39436
rect 312650 39200 312734 39436
rect 312970 39200 313054 39436
rect 313290 39200 313374 39436
rect 313610 39200 313732 39436
rect 0 39158 313732 39200
rect 0 24118 313732 24160
rect 0 23882 5122 24118
rect 5358 23882 5442 24118
rect 5678 23882 5762 24118
rect 5998 23882 6082 24118
rect 6318 23882 6402 24118
rect 6638 23882 6722 24118
rect 6958 23882 7042 24118
rect 7278 23882 7362 24118
rect 7598 23882 7682 24118
rect 7918 23882 8002 24118
rect 8238 23882 8322 24118
rect 8558 23882 8642 24118
rect 8878 23882 304854 24118
rect 305090 23882 305174 24118
rect 305410 23882 305494 24118
rect 305730 23882 305814 24118
rect 306050 23882 306134 24118
rect 306370 23882 306454 24118
rect 306690 23882 306774 24118
rect 307010 23882 307094 24118
rect 307330 23882 307414 24118
rect 307650 23882 307734 24118
rect 307970 23882 308054 24118
rect 308290 23882 308374 24118
rect 308610 23882 313732 24118
rect 0 23840 313732 23882
rect 5000 8878 308732 9000
rect 5000 8642 5122 8878
rect 5358 8642 5442 8878
rect 5678 8642 5762 8878
rect 5998 8642 6082 8878
rect 6318 8642 6402 8878
rect 6638 8642 6722 8878
rect 6958 8642 7042 8878
rect 7278 8642 7362 8878
rect 7598 8642 7682 8878
rect 7918 8642 8002 8878
rect 8238 8642 8322 8878
rect 8558 8642 8642 8878
rect 8878 8642 304854 8878
rect 305090 8642 305174 8878
rect 305410 8642 305494 8878
rect 305730 8642 305814 8878
rect 306050 8642 306134 8878
rect 306370 8642 306454 8878
rect 306690 8642 306774 8878
rect 307010 8642 307094 8878
rect 307330 8642 307414 8878
rect 307650 8642 307734 8878
rect 307970 8642 308054 8878
rect 308290 8642 308374 8878
rect 308610 8642 308732 8878
rect 5000 8558 308732 8642
rect 5000 8322 5122 8558
rect 5358 8322 5442 8558
rect 5678 8322 5762 8558
rect 5998 8322 6082 8558
rect 6318 8322 6402 8558
rect 6638 8322 6722 8558
rect 6958 8322 7042 8558
rect 7278 8322 7362 8558
rect 7598 8322 7682 8558
rect 7918 8322 8002 8558
rect 8238 8322 8322 8558
rect 8558 8322 8642 8558
rect 8878 8322 304854 8558
rect 305090 8322 305174 8558
rect 305410 8322 305494 8558
rect 305730 8322 305814 8558
rect 306050 8322 306134 8558
rect 306370 8322 306454 8558
rect 306690 8322 306774 8558
rect 307010 8322 307094 8558
rect 307330 8322 307414 8558
rect 307650 8322 307734 8558
rect 307970 8322 308054 8558
rect 308290 8322 308374 8558
rect 308610 8322 308732 8558
rect 5000 8238 308732 8322
rect 5000 8002 5122 8238
rect 5358 8002 5442 8238
rect 5678 8002 5762 8238
rect 5998 8002 6082 8238
rect 6318 8002 6402 8238
rect 6638 8002 6722 8238
rect 6958 8002 7042 8238
rect 7278 8002 7362 8238
rect 7598 8002 7682 8238
rect 7918 8002 8002 8238
rect 8238 8002 8322 8238
rect 8558 8002 8642 8238
rect 8878 8002 304854 8238
rect 305090 8002 305174 8238
rect 305410 8002 305494 8238
rect 305730 8002 305814 8238
rect 306050 8002 306134 8238
rect 306370 8002 306454 8238
rect 306690 8002 306774 8238
rect 307010 8002 307094 8238
rect 307330 8002 307414 8238
rect 307650 8002 307734 8238
rect 307970 8002 308054 8238
rect 308290 8002 308374 8238
rect 308610 8002 308732 8238
rect 5000 7918 308732 8002
rect 5000 7682 5122 7918
rect 5358 7682 5442 7918
rect 5678 7682 5762 7918
rect 5998 7682 6082 7918
rect 6318 7682 6402 7918
rect 6638 7682 6722 7918
rect 6958 7682 7042 7918
rect 7278 7682 7362 7918
rect 7598 7682 7682 7918
rect 7918 7682 8002 7918
rect 8238 7682 8322 7918
rect 8558 7682 8642 7918
rect 8878 7682 304854 7918
rect 305090 7682 305174 7918
rect 305410 7682 305494 7918
rect 305730 7682 305814 7918
rect 306050 7682 306134 7918
rect 306370 7682 306454 7918
rect 306690 7682 306774 7918
rect 307010 7682 307094 7918
rect 307330 7682 307414 7918
rect 307650 7682 307734 7918
rect 307970 7682 308054 7918
rect 308290 7682 308374 7918
rect 308610 7682 308732 7918
rect 5000 7598 308732 7682
rect 5000 7362 5122 7598
rect 5358 7362 5442 7598
rect 5678 7362 5762 7598
rect 5998 7362 6082 7598
rect 6318 7362 6402 7598
rect 6638 7362 6722 7598
rect 6958 7362 7042 7598
rect 7278 7362 7362 7598
rect 7598 7362 7682 7598
rect 7918 7362 8002 7598
rect 8238 7362 8322 7598
rect 8558 7362 8642 7598
rect 8878 7362 304854 7598
rect 305090 7362 305174 7598
rect 305410 7362 305494 7598
rect 305730 7362 305814 7598
rect 306050 7362 306134 7598
rect 306370 7362 306454 7598
rect 306690 7362 306774 7598
rect 307010 7362 307094 7598
rect 307330 7362 307414 7598
rect 307650 7362 307734 7598
rect 307970 7362 308054 7598
rect 308290 7362 308374 7598
rect 308610 7362 308732 7598
rect 5000 7278 308732 7362
rect 5000 7042 5122 7278
rect 5358 7042 5442 7278
rect 5678 7042 5762 7278
rect 5998 7042 6082 7278
rect 6318 7042 6402 7278
rect 6638 7042 6722 7278
rect 6958 7042 7042 7278
rect 7278 7042 7362 7278
rect 7598 7042 7682 7278
rect 7918 7042 8002 7278
rect 8238 7042 8322 7278
rect 8558 7042 8642 7278
rect 8878 7042 304854 7278
rect 305090 7042 305174 7278
rect 305410 7042 305494 7278
rect 305730 7042 305814 7278
rect 306050 7042 306134 7278
rect 306370 7042 306454 7278
rect 306690 7042 306774 7278
rect 307010 7042 307094 7278
rect 307330 7042 307414 7278
rect 307650 7042 307734 7278
rect 307970 7042 308054 7278
rect 308290 7042 308374 7278
rect 308610 7042 308732 7278
rect 5000 6958 308732 7042
rect 5000 6722 5122 6958
rect 5358 6722 5442 6958
rect 5678 6722 5762 6958
rect 5998 6722 6082 6958
rect 6318 6722 6402 6958
rect 6638 6722 6722 6958
rect 6958 6722 7042 6958
rect 7278 6722 7362 6958
rect 7598 6722 7682 6958
rect 7918 6722 8002 6958
rect 8238 6722 8322 6958
rect 8558 6722 8642 6958
rect 8878 6722 304854 6958
rect 305090 6722 305174 6958
rect 305410 6722 305494 6958
rect 305730 6722 305814 6958
rect 306050 6722 306134 6958
rect 306370 6722 306454 6958
rect 306690 6722 306774 6958
rect 307010 6722 307094 6958
rect 307330 6722 307414 6958
rect 307650 6722 307734 6958
rect 307970 6722 308054 6958
rect 308290 6722 308374 6958
rect 308610 6722 308732 6958
rect 5000 6638 308732 6722
rect 5000 6402 5122 6638
rect 5358 6402 5442 6638
rect 5678 6402 5762 6638
rect 5998 6402 6082 6638
rect 6318 6402 6402 6638
rect 6638 6402 6722 6638
rect 6958 6402 7042 6638
rect 7278 6402 7362 6638
rect 7598 6402 7682 6638
rect 7918 6402 8002 6638
rect 8238 6402 8322 6638
rect 8558 6402 8642 6638
rect 8878 6402 304854 6638
rect 305090 6402 305174 6638
rect 305410 6402 305494 6638
rect 305730 6402 305814 6638
rect 306050 6402 306134 6638
rect 306370 6402 306454 6638
rect 306690 6402 306774 6638
rect 307010 6402 307094 6638
rect 307330 6402 307414 6638
rect 307650 6402 307734 6638
rect 307970 6402 308054 6638
rect 308290 6402 308374 6638
rect 308610 6402 308732 6638
rect 5000 6318 308732 6402
rect 5000 6082 5122 6318
rect 5358 6082 5442 6318
rect 5678 6082 5762 6318
rect 5998 6082 6082 6318
rect 6318 6082 6402 6318
rect 6638 6082 6722 6318
rect 6958 6082 7042 6318
rect 7278 6082 7362 6318
rect 7598 6082 7682 6318
rect 7918 6082 8002 6318
rect 8238 6082 8322 6318
rect 8558 6082 8642 6318
rect 8878 6082 304854 6318
rect 305090 6082 305174 6318
rect 305410 6082 305494 6318
rect 305730 6082 305814 6318
rect 306050 6082 306134 6318
rect 306370 6082 306454 6318
rect 306690 6082 306774 6318
rect 307010 6082 307094 6318
rect 307330 6082 307414 6318
rect 307650 6082 307734 6318
rect 307970 6082 308054 6318
rect 308290 6082 308374 6318
rect 308610 6082 308732 6318
rect 5000 5998 308732 6082
rect 5000 5762 5122 5998
rect 5358 5762 5442 5998
rect 5678 5762 5762 5998
rect 5998 5762 6082 5998
rect 6318 5762 6402 5998
rect 6638 5762 6722 5998
rect 6958 5762 7042 5998
rect 7278 5762 7362 5998
rect 7598 5762 7682 5998
rect 7918 5762 8002 5998
rect 8238 5762 8322 5998
rect 8558 5762 8642 5998
rect 8878 5762 304854 5998
rect 305090 5762 305174 5998
rect 305410 5762 305494 5998
rect 305730 5762 305814 5998
rect 306050 5762 306134 5998
rect 306370 5762 306454 5998
rect 306690 5762 306774 5998
rect 307010 5762 307094 5998
rect 307330 5762 307414 5998
rect 307650 5762 307734 5998
rect 307970 5762 308054 5998
rect 308290 5762 308374 5998
rect 308610 5762 308732 5998
rect 5000 5678 308732 5762
rect 5000 5442 5122 5678
rect 5358 5442 5442 5678
rect 5678 5442 5762 5678
rect 5998 5442 6082 5678
rect 6318 5442 6402 5678
rect 6638 5442 6722 5678
rect 6958 5442 7042 5678
rect 7278 5442 7362 5678
rect 7598 5442 7682 5678
rect 7918 5442 8002 5678
rect 8238 5442 8322 5678
rect 8558 5442 8642 5678
rect 8878 5442 304854 5678
rect 305090 5442 305174 5678
rect 305410 5442 305494 5678
rect 305730 5442 305814 5678
rect 306050 5442 306134 5678
rect 306370 5442 306454 5678
rect 306690 5442 306774 5678
rect 307010 5442 307094 5678
rect 307330 5442 307414 5678
rect 307650 5442 307734 5678
rect 307970 5442 308054 5678
rect 308290 5442 308374 5678
rect 308610 5442 308732 5678
rect 5000 5358 308732 5442
rect 5000 5122 5122 5358
rect 5358 5122 5442 5358
rect 5678 5122 5762 5358
rect 5998 5122 6082 5358
rect 6318 5122 6402 5358
rect 6638 5122 6722 5358
rect 6958 5122 7042 5358
rect 7278 5122 7362 5358
rect 7598 5122 7682 5358
rect 7918 5122 8002 5358
rect 8238 5122 8322 5358
rect 8558 5122 8642 5358
rect 8878 5122 304854 5358
rect 305090 5122 305174 5358
rect 305410 5122 305494 5358
rect 305730 5122 305814 5358
rect 306050 5122 306134 5358
rect 306370 5122 306454 5358
rect 306690 5122 306774 5358
rect 307010 5122 307094 5358
rect 307330 5122 307414 5358
rect 307650 5122 307734 5358
rect 307970 5122 308054 5358
rect 308290 5122 308374 5358
rect 308610 5122 308732 5358
rect 5000 5000 308732 5122
rect 0 3878 313732 4000
rect 0 3642 122 3878
rect 358 3642 442 3878
rect 678 3642 762 3878
rect 998 3642 1082 3878
rect 1318 3642 1402 3878
rect 1638 3642 1722 3878
rect 1958 3642 2042 3878
rect 2278 3642 2362 3878
rect 2598 3642 2682 3878
rect 2918 3642 3002 3878
rect 3238 3642 3322 3878
rect 3558 3642 3642 3878
rect 3878 3642 309854 3878
rect 310090 3642 310174 3878
rect 310410 3642 310494 3878
rect 310730 3642 310814 3878
rect 311050 3642 311134 3878
rect 311370 3642 311454 3878
rect 311690 3642 311774 3878
rect 312010 3642 312094 3878
rect 312330 3642 312414 3878
rect 312650 3642 312734 3878
rect 312970 3642 313054 3878
rect 313290 3642 313374 3878
rect 313610 3642 313732 3878
rect 0 3558 313732 3642
rect 0 3322 122 3558
rect 358 3322 442 3558
rect 678 3322 762 3558
rect 998 3322 1082 3558
rect 1318 3322 1402 3558
rect 1638 3322 1722 3558
rect 1958 3322 2042 3558
rect 2278 3322 2362 3558
rect 2598 3322 2682 3558
rect 2918 3322 3002 3558
rect 3238 3322 3322 3558
rect 3558 3322 3642 3558
rect 3878 3322 309854 3558
rect 310090 3322 310174 3558
rect 310410 3322 310494 3558
rect 310730 3322 310814 3558
rect 311050 3322 311134 3558
rect 311370 3322 311454 3558
rect 311690 3322 311774 3558
rect 312010 3322 312094 3558
rect 312330 3322 312414 3558
rect 312650 3322 312734 3558
rect 312970 3322 313054 3558
rect 313290 3322 313374 3558
rect 313610 3322 313732 3558
rect 0 3238 313732 3322
rect 0 3002 122 3238
rect 358 3002 442 3238
rect 678 3002 762 3238
rect 998 3002 1082 3238
rect 1318 3002 1402 3238
rect 1638 3002 1722 3238
rect 1958 3002 2042 3238
rect 2278 3002 2362 3238
rect 2598 3002 2682 3238
rect 2918 3002 3002 3238
rect 3238 3002 3322 3238
rect 3558 3002 3642 3238
rect 3878 3002 309854 3238
rect 310090 3002 310174 3238
rect 310410 3002 310494 3238
rect 310730 3002 310814 3238
rect 311050 3002 311134 3238
rect 311370 3002 311454 3238
rect 311690 3002 311774 3238
rect 312010 3002 312094 3238
rect 312330 3002 312414 3238
rect 312650 3002 312734 3238
rect 312970 3002 313054 3238
rect 313290 3002 313374 3238
rect 313610 3002 313732 3238
rect 0 2918 313732 3002
rect 0 2682 122 2918
rect 358 2682 442 2918
rect 678 2682 762 2918
rect 998 2682 1082 2918
rect 1318 2682 1402 2918
rect 1638 2682 1722 2918
rect 1958 2682 2042 2918
rect 2278 2682 2362 2918
rect 2598 2682 2682 2918
rect 2918 2682 3002 2918
rect 3238 2682 3322 2918
rect 3558 2682 3642 2918
rect 3878 2682 309854 2918
rect 310090 2682 310174 2918
rect 310410 2682 310494 2918
rect 310730 2682 310814 2918
rect 311050 2682 311134 2918
rect 311370 2682 311454 2918
rect 311690 2682 311774 2918
rect 312010 2682 312094 2918
rect 312330 2682 312414 2918
rect 312650 2682 312734 2918
rect 312970 2682 313054 2918
rect 313290 2682 313374 2918
rect 313610 2682 313732 2918
rect 0 2598 313732 2682
rect 0 2362 122 2598
rect 358 2362 442 2598
rect 678 2362 762 2598
rect 998 2362 1082 2598
rect 1318 2362 1402 2598
rect 1638 2362 1722 2598
rect 1958 2362 2042 2598
rect 2278 2362 2362 2598
rect 2598 2362 2682 2598
rect 2918 2362 3002 2598
rect 3238 2362 3322 2598
rect 3558 2362 3642 2598
rect 3878 2362 309854 2598
rect 310090 2362 310174 2598
rect 310410 2362 310494 2598
rect 310730 2362 310814 2598
rect 311050 2362 311134 2598
rect 311370 2362 311454 2598
rect 311690 2362 311774 2598
rect 312010 2362 312094 2598
rect 312330 2362 312414 2598
rect 312650 2362 312734 2598
rect 312970 2362 313054 2598
rect 313290 2362 313374 2598
rect 313610 2362 313732 2598
rect 0 2278 313732 2362
rect 0 2042 122 2278
rect 358 2042 442 2278
rect 678 2042 762 2278
rect 998 2042 1082 2278
rect 1318 2042 1402 2278
rect 1638 2042 1722 2278
rect 1958 2042 2042 2278
rect 2278 2042 2362 2278
rect 2598 2042 2682 2278
rect 2918 2042 3002 2278
rect 3238 2042 3322 2278
rect 3558 2042 3642 2278
rect 3878 2042 309854 2278
rect 310090 2042 310174 2278
rect 310410 2042 310494 2278
rect 310730 2042 310814 2278
rect 311050 2042 311134 2278
rect 311370 2042 311454 2278
rect 311690 2042 311774 2278
rect 312010 2042 312094 2278
rect 312330 2042 312414 2278
rect 312650 2042 312734 2278
rect 312970 2042 313054 2278
rect 313290 2042 313374 2278
rect 313610 2042 313732 2278
rect 0 1958 313732 2042
rect 0 1722 122 1958
rect 358 1722 442 1958
rect 678 1722 762 1958
rect 998 1722 1082 1958
rect 1318 1722 1402 1958
rect 1638 1722 1722 1958
rect 1958 1722 2042 1958
rect 2278 1722 2362 1958
rect 2598 1722 2682 1958
rect 2918 1722 3002 1958
rect 3238 1722 3322 1958
rect 3558 1722 3642 1958
rect 3878 1722 309854 1958
rect 310090 1722 310174 1958
rect 310410 1722 310494 1958
rect 310730 1722 310814 1958
rect 311050 1722 311134 1958
rect 311370 1722 311454 1958
rect 311690 1722 311774 1958
rect 312010 1722 312094 1958
rect 312330 1722 312414 1958
rect 312650 1722 312734 1958
rect 312970 1722 313054 1958
rect 313290 1722 313374 1958
rect 313610 1722 313732 1958
rect 0 1638 313732 1722
rect 0 1402 122 1638
rect 358 1402 442 1638
rect 678 1402 762 1638
rect 998 1402 1082 1638
rect 1318 1402 1402 1638
rect 1638 1402 1722 1638
rect 1958 1402 2042 1638
rect 2278 1402 2362 1638
rect 2598 1402 2682 1638
rect 2918 1402 3002 1638
rect 3238 1402 3322 1638
rect 3558 1402 3642 1638
rect 3878 1402 309854 1638
rect 310090 1402 310174 1638
rect 310410 1402 310494 1638
rect 310730 1402 310814 1638
rect 311050 1402 311134 1638
rect 311370 1402 311454 1638
rect 311690 1402 311774 1638
rect 312010 1402 312094 1638
rect 312330 1402 312414 1638
rect 312650 1402 312734 1638
rect 312970 1402 313054 1638
rect 313290 1402 313374 1638
rect 313610 1402 313732 1638
rect 0 1318 313732 1402
rect 0 1082 122 1318
rect 358 1082 442 1318
rect 678 1082 762 1318
rect 998 1082 1082 1318
rect 1318 1082 1402 1318
rect 1638 1082 1722 1318
rect 1958 1082 2042 1318
rect 2278 1082 2362 1318
rect 2598 1082 2682 1318
rect 2918 1082 3002 1318
rect 3238 1082 3322 1318
rect 3558 1082 3642 1318
rect 3878 1082 309854 1318
rect 310090 1082 310174 1318
rect 310410 1082 310494 1318
rect 310730 1082 310814 1318
rect 311050 1082 311134 1318
rect 311370 1082 311454 1318
rect 311690 1082 311774 1318
rect 312010 1082 312094 1318
rect 312330 1082 312414 1318
rect 312650 1082 312734 1318
rect 312970 1082 313054 1318
rect 313290 1082 313374 1318
rect 313610 1082 313732 1318
rect 0 998 313732 1082
rect 0 762 122 998
rect 358 762 442 998
rect 678 762 762 998
rect 998 762 1082 998
rect 1318 762 1402 998
rect 1638 762 1722 998
rect 1958 762 2042 998
rect 2278 762 2362 998
rect 2598 762 2682 998
rect 2918 762 3002 998
rect 3238 762 3322 998
rect 3558 762 3642 998
rect 3878 762 309854 998
rect 310090 762 310174 998
rect 310410 762 310494 998
rect 310730 762 310814 998
rect 311050 762 311134 998
rect 311370 762 311454 998
rect 311690 762 311774 998
rect 312010 762 312094 998
rect 312330 762 312414 998
rect 312650 762 312734 998
rect 312970 762 313054 998
rect 313290 762 313374 998
rect 313610 762 313732 998
rect 0 678 313732 762
rect 0 442 122 678
rect 358 442 442 678
rect 678 442 762 678
rect 998 442 1082 678
rect 1318 442 1402 678
rect 1638 442 1722 678
rect 1958 442 2042 678
rect 2278 442 2362 678
rect 2598 442 2682 678
rect 2918 442 3002 678
rect 3238 442 3322 678
rect 3558 442 3642 678
rect 3878 442 309854 678
rect 310090 442 310174 678
rect 310410 442 310494 678
rect 310730 442 310814 678
rect 311050 442 311134 678
rect 311370 442 311454 678
rect 311690 442 311774 678
rect 312010 442 312094 678
rect 312330 442 312414 678
rect 312650 442 312734 678
rect 312970 442 313054 678
rect 313290 442 313374 678
rect 313610 442 313732 678
rect 0 358 313732 442
rect 0 122 122 358
rect 358 122 442 358
rect 678 122 762 358
rect 998 122 1082 358
rect 1318 122 1402 358
rect 1638 122 1722 358
rect 1958 122 2042 358
rect 2278 122 2362 358
rect 2598 122 2682 358
rect 2918 122 3002 358
rect 3238 122 3322 358
rect 3558 122 3642 358
rect 3878 122 309854 358
rect 310090 122 310174 358
rect 310410 122 310494 358
rect 310730 122 310814 358
rect 311050 122 311134 358
rect 311370 122 311454 358
rect 311690 122 311774 358
rect 312010 122 312094 358
rect 312330 122 312414 358
rect 312650 122 312734 358
rect 312970 122 313054 358
rect 313290 122 313374 358
rect 313610 122 313732 358
rect 0 0 313732 122
use sb_0__0_  sb_0__0_
timestamp 1604349425
transform 1 0 48896 0 1 47824
box 0 0 28000 28000
use grid_io_bottom  grid_io_bottom_1__0_
timestamp 1604349425
transform 1 0 89896 0 1 18824
box 0 0 40000 16000
use cbx_1__0_  cbx_1__0_
timestamp 1604349425
transform 1 0 89896 0 1 53824
box 0 0 40000 16000
use sb_1__0_  sb_1__0_
timestamp 1604349425
transform 1 0 142896 0 1 47824
box 0 0 28000 28000
use grid_io_bottom  grid_io_bottom_2__0_
timestamp 1604349425
transform 1 0 183896 0 1 18824
box 0 0 40000 16000
use cbx_1__0_  cbx_2__0_
timestamp 1604349425
transform 1 0 183896 0 1 53824
box 0 0 40000 16000
use sb_2__0_  sb_2__0_
timestamp 1604349425
transform 1 0 236896 0 1 47824
box 0 0 28000 28000
use grid_io_left  grid_io_left_0__1_
timestamp 1604349425
transform 1 0 19896 0 1 88824
box 0 0 16000 40000
use cby_0__1_  cby_0__1_
timestamp 1604349425
transform 1 0 54896 0 1 88824
box 0 0 16000 40000
use grid_clb  grid_clb_1__1_
timestamp 1604349425
transform 1 0 84896 0 1 83824
box 0 0 50000 50000
use cby_1__1_  cby_1__1_
timestamp 1604349425
transform 1 0 148896 0 1 88824
box 0 0 16000 40000
use grid_clb  grid_clb_2__1_
timestamp 1604349425
transform 1 0 178896 0 1 83824
box 0 0 50000 50000
use cby_1__1_  cby_2__1_
timestamp 1604349425
transform 1 0 242896 0 1 88824
box 0 0 16000 40000
use grid_io_right  grid_io_right_3__1_
timestamp 1604349425
transform 1 0 277896 0 1 88824
box 0 0 16000 40000
use grid_io_left  grid_io_left_0__2_
timestamp 1604349425
transform 1 0 19896 0 1 182824
box 0 0 16000 40000
use sb_0__1_  sb_0__1_
timestamp 1604349425
transform 1 0 48896 0 1 141824
box 0 0 28000 28000
use cby_0__1_  cby_0__2_
timestamp 1604349425
transform 1 0 54896 0 1 182824
box 0 0 16000 40000
use grid_clb  grid_clb_1__2_
timestamp 1604349425
transform 1 0 84896 0 1 177824
box 0 0 50000 50000
use cbx_1__1_  cbx_1__1_
timestamp 1604349425
transform 1 0 89896 0 1 147824
box 0 0 40000 16000
use sb_1__1_  sb_1__1_
timestamp 1604349425
transform 1 0 142896 0 1 141824
box 0 0 28000 28000
use cby_1__1_  cby_1__2_
timestamp 1604349425
transform 1 0 148896 0 1 182824
box 0 0 16000 40000
use grid_clb  grid_clb_2__2_
timestamp 1604349425
transform 1 0 178896 0 1 177824
box 0 0 50000 50000
use cbx_1__1_  cbx_2__1_
timestamp 1604349425
transform 1 0 183896 0 1 147824
box 0 0 40000 16000
use sb_2__1_  sb_2__1_
timestamp 1604349425
transform 1 0 236896 0 1 141824
box 0 0 28000 28000
use cby_1__1_  cby_2__2_
timestamp 1604349425
transform 1 0 242896 0 1 182824
box 0 0 16000 40000
use grid_io_right  grid_io_right_3__2_
timestamp 1604349425
transform 1 0 277896 0 1 182824
box 0 0 16000 40000
use sb_0__2_  sb_0__2_
timestamp 1604349425
transform 1 0 48896 0 1 235824
box 0 0 28000 28000
use sb_1__2_  sb_1__2_
timestamp 1604349425
transform 1 0 142896 0 1 235824
box 0 0 28000 27736
use sb_2__2_  sb_2__2_
timestamp 1604349425
transform 1 0 236896 0 1 235824
box 0 0 28000 27600
use grid_io_top  grid_io_top_1__3_
timestamp 1604349425
transform 1 0 89896 0 1 276824
box 0 0 40000 16000
use cbx_1__2_  cbx_1__2_
timestamp 1604349425
transform 1 0 89896 0 1 241824
box 0 0 40000 16000
use grid_io_top  grid_io_top_2__3_
timestamp 1604349425
transform 1 0 183896 0 1 276824
box 0 0 40000 16000
use cbx_1__2_  cbx_2__2_
timestamp 1604349425
transform 1 0 183896 0 1 241824
box 0 0 40000 16000
<< labels >>
rlabel metal2 s 28222 8824 28278 9304 6 Test_en
port 0 nsew default input
rlabel metal2 s 64930 8824 64986 9304 6 ccff_head
port 1 nsew default input
rlabel metal3 s 303416 21072 303896 21192 6 ccff_tail
port 2 nsew default tristate
rlabel metal3 s 9896 25152 10376 25272 6 clk
port 3 nsew default input
rlabel metal2 s 101730 8824 101786 9304 6 gfpga_pad_GPIO_A[0]
port 4 nsew default tristate
rlabel metal3 s 9896 57792 10376 57912 6 gfpga_pad_GPIO_A[1]
port 5 nsew default tristate
rlabel metal3 s 303416 45552 303896 45672 6 gfpga_pad_GPIO_A[2]
port 6 nsew default tristate
rlabel metal3 s 303416 70032 303896 70152 6 gfpga_pad_GPIO_A[3]
port 7 nsew default tristate
rlabel metal3 s 303416 94512 303896 94632 6 gfpga_pad_GPIO_A[4]
port 8 nsew default tristate
rlabel metal3 s 303416 118992 303896 119112 6 gfpga_pad_GPIO_A[5]
port 9 nsew default tristate
rlabel metal3 s 9896 90432 10376 90552 6 gfpga_pad_GPIO_A[6]
port 10 nsew default tristate
rlabel metal2 s 28222 302344 28278 302824 6 gfpga_pad_GPIO_A[7]
port 11 nsew default tristate
rlabel metal2 s 64930 302344 64986 302824 6 gfpga_pad_GPIO_IE[0]
port 12 nsew default tristate
rlabel metal3 s 9896 123072 10376 123192 6 gfpga_pad_GPIO_IE[1]
port 13 nsew default tristate
rlabel metal2 s 101730 302344 101786 302824 6 gfpga_pad_GPIO_IE[2]
port 14 nsew default tristate
rlabel metal3 s 303416 143472 303896 143592 6 gfpga_pad_GPIO_IE[3]
port 15 nsew default tristate
rlabel metal3 s 9896 155712 10376 155832 6 gfpga_pad_GPIO_IE[4]
port 16 nsew default tristate
rlabel metal3 s 303416 168088 303896 168208 6 gfpga_pad_GPIO_IE[5]
port 17 nsew default tristate
rlabel metal2 s 138438 8824 138494 9304 6 gfpga_pad_GPIO_IE[6]
port 18 nsew default tristate
rlabel metal3 s 303416 192568 303896 192688 6 gfpga_pad_GPIO_IE[7]
port 19 nsew default tristate
rlabel metal3 s 303416 217048 303896 217168 6 gfpga_pad_GPIO_OE[0]
port 20 nsew default tristate
rlabel metal2 s 138438 302344 138494 302824 6 gfpga_pad_GPIO_OE[1]
port 21 nsew default tristate
rlabel metal2 s 175238 8824 175294 9304 6 gfpga_pad_GPIO_OE[2]
port 22 nsew default tristate
rlabel metal2 s 175238 302344 175294 302824 6 gfpga_pad_GPIO_OE[3]
port 23 nsew default tristate
rlabel metal3 s 9896 188488 10376 188608 6 gfpga_pad_GPIO_OE[4]
port 24 nsew default tristate
rlabel metal2 s 211946 8824 212002 9304 6 gfpga_pad_GPIO_OE[5]
port 25 nsew default tristate
rlabel metal2 s 211946 302344 212002 302824 6 gfpga_pad_GPIO_OE[6]
port 26 nsew default tristate
rlabel metal3 s 9896 221128 10376 221248 6 gfpga_pad_GPIO_OE[7]
port 27 nsew default tristate
rlabel metal3 s 303416 241528 303896 241648 6 gfpga_pad_GPIO_Y[0]
port 28 nsew default bidirectional
rlabel metal3 s 303416 266008 303896 266128 6 gfpga_pad_GPIO_Y[1]
port 29 nsew default bidirectional
rlabel metal3 s 9896 253768 10376 253888 6 gfpga_pad_GPIO_Y[2]
port 30 nsew default bidirectional
rlabel metal2 s 248746 302344 248802 302824 6 gfpga_pad_GPIO_Y[3]
port 31 nsew default bidirectional
rlabel metal2 s 248746 8824 248802 9304 6 gfpga_pad_GPIO_Y[4]
port 32 nsew default bidirectional
rlabel metal3 s 303416 290488 303896 290608 6 gfpga_pad_GPIO_Y[5]
port 33 nsew default bidirectional
rlabel metal2 s 285454 302344 285510 302824 6 gfpga_pad_GPIO_Y[6]
port 34 nsew default bidirectional
rlabel metal3 s 9896 286408 10376 286528 6 gfpga_pad_GPIO_Y[7]
port 35 nsew default bidirectional
rlabel metal2 s 285454 8824 285510 9304 6 prog_clk
port 36 nsew default input
rlabel metal5 s 5000 5000 308732 9000 8 vpwr
port 37 nsew default input
rlabel metal5 s 0 0 313732 4000 8 vgnd
port 38 nsew default input
<< properties >>
string FIXED_BBOX 0 0 313732 311408
<< end >>
