magic
tech EFS8A
magscale 1 2
timestamp 1602874717
<< locali >>
rect 2881 19159 2915 19261
rect 29 16779 63 17425
rect 3617 11067 3651 11305
rect 4721 10455 4755 10693
rect 2973 9503 3007 9605
rect 3893 9027 3927 9129
rect 3617 7871 3651 7973
rect 2421 4063 2455 4165
rect 3709 2431 3743 2533
<< viali >>
rect 1685 21301 1719 21335
rect 1501 21097 1535 21131
rect 4169 21097 4203 21131
rect 1685 20961 1719 20995
rect 1961 20961 1995 20995
rect 4077 20961 4111 20995
rect 4629 20961 4663 20995
rect 2421 20757 2455 20791
rect 3157 20757 3191 20791
rect 5181 20757 5215 20791
rect 3617 20417 3651 20451
rect 1685 20349 1719 20383
rect 1961 20349 1995 20383
rect 3065 20349 3099 20383
rect 3525 20349 3559 20383
rect 4537 20349 4571 20383
rect 4629 20349 4663 20383
rect 5181 20349 5215 20383
rect 1501 20213 1535 20247
rect 2421 20213 2455 20247
rect 2789 20213 2823 20247
rect 4077 20213 4111 20247
rect 4721 20213 4755 20247
rect 1593 20009 1627 20043
rect 4629 20009 4663 20043
rect 6285 20009 6319 20043
rect 4353 19941 4387 19975
rect 1685 19873 1719 19907
rect 2099 19873 2133 19907
rect 4537 19873 4571 19907
rect 5089 19873 5123 19907
rect 6101 19873 6135 19907
rect 3065 19669 3099 19703
rect 2053 19465 2087 19499
rect 4261 19465 4295 19499
rect 4537 19465 4571 19499
rect 7021 19465 7055 19499
rect 3709 19329 3743 19363
rect 1685 19261 1719 19295
rect 2881 19261 2915 19295
rect 3157 19261 3191 19295
rect 3617 19261 3651 19295
rect 4905 19261 4939 19295
rect 5457 19261 5491 19295
rect 6837 19261 6871 19295
rect 7297 19261 7331 19295
rect 2881 19125 2915 19159
rect 2973 19125 3007 19159
rect 4997 19125 5031 19159
rect 5917 19125 5951 19159
rect 6285 19125 6319 19159
rect 1777 18921 1811 18955
rect 3249 18921 3283 18955
rect 3893 18921 3927 18955
rect 4353 18921 4387 18955
rect 5825 18921 5859 18955
rect 1961 18785 1995 18819
rect 2237 18785 2271 18819
rect 2697 18785 2731 18819
rect 4077 18785 4111 18819
rect 4629 18785 4663 18819
rect 5641 18785 5675 18819
rect 5273 18581 5307 18615
rect 6193 18581 6227 18615
rect 5457 18377 5491 18411
rect 5825 18377 5859 18411
rect 2329 18241 2363 18275
rect 4353 18241 4387 18275
rect 5089 18241 5123 18275
rect 5549 18241 5583 18275
rect 1777 18173 1811 18207
rect 2237 18173 2271 18207
rect 3341 18173 3375 18207
rect 3801 18173 3835 18207
rect 5328 18173 5362 18207
rect 6837 18173 6871 18207
rect 7297 18173 7331 18207
rect 5181 18105 5215 18139
rect 6285 18105 6319 18139
rect 1685 18037 1719 18071
rect 2789 18037 2823 18071
rect 3249 18037 3283 18071
rect 3433 18037 3467 18071
rect 6561 18037 6595 18071
rect 7021 18037 7055 18071
rect 1501 17833 1535 17867
rect 2421 17833 2455 17867
rect 3341 17833 3375 17867
rect 3801 17833 3835 17867
rect 6193 17833 6227 17867
rect 6929 17833 6963 17867
rect 5825 17765 5859 17799
rect 1685 17697 1719 17731
rect 1961 17697 1995 17731
rect 2789 17697 2823 17731
rect 4077 17697 4111 17731
rect 5089 17697 5123 17731
rect 6745 17697 6779 17731
rect 5457 17629 5491 17663
rect 6561 17629 6595 17663
rect 5254 17561 5288 17595
rect 4261 17493 4295 17527
rect 4537 17493 4571 17527
rect 4905 17493 4939 17527
rect 5365 17493 5399 17527
rect 29 17425 63 17459
rect 5346 17289 5380 17323
rect 5825 17289 5859 17323
rect 5457 17221 5491 17255
rect 6193 17221 6227 17255
rect 7021 17221 7055 17255
rect 3617 17153 3651 17187
rect 5549 17153 5583 17187
rect 1685 17085 1719 17119
rect 1961 17085 1995 17119
rect 3341 17085 3375 17119
rect 3525 17085 3559 17119
rect 6837 17085 6871 17119
rect 2973 17017 3007 17051
rect 5181 17017 5215 17051
rect 1501 16949 1535 16983
rect 2421 16949 2455 16983
rect 4353 16949 4387 16983
rect 4629 16949 4663 16983
rect 5089 16949 5123 16983
rect 6653 16949 6687 16983
rect 7389 16949 7423 16983
rect 29 16745 63 16779
rect 2145 16745 2179 16779
rect 4261 16745 4295 16779
rect 6929 16745 6963 16779
rect 3065 16677 3099 16711
rect 3433 16677 3467 16711
rect 4813 16677 4847 16711
rect 5917 16677 5951 16711
rect 2329 16609 2363 16643
rect 2513 16609 2547 16643
rect 4077 16609 4111 16643
rect 5181 16609 5215 16643
rect 6193 16609 6227 16643
rect 6745 16609 6779 16643
rect 3893 16541 3927 16575
rect 5549 16541 5583 16575
rect 1685 16405 1719 16439
rect 5328 16405 5362 16439
rect 5457 16405 5491 16439
rect 5181 16201 5215 16235
rect 5733 16201 5767 16235
rect 6469 16201 6503 16235
rect 7757 16201 7791 16235
rect 4629 16133 4663 16167
rect 4997 16133 5031 16167
rect 7021 16133 7055 16167
rect 2973 16065 3007 16099
rect 4261 16065 4295 16099
rect 5089 16065 5123 16099
rect 6101 16065 6135 16099
rect 1593 15997 1627 16031
rect 2145 15997 2179 16031
rect 3157 15997 3191 16031
rect 3709 15997 3743 16031
rect 4868 15997 4902 16031
rect 6837 15997 6871 16031
rect 7849 15997 7883 16031
rect 8309 15997 8343 16031
rect 4721 15929 4755 15963
rect 7389 15929 7423 15963
rect 1685 15861 1719 15895
rect 2697 15861 2731 15895
rect 3249 15861 3283 15895
rect 8033 15861 8067 15895
rect 1869 15657 1903 15691
rect 2881 15657 2915 15691
rect 3893 15657 3927 15691
rect 4629 15657 4663 15691
rect 6469 15657 6503 15691
rect 3249 15589 3283 15623
rect 6193 15589 6227 15623
rect 7389 15589 7423 15623
rect 1869 15521 1903 15555
rect 2329 15521 2363 15555
rect 4721 15521 4755 15555
rect 7297 15521 7331 15555
rect 5089 15453 5123 15487
rect 5181 15385 5215 15419
rect 1593 15317 1627 15351
rect 4859 15317 4893 15351
rect 4997 15317 5031 15351
rect 5733 15317 5767 15351
rect 3341 15113 3375 15147
rect 3801 15113 3835 15147
rect 4077 15113 4111 15147
rect 4721 15113 4755 15147
rect 5089 15113 5123 15147
rect 5346 15113 5380 15147
rect 6653 15113 6687 15147
rect 6975 15113 7009 15147
rect 5457 15045 5491 15079
rect 6285 15045 6319 15079
rect 2881 14977 2915 15011
rect 5549 14977 5583 15011
rect 7205 14977 7239 15011
rect 7297 14977 7331 15011
rect 2237 14909 2271 14943
rect 2605 14909 2639 14943
rect 2789 14909 2823 14943
rect 3893 14909 3927 14943
rect 7067 14909 7101 14943
rect 7849 14909 7883 14943
rect 5181 14841 5215 14875
rect 6837 14841 6871 14875
rect 1869 14773 1903 14807
rect 5825 14773 5859 14807
rect 2329 14569 2363 14603
rect 3893 14569 3927 14603
rect 7573 14569 7607 14603
rect 1869 14501 1903 14535
rect 5089 14501 5123 14535
rect 7113 14501 7147 14535
rect 2237 14433 2271 14467
rect 2789 14433 2823 14467
rect 4077 14433 4111 14467
rect 5236 14433 5270 14467
rect 6101 14433 6135 14467
rect 6653 14433 6687 14467
rect 5457 14365 5491 14399
rect 3341 14297 3375 14331
rect 5365 14297 5399 14331
rect 4261 14229 4295 14263
rect 4721 14229 4755 14263
rect 5733 14229 5767 14263
rect 6837 14229 6871 14263
rect 2513 14025 2547 14059
rect 4629 14025 4663 14059
rect 4905 14025 4939 14059
rect 6101 14025 6135 14059
rect 6561 14025 6595 14059
rect 5365 13957 5399 13991
rect 5457 13889 5491 13923
rect 7849 13889 7883 13923
rect 1685 13821 1719 13855
rect 1961 13821 1995 13855
rect 2973 13821 3007 13855
rect 3525 13821 3559 13855
rect 5089 13821 5123 13855
rect 5236 13821 5270 13855
rect 7021 13821 7055 13855
rect 7297 13821 7331 13855
rect 2881 13753 2915 13787
rect 4261 13753 4295 13787
rect 1501 13685 1535 13719
rect 3065 13685 3099 13719
rect 5733 13685 5767 13719
rect 6929 13685 6963 13719
rect 1593 13481 1627 13515
rect 1961 13481 1995 13515
rect 2513 13481 2547 13515
rect 3893 13481 3927 13515
rect 4353 13481 4387 13515
rect 5457 13481 5491 13515
rect 6561 13481 6595 13515
rect 6929 13481 6963 13515
rect 5825 13413 5859 13447
rect 6193 13413 6227 13447
rect 1409 13345 1443 13379
rect 2421 13345 2455 13379
rect 2881 13345 2915 13379
rect 4813 13345 4847 13379
rect 4960 13345 4994 13379
rect 6377 13345 6411 13379
rect 7573 13345 7607 13379
rect 4721 13277 4755 13311
rect 5181 13277 5215 13311
rect 7297 13277 7331 13311
rect 7389 13277 7423 13311
rect 2329 13209 2363 13243
rect 3433 13141 3467 13175
rect 5089 13141 5123 13175
rect 1685 12937 1719 12971
rect 4813 12937 4847 12971
rect 5917 12937 5951 12971
rect 8125 12937 8159 12971
rect 5181 12869 5215 12903
rect 4077 12801 4111 12835
rect 4445 12801 4479 12835
rect 5273 12801 5307 12835
rect 1501 12733 1535 12767
rect 2789 12733 2823 12767
rect 2973 12733 3007 12767
rect 3617 12733 3651 12767
rect 5052 12733 5086 12767
rect 7389 12733 7423 12767
rect 2053 12665 2087 12699
rect 2421 12665 2455 12699
rect 4905 12665 4939 12699
rect 7113 12665 7147 12699
rect 2605 12597 2639 12631
rect 5549 12597 5583 12631
rect 6377 12597 6411 12631
rect 2513 12393 2547 12427
rect 4169 12393 4203 12427
rect 5457 12393 5491 12427
rect 7205 12393 7239 12427
rect 6101 12325 6135 12359
rect 7665 12325 7699 12359
rect 1409 12257 1443 12291
rect 2421 12257 2455 12291
rect 2881 12257 2915 12291
rect 4261 12257 4295 12291
rect 4537 12257 4571 12291
rect 6248 12257 6282 12291
rect 7812 12257 7846 12291
rect 3433 12189 3467 12223
rect 6469 12189 6503 12223
rect 8033 12189 8067 12223
rect 3801 12121 3835 12155
rect 5917 12121 5951 12155
rect 6377 12121 6411 12155
rect 7481 12121 7515 12155
rect 7941 12121 7975 12155
rect 1593 12053 1627 12087
rect 1961 12053 1995 12087
rect 2329 12053 2363 12087
rect 5181 12053 5215 12087
rect 6745 12053 6779 12087
rect 8125 12053 8159 12087
rect 2513 11849 2547 11883
rect 4169 11849 4203 11883
rect 5089 11849 5123 11883
rect 5825 11849 5859 11883
rect 6193 11849 6227 11883
rect 6653 11849 6687 11883
rect 7002 11849 7036 11883
rect 8217 11849 8251 11883
rect 4813 11781 4847 11815
rect 5549 11781 5583 11815
rect 7113 11781 7147 11815
rect 7849 11781 7883 11815
rect 7205 11713 7239 11747
rect 1685 11645 1719 11679
rect 1869 11645 1903 11679
rect 2973 11645 3007 11679
rect 3341 11645 3375 11679
rect 3525 11645 3559 11679
rect 4629 11645 4663 11679
rect 5641 11645 5675 11679
rect 6837 11645 6871 11679
rect 8401 11645 8435 11679
rect 8861 11645 8895 11679
rect 1501 11509 1535 11543
rect 3157 11509 3191 11543
rect 4537 11509 4571 11543
rect 7481 11509 7515 11543
rect 8585 11509 8619 11543
rect 1501 11305 1535 11339
rect 2789 11305 2823 11339
rect 3433 11305 3467 11339
rect 3617 11305 3651 11339
rect 6377 11305 6411 11339
rect 6837 11305 6871 11339
rect 7757 11305 7791 11339
rect 8125 11305 8159 11339
rect 1685 11169 1719 11203
rect 1961 11169 1995 11203
rect 2513 11169 2547 11203
rect 2973 11169 3007 11203
rect 3801 11237 3835 11271
rect 5273 11237 5307 11271
rect 5641 11237 5675 11271
rect 5733 11237 5767 11271
rect 4629 11169 4663 11203
rect 5880 11169 5914 11203
rect 7297 11169 7331 11203
rect 6101 11101 6135 11135
rect 3617 11033 3651 11067
rect 4813 11033 4847 11067
rect 3157 10965 3191 10999
rect 4261 10965 4295 10999
rect 6009 10965 6043 10999
rect 7481 10965 7515 10999
rect 2421 10761 2455 10795
rect 2789 10761 2823 10795
rect 4077 10761 4111 10795
rect 6101 10761 6135 10795
rect 6377 10761 6411 10795
rect 7297 10761 7331 10795
rect 7665 10761 7699 10795
rect 4721 10693 4755 10727
rect 7021 10693 7055 10727
rect 1685 10557 1719 10591
rect 1961 10557 1995 10591
rect 3249 10557 3283 10591
rect 3525 10557 3559 10591
rect 5365 10557 5399 10591
rect 6837 10557 6871 10591
rect 8033 10557 8067 10591
rect 4997 10489 5031 10523
rect 1501 10421 1535 10455
rect 3065 10421 3099 10455
rect 4537 10421 4571 10455
rect 4721 10421 4755 10455
rect 4905 10421 4939 10455
rect 1593 10217 1627 10251
rect 1869 10217 1903 10251
rect 2329 10217 2363 10251
rect 2513 10217 2547 10251
rect 3801 10217 3835 10251
rect 4261 10217 4295 10251
rect 4537 10217 4571 10251
rect 4997 10217 5031 10251
rect 6469 10217 6503 10251
rect 6193 10149 6227 10183
rect 1409 10081 1443 10115
rect 2697 10081 2731 10115
rect 2973 10081 3007 10115
rect 4077 10081 4111 10115
rect 5089 10081 5123 10115
rect 5365 10081 5399 10115
rect 6653 10081 6687 10115
rect 6929 10081 6963 10115
rect 3525 10013 3559 10047
rect 5549 10013 5583 10047
rect 7113 10013 7147 10047
rect 5181 9945 5215 9979
rect 6745 9945 6779 9979
rect 2697 9673 2731 9707
rect 4629 9673 4663 9707
rect 4997 9673 5031 9707
rect 7021 9673 7055 9707
rect 2973 9605 3007 9639
rect 3157 9537 3191 9571
rect 1961 9469 1995 9503
rect 2237 9469 2271 9503
rect 2973 9469 3007 9503
rect 3249 9469 3283 9503
rect 3801 9469 3835 9503
rect 5089 9469 5123 9503
rect 5181 9469 5215 9503
rect 5365 9469 5399 9503
rect 1777 9333 1811 9367
rect 3341 9333 3375 9367
rect 5549 9333 5583 9367
rect 6193 9333 6227 9367
rect 6561 9333 6595 9367
rect 7389 9333 7423 9367
rect 1685 9129 1719 9163
rect 2605 9129 2639 9163
rect 3065 9129 3099 9163
rect 3709 9129 3743 9163
rect 3893 9129 3927 9163
rect 4261 9129 4295 9163
rect 5641 9129 5675 9163
rect 6653 9129 6687 9163
rect 5089 9061 5123 9095
rect 1869 8993 1903 9027
rect 2053 8993 2087 9027
rect 3433 8993 3467 9027
rect 3893 8993 3927 9027
rect 4077 8993 4111 9027
rect 5181 8993 5215 9027
rect 5457 8993 5491 9027
rect 4537 8925 4571 8959
rect 5273 8857 5307 8891
rect 4813 8585 4847 8619
rect 5365 8585 5399 8619
rect 4445 8517 4479 8551
rect 5917 8449 5951 8483
rect 1777 8381 1811 8415
rect 2053 8381 2087 8415
rect 2605 8381 2639 8415
rect 2973 8381 3007 8415
rect 3617 8381 3651 8415
rect 3893 8381 3927 8415
rect 5181 8381 5215 8415
rect 1593 8245 1627 8279
rect 3433 8245 3467 8279
rect 6285 8245 6319 8279
rect 1593 8041 1627 8075
rect 2513 8041 2547 8075
rect 3433 8041 3467 8075
rect 5273 8041 5307 8075
rect 3617 7973 3651 8007
rect 4905 7973 4939 8007
rect 5549 7973 5583 8007
rect 1593 7905 1627 7939
rect 2053 7905 2087 7939
rect 4077 7905 4111 7939
rect 4629 7905 4663 7939
rect 5089 7905 5123 7939
rect 6101 7905 6135 7939
rect 3617 7837 3651 7871
rect 3709 7837 3743 7871
rect 2973 7769 3007 7803
rect 4261 7769 4295 7803
rect 6285 7769 6319 7803
rect 2513 7497 2547 7531
rect 4353 7497 4387 7531
rect 4905 7497 4939 7531
rect 6101 7497 6135 7531
rect 7297 7497 7331 7531
rect 5365 7429 5399 7463
rect 1777 7293 1811 7327
rect 2053 7293 2087 7327
rect 3617 7293 3651 7327
rect 3893 7293 3927 7327
rect 5457 7293 5491 7327
rect 6653 7293 6687 7327
rect 7481 7293 7515 7327
rect 2973 7225 3007 7259
rect 1593 7157 1627 7191
rect 3433 7157 3467 7191
rect 5641 7157 5675 7191
rect 1501 6953 1535 6987
rect 2421 6953 2455 6987
rect 3709 6953 3743 6987
rect 4169 6953 4203 6987
rect 1685 6817 1719 6851
rect 1961 6817 1995 6851
rect 2881 6817 2915 6851
rect 4353 6817 4387 6851
rect 4629 6817 4663 6851
rect 5641 6817 5675 6851
rect 3433 6613 3467 6647
rect 5825 6613 5859 6647
rect 3249 6409 3283 6443
rect 5641 6409 5675 6443
rect 4353 6273 4387 6307
rect 1685 6205 1719 6239
rect 1961 6205 1995 6239
rect 2513 6205 2547 6239
rect 2881 6205 2915 6239
rect 3617 6205 3651 6239
rect 3985 6205 4019 6239
rect 4261 6205 4295 6239
rect 1501 6069 1535 6103
rect 4721 6069 4755 6103
rect 1685 5865 1719 5899
rect 2697 5865 2731 5899
rect 3065 5865 3099 5899
rect 3893 5865 3927 5899
rect 4169 5865 4203 5899
rect 1869 5729 1903 5763
rect 2053 5729 2087 5763
rect 4077 5729 4111 5763
rect 4537 5729 4571 5763
rect 3433 5661 3467 5695
rect 4445 5321 4479 5355
rect 5181 5321 5215 5355
rect 4813 5253 4847 5287
rect 1685 5117 1719 5151
rect 2053 5117 2087 5151
rect 2513 5117 2547 5151
rect 2881 5117 2915 5151
rect 3065 5117 3099 5151
rect 3525 5117 3559 5151
rect 4629 5117 4663 5151
rect 1593 4981 1627 5015
rect 3157 4981 3191 5015
rect 4077 4981 4111 5015
rect 1685 4777 1719 4811
rect 3065 4777 3099 4811
rect 3525 4777 3559 4811
rect 3893 4777 3927 4811
rect 4169 4777 4203 4811
rect 1869 4641 1903 4675
rect 2145 4641 2179 4675
rect 2697 4641 2731 4675
rect 4077 4641 4111 4675
rect 4537 4641 4571 4675
rect 5365 4233 5399 4267
rect 2421 4165 2455 4199
rect 2697 4165 2731 4199
rect 3065 4165 3099 4199
rect 3525 4165 3559 4199
rect 4629 4165 4663 4199
rect 4169 4097 4203 4131
rect 4997 4097 5031 4131
rect 1593 4029 1627 4063
rect 2145 4029 2179 4063
rect 2421 4029 2455 4063
rect 3801 4029 3835 4063
rect 4077 4029 4111 4063
rect 5181 4029 5215 4063
rect 5641 4029 5675 4063
rect 1685 3893 1719 3927
rect 1777 3689 1811 3723
rect 3525 3689 3559 3723
rect 3893 3689 3927 3723
rect 2697 3621 2731 3655
rect 3065 3621 3099 3655
rect 1685 3553 1719 3587
rect 2237 3553 2271 3587
rect 4077 3553 4111 3587
rect 4629 3553 4663 3587
rect 4537 3485 4571 3519
rect 5089 3145 5123 3179
rect 5825 3145 5859 3179
rect 4813 3077 4847 3111
rect 5457 3077 5491 3111
rect 3617 3009 3651 3043
rect 1777 2941 1811 2975
rect 2145 2941 2179 2975
rect 2605 2941 2639 2975
rect 3893 2941 3927 2975
rect 4261 2941 4295 2975
rect 5273 2941 5307 2975
rect 1685 2805 1719 2839
rect 2973 2805 3007 2839
rect 3801 2805 3835 2839
rect 1777 2601 1811 2635
rect 3157 2601 3191 2635
rect 3433 2533 3467 2567
rect 3709 2533 3743 2567
rect 1777 2465 1811 2499
rect 2237 2465 2271 2499
rect 2697 2465 2731 2499
rect 4077 2465 4111 2499
rect 4629 2465 4663 2499
rect 3709 2397 3743 2431
rect 3801 2397 3835 2431
rect 4537 2397 4571 2431
<< metal1 >>
rect 1946 23536 1952 23588
rect 2004 23576 2010 23588
rect 2590 23576 2596 23588
rect 2004 23548 2596 23576
rect 2004 23536 2010 23548
rect 2590 23536 2596 23548
rect 2648 23536 2654 23588
rect 106 21836 112 21888
rect 164 21876 170 21888
rect 4154 21876 4160 21888
rect 164 21848 4160 21876
rect 164 21836 170 21848
rect 4154 21836 4160 21848
rect 4212 21836 4218 21888
rect 1104 21786 22816 21808
rect 1104 21734 4982 21786
rect 5034 21734 5046 21786
rect 5098 21734 5110 21786
rect 5162 21734 5174 21786
rect 5226 21734 12982 21786
rect 13034 21734 13046 21786
rect 13098 21734 13110 21786
rect 13162 21734 13174 21786
rect 13226 21734 20982 21786
rect 21034 21734 21046 21786
rect 21098 21734 21110 21786
rect 21162 21734 21174 21786
rect 21226 21734 22816 21786
rect 1104 21712 22816 21734
rect 106 21360 112 21412
rect 164 21360 170 21412
rect 124 21128 152 21360
rect 1673 21335 1731 21341
rect 1673 21301 1685 21335
rect 1719 21332 1731 21335
rect 2130 21332 2136 21344
rect 1719 21304 2136 21332
rect 1719 21301 1731 21304
rect 1673 21295 1731 21301
rect 2130 21292 2136 21304
rect 2188 21292 2194 21344
rect 1104 21242 22816 21264
rect 1104 21190 8982 21242
rect 9034 21190 9046 21242
rect 9098 21190 9110 21242
rect 9162 21190 9174 21242
rect 9226 21190 16982 21242
rect 17034 21190 17046 21242
rect 17098 21190 17110 21242
rect 17162 21190 17174 21242
rect 17226 21190 22816 21242
rect 1104 21168 22816 21190
rect 1489 21131 1547 21137
rect 1489 21128 1501 21131
rect 124 21100 1501 21128
rect 1489 21097 1501 21100
rect 1535 21097 1547 21131
rect 4154 21128 4160 21140
rect 4115 21100 4160 21128
rect 1489 21091 1547 21097
rect 4154 21088 4160 21100
rect 4212 21088 4218 21140
rect 1673 20995 1731 21001
rect 1673 20961 1685 20995
rect 1719 20961 1731 20995
rect 1673 20955 1731 20961
rect 1949 20995 2007 21001
rect 1949 20961 1961 20995
rect 1995 20992 2007 20995
rect 2130 20992 2136 21004
rect 1995 20964 2136 20992
rect 1995 20961 2007 20964
rect 1949 20955 2007 20961
rect 1688 20924 1716 20955
rect 2130 20952 2136 20964
rect 2188 20952 2194 21004
rect 4062 20992 4068 21004
rect 4023 20964 4068 20992
rect 4062 20952 4068 20964
rect 4120 20952 4126 21004
rect 4617 20995 4675 21001
rect 4617 20961 4629 20995
rect 4663 20992 4675 20995
rect 4663 20964 5212 20992
rect 4663 20961 4675 20964
rect 4617 20955 4675 20961
rect 2498 20924 2504 20936
rect 1688 20896 2504 20924
rect 2498 20884 2504 20896
rect 2556 20884 2562 20936
rect 2130 20748 2136 20800
rect 2188 20788 2194 20800
rect 2409 20791 2467 20797
rect 2409 20788 2421 20791
rect 2188 20760 2421 20788
rect 2188 20748 2194 20760
rect 2409 20757 2421 20760
rect 2455 20757 2467 20791
rect 2409 20751 2467 20757
rect 3145 20791 3203 20797
rect 3145 20757 3157 20791
rect 3191 20788 3203 20791
rect 3510 20788 3516 20800
rect 3191 20760 3516 20788
rect 3191 20757 3203 20760
rect 3145 20751 3203 20757
rect 3510 20748 3516 20760
rect 3568 20788 3574 20800
rect 5184 20797 5212 20964
rect 5169 20791 5227 20797
rect 5169 20788 5181 20791
rect 3568 20760 5181 20788
rect 3568 20748 3574 20760
rect 5169 20757 5181 20760
rect 5215 20788 5227 20791
rect 5350 20788 5356 20800
rect 5215 20760 5356 20788
rect 5215 20757 5227 20760
rect 5169 20751 5227 20757
rect 5350 20748 5356 20760
rect 5408 20748 5414 20800
rect 1104 20698 22816 20720
rect 1104 20646 4982 20698
rect 5034 20646 5046 20698
rect 5098 20646 5110 20698
rect 5162 20646 5174 20698
rect 5226 20646 12982 20698
rect 13034 20646 13046 20698
rect 13098 20646 13110 20698
rect 13162 20646 13174 20698
rect 13226 20646 20982 20698
rect 21034 20646 21046 20698
rect 21098 20646 21110 20698
rect 21162 20646 21174 20698
rect 21226 20646 22816 20698
rect 1104 20624 22816 20646
rect 14 20408 20 20460
rect 72 20448 78 20460
rect 3605 20451 3663 20457
rect 3605 20448 3617 20451
rect 72 20420 3617 20448
rect 72 20408 78 20420
rect 3605 20417 3617 20420
rect 3651 20417 3663 20451
rect 3605 20411 3663 20417
rect 1673 20383 1731 20389
rect 1673 20349 1685 20383
rect 1719 20349 1731 20383
rect 1673 20343 1731 20349
rect 1949 20383 2007 20389
rect 1949 20349 1961 20383
rect 1995 20380 2007 20383
rect 2130 20380 2136 20392
rect 1995 20352 2136 20380
rect 1995 20349 2007 20352
rect 1949 20343 2007 20349
rect 106 20204 112 20256
rect 164 20244 170 20256
rect 1489 20247 1547 20253
rect 1489 20244 1501 20247
rect 164 20216 1501 20244
rect 164 20204 170 20216
rect 1489 20213 1501 20216
rect 1535 20213 1547 20247
rect 1688 20244 1716 20343
rect 2130 20340 2136 20352
rect 2188 20340 2194 20392
rect 3053 20383 3111 20389
rect 3053 20349 3065 20383
rect 3099 20349 3111 20383
rect 3510 20380 3516 20392
rect 3471 20352 3516 20380
rect 3053 20343 3111 20349
rect 2406 20244 2412 20256
rect 1688 20216 2412 20244
rect 1489 20207 1547 20213
rect 2406 20204 2412 20216
rect 2464 20204 2470 20256
rect 2498 20204 2504 20256
rect 2556 20244 2562 20256
rect 2777 20247 2835 20253
rect 2777 20244 2789 20247
rect 2556 20216 2789 20244
rect 2556 20204 2562 20216
rect 2777 20213 2789 20216
rect 2823 20244 2835 20247
rect 3068 20244 3096 20343
rect 3510 20340 3516 20352
rect 3568 20340 3574 20392
rect 4522 20380 4528 20392
rect 4435 20352 4528 20380
rect 4522 20340 4528 20352
rect 4580 20380 4586 20392
rect 4617 20383 4675 20389
rect 4617 20380 4629 20383
rect 4580 20352 4629 20380
rect 4580 20340 4586 20352
rect 4617 20349 4629 20352
rect 4663 20349 4675 20383
rect 4617 20343 4675 20349
rect 5169 20383 5227 20389
rect 5169 20349 5181 20383
rect 5215 20380 5227 20383
rect 5350 20380 5356 20392
rect 5215 20352 5356 20380
rect 5215 20349 5227 20352
rect 5169 20343 5227 20349
rect 5350 20340 5356 20352
rect 5408 20380 5414 20392
rect 7006 20380 7012 20392
rect 5408 20352 7012 20380
rect 5408 20340 5414 20352
rect 7006 20340 7012 20352
rect 7064 20340 7070 20392
rect 4062 20244 4068 20256
rect 2823 20216 3096 20244
rect 4023 20216 4068 20244
rect 2823 20213 2835 20216
rect 2777 20207 2835 20213
rect 4062 20204 4068 20216
rect 4120 20204 4126 20256
rect 4706 20244 4712 20256
rect 4667 20216 4712 20244
rect 4706 20204 4712 20216
rect 4764 20204 4770 20256
rect 1104 20154 22816 20176
rect 1104 20102 8982 20154
rect 9034 20102 9046 20154
rect 9098 20102 9110 20154
rect 9162 20102 9174 20154
rect 9226 20102 16982 20154
rect 17034 20102 17046 20154
rect 17098 20102 17110 20154
rect 17162 20102 17174 20154
rect 17226 20102 22816 20154
rect 1104 20080 22816 20102
rect 382 20000 388 20052
rect 440 20040 446 20052
rect 1581 20043 1639 20049
rect 1581 20040 1593 20043
rect 440 20012 1593 20040
rect 440 20000 446 20012
rect 1581 20009 1593 20012
rect 1627 20009 1639 20043
rect 4614 20040 4620 20052
rect 4575 20012 4620 20040
rect 1581 20003 1639 20009
rect 4614 20000 4620 20012
rect 4672 20000 4678 20052
rect 6273 20043 6331 20049
rect 6273 20040 6285 20043
rect 5460 20012 6285 20040
rect 4338 19972 4344 19984
rect 4251 19944 4344 19972
rect 4338 19932 4344 19944
rect 4396 19972 4402 19984
rect 5350 19972 5356 19984
rect 4396 19944 5356 19972
rect 4396 19932 4402 19944
rect 5350 19932 5356 19944
rect 5408 19932 5414 19984
rect 1670 19904 1676 19916
rect 1631 19876 1676 19904
rect 1670 19864 1676 19876
rect 1728 19864 1734 19916
rect 2130 19913 2136 19916
rect 2087 19907 2136 19913
rect 2087 19873 2099 19907
rect 2133 19873 2136 19907
rect 2087 19867 2136 19873
rect 2130 19864 2136 19867
rect 2188 19904 2194 19916
rect 4522 19904 4528 19916
rect 2188 19876 4200 19904
rect 4483 19876 4528 19904
rect 2188 19864 2194 19876
rect 4172 19848 4200 19876
rect 4522 19864 4528 19876
rect 4580 19864 4586 19916
rect 5077 19907 5135 19913
rect 5077 19873 5089 19907
rect 5123 19904 5135 19907
rect 5460 19904 5488 20012
rect 6273 20009 6285 20012
rect 6319 20009 6331 20043
rect 6273 20003 6331 20009
rect 5123 19876 5488 19904
rect 6089 19907 6147 19913
rect 5123 19873 5135 19876
rect 5077 19867 5135 19873
rect 6089 19873 6101 19907
rect 6135 19904 6147 19907
rect 6270 19904 6276 19916
rect 6135 19876 6276 19904
rect 6135 19873 6147 19876
rect 6089 19867 6147 19873
rect 4154 19796 4160 19848
rect 4212 19836 4218 19848
rect 5092 19836 5120 19867
rect 6270 19864 6276 19876
rect 6328 19864 6334 19916
rect 4212 19808 5120 19836
rect 4212 19796 4218 19808
rect 2498 19660 2504 19712
rect 2556 19700 2562 19712
rect 3053 19703 3111 19709
rect 3053 19700 3065 19703
rect 2556 19672 3065 19700
rect 2556 19660 2562 19672
rect 3053 19669 3065 19672
rect 3099 19669 3111 19703
rect 3053 19663 3111 19669
rect 1104 19610 22816 19632
rect 1104 19558 4982 19610
rect 5034 19558 5046 19610
rect 5098 19558 5110 19610
rect 5162 19558 5174 19610
rect 5226 19558 12982 19610
rect 13034 19558 13046 19610
rect 13098 19558 13110 19610
rect 13162 19558 13174 19610
rect 13226 19558 20982 19610
rect 21034 19558 21046 19610
rect 21098 19558 21110 19610
rect 21162 19558 21174 19610
rect 21226 19558 22816 19610
rect 1104 19536 22816 19558
rect 2041 19499 2099 19505
rect 2041 19465 2053 19499
rect 2087 19496 2099 19499
rect 2130 19496 2136 19508
rect 2087 19468 2136 19496
rect 2087 19465 2099 19468
rect 2041 19459 2099 19465
rect 2130 19456 2136 19468
rect 2188 19456 2194 19508
rect 4249 19499 4307 19505
rect 4249 19465 4261 19499
rect 4295 19496 4307 19499
rect 4522 19496 4528 19508
rect 4295 19468 4528 19496
rect 4295 19465 4307 19468
rect 4249 19459 4307 19465
rect 4522 19456 4528 19468
rect 4580 19456 4586 19508
rect 7006 19496 7012 19508
rect 6967 19468 7012 19496
rect 7006 19456 7012 19468
rect 7064 19456 7070 19508
rect 198 19320 204 19372
rect 256 19360 262 19372
rect 3697 19363 3755 19369
rect 3697 19360 3709 19363
rect 256 19332 3709 19360
rect 256 19320 262 19332
rect 3697 19329 3709 19332
rect 3743 19329 3755 19363
rect 3697 19323 3755 19329
rect 1670 19292 1676 19304
rect 1583 19264 1676 19292
rect 1670 19252 1676 19264
rect 1728 19292 1734 19304
rect 2682 19292 2688 19304
rect 1728 19264 2688 19292
rect 1728 19252 1734 19264
rect 2682 19252 2688 19264
rect 2740 19252 2746 19304
rect 2869 19295 2927 19301
rect 2869 19261 2881 19295
rect 2915 19292 2927 19295
rect 3145 19295 3203 19301
rect 3145 19292 3157 19295
rect 2915 19264 3157 19292
rect 2915 19261 2927 19264
rect 2869 19255 2927 19261
rect 3145 19261 3157 19264
rect 3191 19261 3203 19295
rect 3602 19292 3608 19304
rect 3563 19264 3608 19292
rect 3145 19255 3203 19261
rect 3602 19252 3608 19264
rect 3660 19292 3666 19304
rect 4338 19292 4344 19304
rect 3660 19264 4344 19292
rect 3660 19252 3666 19264
rect 4338 19252 4344 19264
rect 4396 19252 4402 19304
rect 4522 19252 4528 19304
rect 4580 19292 4586 19304
rect 4798 19292 4804 19304
rect 4580 19264 4804 19292
rect 4580 19252 4586 19264
rect 4798 19252 4804 19264
rect 4856 19292 4862 19304
rect 4893 19295 4951 19301
rect 4893 19292 4905 19295
rect 4856 19264 4905 19292
rect 4856 19252 4862 19264
rect 4893 19261 4905 19264
rect 4939 19261 4951 19295
rect 4893 19255 4951 19261
rect 5445 19295 5503 19301
rect 5445 19261 5457 19295
rect 5491 19292 5503 19295
rect 6822 19292 6828 19304
rect 5491 19264 5948 19292
rect 6783 19264 6828 19292
rect 5491 19261 5503 19264
rect 5445 19255 5503 19261
rect 290 19184 296 19236
rect 348 19224 354 19236
rect 348 19196 4752 19224
rect 348 19184 354 19196
rect 1854 19116 1860 19168
rect 1912 19156 1918 19168
rect 2406 19156 2412 19168
rect 1912 19128 2412 19156
rect 1912 19116 1918 19128
rect 2406 19116 2412 19128
rect 2464 19156 2470 19168
rect 2869 19159 2927 19165
rect 2869 19156 2881 19159
rect 2464 19128 2881 19156
rect 2464 19116 2470 19128
rect 2869 19125 2881 19128
rect 2915 19156 2927 19159
rect 2961 19159 3019 19165
rect 2961 19156 2973 19159
rect 2915 19128 2973 19156
rect 2915 19125 2927 19128
rect 2869 19119 2927 19125
rect 2961 19125 2973 19128
rect 3007 19125 3019 19159
rect 4724 19156 4752 19196
rect 5920 19168 5948 19264
rect 6822 19252 6828 19264
rect 6880 19292 6886 19304
rect 7285 19295 7343 19301
rect 7285 19292 7297 19295
rect 6880 19264 7297 19292
rect 6880 19252 6886 19264
rect 7285 19261 7297 19264
rect 7331 19261 7343 19295
rect 7285 19255 7343 19261
rect 4985 19159 5043 19165
rect 4985 19156 4997 19159
rect 4724 19128 4997 19156
rect 2961 19119 3019 19125
rect 4985 19125 4997 19128
rect 5031 19125 5043 19159
rect 5902 19156 5908 19168
rect 5863 19128 5908 19156
rect 4985 19119 5043 19125
rect 5902 19116 5908 19128
rect 5960 19116 5966 19168
rect 6270 19156 6276 19168
rect 6231 19128 6276 19156
rect 6270 19116 6276 19128
rect 6328 19116 6334 19168
rect 1104 19066 22816 19088
rect 1104 19014 8982 19066
rect 9034 19014 9046 19066
rect 9098 19014 9110 19066
rect 9162 19014 9174 19066
rect 9226 19014 16982 19066
rect 17034 19014 17046 19066
rect 17098 19014 17110 19066
rect 17162 19014 17174 19066
rect 17226 19014 22816 19066
rect 1104 18992 22816 19014
rect 1762 18952 1768 18964
rect 1723 18924 1768 18952
rect 1762 18912 1768 18924
rect 1820 18912 1826 18964
rect 3237 18955 3295 18961
rect 3237 18921 3249 18955
rect 3283 18952 3295 18955
rect 3602 18952 3608 18964
rect 3283 18924 3608 18952
rect 3283 18921 3295 18924
rect 3237 18915 3295 18921
rect 3602 18912 3608 18924
rect 3660 18912 3666 18964
rect 3881 18955 3939 18961
rect 3881 18921 3893 18955
rect 3927 18952 3939 18955
rect 4154 18952 4160 18964
rect 3927 18924 4160 18952
rect 3927 18921 3939 18924
rect 3881 18915 3939 18921
rect 4154 18912 4160 18924
rect 4212 18912 4218 18964
rect 4246 18912 4252 18964
rect 4304 18952 4310 18964
rect 4341 18955 4399 18961
rect 4341 18952 4353 18955
rect 4304 18924 4353 18952
rect 4304 18912 4310 18924
rect 4341 18921 4353 18924
rect 4387 18921 4399 18955
rect 5813 18955 5871 18961
rect 5813 18952 5825 18955
rect 4341 18915 4399 18921
rect 4816 18924 5825 18952
rect 1949 18819 2007 18825
rect 1949 18785 1961 18819
rect 1995 18785 2007 18819
rect 2222 18816 2228 18828
rect 2135 18788 2228 18816
rect 1949 18779 2007 18785
rect 1964 18748 1992 18779
rect 2222 18776 2228 18788
rect 2280 18816 2286 18828
rect 2685 18819 2743 18825
rect 2685 18816 2697 18819
rect 2280 18788 2697 18816
rect 2280 18776 2286 18788
rect 2685 18785 2697 18788
rect 2731 18785 2743 18819
rect 4062 18816 4068 18828
rect 4023 18788 4068 18816
rect 2685 18779 2743 18785
rect 4062 18776 4068 18788
rect 4120 18776 4126 18828
rect 4614 18816 4620 18828
rect 4527 18788 4620 18816
rect 4614 18776 4620 18788
rect 4672 18816 4678 18828
rect 4816 18816 4844 18924
rect 5813 18921 5825 18924
rect 5859 18921 5871 18955
rect 5813 18915 5871 18921
rect 5626 18816 5632 18828
rect 4672 18788 4844 18816
rect 5587 18788 5632 18816
rect 4672 18776 4678 18788
rect 5626 18776 5632 18788
rect 5684 18776 5690 18828
rect 2406 18748 2412 18760
rect 1964 18720 2412 18748
rect 2406 18708 2412 18720
rect 2464 18708 2470 18760
rect 5261 18615 5319 18621
rect 5261 18581 5273 18615
rect 5307 18612 5319 18615
rect 5442 18612 5448 18624
rect 5307 18584 5448 18612
rect 5307 18581 5319 18584
rect 5261 18575 5319 18581
rect 5442 18572 5448 18584
rect 5500 18572 5506 18624
rect 6178 18612 6184 18624
rect 6139 18584 6184 18612
rect 6178 18572 6184 18584
rect 6236 18572 6242 18624
rect 1104 18522 22816 18544
rect 1104 18470 4982 18522
rect 5034 18470 5046 18522
rect 5098 18470 5110 18522
rect 5162 18470 5174 18522
rect 5226 18470 12982 18522
rect 13034 18470 13046 18522
rect 13098 18470 13110 18522
rect 13162 18470 13174 18522
rect 13226 18470 20982 18522
rect 21034 18470 21046 18522
rect 21098 18470 21110 18522
rect 21162 18470 21174 18522
rect 21226 18470 22816 18522
rect 1104 18448 22816 18470
rect 5442 18408 5448 18420
rect 5403 18380 5448 18408
rect 5442 18368 5448 18380
rect 5500 18368 5506 18420
rect 5813 18411 5871 18417
rect 5813 18377 5825 18411
rect 5859 18408 5871 18411
rect 6270 18408 6276 18420
rect 5859 18380 6276 18408
rect 5859 18377 5871 18380
rect 5813 18371 5871 18377
rect 6270 18368 6276 18380
rect 6328 18368 6334 18420
rect 106 18232 112 18284
rect 164 18272 170 18284
rect 2317 18275 2375 18281
rect 2317 18272 2329 18275
rect 164 18244 2329 18272
rect 164 18232 170 18244
rect 2317 18241 2329 18244
rect 2363 18241 2375 18275
rect 2317 18235 2375 18241
rect 2682 18232 2688 18284
rect 2740 18272 2746 18284
rect 4062 18272 4068 18284
rect 2740 18244 4068 18272
rect 2740 18232 2746 18244
rect 4062 18232 4068 18244
rect 4120 18272 4126 18284
rect 4341 18275 4399 18281
rect 4341 18272 4353 18275
rect 4120 18244 4353 18272
rect 4120 18232 4126 18244
rect 4341 18241 4353 18244
rect 4387 18241 4399 18275
rect 4341 18235 4399 18241
rect 5077 18275 5135 18281
rect 5077 18241 5089 18275
rect 5123 18272 5135 18275
rect 5534 18272 5540 18284
rect 5123 18244 5540 18272
rect 5123 18241 5135 18244
rect 5077 18235 5135 18241
rect 5534 18232 5540 18244
rect 5592 18232 5598 18284
rect 1765 18207 1823 18213
rect 1765 18173 1777 18207
rect 1811 18173 1823 18207
rect 2222 18204 2228 18216
rect 2183 18176 2228 18204
rect 1765 18167 1823 18173
rect 1780 18080 1808 18167
rect 2222 18164 2228 18176
rect 2280 18164 2286 18216
rect 3329 18207 3387 18213
rect 3329 18204 3341 18207
rect 3252 18176 3341 18204
rect 3252 18136 3280 18176
rect 3329 18173 3341 18176
rect 3375 18173 3387 18207
rect 3786 18204 3792 18216
rect 3747 18176 3792 18204
rect 3329 18167 3387 18173
rect 3786 18164 3792 18176
rect 3844 18204 3850 18216
rect 4614 18204 4620 18216
rect 3844 18176 4620 18204
rect 3844 18164 3850 18176
rect 4614 18164 4620 18176
rect 4672 18164 4678 18216
rect 5316 18207 5374 18213
rect 5316 18173 5328 18207
rect 5362 18204 5374 18207
rect 6178 18204 6184 18216
rect 5362 18176 6184 18204
rect 5362 18173 5374 18176
rect 5316 18167 5374 18173
rect 6178 18164 6184 18176
rect 6236 18164 6242 18216
rect 6825 18207 6883 18213
rect 6825 18173 6837 18207
rect 6871 18204 6883 18207
rect 6914 18204 6920 18216
rect 6871 18176 6920 18204
rect 6871 18173 6883 18176
rect 6825 18167 6883 18173
rect 6914 18164 6920 18176
rect 6972 18204 6978 18216
rect 7285 18207 7343 18213
rect 7285 18204 7297 18207
rect 6972 18176 7297 18204
rect 6972 18164 6978 18176
rect 7285 18173 7297 18176
rect 7331 18173 7343 18207
rect 7285 18167 7343 18173
rect 4798 18136 4804 18148
rect 3252 18108 4804 18136
rect 3252 18080 3280 18108
rect 4798 18096 4804 18108
rect 4856 18096 4862 18148
rect 5166 18136 5172 18148
rect 5127 18108 5172 18136
rect 5166 18096 5172 18108
rect 5224 18136 5230 18148
rect 6273 18139 6331 18145
rect 6273 18136 6285 18139
rect 5224 18108 6285 18136
rect 5224 18096 5230 18108
rect 6273 18105 6285 18108
rect 6319 18105 6331 18139
rect 6273 18099 6331 18105
rect 1673 18071 1731 18077
rect 1673 18037 1685 18071
rect 1719 18068 1731 18071
rect 1762 18068 1768 18080
rect 1719 18040 1768 18068
rect 1719 18037 1731 18040
rect 1673 18031 1731 18037
rect 1762 18028 1768 18040
rect 1820 18028 1826 18080
rect 2406 18028 2412 18080
rect 2464 18068 2470 18080
rect 2777 18071 2835 18077
rect 2777 18068 2789 18071
rect 2464 18040 2789 18068
rect 2464 18028 2470 18040
rect 2777 18037 2789 18040
rect 2823 18037 2835 18071
rect 3234 18068 3240 18080
rect 3195 18040 3240 18068
rect 2777 18031 2835 18037
rect 3234 18028 3240 18040
rect 3292 18028 3298 18080
rect 3418 18068 3424 18080
rect 3379 18040 3424 18068
rect 3418 18028 3424 18040
rect 3476 18028 3482 18080
rect 6546 18068 6552 18080
rect 6507 18040 6552 18068
rect 6546 18028 6552 18040
rect 6604 18028 6610 18080
rect 7006 18068 7012 18080
rect 6967 18040 7012 18068
rect 7006 18028 7012 18040
rect 7064 18028 7070 18080
rect 1104 17978 22816 18000
rect 1104 17926 8982 17978
rect 9034 17926 9046 17978
rect 9098 17926 9110 17978
rect 9162 17926 9174 17978
rect 9226 17926 16982 17978
rect 17034 17926 17046 17978
rect 17098 17926 17110 17978
rect 17162 17926 17174 17978
rect 17226 17926 22816 17978
rect 1104 17904 22816 17926
rect 14 17824 20 17876
rect 72 17864 78 17876
rect 1489 17867 1547 17873
rect 1489 17864 1501 17867
rect 72 17836 1501 17864
rect 72 17824 78 17836
rect 1489 17833 1501 17836
rect 1535 17833 1547 17867
rect 1489 17827 1547 17833
rect 2222 17824 2228 17876
rect 2280 17864 2286 17876
rect 2409 17867 2467 17873
rect 2409 17864 2421 17867
rect 2280 17836 2421 17864
rect 2280 17824 2286 17836
rect 2409 17833 2421 17836
rect 2455 17864 2467 17867
rect 3329 17867 3387 17873
rect 3329 17864 3341 17867
rect 2455 17836 3341 17864
rect 2455 17833 2467 17836
rect 2409 17827 2467 17833
rect 3329 17833 3341 17836
rect 3375 17864 3387 17867
rect 3786 17864 3792 17876
rect 3375 17836 3792 17864
rect 3375 17833 3387 17836
rect 3329 17827 3387 17833
rect 3786 17824 3792 17836
rect 3844 17824 3850 17876
rect 6178 17864 6184 17876
rect 6091 17836 6184 17864
rect 6178 17824 6184 17836
rect 6236 17864 6242 17876
rect 6914 17864 6920 17876
rect 6236 17836 6920 17864
rect 6236 17824 6242 17836
rect 6914 17824 6920 17836
rect 6972 17824 6978 17876
rect 5626 17756 5632 17808
rect 5684 17796 5690 17808
rect 5813 17799 5871 17805
rect 5813 17796 5825 17799
rect 5684 17768 5825 17796
rect 5684 17756 5690 17768
rect 5813 17765 5825 17768
rect 5859 17796 5871 17799
rect 6546 17796 6552 17808
rect 5859 17768 6552 17796
rect 5859 17765 5871 17768
rect 5813 17759 5871 17765
rect 6546 17756 6552 17768
rect 6604 17756 6610 17808
rect 1673 17731 1731 17737
rect 1673 17697 1685 17731
rect 1719 17697 1731 17731
rect 1946 17728 1952 17740
rect 1907 17700 1952 17728
rect 1673 17691 1731 17697
rect 1688 17660 1716 17691
rect 1946 17688 1952 17700
rect 2004 17728 2010 17740
rect 2777 17731 2835 17737
rect 2777 17728 2789 17731
rect 2004 17700 2789 17728
rect 2004 17688 2010 17700
rect 2777 17697 2789 17700
rect 2823 17697 2835 17731
rect 2777 17691 2835 17697
rect 4065 17731 4123 17737
rect 4065 17697 4077 17731
rect 4111 17728 4123 17731
rect 4430 17728 4436 17740
rect 4111 17700 4436 17728
rect 4111 17697 4123 17700
rect 4065 17691 4123 17697
rect 4430 17688 4436 17700
rect 4488 17688 4494 17740
rect 5077 17731 5135 17737
rect 5077 17728 5089 17731
rect 4908 17700 5089 17728
rect 2406 17660 2412 17672
rect 1688 17632 2412 17660
rect 2406 17620 2412 17632
rect 2464 17620 2470 17672
rect 4246 17524 4252 17536
rect 4207 17496 4252 17524
rect 4246 17484 4252 17496
rect 4304 17484 4310 17536
rect 4522 17524 4528 17536
rect 4483 17496 4528 17524
rect 4522 17484 4528 17496
rect 4580 17524 4586 17536
rect 4908 17533 4936 17700
rect 5077 17697 5089 17700
rect 5123 17728 5135 17731
rect 5166 17728 5172 17740
rect 5123 17700 5172 17728
rect 5123 17697 5135 17700
rect 5077 17691 5135 17697
rect 5166 17688 5172 17700
rect 5224 17688 5230 17740
rect 6638 17688 6644 17740
rect 6696 17728 6702 17740
rect 6733 17731 6791 17737
rect 6733 17728 6745 17731
rect 6696 17700 6745 17728
rect 6696 17688 6702 17700
rect 6733 17697 6745 17700
rect 6779 17697 6791 17731
rect 6733 17691 6791 17697
rect 5445 17663 5503 17669
rect 5445 17629 5457 17663
rect 5491 17660 5503 17663
rect 5626 17660 5632 17672
rect 5491 17632 5632 17660
rect 5491 17629 5503 17632
rect 5445 17623 5503 17629
rect 5626 17620 5632 17632
rect 5684 17620 5690 17672
rect 5718 17620 5724 17672
rect 5776 17660 5782 17672
rect 6549 17663 6607 17669
rect 6549 17660 6561 17663
rect 5776 17632 6561 17660
rect 5776 17620 5782 17632
rect 6549 17629 6561 17632
rect 6595 17660 6607 17663
rect 7006 17660 7012 17672
rect 6595 17632 7012 17660
rect 6595 17629 6607 17632
rect 6549 17623 6607 17629
rect 7006 17620 7012 17632
rect 7064 17620 7070 17672
rect 5242 17595 5300 17601
rect 5242 17561 5254 17595
rect 5288 17592 5300 17595
rect 6178 17592 6184 17604
rect 5288 17564 6184 17592
rect 5288 17561 5300 17564
rect 5242 17555 5300 17561
rect 6178 17552 6184 17564
rect 6236 17552 6242 17604
rect 4893 17527 4951 17533
rect 4893 17524 4905 17527
rect 4580 17496 4905 17524
rect 4580 17484 4586 17496
rect 4893 17493 4905 17496
rect 4939 17493 4951 17527
rect 4893 17487 4951 17493
rect 5353 17527 5411 17533
rect 5353 17493 5365 17527
rect 5399 17524 5411 17527
rect 5442 17524 5448 17536
rect 5399 17496 5448 17524
rect 5399 17493 5411 17496
rect 5353 17487 5411 17493
rect 5442 17484 5448 17496
rect 5500 17524 5506 17536
rect 6086 17524 6092 17536
rect 5500 17496 6092 17524
rect 5500 17484 5506 17496
rect 6086 17484 6092 17496
rect 6144 17484 6150 17536
rect 14 17416 20 17468
rect 72 17456 78 17468
rect 72 17428 117 17456
rect 1104 17434 22816 17456
rect 72 17416 78 17428
rect 1104 17382 4982 17434
rect 5034 17382 5046 17434
rect 5098 17382 5110 17434
rect 5162 17382 5174 17434
rect 5226 17382 12982 17434
rect 13034 17382 13046 17434
rect 13098 17382 13110 17434
rect 13162 17382 13174 17434
rect 13226 17382 20982 17434
rect 21034 17382 21046 17434
rect 21098 17382 21110 17434
rect 21162 17382 21174 17434
rect 21226 17382 22816 17434
rect 1104 17360 22816 17382
rect 5334 17323 5392 17329
rect 5334 17289 5346 17323
rect 5380 17320 5392 17323
rect 5718 17320 5724 17332
rect 5380 17292 5724 17320
rect 5380 17289 5392 17292
rect 5334 17283 5392 17289
rect 5718 17280 5724 17292
rect 5776 17280 5782 17332
rect 5813 17323 5871 17329
rect 5813 17289 5825 17323
rect 5859 17320 5871 17323
rect 6822 17320 6828 17332
rect 5859 17292 6828 17320
rect 5859 17289 5871 17292
rect 5813 17283 5871 17289
rect 6822 17280 6828 17292
rect 6880 17280 6886 17332
rect 5445 17255 5503 17261
rect 5445 17221 5457 17255
rect 5491 17221 5503 17255
rect 5445 17215 5503 17221
rect 14 17144 20 17196
rect 72 17184 78 17196
rect 3605 17187 3663 17193
rect 3605 17184 3617 17187
rect 72 17156 3617 17184
rect 72 17144 78 17156
rect 3605 17153 3617 17156
rect 3651 17153 3663 17187
rect 3605 17147 3663 17153
rect 5350 17144 5356 17196
rect 5408 17184 5414 17196
rect 5460 17184 5488 17215
rect 6086 17212 6092 17264
rect 6144 17252 6150 17264
rect 6181 17255 6239 17261
rect 6181 17252 6193 17255
rect 6144 17224 6193 17252
rect 6144 17212 6150 17224
rect 6181 17221 6193 17224
rect 6227 17252 6239 17255
rect 7009 17255 7067 17261
rect 7009 17252 7021 17255
rect 6227 17224 7021 17252
rect 6227 17221 6239 17224
rect 6181 17215 6239 17221
rect 7009 17221 7021 17224
rect 7055 17221 7067 17255
rect 7009 17215 7067 17221
rect 5408 17156 5488 17184
rect 5537 17187 5595 17193
rect 5408 17144 5414 17156
rect 5537 17153 5549 17187
rect 5583 17184 5595 17187
rect 5626 17184 5632 17196
rect 5583 17156 5632 17184
rect 5583 17153 5595 17156
rect 5537 17147 5595 17153
rect 1673 17119 1731 17125
rect 1673 17085 1685 17119
rect 1719 17116 1731 17119
rect 1762 17116 1768 17128
rect 1719 17088 1768 17116
rect 1719 17085 1731 17088
rect 1673 17079 1731 17085
rect 1762 17076 1768 17088
rect 1820 17076 1826 17128
rect 1946 17116 1952 17128
rect 1907 17088 1952 17116
rect 1946 17076 1952 17088
rect 2004 17076 2010 17128
rect 3329 17119 3387 17125
rect 3329 17085 3341 17119
rect 3375 17085 3387 17119
rect 3510 17116 3516 17128
rect 3471 17088 3516 17116
rect 3329 17079 3387 17085
rect 2961 17051 3019 17057
rect 2961 17017 2973 17051
rect 3007 17048 3019 17051
rect 3234 17048 3240 17060
rect 3007 17020 3240 17048
rect 3007 17017 3019 17020
rect 2961 17011 3019 17017
rect 3234 17008 3240 17020
rect 3292 17048 3298 17060
rect 3344 17048 3372 17079
rect 3510 17076 3516 17088
rect 3568 17076 3574 17128
rect 5552 17116 5580 17147
rect 5626 17144 5632 17156
rect 5684 17184 5690 17196
rect 6914 17184 6920 17196
rect 5684 17156 6920 17184
rect 5684 17144 5690 17156
rect 6914 17144 6920 17156
rect 6972 17144 6978 17196
rect 4632 17088 5580 17116
rect 6825 17119 6883 17125
rect 3694 17048 3700 17060
rect 3292 17020 3700 17048
rect 3292 17008 3298 17020
rect 3694 17008 3700 17020
rect 3752 17008 3758 17060
rect 106 16940 112 16992
rect 164 16980 170 16992
rect 1489 16983 1547 16989
rect 1489 16980 1501 16983
rect 164 16952 1501 16980
rect 164 16940 170 16952
rect 1489 16949 1501 16952
rect 1535 16949 1547 16983
rect 2406 16980 2412 16992
rect 2367 16952 2412 16980
rect 1489 16943 1547 16949
rect 2406 16940 2412 16952
rect 2464 16940 2470 16992
rect 4338 16980 4344 16992
rect 4299 16952 4344 16980
rect 4338 16940 4344 16952
rect 4396 16980 4402 16992
rect 4632 16989 4660 17088
rect 6825 17085 6837 17119
rect 6871 17116 6883 17119
rect 7374 17116 7380 17128
rect 6871 17088 7380 17116
rect 6871 17085 6883 17088
rect 6825 17079 6883 17085
rect 7374 17076 7380 17088
rect 7432 17076 7438 17128
rect 5166 17048 5172 17060
rect 5127 17020 5172 17048
rect 5166 17008 5172 17020
rect 5224 17008 5230 17060
rect 4617 16983 4675 16989
rect 4617 16980 4629 16983
rect 4396 16952 4629 16980
rect 4396 16940 4402 16952
rect 4617 16949 4629 16952
rect 4663 16949 4675 16983
rect 4617 16943 4675 16949
rect 5077 16983 5135 16989
rect 5077 16949 5089 16983
rect 5123 16980 5135 16983
rect 5350 16980 5356 16992
rect 5123 16952 5356 16980
rect 5123 16949 5135 16952
rect 5077 16943 5135 16949
rect 5350 16940 5356 16952
rect 5408 16940 5414 16992
rect 6638 16980 6644 16992
rect 6599 16952 6644 16980
rect 6638 16940 6644 16952
rect 6696 16940 6702 16992
rect 7374 16980 7380 16992
rect 7335 16952 7380 16980
rect 7374 16940 7380 16952
rect 7432 16940 7438 16992
rect 1104 16890 22816 16912
rect 1104 16838 8982 16890
rect 9034 16838 9046 16890
rect 9098 16838 9110 16890
rect 9162 16838 9174 16890
rect 9226 16838 16982 16890
rect 17034 16838 17046 16890
rect 17098 16838 17110 16890
rect 17162 16838 17174 16890
rect 17226 16838 22816 16890
rect 1104 16816 22816 16838
rect 17 16779 75 16785
rect 17 16745 29 16779
rect 63 16776 75 16779
rect 2133 16779 2191 16785
rect 2133 16776 2145 16779
rect 63 16748 2145 16776
rect 63 16745 75 16748
rect 17 16739 75 16745
rect 2133 16745 2145 16748
rect 2179 16745 2191 16779
rect 4249 16779 4307 16785
rect 4249 16776 4261 16779
rect 2133 16739 2191 16745
rect 4126 16748 4261 16776
rect 1946 16668 1952 16720
rect 2004 16708 2010 16720
rect 2866 16708 2872 16720
rect 2004 16680 2872 16708
rect 2004 16668 2010 16680
rect 2516 16649 2544 16680
rect 2866 16668 2872 16680
rect 2924 16708 2930 16720
rect 3053 16711 3111 16717
rect 3053 16708 3065 16711
rect 2924 16680 3065 16708
rect 2924 16668 2930 16680
rect 3053 16677 3065 16680
rect 3099 16708 3111 16711
rect 3421 16711 3479 16717
rect 3421 16708 3433 16711
rect 3099 16680 3433 16708
rect 3099 16677 3111 16680
rect 3053 16671 3111 16677
rect 3421 16677 3433 16680
rect 3467 16708 3479 16711
rect 3510 16708 3516 16720
rect 3467 16680 3516 16708
rect 3467 16677 3479 16680
rect 3421 16671 3479 16677
rect 3510 16668 3516 16680
rect 3568 16708 3574 16720
rect 4126 16708 4154 16748
rect 4249 16745 4261 16748
rect 4295 16745 4307 16779
rect 6914 16776 6920 16788
rect 6875 16748 6920 16776
rect 4249 16739 4307 16745
rect 6914 16736 6920 16748
rect 6972 16736 6978 16788
rect 3568 16680 4154 16708
rect 4801 16711 4859 16717
rect 3568 16668 3574 16680
rect 4801 16677 4813 16711
rect 4847 16708 4859 16711
rect 5626 16708 5632 16720
rect 4847 16680 5632 16708
rect 4847 16677 4859 16680
rect 4801 16671 4859 16677
rect 5626 16668 5632 16680
rect 5684 16668 5690 16720
rect 5902 16708 5908 16720
rect 5863 16680 5908 16708
rect 5902 16668 5908 16680
rect 5960 16668 5966 16720
rect 2317 16643 2375 16649
rect 2317 16609 2329 16643
rect 2363 16609 2375 16643
rect 2317 16603 2375 16609
rect 2501 16643 2559 16649
rect 2501 16609 2513 16643
rect 2547 16609 2559 16643
rect 2501 16603 2559 16609
rect 2332 16572 2360 16603
rect 3970 16600 3976 16652
rect 4028 16640 4034 16652
rect 4065 16643 4123 16649
rect 4065 16640 4077 16643
rect 4028 16612 4077 16640
rect 4028 16600 4034 16612
rect 4065 16609 4077 16612
rect 4111 16609 4123 16643
rect 4065 16603 4123 16609
rect 4522 16600 4528 16652
rect 4580 16640 4586 16652
rect 5166 16640 5172 16652
rect 4580 16612 5172 16640
rect 4580 16600 4586 16612
rect 5166 16600 5172 16612
rect 5224 16640 5230 16652
rect 6181 16643 6239 16649
rect 6181 16640 6193 16643
rect 5224 16612 6193 16640
rect 5224 16600 5230 16612
rect 6181 16609 6193 16612
rect 6227 16640 6239 16643
rect 6362 16640 6368 16652
rect 6227 16612 6368 16640
rect 6227 16609 6239 16612
rect 6181 16603 6239 16609
rect 6362 16600 6368 16612
rect 6420 16600 6426 16652
rect 6730 16640 6736 16652
rect 6691 16612 6736 16640
rect 6730 16600 6736 16612
rect 6788 16600 6794 16652
rect 2682 16572 2688 16584
rect 2332 16544 2688 16572
rect 2682 16532 2688 16544
rect 2740 16532 2746 16584
rect 3881 16575 3939 16581
rect 3881 16541 3893 16575
rect 3927 16572 3939 16575
rect 4430 16572 4436 16584
rect 3927 16544 4436 16572
rect 3927 16541 3939 16544
rect 3881 16535 3939 16541
rect 4430 16532 4436 16544
rect 4488 16532 4494 16584
rect 5534 16572 5540 16584
rect 5495 16544 5540 16572
rect 5534 16532 5540 16544
rect 5592 16532 5598 16584
rect 5718 16504 5724 16516
rect 5331 16476 5724 16504
rect 1673 16439 1731 16445
rect 1673 16405 1685 16439
rect 1719 16436 1731 16439
rect 1762 16436 1768 16448
rect 1719 16408 1768 16436
rect 1719 16405 1731 16408
rect 1673 16399 1731 16405
rect 1762 16396 1768 16408
rect 1820 16396 1826 16448
rect 5331 16445 5359 16476
rect 5718 16464 5724 16476
rect 5776 16464 5782 16516
rect 5316 16439 5374 16445
rect 5316 16405 5328 16439
rect 5362 16405 5374 16439
rect 5442 16436 5448 16448
rect 5403 16408 5448 16436
rect 5316 16399 5374 16405
rect 5442 16396 5448 16408
rect 5500 16396 5506 16448
rect 1104 16346 22816 16368
rect 1104 16294 4982 16346
rect 5034 16294 5046 16346
rect 5098 16294 5110 16346
rect 5162 16294 5174 16346
rect 5226 16294 12982 16346
rect 13034 16294 13046 16346
rect 13098 16294 13110 16346
rect 13162 16294 13174 16346
rect 13226 16294 20982 16346
rect 21034 16294 21046 16346
rect 21098 16294 21110 16346
rect 21162 16294 21174 16346
rect 21226 16294 22816 16346
rect 1104 16272 22816 16294
rect 4430 16192 4436 16244
rect 4488 16232 4494 16244
rect 5169 16235 5227 16241
rect 5169 16232 5181 16235
rect 4488 16204 5181 16232
rect 4488 16192 4494 16204
rect 5169 16201 5181 16204
rect 5215 16201 5227 16235
rect 5169 16195 5227 16201
rect 5534 16192 5540 16244
rect 5592 16232 5598 16244
rect 5721 16235 5779 16241
rect 5721 16232 5733 16235
rect 5592 16204 5733 16232
rect 5592 16192 5598 16204
rect 5721 16201 5733 16204
rect 5767 16201 5779 16235
rect 5721 16195 5779 16201
rect 6362 16192 6368 16244
rect 6420 16232 6426 16244
rect 6457 16235 6515 16241
rect 6457 16232 6469 16235
rect 6420 16204 6469 16232
rect 6420 16192 6426 16204
rect 6457 16201 6469 16204
rect 6503 16201 6515 16235
rect 7742 16232 7748 16244
rect 7703 16204 7748 16232
rect 6457 16195 6515 16201
rect 7742 16192 7748 16204
rect 7800 16192 7806 16244
rect 4617 16167 4675 16173
rect 4617 16133 4629 16167
rect 4663 16164 4675 16167
rect 4985 16167 5043 16173
rect 4985 16164 4997 16167
rect 4663 16136 4997 16164
rect 4663 16133 4675 16136
rect 4617 16127 4675 16133
rect 4985 16133 4997 16136
rect 5031 16164 5043 16167
rect 5350 16164 5356 16176
rect 5031 16136 5356 16164
rect 5031 16133 5043 16136
rect 4985 16127 5043 16133
rect 5350 16124 5356 16136
rect 5408 16124 5414 16176
rect 5626 16124 5632 16176
rect 5684 16164 5690 16176
rect 7009 16167 7067 16173
rect 7009 16164 7021 16167
rect 5684 16136 7021 16164
rect 5684 16124 5690 16136
rect 7009 16133 7021 16136
rect 7055 16133 7067 16167
rect 7009 16127 7067 16133
rect 2406 16096 2412 16108
rect 1596 16068 2412 16096
rect 1596 16040 1624 16068
rect 2406 16056 2412 16068
rect 2464 16096 2470 16108
rect 2961 16099 3019 16105
rect 2961 16096 2973 16099
rect 2464 16068 2973 16096
rect 2464 16056 2470 16068
rect 2961 16065 2973 16068
rect 3007 16065 3019 16099
rect 2961 16059 3019 16065
rect 4249 16099 4307 16105
rect 4249 16065 4261 16099
rect 4295 16096 4307 16099
rect 4338 16096 4344 16108
rect 4295 16068 4344 16096
rect 4295 16065 4307 16068
rect 4249 16059 4307 16065
rect 1578 16028 1584 16040
rect 1539 16000 1584 16028
rect 1578 15988 1584 16000
rect 1636 15988 1642 16040
rect 2130 16028 2136 16040
rect 2091 16000 2136 16028
rect 2130 15988 2136 16000
rect 2188 15988 2194 16040
rect 2976 16028 3004 16059
rect 4338 16056 4344 16068
rect 4396 16096 4402 16108
rect 5077 16099 5135 16105
rect 5077 16096 5089 16099
rect 4396 16068 5089 16096
rect 4396 16056 4402 16068
rect 5077 16065 5089 16068
rect 5123 16065 5135 16099
rect 5368 16096 5396 16124
rect 6089 16099 6147 16105
rect 6089 16096 6101 16099
rect 5368 16068 6101 16096
rect 5077 16059 5135 16065
rect 6089 16065 6101 16068
rect 6135 16065 6147 16099
rect 6089 16059 6147 16065
rect 3145 16031 3203 16037
rect 3145 16028 3157 16031
rect 2976 16000 3157 16028
rect 3145 15997 3157 16000
rect 3191 15997 3203 16031
rect 3145 15991 3203 15997
rect 3697 16031 3755 16037
rect 3697 15997 3709 16031
rect 3743 16028 3755 16031
rect 4062 16028 4068 16040
rect 3743 16000 4068 16028
rect 3743 15997 3755 16000
rect 3697 15991 3755 15997
rect 4062 15988 4068 16000
rect 4120 15988 4126 16040
rect 4853 16028 4859 16040
rect 4814 16000 4859 16028
rect 4853 15988 4859 16000
rect 4911 15988 4917 16040
rect 5092 16028 5120 16059
rect 6638 16056 6644 16108
rect 6696 16096 6702 16108
rect 7760 16096 7788 16192
rect 6696 16068 7788 16096
rect 6696 16056 6702 16068
rect 5442 16028 5448 16040
rect 5092 16000 5448 16028
rect 5442 15988 5448 16000
rect 5500 15988 5506 16040
rect 6840 16037 6868 16068
rect 6825 16031 6883 16037
rect 6825 15997 6837 16031
rect 6871 15997 6883 16031
rect 7834 16028 7840 16040
rect 7747 16000 7840 16028
rect 6825 15991 6883 15997
rect 7834 15988 7840 16000
rect 7892 16028 7898 16040
rect 8297 16031 8355 16037
rect 8297 16028 8309 16031
rect 7892 16000 8309 16028
rect 7892 15988 7898 16000
rect 8297 15997 8309 16000
rect 8343 15997 8355 16031
rect 8297 15991 8355 15997
rect 14 15920 20 15972
rect 72 15920 78 15972
rect 4522 15920 4528 15972
rect 4580 15960 4586 15972
rect 4709 15963 4767 15969
rect 4709 15960 4721 15963
rect 4580 15932 4721 15960
rect 4580 15920 4586 15932
rect 4709 15929 4721 15932
rect 4755 15929 4767 15963
rect 4709 15923 4767 15929
rect 6730 15920 6736 15972
rect 6788 15960 6794 15972
rect 7377 15963 7435 15969
rect 7377 15960 7389 15963
rect 6788 15932 7389 15960
rect 6788 15920 6794 15932
rect 7377 15929 7389 15932
rect 7423 15960 7435 15963
rect 7558 15960 7564 15972
rect 7423 15932 7564 15960
rect 7423 15929 7435 15932
rect 7377 15923 7435 15929
rect 7558 15920 7564 15932
rect 7616 15960 7622 15972
rect 9582 15960 9588 15972
rect 7616 15932 9588 15960
rect 7616 15920 7622 15932
rect 9582 15920 9588 15932
rect 9640 15920 9646 15972
rect 32 15892 60 15920
rect 1673 15895 1731 15901
rect 1673 15892 1685 15895
rect 32 15864 1685 15892
rect 1673 15861 1685 15864
rect 1719 15861 1731 15895
rect 2682 15892 2688 15904
rect 2643 15864 2688 15892
rect 1673 15855 1731 15861
rect 2682 15852 2688 15864
rect 2740 15852 2746 15904
rect 3234 15892 3240 15904
rect 3195 15864 3240 15892
rect 3234 15852 3240 15864
rect 3292 15852 3298 15904
rect 6362 15852 6368 15904
rect 6420 15892 6426 15904
rect 8021 15895 8079 15901
rect 8021 15892 8033 15895
rect 6420 15864 8033 15892
rect 6420 15852 6426 15864
rect 8021 15861 8033 15864
rect 8067 15861 8079 15895
rect 8021 15855 8079 15861
rect 1104 15802 22816 15824
rect 1104 15750 8982 15802
rect 9034 15750 9046 15802
rect 9098 15750 9110 15802
rect 9162 15750 9174 15802
rect 9226 15750 16982 15802
rect 17034 15750 17046 15802
rect 17098 15750 17110 15802
rect 17162 15750 17174 15802
rect 17226 15750 22816 15802
rect 1104 15728 22816 15750
rect 198 15648 204 15700
rect 256 15688 262 15700
rect 1857 15691 1915 15697
rect 1857 15688 1869 15691
rect 256 15660 1869 15688
rect 256 15648 262 15660
rect 1857 15657 1869 15660
rect 1903 15657 1915 15691
rect 2866 15688 2872 15700
rect 2827 15660 2872 15688
rect 1857 15651 1915 15657
rect 2866 15648 2872 15660
rect 2924 15648 2930 15700
rect 3881 15691 3939 15697
rect 3881 15657 3893 15691
rect 3927 15688 3939 15691
rect 3970 15688 3976 15700
rect 3927 15660 3976 15688
rect 3927 15657 3939 15660
rect 3881 15651 3939 15657
rect 3970 15648 3976 15660
rect 4028 15648 4034 15700
rect 4617 15691 4675 15697
rect 4617 15657 4629 15691
rect 4663 15688 4675 15691
rect 4706 15688 4712 15700
rect 4663 15660 4712 15688
rect 4663 15657 4675 15660
rect 4617 15651 4675 15657
rect 4706 15648 4712 15660
rect 4764 15688 4770 15700
rect 5626 15688 5632 15700
rect 4764 15660 5632 15688
rect 4764 15648 4770 15660
rect 5626 15648 5632 15660
rect 5684 15648 5690 15700
rect 5718 15648 5724 15700
rect 5776 15688 5782 15700
rect 6454 15688 6460 15700
rect 5776 15660 6460 15688
rect 5776 15648 5782 15660
rect 6454 15648 6460 15660
rect 6512 15648 6518 15700
rect 2130 15580 2136 15632
rect 2188 15620 2194 15632
rect 3237 15623 3295 15629
rect 3237 15620 3249 15623
rect 2188 15592 3249 15620
rect 2188 15580 2194 15592
rect 1854 15552 1860 15564
rect 1815 15524 1860 15552
rect 1854 15512 1860 15524
rect 1912 15512 1918 15564
rect 2332 15561 2360 15592
rect 3237 15589 3249 15592
rect 3283 15620 3295 15623
rect 3326 15620 3332 15632
rect 3283 15592 3332 15620
rect 3283 15589 3295 15592
rect 3237 15583 3295 15589
rect 3326 15580 3332 15592
rect 3384 15620 3390 15632
rect 4246 15620 4252 15632
rect 3384 15592 4252 15620
rect 3384 15580 3390 15592
rect 4246 15580 4252 15592
rect 4304 15580 4310 15632
rect 6181 15623 6239 15629
rect 6181 15589 6193 15623
rect 6227 15620 6239 15623
rect 7377 15623 7435 15629
rect 7377 15620 7389 15623
rect 6227 15592 7389 15620
rect 6227 15589 6239 15592
rect 6181 15583 6239 15589
rect 7377 15589 7389 15592
rect 7423 15620 7435 15623
rect 7834 15620 7840 15632
rect 7423 15592 7840 15620
rect 7423 15589 7435 15592
rect 7377 15583 7435 15589
rect 7834 15580 7840 15592
rect 7892 15580 7898 15632
rect 2317 15555 2375 15561
rect 2317 15521 2329 15555
rect 2363 15521 2375 15555
rect 2317 15515 2375 15521
rect 3786 15512 3792 15564
rect 3844 15552 3850 15564
rect 4522 15552 4528 15564
rect 3844 15524 4528 15552
rect 3844 15512 3850 15524
rect 4522 15512 4528 15524
rect 4580 15552 4586 15564
rect 4709 15555 4767 15561
rect 4709 15552 4721 15555
rect 4580 15524 4721 15552
rect 4580 15512 4586 15524
rect 4709 15521 4721 15524
rect 4755 15521 4767 15555
rect 4709 15515 4767 15521
rect 6270 15512 6276 15564
rect 6328 15552 6334 15564
rect 7285 15555 7343 15561
rect 7285 15552 7297 15555
rect 6328 15524 7297 15552
rect 6328 15512 6334 15524
rect 7285 15521 7297 15524
rect 7331 15552 7343 15555
rect 7331 15524 7696 15552
rect 7331 15521 7343 15524
rect 7285 15515 7343 15521
rect 7668 15496 7696 15524
rect 4798 15444 4804 15496
rect 4856 15484 4862 15496
rect 5077 15487 5135 15493
rect 5077 15484 5089 15487
rect 4856 15456 5089 15484
rect 4856 15444 4862 15456
rect 5077 15453 5089 15456
rect 5123 15484 5135 15487
rect 5534 15484 5540 15496
rect 5123 15456 5540 15484
rect 5123 15453 5135 15456
rect 5077 15447 5135 15453
rect 5534 15444 5540 15456
rect 5592 15444 5598 15496
rect 7650 15444 7656 15496
rect 7708 15444 7714 15496
rect 3970 15376 3976 15428
rect 4028 15416 4034 15428
rect 5169 15419 5227 15425
rect 5169 15416 5181 15419
rect 4028 15388 5181 15416
rect 4028 15376 4034 15388
rect 5169 15385 5181 15388
rect 5215 15385 5227 15419
rect 5169 15379 5227 15385
rect 1578 15348 1584 15360
rect 1539 15320 1584 15348
rect 1578 15308 1584 15320
rect 1636 15308 1642 15360
rect 4706 15308 4712 15360
rect 4764 15348 4770 15360
rect 4847 15351 4905 15357
rect 4847 15348 4859 15351
rect 4764 15320 4859 15348
rect 4764 15308 4770 15320
rect 4847 15317 4859 15320
rect 4893 15317 4905 15351
rect 4847 15311 4905 15317
rect 4985 15351 5043 15357
rect 4985 15317 4997 15351
rect 5031 15348 5043 15351
rect 5350 15348 5356 15360
rect 5031 15320 5356 15348
rect 5031 15317 5043 15320
rect 4985 15311 5043 15317
rect 5350 15308 5356 15320
rect 5408 15308 5414 15360
rect 5442 15308 5448 15360
rect 5500 15348 5506 15360
rect 5721 15351 5779 15357
rect 5721 15348 5733 15351
rect 5500 15320 5733 15348
rect 5500 15308 5506 15320
rect 5721 15317 5733 15320
rect 5767 15317 5779 15351
rect 5721 15311 5779 15317
rect 1104 15258 22816 15280
rect 1104 15206 4982 15258
rect 5034 15206 5046 15258
rect 5098 15206 5110 15258
rect 5162 15206 5174 15258
rect 5226 15206 12982 15258
rect 13034 15206 13046 15258
rect 13098 15206 13110 15258
rect 13162 15206 13174 15258
rect 13226 15206 20982 15258
rect 21034 15206 21046 15258
rect 21098 15206 21110 15258
rect 21162 15206 21174 15258
rect 21226 15206 22816 15258
rect 1104 15184 22816 15206
rect 106 15104 112 15156
rect 164 15144 170 15156
rect 3326 15144 3332 15156
rect 164 15116 2912 15144
rect 3287 15116 3332 15144
rect 164 15104 170 15116
rect 2884 15017 2912 15116
rect 3326 15104 3332 15116
rect 3384 15104 3390 15156
rect 3786 15144 3792 15156
rect 3747 15116 3792 15144
rect 3786 15104 3792 15116
rect 3844 15104 3850 15156
rect 4062 15144 4068 15156
rect 4023 15116 4068 15144
rect 4062 15104 4068 15116
rect 4120 15104 4126 15156
rect 4709 15147 4767 15153
rect 4709 15113 4721 15147
rect 4755 15144 4767 15147
rect 4798 15144 4804 15156
rect 4755 15116 4804 15144
rect 4755 15113 4767 15116
rect 4709 15107 4767 15113
rect 4798 15104 4804 15116
rect 4856 15104 4862 15156
rect 5077 15147 5135 15153
rect 5077 15113 5089 15147
rect 5123 15144 5135 15147
rect 5334 15147 5392 15153
rect 5334 15144 5346 15147
rect 5123 15116 5346 15144
rect 5123 15113 5135 15116
rect 5077 15107 5135 15113
rect 5334 15113 5346 15116
rect 5380 15144 5392 15147
rect 6638 15144 6644 15156
rect 5380 15116 6644 15144
rect 5380 15113 5392 15116
rect 5334 15107 5392 15113
rect 6638 15104 6644 15116
rect 6696 15144 6702 15156
rect 6963 15147 7021 15153
rect 6963 15144 6975 15147
rect 6696 15116 6975 15144
rect 6696 15104 6702 15116
rect 6963 15113 6975 15116
rect 7009 15113 7021 15147
rect 6963 15107 7021 15113
rect 5445 15079 5503 15085
rect 5445 15045 5457 15079
rect 5491 15076 5503 15079
rect 6086 15076 6092 15088
rect 5491 15048 6092 15076
rect 5491 15045 5503 15048
rect 5445 15039 5503 15045
rect 2869 15011 2927 15017
rect 2869 14977 2881 15011
rect 2915 14977 2927 15011
rect 2869 14971 2927 14977
rect 5258 14968 5264 15020
rect 5316 15008 5322 15020
rect 5460 15008 5488 15039
rect 6086 15036 6092 15048
rect 6144 15036 6150 15088
rect 6270 15076 6276 15088
rect 6231 15048 6276 15076
rect 6270 15036 6276 15048
rect 6328 15036 6334 15088
rect 5316 14980 5488 15008
rect 5537 15011 5595 15017
rect 5316 14968 5322 14980
rect 5537 14977 5549 15011
rect 5583 14977 5595 15011
rect 5537 14971 5595 14977
rect 2225 14943 2283 14949
rect 2225 14909 2237 14943
rect 2271 14940 2283 14943
rect 2593 14943 2651 14949
rect 2593 14940 2605 14943
rect 2271 14912 2605 14940
rect 2271 14909 2283 14912
rect 2225 14903 2283 14909
rect 2593 14909 2605 14912
rect 2639 14909 2651 14943
rect 2774 14940 2780 14952
rect 2687 14912 2780 14940
rect 2593 14903 2651 14909
rect 2608 14872 2636 14903
rect 2774 14900 2780 14912
rect 2832 14940 2838 14952
rect 3326 14940 3332 14952
rect 2832 14912 3332 14940
rect 2832 14900 2838 14912
rect 3326 14900 3332 14912
rect 3384 14900 3390 14952
rect 3881 14943 3939 14949
rect 3881 14909 3893 14943
rect 3927 14940 3939 14943
rect 4246 14940 4252 14952
rect 3927 14912 4252 14940
rect 3927 14909 3939 14912
rect 3881 14903 3939 14909
rect 4246 14900 4252 14912
rect 4304 14900 4310 14952
rect 5442 14900 5448 14952
rect 5500 14940 5506 14952
rect 5552 14940 5580 14971
rect 5500 14912 5580 14940
rect 6104 14940 6132 15036
rect 7190 15008 7196 15020
rect 7151 14980 7196 15008
rect 7190 14968 7196 14980
rect 7248 14968 7254 15020
rect 7282 14968 7288 15020
rect 7340 15008 7346 15020
rect 7340 14980 7385 15008
rect 7340 14968 7346 14980
rect 7055 14943 7113 14949
rect 7055 14940 7067 14943
rect 6104 14912 7067 14940
rect 5500 14900 5506 14912
rect 7055 14909 7067 14912
rect 7101 14940 7113 14943
rect 7837 14943 7895 14949
rect 7837 14940 7849 14943
rect 7101 14912 7849 14940
rect 7101 14909 7113 14912
rect 7055 14903 7113 14909
rect 7837 14909 7849 14912
rect 7883 14909 7895 14943
rect 7837 14903 7895 14909
rect 2682 14872 2688 14884
rect 2595 14844 2688 14872
rect 2682 14832 2688 14844
rect 2740 14872 2746 14884
rect 3602 14872 3608 14884
rect 2740 14844 3608 14872
rect 2740 14832 2746 14844
rect 3602 14832 3608 14844
rect 3660 14832 3666 14884
rect 5169 14875 5227 14881
rect 5169 14841 5181 14875
rect 5215 14872 5227 14875
rect 6822 14872 6828 14884
rect 5215 14844 6828 14872
rect 5215 14841 5227 14844
rect 5169 14835 5227 14841
rect 6822 14832 6828 14844
rect 6880 14832 6886 14884
rect 1854 14804 1860 14816
rect 1815 14776 1860 14804
rect 1854 14764 1860 14776
rect 1912 14764 1918 14816
rect 4062 14764 4068 14816
rect 4120 14804 4126 14816
rect 4430 14804 4436 14816
rect 4120 14776 4436 14804
rect 4120 14764 4126 14776
rect 4430 14764 4436 14776
rect 4488 14764 4494 14816
rect 4522 14764 4528 14816
rect 4580 14804 4586 14816
rect 5813 14807 5871 14813
rect 5813 14804 5825 14807
rect 4580 14776 5825 14804
rect 4580 14764 4586 14776
rect 5813 14773 5825 14776
rect 5859 14773 5871 14807
rect 5813 14767 5871 14773
rect 1104 14714 22816 14736
rect 1104 14662 8982 14714
rect 9034 14662 9046 14714
rect 9098 14662 9110 14714
rect 9162 14662 9174 14714
rect 9226 14662 16982 14714
rect 17034 14662 17046 14714
rect 17098 14662 17110 14714
rect 17162 14662 17174 14714
rect 17226 14662 22816 14714
rect 1104 14640 22816 14662
rect 14 14560 20 14612
rect 72 14600 78 14612
rect 2317 14603 2375 14609
rect 2317 14600 2329 14603
rect 72 14572 2329 14600
rect 72 14560 78 14572
rect 2317 14569 2329 14572
rect 2363 14569 2375 14603
rect 2317 14563 2375 14569
rect 3881 14603 3939 14609
rect 3881 14569 3893 14603
rect 3927 14600 3939 14603
rect 4246 14600 4252 14612
rect 3927 14572 4252 14600
rect 3927 14569 3939 14572
rect 3881 14563 3939 14569
rect 4246 14560 4252 14572
rect 4304 14560 4310 14612
rect 6270 14600 6276 14612
rect 5092 14572 6276 14600
rect 1857 14535 1915 14541
rect 1857 14501 1869 14535
rect 1903 14532 1915 14535
rect 1903 14504 2820 14532
rect 1903 14501 1915 14504
rect 1857 14495 1915 14501
rect 2792 14476 2820 14504
rect 4798 14492 4804 14544
rect 4856 14532 4862 14544
rect 5092 14541 5120 14572
rect 6270 14560 6276 14572
rect 6328 14560 6334 14612
rect 6822 14560 6828 14612
rect 6880 14600 6886 14612
rect 7561 14603 7619 14609
rect 7561 14600 7573 14603
rect 6880 14572 7573 14600
rect 6880 14560 6886 14572
rect 7561 14569 7573 14572
rect 7607 14600 7619 14603
rect 7834 14600 7840 14612
rect 7607 14572 7840 14600
rect 7607 14569 7619 14572
rect 7561 14563 7619 14569
rect 7834 14560 7840 14572
rect 7892 14560 7898 14612
rect 5077 14535 5135 14541
rect 5077 14532 5089 14535
rect 4856 14504 5089 14532
rect 4856 14492 4862 14504
rect 5077 14501 5089 14504
rect 5123 14501 5135 14535
rect 5077 14495 5135 14501
rect 5534 14492 5540 14544
rect 5592 14532 5598 14544
rect 7101 14535 7159 14541
rect 7101 14532 7113 14535
rect 5592 14504 7113 14532
rect 5592 14492 5598 14504
rect 7101 14501 7113 14504
rect 7147 14532 7159 14535
rect 7190 14532 7196 14544
rect 7147 14504 7196 14532
rect 7147 14501 7159 14504
rect 7101 14495 7159 14501
rect 7190 14492 7196 14504
rect 7248 14492 7254 14544
rect 1670 14424 1676 14476
rect 1728 14464 1734 14476
rect 2225 14467 2283 14473
rect 2225 14464 2237 14467
rect 1728 14436 2237 14464
rect 1728 14424 1734 14436
rect 2225 14433 2237 14436
rect 2271 14433 2283 14467
rect 2774 14464 2780 14476
rect 2735 14436 2780 14464
rect 2225 14427 2283 14433
rect 2774 14424 2780 14436
rect 2832 14424 2838 14476
rect 3878 14424 3884 14476
rect 3936 14464 3942 14476
rect 4065 14467 4123 14473
rect 4065 14464 4077 14467
rect 3936 14436 4077 14464
rect 3936 14424 3942 14436
rect 4065 14433 4077 14436
rect 4111 14464 4123 14467
rect 4522 14464 4528 14476
rect 4111 14436 4528 14464
rect 4111 14433 4123 14436
rect 4065 14427 4123 14433
rect 4522 14424 4528 14436
rect 4580 14424 4586 14476
rect 4706 14424 4712 14476
rect 4764 14464 4770 14476
rect 5224 14467 5282 14473
rect 5224 14464 5236 14467
rect 4764 14436 5236 14464
rect 4764 14424 4770 14436
rect 5224 14433 5236 14436
rect 5270 14433 5282 14467
rect 6086 14464 6092 14476
rect 6047 14436 6092 14464
rect 5224 14427 5282 14433
rect 6086 14424 6092 14436
rect 6144 14424 6150 14476
rect 6270 14424 6276 14476
rect 6328 14464 6334 14476
rect 6641 14467 6699 14473
rect 6641 14464 6653 14467
rect 6328 14436 6653 14464
rect 6328 14424 6334 14436
rect 6641 14433 6653 14436
rect 6687 14433 6699 14467
rect 6641 14427 6699 14433
rect 5442 14396 5448 14408
rect 5403 14368 5448 14396
rect 5442 14356 5448 14368
rect 5500 14356 5506 14408
rect 1946 14288 1952 14340
rect 2004 14328 2010 14340
rect 3329 14331 3387 14337
rect 3329 14328 3341 14331
rect 2004 14300 3341 14328
rect 2004 14288 2010 14300
rect 3329 14297 3341 14300
rect 3375 14328 3387 14331
rect 4430 14328 4436 14340
rect 3375 14300 4436 14328
rect 3375 14297 3387 14300
rect 3329 14291 3387 14297
rect 4430 14288 4436 14300
rect 4488 14288 4494 14340
rect 5258 14328 5264 14340
rect 4540 14300 5264 14328
rect 4246 14260 4252 14272
rect 4207 14232 4252 14260
rect 4246 14220 4252 14232
rect 4304 14220 4310 14272
rect 4338 14220 4344 14272
rect 4396 14260 4402 14272
rect 4540 14260 4568 14300
rect 5258 14288 5264 14300
rect 5316 14328 5322 14340
rect 5353 14331 5411 14337
rect 5353 14328 5365 14331
rect 5316 14300 5365 14328
rect 5316 14288 5322 14300
rect 5353 14297 5365 14300
rect 5399 14297 5411 14331
rect 5353 14291 5411 14297
rect 4706 14260 4712 14272
rect 4396 14232 4568 14260
rect 4667 14232 4712 14260
rect 4396 14220 4402 14232
rect 4706 14220 4712 14232
rect 4764 14220 4770 14272
rect 5718 14260 5724 14272
rect 5679 14232 5724 14260
rect 5718 14220 5724 14232
rect 5776 14220 5782 14272
rect 6362 14220 6368 14272
rect 6420 14260 6426 14272
rect 6825 14263 6883 14269
rect 6825 14260 6837 14263
rect 6420 14232 6837 14260
rect 6420 14220 6426 14232
rect 6825 14229 6837 14232
rect 6871 14229 6883 14263
rect 6825 14223 6883 14229
rect 1104 14170 22816 14192
rect 1104 14118 4982 14170
rect 5034 14118 5046 14170
rect 5098 14118 5110 14170
rect 5162 14118 5174 14170
rect 5226 14118 12982 14170
rect 13034 14118 13046 14170
rect 13098 14118 13110 14170
rect 13162 14118 13174 14170
rect 13226 14118 20982 14170
rect 21034 14118 21046 14170
rect 21098 14118 21110 14170
rect 21162 14118 21174 14170
rect 21226 14118 22816 14170
rect 1104 14096 22816 14118
rect 2501 14059 2559 14065
rect 2501 14025 2513 14059
rect 2547 14056 2559 14059
rect 2774 14056 2780 14068
rect 2547 14028 2780 14056
rect 2547 14025 2559 14028
rect 2501 14019 2559 14025
rect 2774 14016 2780 14028
rect 2832 14016 2838 14068
rect 4617 14059 4675 14065
rect 4617 14025 4629 14059
rect 4663 14056 4675 14059
rect 4798 14056 4804 14068
rect 4663 14028 4804 14056
rect 4663 14025 4675 14028
rect 4617 14019 4675 14025
rect 4798 14016 4804 14028
rect 4856 14056 4862 14068
rect 4893 14059 4951 14065
rect 4893 14056 4905 14059
rect 4856 14028 4905 14056
rect 4856 14016 4862 14028
rect 4893 14025 4905 14028
rect 4939 14025 4951 14059
rect 4893 14019 4951 14025
rect 2130 13948 2136 14000
rect 2188 13988 2194 14000
rect 2188 13960 3004 13988
rect 2188 13948 2194 13960
rect 1670 13852 1676 13864
rect 1631 13824 1676 13852
rect 1670 13812 1676 13824
rect 1728 13812 1734 13864
rect 1946 13852 1952 13864
rect 1907 13824 1952 13852
rect 1946 13812 1952 13824
rect 2004 13812 2010 13864
rect 2976 13861 3004 13960
rect 4246 13920 4252 13932
rect 4126 13892 4252 13920
rect 2961 13855 3019 13861
rect 2961 13821 2973 13855
rect 3007 13821 3019 13855
rect 3513 13855 3571 13861
rect 3513 13852 3525 13855
rect 3423 13824 3525 13852
rect 2961 13815 3019 13821
rect 3513 13821 3525 13824
rect 3559 13852 3571 13855
rect 4126 13852 4154 13892
rect 4246 13880 4252 13892
rect 4304 13880 4310 13932
rect 3559 13824 4154 13852
rect 4908 13852 4936 14019
rect 5626 14016 5632 14068
rect 5684 14056 5690 14068
rect 6089 14059 6147 14065
rect 6089 14056 6101 14059
rect 5684 14028 6101 14056
rect 5684 14016 5690 14028
rect 6089 14025 6101 14028
rect 6135 14025 6147 14059
rect 6089 14019 6147 14025
rect 6270 14016 6276 14068
rect 6328 14056 6334 14068
rect 6549 14059 6607 14065
rect 6549 14056 6561 14059
rect 6328 14028 6561 14056
rect 6328 14016 6334 14028
rect 6549 14025 6561 14028
rect 6595 14025 6607 14059
rect 6549 14019 6607 14025
rect 5353 13991 5411 13997
rect 5353 13957 5365 13991
rect 5399 13988 5411 13991
rect 5399 13960 6132 13988
rect 5399 13957 5411 13960
rect 5353 13951 5411 13957
rect 6104 13932 6132 13960
rect 5445 13923 5503 13929
rect 5445 13920 5457 13923
rect 5368 13892 5457 13920
rect 5258 13861 5264 13864
rect 5077 13855 5135 13861
rect 5077 13852 5089 13855
rect 4908 13824 5089 13852
rect 3559 13821 3571 13824
rect 3513 13815 3571 13821
rect 5077 13821 5089 13824
rect 5123 13821 5135 13855
rect 5077 13815 5135 13821
rect 5224 13855 5264 13861
rect 5224 13821 5236 13855
rect 5224 13815 5264 13821
rect 2866 13784 2872 13796
rect 2779 13756 2872 13784
rect 2866 13744 2872 13756
rect 2924 13784 2930 13796
rect 3528 13784 3556 13815
rect 5258 13812 5264 13815
rect 5316 13812 5322 13864
rect 2924 13756 3556 13784
rect 4249 13787 4307 13793
rect 2924 13744 2930 13756
rect 4249 13753 4261 13787
rect 4295 13784 4307 13787
rect 4798 13784 4804 13796
rect 4295 13756 4804 13784
rect 4295 13753 4307 13756
rect 4249 13747 4307 13753
rect 4798 13744 4804 13756
rect 4856 13784 4862 13796
rect 5368 13784 5396 13892
rect 5445 13889 5457 13892
rect 5491 13920 5503 13923
rect 5534 13920 5540 13932
rect 5491 13892 5540 13920
rect 5491 13889 5503 13892
rect 5445 13883 5503 13889
rect 5534 13880 5540 13892
rect 5592 13880 5598 13932
rect 6086 13880 6092 13932
rect 6144 13880 6150 13932
rect 7466 13920 7472 13932
rect 7024 13892 7472 13920
rect 7024 13861 7052 13892
rect 7466 13880 7472 13892
rect 7524 13920 7530 13932
rect 7837 13923 7895 13929
rect 7837 13920 7849 13923
rect 7524 13892 7849 13920
rect 7524 13880 7530 13892
rect 7837 13889 7849 13892
rect 7883 13889 7895 13923
rect 7837 13883 7895 13889
rect 7009 13855 7067 13861
rect 7009 13821 7021 13855
rect 7055 13821 7067 13855
rect 7282 13852 7288 13864
rect 7243 13824 7288 13852
rect 7009 13815 7067 13821
rect 7282 13812 7288 13824
rect 7340 13812 7346 13864
rect 4856 13756 5396 13784
rect 4856 13744 4862 13756
rect 106 13676 112 13728
rect 164 13716 170 13728
rect 1489 13719 1547 13725
rect 1489 13716 1501 13719
rect 164 13688 1501 13716
rect 164 13676 170 13688
rect 1489 13685 1501 13688
rect 1535 13685 1547 13719
rect 3050 13716 3056 13728
rect 3011 13688 3056 13716
rect 1489 13679 1547 13685
rect 3050 13676 3056 13688
rect 3108 13676 3114 13728
rect 5721 13719 5779 13725
rect 5721 13685 5733 13719
rect 5767 13716 5779 13719
rect 5902 13716 5908 13728
rect 5767 13688 5908 13716
rect 5767 13685 5779 13688
rect 5721 13679 5779 13685
rect 5902 13676 5908 13688
rect 5960 13676 5966 13728
rect 6914 13716 6920 13728
rect 6875 13688 6920 13716
rect 6914 13676 6920 13688
rect 6972 13676 6978 13728
rect 1104 13626 22816 13648
rect 1104 13574 8982 13626
rect 9034 13574 9046 13626
rect 9098 13574 9110 13626
rect 9162 13574 9174 13626
rect 9226 13574 16982 13626
rect 17034 13574 17046 13626
rect 17098 13574 17110 13626
rect 17162 13574 17174 13626
rect 17226 13574 22816 13626
rect 1104 13552 22816 13574
rect 1578 13512 1584 13524
rect 1539 13484 1584 13512
rect 1578 13472 1584 13484
rect 1636 13472 1642 13524
rect 1946 13512 1952 13524
rect 1907 13484 1952 13512
rect 1946 13472 1952 13484
rect 2004 13472 2010 13524
rect 2501 13515 2559 13521
rect 2501 13481 2513 13515
rect 2547 13481 2559 13515
rect 3878 13512 3884 13524
rect 3839 13484 3884 13512
rect 2501 13475 2559 13481
rect 106 13404 112 13456
rect 164 13444 170 13456
rect 2516 13444 2544 13475
rect 3878 13472 3884 13484
rect 3936 13472 3942 13524
rect 4338 13512 4344 13524
rect 4299 13484 4344 13512
rect 4338 13472 4344 13484
rect 4396 13472 4402 13524
rect 4430 13472 4436 13524
rect 4488 13512 4494 13524
rect 5445 13515 5503 13521
rect 5445 13512 5457 13515
rect 4488 13484 5457 13512
rect 4488 13472 4494 13484
rect 5445 13481 5457 13484
rect 5491 13481 5503 13515
rect 5445 13475 5503 13481
rect 5534 13472 5540 13524
rect 5592 13512 5598 13524
rect 6549 13515 6607 13521
rect 6549 13512 6561 13515
rect 5592 13484 6561 13512
rect 5592 13472 5598 13484
rect 6549 13481 6561 13484
rect 6595 13481 6607 13515
rect 6549 13475 6607 13481
rect 6917 13515 6975 13521
rect 6917 13481 6929 13515
rect 6963 13512 6975 13515
rect 7282 13512 7288 13524
rect 6963 13484 7288 13512
rect 6963 13481 6975 13484
rect 6917 13475 6975 13481
rect 7282 13472 7288 13484
rect 7340 13472 7346 13524
rect 164 13416 2544 13444
rect 164 13404 170 13416
rect 5626 13404 5632 13456
rect 5684 13444 5690 13456
rect 5813 13447 5871 13453
rect 5813 13444 5825 13447
rect 5684 13416 5825 13444
rect 5684 13404 5690 13416
rect 5813 13413 5825 13416
rect 5859 13413 5871 13447
rect 5813 13407 5871 13413
rect 6086 13404 6092 13456
rect 6144 13444 6150 13456
rect 6181 13447 6239 13453
rect 6181 13444 6193 13447
rect 6144 13416 6193 13444
rect 6144 13404 6150 13416
rect 6181 13413 6193 13416
rect 6227 13413 6239 13447
rect 6181 13407 6239 13413
rect 1397 13379 1455 13385
rect 1397 13345 1409 13379
rect 1443 13376 1455 13379
rect 2130 13376 2136 13388
rect 1443 13348 2136 13376
rect 1443 13345 1455 13348
rect 1397 13339 1455 13345
rect 2130 13336 2136 13348
rect 2188 13336 2194 13388
rect 2222 13336 2228 13388
rect 2280 13376 2286 13388
rect 2409 13379 2467 13385
rect 2409 13376 2421 13379
rect 2280 13348 2421 13376
rect 2280 13336 2286 13348
rect 2409 13345 2421 13348
rect 2455 13345 2467 13379
rect 2866 13376 2872 13388
rect 2827 13348 2872 13376
rect 2409 13339 2467 13345
rect 2866 13336 2872 13348
rect 2924 13336 2930 13388
rect 4614 13336 4620 13388
rect 4672 13376 4678 13388
rect 4801 13379 4859 13385
rect 4801 13376 4813 13379
rect 4672 13348 4813 13376
rect 4672 13336 4678 13348
rect 4801 13345 4813 13348
rect 4847 13345 4859 13379
rect 4801 13339 4859 13345
rect 4948 13379 5006 13385
rect 4948 13345 4960 13379
rect 4994 13376 5006 13379
rect 5258 13376 5264 13388
rect 4994 13348 5264 13376
rect 4994 13345 5006 13348
rect 4948 13339 5006 13345
rect 5258 13336 5264 13348
rect 5316 13376 5322 13388
rect 5644 13376 5672 13404
rect 5316 13348 5672 13376
rect 6365 13379 6423 13385
rect 5316 13336 5322 13348
rect 6365 13345 6377 13379
rect 6411 13376 6423 13379
rect 7558 13376 7564 13388
rect 6411 13348 7328 13376
rect 7519 13348 7564 13376
rect 6411 13345 6423 13348
rect 6365 13339 6423 13345
rect 7300 13320 7328 13348
rect 7558 13336 7564 13348
rect 7616 13336 7622 13388
rect 4709 13311 4767 13317
rect 4709 13277 4721 13311
rect 4755 13308 4767 13311
rect 5169 13311 5227 13317
rect 5169 13308 5181 13311
rect 4755 13280 5181 13308
rect 4755 13277 4767 13280
rect 4709 13271 4767 13277
rect 5169 13277 5181 13280
rect 5215 13308 5227 13311
rect 5442 13308 5448 13320
rect 5215 13280 5448 13308
rect 5215 13277 5227 13280
rect 5169 13271 5227 13277
rect 5442 13268 5448 13280
rect 5500 13268 5506 13320
rect 7282 13308 7288 13320
rect 7195 13280 7288 13308
rect 7282 13268 7288 13280
rect 7340 13308 7346 13320
rect 7377 13311 7435 13317
rect 7377 13308 7389 13311
rect 7340 13280 7389 13308
rect 7340 13268 7346 13280
rect 7377 13277 7389 13280
rect 7423 13277 7435 13311
rect 7377 13271 7435 13277
rect 2317 13243 2375 13249
rect 2317 13209 2329 13243
rect 2363 13240 2375 13243
rect 2774 13240 2780 13252
rect 2363 13212 2780 13240
rect 2363 13209 2375 13212
rect 2317 13203 2375 13209
rect 2774 13200 2780 13212
rect 2832 13240 2838 13252
rect 7466 13240 7472 13252
rect 2832 13212 7472 13240
rect 2832 13200 2838 13212
rect 7466 13200 7472 13212
rect 7524 13200 7530 13252
rect 3418 13172 3424 13184
rect 3379 13144 3424 13172
rect 3418 13132 3424 13144
rect 3476 13132 3482 13184
rect 5077 13175 5135 13181
rect 5077 13141 5089 13175
rect 5123 13172 5135 13175
rect 5350 13172 5356 13184
rect 5123 13144 5356 13172
rect 5123 13141 5135 13144
rect 5077 13135 5135 13141
rect 5350 13132 5356 13144
rect 5408 13132 5414 13184
rect 1104 13082 22816 13104
rect 1104 13030 4982 13082
rect 5034 13030 5046 13082
rect 5098 13030 5110 13082
rect 5162 13030 5174 13082
rect 5226 13030 12982 13082
rect 13034 13030 13046 13082
rect 13098 13030 13110 13082
rect 13162 13030 13174 13082
rect 13226 13030 20982 13082
rect 21034 13030 21046 13082
rect 21098 13030 21110 13082
rect 21162 13030 21174 13082
rect 21226 13030 22816 13082
rect 1104 13008 22816 13030
rect 1673 12971 1731 12977
rect 1673 12937 1685 12971
rect 1719 12968 1731 12971
rect 1854 12968 1860 12980
rect 1719 12940 1860 12968
rect 1719 12937 1731 12940
rect 1673 12931 1731 12937
rect 1854 12928 1860 12940
rect 1912 12968 1918 12980
rect 3234 12968 3240 12980
rect 1912 12940 3240 12968
rect 1912 12928 1918 12940
rect 3234 12928 3240 12940
rect 3292 12928 3298 12980
rect 4798 12968 4804 12980
rect 4759 12940 4804 12968
rect 4798 12928 4804 12940
rect 4856 12968 4862 12980
rect 4856 12940 5304 12968
rect 4856 12928 4862 12940
rect 5169 12903 5227 12909
rect 5169 12869 5181 12903
rect 5215 12869 5227 12903
rect 5169 12863 5227 12869
rect 4065 12835 4123 12841
rect 4065 12801 4077 12835
rect 4111 12832 4123 12835
rect 4433 12835 4491 12841
rect 4111 12804 4384 12832
rect 4111 12801 4123 12804
rect 4065 12795 4123 12801
rect 1489 12767 1547 12773
rect 1489 12733 1501 12767
rect 1535 12764 1547 12767
rect 2222 12764 2228 12776
rect 1535 12736 2228 12764
rect 1535 12733 1547 12736
rect 1489 12727 1547 12733
rect 2222 12724 2228 12736
rect 2280 12724 2286 12776
rect 2774 12764 2780 12776
rect 2735 12736 2780 12764
rect 2774 12724 2780 12736
rect 2832 12724 2838 12776
rect 2866 12724 2872 12776
rect 2924 12764 2930 12776
rect 2961 12767 3019 12773
rect 2961 12764 2973 12767
rect 2924 12736 2973 12764
rect 2924 12724 2930 12736
rect 2961 12733 2973 12736
rect 3007 12733 3019 12767
rect 2961 12727 3019 12733
rect 3605 12767 3663 12773
rect 3605 12733 3617 12767
rect 3651 12764 3663 12767
rect 4246 12764 4252 12776
rect 3651 12736 4252 12764
rect 3651 12733 3663 12736
rect 3605 12727 3663 12733
rect 4246 12724 4252 12736
rect 4304 12724 4310 12776
rect 4356 12764 4384 12804
rect 4433 12801 4445 12835
rect 4479 12832 4491 12835
rect 4706 12832 4712 12844
rect 4479 12804 4712 12832
rect 4479 12801 4491 12804
rect 4433 12795 4491 12801
rect 4706 12792 4712 12804
rect 4764 12832 4770 12844
rect 5184 12832 5212 12863
rect 5276 12841 5304 12940
rect 5626 12928 5632 12980
rect 5684 12968 5690 12980
rect 5905 12971 5963 12977
rect 5905 12968 5917 12971
rect 5684 12940 5917 12968
rect 5684 12928 5690 12940
rect 5905 12937 5917 12940
rect 5951 12937 5963 12971
rect 5905 12931 5963 12937
rect 7558 12928 7564 12980
rect 7616 12968 7622 12980
rect 8113 12971 8171 12977
rect 8113 12968 8125 12971
rect 7616 12940 8125 12968
rect 7616 12928 7622 12940
rect 8113 12937 8125 12940
rect 8159 12937 8171 12971
rect 8113 12931 8171 12937
rect 4764 12804 5212 12832
rect 4764 12792 4770 12804
rect 5040 12767 5098 12773
rect 5040 12764 5052 12767
rect 4356 12736 5052 12764
rect 5040 12733 5052 12736
rect 5086 12764 5098 12767
rect 5184 12764 5212 12804
rect 5261 12835 5319 12841
rect 5261 12801 5273 12835
rect 5307 12801 5319 12835
rect 5261 12795 5319 12801
rect 5350 12764 5356 12776
rect 5086 12733 5120 12764
rect 5184 12736 5356 12764
rect 5040 12727 5120 12733
rect 2041 12699 2099 12705
rect 2041 12665 2053 12699
rect 2087 12696 2099 12699
rect 2409 12699 2467 12705
rect 2409 12696 2421 12699
rect 2087 12668 2421 12696
rect 2087 12665 2099 12668
rect 2041 12659 2099 12665
rect 2409 12665 2421 12668
rect 2455 12696 2467 12699
rect 2884 12696 2912 12724
rect 2455 12668 2912 12696
rect 2455 12665 2467 12668
rect 2409 12659 2467 12665
rect 4614 12656 4620 12708
rect 4672 12696 4678 12708
rect 4893 12699 4951 12705
rect 4893 12696 4905 12699
rect 4672 12668 4905 12696
rect 4672 12656 4678 12668
rect 4893 12665 4905 12668
rect 4939 12665 4951 12699
rect 5092 12696 5120 12727
rect 5350 12724 5356 12736
rect 5408 12724 5414 12776
rect 7374 12764 7380 12776
rect 7335 12736 7380 12764
rect 7374 12724 7380 12736
rect 7432 12724 7438 12776
rect 5626 12696 5632 12708
rect 5092 12668 5632 12696
rect 4893 12659 4951 12665
rect 5626 12656 5632 12668
rect 5684 12656 5690 12708
rect 6086 12656 6092 12708
rect 6144 12696 6150 12708
rect 7101 12699 7159 12705
rect 7101 12696 7113 12699
rect 6144 12668 7113 12696
rect 6144 12656 6150 12668
rect 7101 12665 7113 12668
rect 7147 12665 7159 12699
rect 7101 12659 7159 12665
rect 14 12588 20 12640
rect 72 12628 78 12640
rect 2593 12631 2651 12637
rect 2593 12628 2605 12631
rect 72 12600 2605 12628
rect 72 12588 78 12600
rect 2593 12597 2605 12600
rect 2639 12597 2651 12631
rect 5534 12628 5540 12640
rect 5495 12600 5540 12628
rect 2593 12591 2651 12597
rect 5534 12588 5540 12600
rect 5592 12588 5598 12640
rect 6362 12628 6368 12640
rect 6323 12600 6368 12628
rect 6362 12588 6368 12600
rect 6420 12588 6426 12640
rect 1104 12538 22816 12560
rect 1104 12486 8982 12538
rect 9034 12486 9046 12538
rect 9098 12486 9110 12538
rect 9162 12486 9174 12538
rect 9226 12486 16982 12538
rect 17034 12486 17046 12538
rect 17098 12486 17110 12538
rect 17162 12486 17174 12538
rect 17226 12486 22816 12538
rect 1104 12464 22816 12486
rect 106 12384 112 12436
rect 164 12424 170 12436
rect 2501 12427 2559 12433
rect 2501 12424 2513 12427
rect 164 12396 2513 12424
rect 164 12384 170 12396
rect 2501 12393 2513 12396
rect 2547 12393 2559 12427
rect 4157 12427 4215 12433
rect 4157 12424 4169 12427
rect 2501 12387 2559 12393
rect 2976 12396 4169 12424
rect 198 12316 204 12368
rect 256 12356 262 12368
rect 2976 12356 3004 12396
rect 4157 12393 4169 12396
rect 4203 12393 4215 12427
rect 5442 12424 5448 12436
rect 5403 12396 5448 12424
rect 4157 12387 4215 12393
rect 5442 12384 5448 12396
rect 5500 12384 5506 12436
rect 6638 12384 6644 12436
rect 6696 12424 6702 12436
rect 7193 12427 7251 12433
rect 7193 12424 7205 12427
rect 6696 12396 7205 12424
rect 6696 12384 6702 12396
rect 7193 12393 7205 12396
rect 7239 12424 7251 12427
rect 7374 12424 7380 12436
rect 7239 12396 7380 12424
rect 7239 12393 7251 12396
rect 7193 12387 7251 12393
rect 7374 12384 7380 12396
rect 7432 12384 7438 12436
rect 256 12328 3004 12356
rect 256 12316 262 12328
rect 3694 12316 3700 12368
rect 3752 12356 3758 12368
rect 4798 12356 4804 12368
rect 3752 12328 4804 12356
rect 3752 12316 3758 12328
rect 4798 12316 4804 12328
rect 4856 12316 4862 12368
rect 6086 12356 6092 12368
rect 6047 12328 6092 12356
rect 6086 12316 6092 12328
rect 6144 12316 6150 12368
rect 7392 12356 7420 12384
rect 7653 12359 7711 12365
rect 7653 12356 7665 12359
rect 7392 12328 7665 12356
rect 7653 12325 7665 12328
rect 7699 12325 7711 12359
rect 7653 12319 7711 12325
rect 1397 12291 1455 12297
rect 1397 12257 1409 12291
rect 1443 12288 1455 12291
rect 1670 12288 1676 12300
rect 1443 12260 1676 12288
rect 1443 12257 1455 12260
rect 1397 12251 1455 12257
rect 1670 12248 1676 12260
rect 1728 12288 1734 12300
rect 2409 12291 2467 12297
rect 2409 12288 2421 12291
rect 1728 12260 2421 12288
rect 1728 12248 1734 12260
rect 2409 12257 2421 12260
rect 2455 12257 2467 12291
rect 2866 12288 2872 12300
rect 2827 12260 2872 12288
rect 2409 12251 2467 12257
rect 2424 12220 2452 12251
rect 2866 12248 2872 12260
rect 2924 12248 2930 12300
rect 4246 12288 4252 12300
rect 4207 12260 4252 12288
rect 4246 12248 4252 12260
rect 4304 12248 4310 12300
rect 4522 12288 4528 12300
rect 4483 12260 4528 12288
rect 4522 12248 4528 12260
rect 4580 12248 4586 12300
rect 6178 12288 6184 12300
rect 6146 12260 6184 12288
rect 6178 12248 6184 12260
rect 6236 12297 6242 12300
rect 6236 12291 6294 12297
rect 6236 12257 6248 12291
rect 6282 12288 6294 12291
rect 7558 12288 7564 12300
rect 6282 12260 7564 12288
rect 6282 12257 6294 12260
rect 6236 12251 6294 12257
rect 6236 12248 6242 12251
rect 7558 12248 7564 12260
rect 7616 12288 7622 12300
rect 7800 12291 7858 12297
rect 7800 12288 7812 12291
rect 7616 12260 7812 12288
rect 7616 12248 7622 12260
rect 7800 12257 7812 12260
rect 7846 12257 7858 12291
rect 7800 12251 7858 12257
rect 2682 12220 2688 12232
rect 2424 12192 2688 12220
rect 2682 12180 2688 12192
rect 2740 12220 2746 12232
rect 3418 12220 3424 12232
rect 2740 12192 3424 12220
rect 2740 12180 2746 12192
rect 3418 12180 3424 12192
rect 3476 12180 3482 12232
rect 6454 12220 6460 12232
rect 6415 12192 6460 12220
rect 6454 12180 6460 12192
rect 6512 12220 6518 12232
rect 8021 12223 8079 12229
rect 8021 12220 8033 12223
rect 6512 12192 8033 12220
rect 6512 12180 6518 12192
rect 8021 12189 8033 12192
rect 8067 12189 8079 12223
rect 8021 12183 8079 12189
rect 2130 12112 2136 12164
rect 2188 12152 2194 12164
rect 3510 12152 3516 12164
rect 2188 12124 3516 12152
rect 2188 12112 2194 12124
rect 3510 12112 3516 12124
rect 3568 12152 3574 12164
rect 3789 12155 3847 12161
rect 3789 12152 3801 12155
rect 3568 12124 3801 12152
rect 3568 12112 3574 12124
rect 3789 12121 3801 12124
rect 3835 12121 3847 12155
rect 3789 12115 3847 12121
rect 4614 12112 4620 12164
rect 4672 12152 4678 12164
rect 5905 12155 5963 12161
rect 5905 12152 5917 12155
rect 4672 12124 5917 12152
rect 4672 12112 4678 12124
rect 5905 12121 5917 12124
rect 5951 12152 5963 12155
rect 6362 12152 6368 12164
rect 5951 12124 6368 12152
rect 5951 12121 5963 12124
rect 5905 12115 5963 12121
rect 6362 12112 6368 12124
rect 6420 12152 6426 12164
rect 7098 12152 7104 12164
rect 6420 12124 7104 12152
rect 6420 12112 6426 12124
rect 7098 12112 7104 12124
rect 7156 12152 7162 12164
rect 7469 12155 7527 12161
rect 7469 12152 7481 12155
rect 7156 12124 7481 12152
rect 7156 12112 7162 12124
rect 7469 12121 7481 12124
rect 7515 12152 7527 12155
rect 7926 12152 7932 12164
rect 7515 12124 7932 12152
rect 7515 12121 7527 12124
rect 7469 12115 7527 12121
rect 7926 12112 7932 12124
rect 7984 12112 7990 12164
rect 1578 12084 1584 12096
rect 1539 12056 1584 12084
rect 1578 12044 1584 12056
rect 1636 12044 1642 12096
rect 1946 12084 1952 12096
rect 1907 12056 1952 12084
rect 1946 12044 1952 12056
rect 2004 12044 2010 12096
rect 2314 12084 2320 12096
rect 2275 12056 2320 12084
rect 2314 12044 2320 12056
rect 2372 12044 2378 12096
rect 5169 12087 5227 12093
rect 5169 12053 5181 12087
rect 5215 12084 5227 12087
rect 5350 12084 5356 12096
rect 5215 12056 5356 12084
rect 5215 12053 5227 12056
rect 5169 12047 5227 12053
rect 5350 12044 5356 12056
rect 5408 12044 5414 12096
rect 6730 12084 6736 12096
rect 6691 12056 6736 12084
rect 6730 12044 6736 12056
rect 6788 12044 6794 12096
rect 8018 12044 8024 12096
rect 8076 12084 8082 12096
rect 8113 12087 8171 12093
rect 8113 12084 8125 12087
rect 8076 12056 8125 12084
rect 8076 12044 8082 12056
rect 8113 12053 8125 12056
rect 8159 12053 8171 12087
rect 8113 12047 8171 12053
rect 1104 11994 22816 12016
rect 1104 11942 4982 11994
rect 5034 11942 5046 11994
rect 5098 11942 5110 11994
rect 5162 11942 5174 11994
rect 5226 11942 12982 11994
rect 13034 11942 13046 11994
rect 13098 11942 13110 11994
rect 13162 11942 13174 11994
rect 13226 11942 20982 11994
rect 21034 11942 21046 11994
rect 21098 11942 21110 11994
rect 21162 11942 21174 11994
rect 21226 11942 22816 11994
rect 1104 11920 22816 11942
rect 2501 11883 2559 11889
rect 2501 11849 2513 11883
rect 2547 11880 2559 11883
rect 2866 11880 2872 11892
rect 2547 11852 2872 11880
rect 2547 11849 2559 11852
rect 2501 11843 2559 11849
rect 2866 11840 2872 11852
rect 2924 11840 2930 11892
rect 4157 11883 4215 11889
rect 4157 11849 4169 11883
rect 4203 11880 4215 11883
rect 4522 11880 4528 11892
rect 4203 11852 4528 11880
rect 4203 11849 4215 11852
rect 4157 11843 4215 11849
rect 4522 11840 4528 11852
rect 4580 11840 4586 11892
rect 4614 11840 4620 11892
rect 4672 11880 4678 11892
rect 5077 11883 5135 11889
rect 5077 11880 5089 11883
rect 4672 11852 5089 11880
rect 4672 11840 4678 11852
rect 5077 11849 5089 11852
rect 5123 11849 5135 11883
rect 5077 11843 5135 11849
rect 5350 11840 5356 11892
rect 5408 11880 5414 11892
rect 5813 11883 5871 11889
rect 5813 11880 5825 11883
rect 5408 11852 5825 11880
rect 5408 11840 5414 11852
rect 5813 11849 5825 11852
rect 5859 11849 5871 11883
rect 6178 11880 6184 11892
rect 6139 11852 6184 11880
rect 5813 11843 5871 11849
rect 6178 11840 6184 11852
rect 6236 11840 6242 11892
rect 6638 11880 6644 11892
rect 6599 11852 6644 11880
rect 6638 11840 6644 11852
rect 6696 11840 6702 11892
rect 6990 11883 7048 11889
rect 6990 11849 7002 11883
rect 7036 11880 7048 11883
rect 7282 11880 7288 11892
rect 7036 11852 7288 11880
rect 7036 11849 7048 11852
rect 6990 11843 7048 11849
rect 7282 11840 7288 11852
rect 7340 11840 7346 11892
rect 7374 11840 7380 11892
rect 7432 11880 7438 11892
rect 8205 11883 8263 11889
rect 8205 11880 8217 11883
rect 7432 11852 8217 11880
rect 7432 11840 7438 11852
rect 8205 11849 8217 11852
rect 8251 11849 8263 11883
rect 8205 11843 8263 11849
rect 4801 11815 4859 11821
rect 4801 11812 4813 11815
rect 4126 11784 4813 11812
rect 1946 11744 1952 11756
rect 1688 11716 1952 11744
rect 1688 11688 1716 11716
rect 1946 11704 1952 11716
rect 2004 11744 2010 11756
rect 4126 11744 4154 11784
rect 4801 11781 4813 11784
rect 4847 11781 4859 11815
rect 4801 11775 4859 11781
rect 5537 11815 5595 11821
rect 5537 11781 5549 11815
rect 5583 11812 5595 11815
rect 6454 11812 6460 11824
rect 5583 11784 6460 11812
rect 5583 11781 5595 11784
rect 5537 11775 5595 11781
rect 6454 11772 6460 11784
rect 6512 11772 6518 11824
rect 7098 11812 7104 11824
rect 7059 11784 7104 11812
rect 7098 11772 7104 11784
rect 7156 11772 7162 11824
rect 7558 11772 7564 11824
rect 7616 11812 7622 11824
rect 7837 11815 7895 11821
rect 7837 11812 7849 11815
rect 7616 11784 7849 11812
rect 7616 11772 7622 11784
rect 7837 11781 7849 11784
rect 7883 11781 7895 11815
rect 7837 11775 7895 11781
rect 2004 11716 3004 11744
rect 2004 11704 2010 11716
rect 1670 11676 1676 11688
rect 1583 11648 1676 11676
rect 1670 11636 1676 11648
rect 1728 11636 1734 11688
rect 1857 11679 1915 11685
rect 1857 11645 1869 11679
rect 1903 11676 1915 11679
rect 2314 11676 2320 11688
rect 1903 11648 2320 11676
rect 1903 11645 1915 11648
rect 1857 11639 1915 11645
rect 2314 11636 2320 11648
rect 2372 11676 2378 11688
rect 2774 11676 2780 11688
rect 2372 11648 2780 11676
rect 2372 11636 2378 11648
rect 2774 11636 2780 11648
rect 2832 11636 2838 11688
rect 2976 11685 3004 11716
rect 3344 11716 4154 11744
rect 6472 11744 6500 11772
rect 7193 11747 7251 11753
rect 7193 11744 7205 11747
rect 6472 11716 7205 11744
rect 3344 11685 3372 11716
rect 7193 11713 7205 11716
rect 7239 11713 7251 11747
rect 7193 11707 7251 11713
rect 2961 11679 3019 11685
rect 2961 11645 2973 11679
rect 3007 11676 3019 11679
rect 3329 11679 3387 11685
rect 3329 11676 3341 11679
rect 3007 11648 3341 11676
rect 3007 11645 3019 11648
rect 2961 11639 3019 11645
rect 3329 11645 3341 11648
rect 3375 11645 3387 11679
rect 3510 11676 3516 11688
rect 3471 11648 3516 11676
rect 3329 11639 3387 11645
rect 3510 11636 3516 11648
rect 3568 11636 3574 11688
rect 4617 11679 4675 11685
rect 4617 11676 4629 11679
rect 4540 11648 4629 11676
rect 14 11568 20 11620
rect 72 11608 78 11620
rect 72 11580 3004 11608
rect 72 11568 78 11580
rect 106 11500 112 11552
rect 164 11540 170 11552
rect 1489 11543 1547 11549
rect 1489 11540 1501 11543
rect 164 11512 1501 11540
rect 164 11500 170 11512
rect 1489 11509 1501 11512
rect 1535 11509 1547 11543
rect 2976 11540 3004 11580
rect 4540 11552 4568 11648
rect 4617 11645 4629 11648
rect 4663 11645 4675 11679
rect 4617 11639 4675 11645
rect 5629 11679 5687 11685
rect 5629 11645 5641 11679
rect 5675 11676 5687 11679
rect 5718 11676 5724 11688
rect 5675 11648 5724 11676
rect 5675 11645 5687 11648
rect 5629 11639 5687 11645
rect 5718 11636 5724 11648
rect 5776 11676 5782 11688
rect 6086 11676 6092 11688
rect 5776 11648 6092 11676
rect 5776 11636 5782 11648
rect 6086 11636 6092 11648
rect 6144 11636 6150 11688
rect 6638 11636 6644 11688
rect 6696 11676 6702 11688
rect 6825 11679 6883 11685
rect 6825 11676 6837 11679
rect 6696 11648 6837 11676
rect 6696 11636 6702 11648
rect 6825 11645 6837 11648
rect 6871 11645 6883 11679
rect 6825 11639 6883 11645
rect 7006 11636 7012 11688
rect 7064 11676 7070 11688
rect 8389 11679 8447 11685
rect 8389 11676 8401 11679
rect 7064 11648 8401 11676
rect 7064 11636 7070 11648
rect 8389 11645 8401 11648
rect 8435 11676 8447 11679
rect 8849 11679 8907 11685
rect 8849 11676 8861 11679
rect 8435 11648 8861 11676
rect 8435 11645 8447 11648
rect 8389 11639 8447 11645
rect 8849 11645 8861 11648
rect 8895 11645 8907 11679
rect 8849 11639 8907 11645
rect 4798 11568 4804 11620
rect 4856 11608 4862 11620
rect 4856 11580 7696 11608
rect 4856 11568 4862 11580
rect 3145 11543 3203 11549
rect 3145 11540 3157 11543
rect 2976 11512 3157 11540
rect 1489 11503 1547 11509
rect 3145 11509 3157 11512
rect 3191 11509 3203 11543
rect 4522 11540 4528 11552
rect 4483 11512 4528 11540
rect 3145 11503 3203 11509
rect 4522 11500 4528 11512
rect 4580 11500 4586 11552
rect 6914 11500 6920 11552
rect 6972 11540 6978 11552
rect 7469 11543 7527 11549
rect 7469 11540 7481 11543
rect 6972 11512 7481 11540
rect 6972 11500 6978 11512
rect 7469 11509 7481 11512
rect 7515 11509 7527 11543
rect 7668 11540 7696 11580
rect 8573 11543 8631 11549
rect 8573 11540 8585 11543
rect 7668 11512 8585 11540
rect 7469 11503 7527 11509
rect 8573 11509 8585 11512
rect 8619 11509 8631 11543
rect 8573 11503 8631 11509
rect 1104 11450 22816 11472
rect 1104 11398 8982 11450
rect 9034 11398 9046 11450
rect 9098 11398 9110 11450
rect 9162 11398 9174 11450
rect 9226 11398 16982 11450
rect 17034 11398 17046 11450
rect 17098 11398 17110 11450
rect 17162 11398 17174 11450
rect 17226 11398 22816 11450
rect 1104 11376 22816 11398
rect 106 11296 112 11348
rect 164 11336 170 11348
rect 1489 11339 1547 11345
rect 1489 11336 1501 11339
rect 164 11308 1501 11336
rect 164 11296 170 11308
rect 1489 11305 1501 11308
rect 1535 11305 1547 11339
rect 1489 11299 1547 11305
rect 2682 11296 2688 11348
rect 2740 11336 2746 11348
rect 2777 11339 2835 11345
rect 2777 11336 2789 11339
rect 2740 11308 2789 11336
rect 2740 11296 2746 11308
rect 2777 11305 2789 11308
rect 2823 11336 2835 11339
rect 3421 11339 3479 11345
rect 3421 11336 3433 11339
rect 2823 11308 3433 11336
rect 2823 11305 2835 11308
rect 2777 11299 2835 11305
rect 3421 11305 3433 11308
rect 3467 11336 3479 11339
rect 3605 11339 3663 11345
rect 3605 11336 3617 11339
rect 3467 11308 3617 11336
rect 3467 11305 3479 11308
rect 3421 11299 3479 11305
rect 3605 11305 3617 11308
rect 3651 11305 3663 11339
rect 3605 11299 3663 11305
rect 4522 11296 4528 11348
rect 4580 11336 4586 11348
rect 6365 11339 6423 11345
rect 6365 11336 6377 11339
rect 4580 11308 6377 11336
rect 4580 11296 4586 11308
rect 6365 11305 6377 11308
rect 6411 11305 6423 11339
rect 6365 11299 6423 11305
rect 6454 11296 6460 11348
rect 6512 11336 6518 11348
rect 6825 11339 6883 11345
rect 6825 11336 6837 11339
rect 6512 11308 6837 11336
rect 6512 11296 6518 11308
rect 6825 11305 6837 11308
rect 6871 11336 6883 11339
rect 7745 11339 7803 11345
rect 7745 11336 7757 11339
rect 6871 11308 7757 11336
rect 6871 11305 6883 11308
rect 6825 11299 6883 11305
rect 7745 11305 7757 11308
rect 7791 11305 7803 11339
rect 7745 11299 7803 11305
rect 7926 11296 7932 11348
rect 7984 11336 7990 11348
rect 8113 11339 8171 11345
rect 8113 11336 8125 11339
rect 7984 11308 8125 11336
rect 7984 11296 7990 11308
rect 8113 11305 8125 11308
rect 8159 11305 8171 11339
rect 8113 11299 8171 11305
rect 2700 11268 2728 11296
rect 1964 11240 2728 11268
rect 1670 11200 1676 11212
rect 1631 11172 1676 11200
rect 1670 11160 1676 11172
rect 1728 11160 1734 11212
rect 1964 11209 1992 11240
rect 3510 11228 3516 11280
rect 3568 11268 3574 11280
rect 3789 11271 3847 11277
rect 3789 11268 3801 11271
rect 3568 11240 3801 11268
rect 3568 11228 3574 11240
rect 3789 11237 3801 11240
rect 3835 11237 3847 11271
rect 3789 11231 3847 11237
rect 5261 11271 5319 11277
rect 5261 11237 5273 11271
rect 5307 11268 5319 11271
rect 5629 11271 5687 11277
rect 5629 11268 5641 11271
rect 5307 11240 5641 11268
rect 5307 11237 5319 11240
rect 5261 11231 5319 11237
rect 5629 11237 5641 11240
rect 5675 11268 5687 11271
rect 5718 11268 5724 11280
rect 5675 11240 5724 11268
rect 5675 11237 5687 11240
rect 5629 11231 5687 11237
rect 5718 11228 5724 11240
rect 5776 11228 5782 11280
rect 1949 11203 2007 11209
rect 1949 11169 1961 11203
rect 1995 11169 2007 11203
rect 1949 11163 2007 11169
rect 2501 11203 2559 11209
rect 2501 11169 2513 11203
rect 2547 11200 2559 11203
rect 2774 11200 2780 11212
rect 2547 11172 2780 11200
rect 2547 11169 2559 11172
rect 2501 11163 2559 11169
rect 2774 11160 2780 11172
rect 2832 11200 2838 11212
rect 2961 11203 3019 11209
rect 2961 11200 2973 11203
rect 2832 11172 2973 11200
rect 2832 11160 2838 11172
rect 2961 11169 2973 11172
rect 3007 11200 3019 11203
rect 4246 11200 4252 11212
rect 3007 11172 4252 11200
rect 3007 11169 3019 11172
rect 2961 11163 3019 11169
rect 4246 11160 4252 11172
rect 4304 11160 4310 11212
rect 4614 11200 4620 11212
rect 4575 11172 4620 11200
rect 4614 11160 4620 11172
rect 4672 11160 4678 11212
rect 5868 11203 5926 11209
rect 5868 11169 5880 11203
rect 5914 11200 5926 11203
rect 6178 11200 6184 11212
rect 5914 11172 6184 11200
rect 5914 11169 5926 11172
rect 5868 11163 5926 11169
rect 6178 11160 6184 11172
rect 6236 11200 6242 11212
rect 7190 11200 7196 11212
rect 6236 11172 7196 11200
rect 6236 11160 6242 11172
rect 7190 11160 7196 11172
rect 7248 11160 7254 11212
rect 7285 11203 7343 11209
rect 7285 11169 7297 11203
rect 7331 11200 7343 11203
rect 7466 11200 7472 11212
rect 7331 11172 7472 11200
rect 7331 11169 7343 11172
rect 7285 11163 7343 11169
rect 7466 11160 7472 11172
rect 7524 11160 7530 11212
rect 6086 11132 6092 11144
rect 5999 11104 6092 11132
rect 6086 11092 6092 11104
rect 6144 11132 6150 11144
rect 6454 11132 6460 11144
rect 6144 11104 6460 11132
rect 6144 11092 6150 11104
rect 6454 11092 6460 11104
rect 6512 11092 6518 11144
rect 3605 11067 3663 11073
rect 3605 11033 3617 11067
rect 3651 11064 3663 11067
rect 4154 11064 4160 11076
rect 3651 11036 4160 11064
rect 3651 11033 3663 11036
rect 3605 11027 3663 11033
rect 4154 11024 4160 11036
rect 4212 11064 4218 11076
rect 4801 11067 4859 11073
rect 4801 11064 4813 11067
rect 4212 11036 4813 11064
rect 4212 11024 4218 11036
rect 4801 11033 4813 11036
rect 4847 11064 4859 11067
rect 7006 11064 7012 11076
rect 4847 11036 7012 11064
rect 4847 11033 4859 11036
rect 4801 11027 4859 11033
rect 7006 11024 7012 11036
rect 7064 11024 7070 11076
rect 3142 10996 3148 11008
rect 3103 10968 3148 10996
rect 3142 10956 3148 10968
rect 3200 10956 3206 11008
rect 4246 10996 4252 11008
rect 4207 10968 4252 10996
rect 4246 10956 4252 10968
rect 4304 10956 4310 11008
rect 5997 10999 6055 11005
rect 5997 10965 6009 10999
rect 6043 10996 6055 10999
rect 6362 10996 6368 11008
rect 6043 10968 6368 10996
rect 6043 10965 6055 10968
rect 5997 10959 6055 10965
rect 6362 10956 6368 10968
rect 6420 10956 6426 11008
rect 7466 10996 7472 11008
rect 7427 10968 7472 10996
rect 7466 10956 7472 10968
rect 7524 10956 7530 11008
rect 1104 10906 22816 10928
rect 1104 10854 4982 10906
rect 5034 10854 5046 10906
rect 5098 10854 5110 10906
rect 5162 10854 5174 10906
rect 5226 10854 12982 10906
rect 13034 10854 13046 10906
rect 13098 10854 13110 10906
rect 13162 10854 13174 10906
rect 13226 10854 20982 10906
rect 21034 10854 21046 10906
rect 21098 10854 21110 10906
rect 21162 10854 21174 10906
rect 21226 10854 22816 10906
rect 1104 10832 22816 10854
rect 1670 10752 1676 10804
rect 1728 10792 1734 10804
rect 2409 10795 2467 10801
rect 2409 10792 2421 10795
rect 1728 10764 2421 10792
rect 1728 10752 1734 10764
rect 2409 10761 2421 10764
rect 2455 10761 2467 10795
rect 2774 10792 2780 10804
rect 2735 10764 2780 10792
rect 2409 10755 2467 10761
rect 2774 10752 2780 10764
rect 2832 10752 2838 10804
rect 4065 10795 4123 10801
rect 4065 10761 4077 10795
rect 4111 10792 4123 10795
rect 4154 10792 4160 10804
rect 4111 10764 4160 10792
rect 4111 10761 4123 10764
rect 4065 10755 4123 10761
rect 4154 10752 4160 10764
rect 4212 10752 4218 10804
rect 6086 10792 6092 10804
rect 6047 10764 6092 10792
rect 6086 10752 6092 10764
rect 6144 10752 6150 10804
rect 6362 10792 6368 10804
rect 6323 10764 6368 10792
rect 6362 10752 6368 10764
rect 6420 10752 6426 10804
rect 7282 10792 7288 10804
rect 7243 10764 7288 10792
rect 7282 10752 7288 10764
rect 7340 10752 7346 10804
rect 7558 10752 7564 10804
rect 7616 10792 7622 10804
rect 7653 10795 7711 10801
rect 7653 10792 7665 10795
rect 7616 10764 7665 10792
rect 7616 10752 7622 10764
rect 7653 10761 7665 10764
rect 7699 10761 7711 10795
rect 7653 10755 7711 10761
rect 2590 10684 2596 10736
rect 2648 10724 2654 10736
rect 4709 10727 4767 10733
rect 4709 10724 4721 10727
rect 2648 10696 4721 10724
rect 2648 10684 2654 10696
rect 4709 10693 4721 10696
rect 4755 10693 4767 10727
rect 7009 10727 7067 10733
rect 7009 10724 7021 10727
rect 4709 10687 4767 10693
rect 4908 10696 7021 10724
rect 198 10616 204 10668
rect 256 10656 262 10668
rect 2498 10656 2504 10668
rect 256 10628 2504 10656
rect 256 10616 262 10628
rect 2498 10616 2504 10628
rect 2556 10616 2562 10668
rect 3878 10656 3884 10668
rect 3252 10628 3884 10656
rect 1670 10588 1676 10600
rect 1631 10560 1676 10588
rect 1670 10548 1676 10560
rect 1728 10548 1734 10600
rect 1949 10591 2007 10597
rect 1949 10557 1961 10591
rect 1995 10588 2007 10591
rect 2314 10588 2320 10600
rect 1995 10560 2320 10588
rect 1995 10557 2007 10560
rect 1949 10551 2007 10557
rect 2314 10548 2320 10560
rect 2372 10588 2378 10600
rect 2866 10588 2872 10600
rect 2372 10560 2872 10588
rect 2372 10548 2378 10560
rect 2866 10548 2872 10560
rect 2924 10548 2930 10600
rect 3252 10597 3280 10628
rect 3878 10616 3884 10628
rect 3936 10656 3942 10668
rect 4522 10656 4528 10668
rect 3936 10628 4528 10656
rect 3936 10616 3942 10628
rect 4522 10616 4528 10628
rect 4580 10616 4586 10668
rect 3237 10591 3295 10597
rect 3237 10557 3249 10591
rect 3283 10557 3295 10591
rect 3237 10551 3295 10557
rect 3513 10591 3571 10597
rect 3513 10557 3525 10591
rect 3559 10588 3571 10591
rect 3786 10588 3792 10600
rect 3559 10560 3792 10588
rect 3559 10557 3571 10560
rect 3513 10551 3571 10557
rect 3786 10548 3792 10560
rect 3844 10588 3850 10600
rect 4908 10588 4936 10696
rect 7009 10693 7021 10696
rect 7055 10693 7067 10727
rect 7009 10687 7067 10693
rect 3844 10560 4936 10588
rect 5353 10591 5411 10597
rect 3844 10548 3850 10560
rect 5353 10557 5365 10591
rect 5399 10557 5411 10591
rect 5353 10551 5411 10557
rect 14 10480 20 10532
rect 72 10480 78 10532
rect 106 10480 112 10532
rect 164 10520 170 10532
rect 4982 10520 4988 10532
rect 164 10492 3004 10520
rect 4943 10492 4988 10520
rect 164 10480 170 10492
rect 32 10452 60 10480
rect 1489 10455 1547 10461
rect 1489 10452 1501 10455
rect 32 10424 1501 10452
rect 1489 10421 1501 10424
rect 1535 10421 1547 10455
rect 2976 10452 3004 10492
rect 4982 10480 4988 10492
rect 5040 10480 5046 10532
rect 5368 10464 5396 10551
rect 6730 10548 6736 10600
rect 6788 10588 6794 10600
rect 6825 10591 6883 10597
rect 6825 10588 6837 10591
rect 6788 10560 6837 10588
rect 6788 10548 6794 10560
rect 6825 10557 6837 10560
rect 6871 10588 6883 10591
rect 8021 10591 8079 10597
rect 8021 10588 8033 10591
rect 6871 10560 8033 10588
rect 6871 10557 6883 10560
rect 6825 10551 6883 10557
rect 8021 10557 8033 10560
rect 8067 10557 8079 10591
rect 8021 10551 8079 10557
rect 3053 10455 3111 10461
rect 3053 10452 3065 10455
rect 2976 10424 3065 10452
rect 1489 10415 1547 10421
rect 3053 10421 3065 10424
rect 3099 10421 3111 10455
rect 3053 10415 3111 10421
rect 4525 10455 4583 10461
rect 4525 10421 4537 10455
rect 4571 10452 4583 10455
rect 4614 10452 4620 10464
rect 4571 10424 4620 10452
rect 4571 10421 4583 10424
rect 4525 10415 4583 10421
rect 4614 10412 4620 10424
rect 4672 10412 4678 10464
rect 4709 10455 4767 10461
rect 4709 10421 4721 10455
rect 4755 10452 4767 10455
rect 4893 10455 4951 10461
rect 4893 10452 4905 10455
rect 4755 10424 4905 10452
rect 4755 10421 4767 10424
rect 4709 10415 4767 10421
rect 4893 10421 4905 10424
rect 4939 10452 4951 10455
rect 5350 10452 5356 10464
rect 4939 10424 5356 10452
rect 4939 10421 4951 10424
rect 4893 10415 4951 10421
rect 5350 10412 5356 10424
rect 5408 10412 5414 10464
rect 1104 10362 22816 10384
rect 1104 10310 8982 10362
rect 9034 10310 9046 10362
rect 9098 10310 9110 10362
rect 9162 10310 9174 10362
rect 9226 10310 16982 10362
rect 17034 10310 17046 10362
rect 17098 10310 17110 10362
rect 17162 10310 17174 10362
rect 17226 10310 22816 10362
rect 1104 10288 22816 10310
rect 1581 10251 1639 10257
rect 1581 10217 1593 10251
rect 1627 10217 1639 10251
rect 1581 10211 1639 10217
rect 1596 10180 1624 10211
rect 1670 10208 1676 10260
rect 1728 10248 1734 10260
rect 1857 10251 1915 10257
rect 1857 10248 1869 10251
rect 1728 10220 1869 10248
rect 1728 10208 1734 10220
rect 1857 10217 1869 10220
rect 1903 10217 1915 10251
rect 2314 10248 2320 10260
rect 2275 10220 2320 10248
rect 1857 10211 1915 10217
rect 2314 10208 2320 10220
rect 2372 10208 2378 10260
rect 2498 10248 2504 10260
rect 2459 10220 2504 10248
rect 2498 10208 2504 10220
rect 2556 10208 2562 10260
rect 3510 10208 3516 10260
rect 3568 10248 3574 10260
rect 3789 10251 3847 10257
rect 3789 10248 3801 10251
rect 3568 10220 3801 10248
rect 3568 10208 3574 10220
rect 3789 10217 3801 10220
rect 3835 10217 3847 10251
rect 4246 10248 4252 10260
rect 4207 10220 4252 10248
rect 3789 10211 3847 10217
rect 4246 10208 4252 10220
rect 4304 10208 4310 10260
rect 4522 10248 4528 10260
rect 4483 10220 4528 10248
rect 4522 10208 4528 10220
rect 4580 10208 4586 10260
rect 4982 10248 4988 10260
rect 4943 10220 4988 10248
rect 4982 10208 4988 10220
rect 5040 10208 5046 10260
rect 5718 10208 5724 10260
rect 5776 10248 5782 10260
rect 6457 10251 6515 10257
rect 6457 10248 6469 10251
rect 5776 10220 6469 10248
rect 5776 10208 5782 10220
rect 6457 10217 6469 10220
rect 6503 10217 6515 10251
rect 6457 10211 6515 10217
rect 2332 10180 2360 10208
rect 1596 10152 2360 10180
rect 1394 10112 1400 10124
rect 1355 10084 1400 10112
rect 1394 10072 1400 10084
rect 1452 10072 1458 10124
rect 2685 10115 2743 10121
rect 2685 10081 2697 10115
rect 2731 10081 2743 10115
rect 2685 10075 2743 10081
rect 2961 10115 3019 10121
rect 2961 10081 2973 10115
rect 3007 10112 3019 10115
rect 3528 10112 3556 10208
rect 4154 10140 4160 10192
rect 4212 10180 4218 10192
rect 5000 10180 5028 10208
rect 5994 10180 6000 10192
rect 4212 10152 5028 10180
rect 5092 10152 6000 10180
rect 4212 10140 4218 10152
rect 3007 10084 3556 10112
rect 4065 10115 4123 10121
rect 3007 10081 3019 10084
rect 2961 10075 3019 10081
rect 4065 10081 4077 10115
rect 4111 10081 4123 10115
rect 4065 10075 4123 10081
rect 2700 10044 2728 10075
rect 3513 10047 3571 10053
rect 3513 10044 3525 10047
rect 2700 10016 3525 10044
rect 3513 10013 3525 10016
rect 3559 10044 3571 10047
rect 3786 10044 3792 10056
rect 3559 10016 3792 10044
rect 3559 10013 3571 10016
rect 3513 10007 3571 10013
rect 3786 10004 3792 10016
rect 3844 10004 3850 10056
rect 4080 10044 4108 10075
rect 4706 10072 4712 10124
rect 4764 10112 4770 10124
rect 5092 10121 5120 10152
rect 5994 10140 6000 10152
rect 6052 10140 6058 10192
rect 6178 10180 6184 10192
rect 6139 10152 6184 10180
rect 6178 10140 6184 10152
rect 6236 10140 6242 10192
rect 5077 10115 5135 10121
rect 5077 10112 5089 10115
rect 4764 10084 5089 10112
rect 4764 10072 4770 10084
rect 5077 10081 5089 10084
rect 5123 10081 5135 10115
rect 5077 10075 5135 10081
rect 5353 10115 5411 10121
rect 5353 10081 5365 10115
rect 5399 10112 5411 10115
rect 5718 10112 5724 10124
rect 5399 10084 5724 10112
rect 5399 10081 5411 10084
rect 5353 10075 5411 10081
rect 5718 10072 5724 10084
rect 5776 10072 5782 10124
rect 6638 10112 6644 10124
rect 6599 10084 6644 10112
rect 6638 10072 6644 10084
rect 6696 10072 6702 10124
rect 6917 10115 6975 10121
rect 6917 10081 6929 10115
rect 6963 10112 6975 10115
rect 7282 10112 7288 10124
rect 6963 10084 7288 10112
rect 6963 10081 6975 10084
rect 6917 10075 6975 10081
rect 7282 10072 7288 10084
rect 7340 10072 7346 10124
rect 4043 10016 4154 10044
rect 4126 9908 4154 10016
rect 4614 10004 4620 10056
rect 4672 10044 4678 10056
rect 5537 10047 5595 10053
rect 5537 10044 5549 10047
rect 4672 10016 5549 10044
rect 4672 10004 4678 10016
rect 5537 10013 5549 10016
rect 5583 10013 5595 10047
rect 7101 10047 7159 10053
rect 7101 10044 7113 10047
rect 5537 10007 5595 10013
rect 5736 10016 7113 10044
rect 4522 9936 4528 9988
rect 4580 9976 4586 9988
rect 4798 9976 4804 9988
rect 4580 9948 4804 9976
rect 4580 9936 4586 9948
rect 4798 9936 4804 9948
rect 4856 9936 4862 9988
rect 5169 9979 5227 9985
rect 5169 9945 5181 9979
rect 5215 9976 5227 9979
rect 5350 9976 5356 9988
rect 5215 9948 5356 9976
rect 5215 9945 5227 9948
rect 5169 9939 5227 9945
rect 5350 9936 5356 9948
rect 5408 9936 5414 9988
rect 4246 9908 4252 9920
rect 4126 9880 4252 9908
rect 4246 9868 4252 9880
rect 4304 9908 4310 9920
rect 5736 9908 5764 10016
rect 7101 10013 7113 10016
rect 7147 10013 7159 10047
rect 7101 10007 7159 10013
rect 6730 9976 6736 9988
rect 6691 9948 6736 9976
rect 6730 9936 6736 9948
rect 6788 9936 6794 9988
rect 4304 9880 5764 9908
rect 4304 9868 4310 9880
rect 1104 9818 22816 9840
rect 1104 9766 4982 9818
rect 5034 9766 5046 9818
rect 5098 9766 5110 9818
rect 5162 9766 5174 9818
rect 5226 9766 12982 9818
rect 13034 9766 13046 9818
rect 13098 9766 13110 9818
rect 13162 9766 13174 9818
rect 13226 9766 20982 9818
rect 21034 9766 21046 9818
rect 21098 9766 21110 9818
rect 21162 9766 21174 9818
rect 21226 9766 22816 9818
rect 1104 9744 22816 9766
rect 1394 9664 1400 9716
rect 1452 9704 1458 9716
rect 2682 9704 2688 9716
rect 1452 9676 2688 9704
rect 1452 9664 1458 9676
rect 2682 9664 2688 9676
rect 2740 9664 2746 9716
rect 4617 9707 4675 9713
rect 4617 9673 4629 9707
rect 4663 9704 4675 9707
rect 4706 9704 4712 9716
rect 4663 9676 4712 9704
rect 4663 9673 4675 9676
rect 4617 9667 4675 9673
rect 4706 9664 4712 9676
rect 4764 9664 4770 9716
rect 4985 9707 5043 9713
rect 4985 9673 4997 9707
rect 5031 9704 5043 9707
rect 5350 9704 5356 9716
rect 5031 9676 5356 9704
rect 5031 9673 5043 9676
rect 4985 9667 5043 9673
rect 5350 9664 5356 9676
rect 5408 9704 5414 9716
rect 6730 9704 6736 9716
rect 5408 9676 6736 9704
rect 5408 9664 5414 9676
rect 6730 9664 6736 9676
rect 6788 9704 6794 9716
rect 7009 9707 7067 9713
rect 7009 9704 7021 9707
rect 6788 9676 7021 9704
rect 6788 9664 6794 9676
rect 7009 9673 7021 9676
rect 7055 9673 7067 9707
rect 7009 9667 7067 9673
rect 1578 9596 1584 9648
rect 1636 9636 1642 9648
rect 2961 9639 3019 9645
rect 2961 9636 2973 9639
rect 1636 9608 2973 9636
rect 1636 9596 1642 9608
rect 2961 9605 2973 9608
rect 3007 9605 3019 9639
rect 2961 9599 3019 9605
rect 4062 9596 4068 9648
rect 4120 9636 4126 9648
rect 5166 9636 5172 9648
rect 4120 9608 5172 9636
rect 4120 9596 4126 9608
rect 5166 9596 5172 9608
rect 5224 9596 5230 9648
rect 3050 9568 3056 9580
rect 2240 9540 3056 9568
rect 2240 9509 2268 9540
rect 3050 9528 3056 9540
rect 3108 9568 3114 9580
rect 3145 9571 3203 9577
rect 3145 9568 3157 9571
rect 3108 9540 3157 9568
rect 3108 9528 3114 9540
rect 3145 9537 3157 9540
rect 3191 9568 3203 9571
rect 6638 9568 6644 9580
rect 3191 9540 3832 9568
rect 3191 9537 3203 9540
rect 3145 9531 3203 9537
rect 3804 9512 3832 9540
rect 5092 9540 6644 9568
rect 5092 9512 5120 9540
rect 6638 9528 6644 9540
rect 6696 9528 6702 9580
rect 1949 9503 2007 9509
rect 1949 9469 1961 9503
rect 1995 9469 2007 9503
rect 1949 9463 2007 9469
rect 2225 9503 2283 9509
rect 2225 9469 2237 9503
rect 2271 9469 2283 9503
rect 2225 9463 2283 9469
rect 2961 9503 3019 9509
rect 2961 9469 2973 9503
rect 3007 9500 3019 9503
rect 3237 9503 3295 9509
rect 3237 9500 3249 9503
rect 3007 9472 3249 9500
rect 3007 9469 3019 9472
rect 2961 9463 3019 9469
rect 3237 9469 3249 9472
rect 3283 9469 3295 9503
rect 3786 9500 3792 9512
rect 3747 9472 3792 9500
rect 3237 9463 3295 9469
rect 1854 9392 1860 9444
rect 1912 9432 1918 9444
rect 1964 9432 1992 9463
rect 3786 9460 3792 9472
rect 3844 9460 3850 9512
rect 5074 9500 5080 9512
rect 4987 9472 5080 9500
rect 5074 9460 5080 9472
rect 5132 9460 5138 9512
rect 5166 9460 5172 9512
rect 5224 9500 5230 9512
rect 5353 9503 5411 9509
rect 5224 9472 5269 9500
rect 5224 9460 5230 9472
rect 5353 9469 5365 9503
rect 5399 9500 5411 9503
rect 5718 9500 5724 9512
rect 5399 9472 5724 9500
rect 5399 9469 5411 9472
rect 5353 9463 5411 9469
rect 5718 9460 5724 9472
rect 5776 9500 5782 9512
rect 5776 9472 6224 9500
rect 5776 9460 5782 9472
rect 3142 9432 3148 9444
rect 1912 9404 3148 9432
rect 1912 9392 1918 9404
rect 3142 9392 3148 9404
rect 3200 9392 3206 9444
rect 106 9324 112 9376
rect 164 9364 170 9376
rect 1765 9367 1823 9373
rect 1765 9364 1777 9367
rect 164 9336 1777 9364
rect 164 9324 170 9336
rect 1765 9333 1777 9336
rect 1811 9333 1823 9367
rect 3326 9364 3332 9376
rect 3287 9336 3332 9364
rect 1765 9327 1823 9333
rect 3326 9324 3332 9336
rect 3384 9324 3390 9376
rect 4982 9324 4988 9376
rect 5040 9364 5046 9376
rect 6196 9373 6224 9472
rect 5537 9367 5595 9373
rect 5537 9364 5549 9367
rect 5040 9336 5549 9364
rect 5040 9324 5046 9336
rect 5537 9333 5549 9336
rect 5583 9333 5595 9367
rect 5537 9327 5595 9333
rect 6181 9367 6239 9373
rect 6181 9333 6193 9367
rect 6227 9364 6239 9367
rect 6549 9367 6607 9373
rect 6549 9364 6561 9367
rect 6227 9336 6561 9364
rect 6227 9333 6239 9336
rect 6181 9327 6239 9333
rect 6549 9333 6561 9336
rect 6595 9364 6607 9367
rect 7282 9364 7288 9376
rect 6595 9336 7288 9364
rect 6595 9333 6607 9336
rect 6549 9327 6607 9333
rect 7282 9324 7288 9336
rect 7340 9364 7346 9376
rect 7377 9367 7435 9373
rect 7377 9364 7389 9367
rect 7340 9336 7389 9364
rect 7340 9324 7346 9336
rect 7377 9333 7389 9336
rect 7423 9333 7435 9367
rect 7377 9327 7435 9333
rect 1104 9274 22816 9296
rect 1104 9222 8982 9274
rect 9034 9222 9046 9274
rect 9098 9222 9110 9274
rect 9162 9222 9174 9274
rect 9226 9222 16982 9274
rect 17034 9222 17046 9274
rect 17098 9222 17110 9274
rect 17162 9222 17174 9274
rect 17226 9222 22816 9274
rect 1104 9200 22816 9222
rect 106 9120 112 9172
rect 164 9160 170 9172
rect 1673 9163 1731 9169
rect 1673 9160 1685 9163
rect 164 9132 1685 9160
rect 164 9120 170 9132
rect 1673 9129 1685 9132
rect 1719 9129 1731 9163
rect 1673 9123 1731 9129
rect 2593 9163 2651 9169
rect 2593 9129 2605 9163
rect 2639 9160 2651 9163
rect 3050 9160 3056 9172
rect 2639 9132 3056 9160
rect 2639 9129 2651 9132
rect 2593 9123 2651 9129
rect 3050 9120 3056 9132
rect 3108 9120 3114 9172
rect 3142 9120 3148 9172
rect 3200 9160 3206 9172
rect 3697 9163 3755 9169
rect 3697 9160 3709 9163
rect 3200 9132 3709 9160
rect 3200 9120 3206 9132
rect 3697 9129 3709 9132
rect 3743 9129 3755 9163
rect 3697 9123 3755 9129
rect 3881 9163 3939 9169
rect 3881 9129 3893 9163
rect 3927 9160 3939 9163
rect 4249 9163 4307 9169
rect 4249 9160 4261 9163
rect 3927 9132 4261 9160
rect 3927 9129 3939 9132
rect 3881 9123 3939 9129
rect 4249 9129 4261 9132
rect 4295 9160 4307 9163
rect 4706 9160 4712 9172
rect 4295 9132 4712 9160
rect 4295 9129 4307 9132
rect 4249 9123 4307 9129
rect 4706 9120 4712 9132
rect 4764 9120 4770 9172
rect 5629 9163 5687 9169
rect 5629 9160 5641 9163
rect 4816 9132 5641 9160
rect 2682 9052 2688 9104
rect 2740 9092 2746 9104
rect 4816 9092 4844 9132
rect 5629 9129 5641 9132
rect 5675 9129 5687 9163
rect 6638 9160 6644 9172
rect 6599 9132 6644 9160
rect 5629 9123 5687 9129
rect 6638 9120 6644 9132
rect 6696 9120 6702 9172
rect 5074 9092 5080 9104
rect 2740 9064 4844 9092
rect 5035 9064 5080 9092
rect 2740 9052 2746 9064
rect 5074 9052 5080 9064
rect 5132 9092 5138 9104
rect 5350 9092 5356 9104
rect 5132 9064 5356 9092
rect 5132 9052 5138 9064
rect 5350 9052 5356 9064
rect 5408 9052 5414 9104
rect 1854 9024 1860 9036
rect 1815 8996 1860 9024
rect 1854 8984 1860 8996
rect 1912 8984 1918 9036
rect 2038 9024 2044 9036
rect 1999 8996 2044 9024
rect 2038 8984 2044 8996
rect 2096 8984 2102 9036
rect 3421 9027 3479 9033
rect 3421 8993 3433 9027
rect 3467 9024 3479 9027
rect 3510 9024 3516 9036
rect 3467 8996 3516 9024
rect 3467 8993 3479 8996
rect 3421 8987 3479 8993
rect 3510 8984 3516 8996
rect 3568 9024 3574 9036
rect 3881 9027 3939 9033
rect 3881 9024 3893 9027
rect 3568 8996 3893 9024
rect 3568 8984 3574 8996
rect 3881 8993 3893 8996
rect 3927 8993 3939 9027
rect 3881 8987 3939 8993
rect 4065 9027 4123 9033
rect 4065 8993 4077 9027
rect 4111 9024 4123 9027
rect 4614 9024 4620 9036
rect 4111 8996 4620 9024
rect 4111 8993 4123 8996
rect 4065 8987 4123 8993
rect 4614 8984 4620 8996
rect 4672 9024 4678 9036
rect 4982 9024 4988 9036
rect 4672 8996 4988 9024
rect 4672 8984 4678 8996
rect 4982 8984 4988 8996
rect 5040 8984 5046 9036
rect 5169 9027 5227 9033
rect 5169 8993 5181 9027
rect 5215 8993 5227 9027
rect 5169 8987 5227 8993
rect 5445 9027 5503 9033
rect 5445 8993 5457 9027
rect 5491 9024 5503 9027
rect 5718 9024 5724 9036
rect 5491 8996 5724 9024
rect 5491 8993 5503 8996
rect 5445 8987 5503 8993
rect 4246 8916 4252 8968
rect 4304 8956 4310 8968
rect 4525 8959 4583 8965
rect 4525 8956 4537 8959
rect 4304 8928 4537 8956
rect 4304 8916 4310 8928
rect 4525 8925 4537 8928
rect 4571 8925 4583 8959
rect 4525 8919 4583 8925
rect 4798 8916 4804 8968
rect 4856 8956 4862 8968
rect 5184 8956 5212 8987
rect 5718 8984 5724 8996
rect 5776 8984 5782 9036
rect 4856 8928 5212 8956
rect 4856 8916 4862 8928
rect 5166 8848 5172 8900
rect 5224 8888 5230 8900
rect 5261 8891 5319 8897
rect 5261 8888 5273 8891
rect 5224 8860 5273 8888
rect 5224 8848 5230 8860
rect 5261 8857 5273 8860
rect 5307 8888 5319 8891
rect 5534 8888 5540 8900
rect 5307 8860 5540 8888
rect 5307 8857 5319 8860
rect 5261 8851 5319 8857
rect 5534 8848 5540 8860
rect 5592 8848 5598 8900
rect 1104 8730 22816 8752
rect 1104 8678 4982 8730
rect 5034 8678 5046 8730
rect 5098 8678 5110 8730
rect 5162 8678 5174 8730
rect 5226 8678 12982 8730
rect 13034 8678 13046 8730
rect 13098 8678 13110 8730
rect 13162 8678 13174 8730
rect 13226 8678 20982 8730
rect 21034 8678 21046 8730
rect 21098 8678 21110 8730
rect 21162 8678 21174 8730
rect 21226 8678 22816 8730
rect 1104 8656 22816 8678
rect 4798 8616 4804 8628
rect 4759 8588 4804 8616
rect 4798 8576 4804 8588
rect 4856 8576 4862 8628
rect 5350 8616 5356 8628
rect 5311 8588 5356 8616
rect 5350 8576 5356 8588
rect 5408 8576 5414 8628
rect 4433 8551 4491 8557
rect 4433 8517 4445 8551
rect 4479 8548 4491 8551
rect 5718 8548 5724 8560
rect 4479 8520 5724 8548
rect 4479 8517 4491 8520
rect 4433 8511 4491 8517
rect 5718 8508 5724 8520
rect 5776 8508 5782 8560
rect 2866 8480 2872 8492
rect 1780 8452 2872 8480
rect 1780 8421 1808 8452
rect 2866 8440 2872 8452
rect 2924 8440 2930 8492
rect 4798 8440 4804 8492
rect 4856 8480 4862 8492
rect 5905 8483 5963 8489
rect 5905 8480 5917 8483
rect 4856 8452 5917 8480
rect 4856 8440 4862 8452
rect 1765 8415 1823 8421
rect 1765 8381 1777 8415
rect 1811 8381 1823 8415
rect 2038 8412 2044 8424
rect 1951 8384 2044 8412
rect 1765 8375 1823 8381
rect 2038 8372 2044 8384
rect 2096 8412 2102 8424
rect 2593 8415 2651 8421
rect 2593 8412 2605 8415
rect 2096 8384 2605 8412
rect 2096 8372 2102 8384
rect 2593 8381 2605 8384
rect 2639 8412 2651 8415
rect 2961 8415 3019 8421
rect 2961 8412 2973 8415
rect 2639 8384 2973 8412
rect 2639 8381 2651 8384
rect 2593 8375 2651 8381
rect 2961 8381 2973 8384
rect 3007 8412 3019 8415
rect 3602 8412 3608 8424
rect 3007 8384 3096 8412
rect 3563 8384 3608 8412
rect 3007 8381 3019 8384
rect 2961 8375 3019 8381
rect 14 8304 20 8356
rect 72 8344 78 8356
rect 3068 8344 3096 8384
rect 3602 8372 3608 8384
rect 3660 8372 3666 8424
rect 5184 8421 5212 8452
rect 5905 8449 5917 8452
rect 5951 8449 5963 8483
rect 5905 8443 5963 8449
rect 3881 8415 3939 8421
rect 3881 8381 3893 8415
rect 3927 8381 3939 8415
rect 5169 8415 5227 8421
rect 5169 8412 5181 8415
rect 5147 8384 5181 8412
rect 3881 8375 3939 8381
rect 5169 8381 5181 8384
rect 5215 8381 5227 8415
rect 5169 8375 5227 8381
rect 3510 8344 3516 8356
rect 72 8316 3004 8344
rect 3068 8316 3516 8344
rect 72 8304 78 8316
rect 106 8236 112 8288
rect 164 8276 170 8288
rect 1581 8279 1639 8285
rect 1581 8276 1593 8279
rect 164 8248 1593 8276
rect 164 8236 170 8248
rect 1581 8245 1593 8248
rect 1627 8245 1639 8279
rect 2976 8276 3004 8316
rect 3510 8304 3516 8316
rect 3568 8344 3574 8356
rect 3896 8344 3924 8375
rect 6178 8344 6184 8356
rect 3568 8316 6184 8344
rect 3568 8304 3574 8316
rect 6178 8304 6184 8316
rect 6236 8304 6242 8356
rect 3421 8279 3479 8285
rect 3421 8276 3433 8279
rect 2976 8248 3433 8276
rect 1581 8239 1639 8245
rect 3421 8245 3433 8248
rect 3467 8245 3479 8279
rect 3421 8239 3479 8245
rect 3602 8236 3608 8288
rect 3660 8276 3666 8288
rect 3970 8276 3976 8288
rect 3660 8248 3976 8276
rect 3660 8236 3666 8248
rect 3970 8236 3976 8248
rect 4028 8276 4034 8288
rect 5258 8276 5264 8288
rect 4028 8248 5264 8276
rect 4028 8236 4034 8248
rect 5258 8236 5264 8248
rect 5316 8276 5322 8288
rect 6273 8279 6331 8285
rect 6273 8276 6285 8279
rect 5316 8248 6285 8276
rect 5316 8236 5322 8248
rect 6273 8245 6285 8248
rect 6319 8245 6331 8279
rect 6273 8239 6331 8245
rect 1104 8186 22816 8208
rect 1104 8134 8982 8186
rect 9034 8134 9046 8186
rect 9098 8134 9110 8186
rect 9162 8134 9174 8186
rect 9226 8134 16982 8186
rect 17034 8134 17046 8186
rect 17098 8134 17110 8186
rect 17162 8134 17174 8186
rect 17226 8134 22816 8186
rect 1104 8112 22816 8134
rect 106 8032 112 8084
rect 164 8072 170 8084
rect 1581 8075 1639 8081
rect 1581 8072 1593 8075
rect 164 8044 1593 8072
rect 164 8032 170 8044
rect 1581 8041 1593 8044
rect 1627 8041 1639 8075
rect 1581 8035 1639 8041
rect 1854 8032 1860 8084
rect 1912 8072 1918 8084
rect 2501 8075 2559 8081
rect 2501 8072 2513 8075
rect 1912 8044 2513 8072
rect 1912 8032 1918 8044
rect 2501 8041 2513 8044
rect 2547 8041 2559 8075
rect 2501 8035 2559 8041
rect 3421 8075 3479 8081
rect 3421 8041 3433 8075
rect 3467 8072 3479 8075
rect 3510 8072 3516 8084
rect 3467 8044 3516 8072
rect 3467 8041 3479 8044
rect 3421 8035 3479 8041
rect 3510 8032 3516 8044
rect 3568 8032 3574 8084
rect 5258 8072 5264 8084
rect 5219 8044 5264 8072
rect 5258 8032 5264 8044
rect 5316 8032 5322 8084
rect 3605 8007 3663 8013
rect 3605 7973 3617 8007
rect 3651 8004 3663 8007
rect 4893 8007 4951 8013
rect 4893 8004 4905 8007
rect 3651 7976 4905 8004
rect 3651 7973 3663 7976
rect 3605 7967 3663 7973
rect 4893 7973 4905 7976
rect 4939 7973 4951 8007
rect 5534 8004 5540 8016
rect 5495 7976 5540 8004
rect 4893 7967 4951 7973
rect 5534 7964 5540 7976
rect 5592 7964 5598 8016
rect 1578 7936 1584 7948
rect 1539 7908 1584 7936
rect 1578 7896 1584 7908
rect 1636 7896 1642 7948
rect 2038 7936 2044 7948
rect 1999 7908 2044 7936
rect 2038 7896 2044 7908
rect 2096 7896 2102 7948
rect 2314 7896 2320 7948
rect 2372 7936 2378 7948
rect 4065 7939 4123 7945
rect 4065 7936 4077 7939
rect 2372 7908 4077 7936
rect 2372 7896 2378 7908
rect 4065 7905 4077 7908
rect 4111 7936 4123 7939
rect 4338 7936 4344 7948
rect 4111 7908 4344 7936
rect 4111 7905 4123 7908
rect 4065 7899 4123 7905
rect 4338 7896 4344 7908
rect 4396 7896 4402 7948
rect 4614 7936 4620 7948
rect 4575 7908 4620 7936
rect 4614 7896 4620 7908
rect 4672 7896 4678 7948
rect 4706 7896 4712 7948
rect 4764 7936 4770 7948
rect 5077 7939 5135 7945
rect 5077 7936 5089 7939
rect 4764 7908 5089 7936
rect 4764 7896 4770 7908
rect 5077 7905 5089 7908
rect 5123 7905 5135 7939
rect 6086 7936 6092 7948
rect 5999 7908 6092 7936
rect 5077 7899 5135 7905
rect 6086 7896 6092 7908
rect 6144 7936 6150 7948
rect 6914 7936 6920 7948
rect 6144 7908 6920 7936
rect 6144 7896 6150 7908
rect 6914 7896 6920 7908
rect 6972 7896 6978 7948
rect 1596 7868 1624 7896
rect 3605 7871 3663 7877
rect 3605 7868 3617 7871
rect 1596 7840 3617 7868
rect 3605 7837 3617 7840
rect 3651 7868 3663 7871
rect 3697 7871 3755 7877
rect 3697 7868 3709 7871
rect 3651 7840 3709 7868
rect 3651 7837 3663 7840
rect 3605 7831 3663 7837
rect 3697 7837 3709 7840
rect 3743 7837 3755 7871
rect 3697 7831 3755 7837
rect 2866 7760 2872 7812
rect 2924 7800 2930 7812
rect 2961 7803 3019 7809
rect 2961 7800 2973 7803
rect 2924 7772 2973 7800
rect 2924 7760 2930 7772
rect 2961 7769 2973 7772
rect 3007 7800 3019 7803
rect 3878 7800 3884 7812
rect 3007 7772 3884 7800
rect 3007 7769 3019 7772
rect 2961 7763 3019 7769
rect 3878 7760 3884 7772
rect 3936 7800 3942 7812
rect 4249 7803 4307 7809
rect 4249 7800 4261 7803
rect 3936 7772 4261 7800
rect 3936 7760 3942 7772
rect 4249 7769 4261 7772
rect 4295 7769 4307 7803
rect 4249 7763 4307 7769
rect 6178 7760 6184 7812
rect 6236 7800 6242 7812
rect 6273 7803 6331 7809
rect 6273 7800 6285 7803
rect 6236 7772 6285 7800
rect 6236 7760 6242 7772
rect 6273 7769 6285 7772
rect 6319 7769 6331 7803
rect 6273 7763 6331 7769
rect 1104 7642 22816 7664
rect 1104 7590 4982 7642
rect 5034 7590 5046 7642
rect 5098 7590 5110 7642
rect 5162 7590 5174 7642
rect 5226 7590 12982 7642
rect 13034 7590 13046 7642
rect 13098 7590 13110 7642
rect 13162 7590 13174 7642
rect 13226 7590 20982 7642
rect 21034 7590 21046 7642
rect 21098 7590 21110 7642
rect 21162 7590 21174 7642
rect 21226 7590 22816 7642
rect 1104 7568 22816 7590
rect 2038 7488 2044 7540
rect 2096 7528 2102 7540
rect 2501 7531 2559 7537
rect 2501 7528 2513 7531
rect 2096 7500 2513 7528
rect 2096 7488 2102 7500
rect 2501 7497 2513 7500
rect 2547 7497 2559 7531
rect 4338 7528 4344 7540
rect 4299 7500 4344 7528
rect 2501 7491 2559 7497
rect 4338 7488 4344 7500
rect 4396 7488 4402 7540
rect 4706 7488 4712 7540
rect 4764 7528 4770 7540
rect 4893 7531 4951 7537
rect 4893 7528 4905 7531
rect 4764 7500 4905 7528
rect 4764 7488 4770 7500
rect 4893 7497 4905 7500
rect 4939 7497 4951 7531
rect 6086 7528 6092 7540
rect 6047 7500 6092 7528
rect 4893 7491 4951 7497
rect 6086 7488 6092 7500
rect 6144 7488 6150 7540
rect 7282 7528 7288 7540
rect 7243 7500 7288 7528
rect 7282 7488 7288 7500
rect 7340 7488 7346 7540
rect 5353 7463 5411 7469
rect 5353 7429 5365 7463
rect 5399 7460 5411 7463
rect 8018 7460 8024 7472
rect 5399 7432 8024 7460
rect 5399 7429 5411 7432
rect 5353 7423 5411 7429
rect 1765 7327 1823 7333
rect 1765 7293 1777 7327
rect 1811 7324 1823 7327
rect 1854 7324 1860 7336
rect 1811 7296 1860 7324
rect 1811 7293 1823 7296
rect 1765 7287 1823 7293
rect 1854 7284 1860 7296
rect 1912 7284 1918 7336
rect 1946 7284 1952 7336
rect 2004 7324 2010 7336
rect 2041 7327 2099 7333
rect 2041 7324 2053 7327
rect 2004 7296 2053 7324
rect 2004 7284 2010 7296
rect 2041 7293 2053 7296
rect 2087 7324 2099 7327
rect 3605 7327 3663 7333
rect 2087 7296 3004 7324
rect 2087 7293 2099 7296
rect 2041 7287 2099 7293
rect 2976 7265 3004 7296
rect 3605 7293 3617 7327
rect 3651 7324 3663 7327
rect 3694 7324 3700 7336
rect 3651 7296 3700 7324
rect 3651 7293 3663 7296
rect 3605 7287 3663 7293
rect 3694 7284 3700 7296
rect 3752 7284 3758 7336
rect 3878 7324 3884 7336
rect 3839 7296 3884 7324
rect 3878 7284 3884 7296
rect 3936 7284 3942 7336
rect 5460 7333 5488 7432
rect 8018 7420 8024 7432
rect 8076 7420 8082 7472
rect 5445 7327 5503 7333
rect 5445 7293 5457 7327
rect 5491 7293 5503 7327
rect 5445 7287 5503 7293
rect 6641 7327 6699 7333
rect 6641 7293 6653 7327
rect 6687 7324 6699 7327
rect 7469 7327 7527 7333
rect 7469 7324 7481 7327
rect 6687 7296 7481 7324
rect 6687 7293 6699 7296
rect 6641 7287 6699 7293
rect 7469 7293 7481 7296
rect 7515 7324 7527 7327
rect 12066 7324 12072 7336
rect 7515 7296 12072 7324
rect 7515 7293 7527 7296
rect 7469 7287 7527 7293
rect 12066 7284 12072 7296
rect 12124 7284 12130 7336
rect 2961 7259 3019 7265
rect 2961 7225 2973 7259
rect 3007 7256 3019 7259
rect 3007 7228 3648 7256
rect 3007 7225 3019 7228
rect 2961 7219 3019 7225
rect 3620 7200 3648 7228
rect 1578 7188 1584 7200
rect 1539 7160 1584 7188
rect 1578 7148 1584 7160
rect 1636 7148 1642 7200
rect 3418 7188 3424 7200
rect 3379 7160 3424 7188
rect 3418 7148 3424 7160
rect 3476 7148 3482 7200
rect 3602 7148 3608 7200
rect 3660 7188 3666 7200
rect 5629 7191 5687 7197
rect 5629 7188 5641 7191
rect 3660 7160 5641 7188
rect 3660 7148 3666 7160
rect 5629 7157 5641 7160
rect 5675 7157 5687 7191
rect 5629 7151 5687 7157
rect 1104 7098 22816 7120
rect 1104 7046 8982 7098
rect 9034 7046 9046 7098
rect 9098 7046 9110 7098
rect 9162 7046 9174 7098
rect 9226 7046 16982 7098
rect 17034 7046 17046 7098
rect 17098 7046 17110 7098
rect 17162 7046 17174 7098
rect 17226 7046 22816 7098
rect 1104 7024 22816 7046
rect 106 6944 112 6996
rect 164 6984 170 6996
rect 1489 6987 1547 6993
rect 1489 6984 1501 6987
rect 164 6956 1501 6984
rect 164 6944 170 6956
rect 1489 6953 1501 6956
rect 1535 6953 1547 6987
rect 1489 6947 1547 6953
rect 1854 6944 1860 6996
rect 1912 6984 1918 6996
rect 2409 6987 2467 6993
rect 2409 6984 2421 6987
rect 1912 6956 2421 6984
rect 1912 6944 1918 6956
rect 2409 6953 2421 6956
rect 2455 6984 2467 6987
rect 3050 6984 3056 6996
rect 2455 6956 3056 6984
rect 2455 6953 2467 6956
rect 2409 6947 2467 6953
rect 3050 6944 3056 6956
rect 3108 6944 3114 6996
rect 3694 6984 3700 6996
rect 3655 6956 3700 6984
rect 3694 6944 3700 6956
rect 3752 6944 3758 6996
rect 4157 6987 4215 6993
rect 4157 6953 4169 6987
rect 4203 6953 4215 6987
rect 4157 6947 4215 6953
rect 290 6876 296 6928
rect 348 6916 354 6928
rect 4172 6916 4200 6947
rect 348 6888 4200 6916
rect 348 6876 354 6888
rect 1673 6851 1731 6857
rect 1673 6817 1685 6851
rect 1719 6817 1731 6851
rect 1946 6848 1952 6860
rect 1907 6820 1952 6848
rect 1673 6811 1731 6817
rect 1688 6780 1716 6811
rect 1946 6808 1952 6820
rect 2004 6808 2010 6860
rect 2866 6848 2872 6860
rect 2827 6820 2872 6848
rect 2866 6808 2872 6820
rect 2924 6808 2930 6860
rect 4341 6851 4399 6857
rect 4341 6817 4353 6851
rect 4387 6848 4399 6851
rect 4522 6848 4528 6860
rect 4387 6820 4528 6848
rect 4387 6817 4399 6820
rect 4341 6811 4399 6817
rect 4522 6808 4528 6820
rect 4580 6808 4586 6860
rect 4617 6851 4675 6857
rect 4617 6817 4629 6851
rect 4663 6817 4675 6851
rect 5626 6848 5632 6860
rect 5587 6820 5632 6848
rect 4617 6811 4675 6817
rect 2884 6780 2912 6808
rect 1688 6752 2912 6780
rect 3421 6647 3479 6653
rect 3421 6613 3433 6647
rect 3467 6644 3479 6647
rect 3878 6644 3884 6656
rect 3467 6616 3884 6644
rect 3467 6613 3479 6616
rect 3421 6607 3479 6613
rect 3878 6604 3884 6616
rect 3936 6644 3942 6656
rect 4632 6644 4660 6811
rect 5626 6808 5632 6820
rect 5684 6808 5690 6860
rect 4706 6644 4712 6656
rect 3936 6616 4712 6644
rect 3936 6604 3942 6616
rect 4706 6604 4712 6616
rect 4764 6644 4770 6656
rect 5813 6647 5871 6653
rect 5813 6644 5825 6647
rect 4764 6616 5825 6644
rect 4764 6604 4770 6616
rect 5813 6613 5825 6616
rect 5859 6613 5871 6647
rect 5813 6607 5871 6613
rect 1104 6554 22816 6576
rect 1104 6502 4982 6554
rect 5034 6502 5046 6554
rect 5098 6502 5110 6554
rect 5162 6502 5174 6554
rect 5226 6502 12982 6554
rect 13034 6502 13046 6554
rect 13098 6502 13110 6554
rect 13162 6502 13174 6554
rect 13226 6502 20982 6554
rect 21034 6502 21046 6554
rect 21098 6502 21110 6554
rect 21162 6502 21174 6554
rect 21226 6502 22816 6554
rect 1104 6480 22816 6502
rect 3237 6443 3295 6449
rect 3237 6409 3249 6443
rect 3283 6440 3295 6443
rect 4522 6440 4528 6452
rect 3283 6412 4528 6440
rect 3283 6409 3295 6412
rect 3237 6403 3295 6409
rect 4522 6400 4528 6412
rect 4580 6400 4586 6452
rect 5626 6440 5632 6452
rect 5587 6412 5632 6440
rect 5626 6400 5632 6412
rect 5684 6400 5690 6452
rect 14 6264 20 6316
rect 72 6304 78 6316
rect 4341 6307 4399 6313
rect 4341 6304 4353 6307
rect 72 6276 4353 6304
rect 72 6264 78 6276
rect 4341 6273 4353 6276
rect 4387 6273 4399 6307
rect 4341 6267 4399 6273
rect 1670 6236 1676 6248
rect 1631 6208 1676 6236
rect 1670 6196 1676 6208
rect 1728 6196 1734 6248
rect 1949 6239 2007 6245
rect 1949 6205 1961 6239
rect 1995 6236 2007 6239
rect 2501 6239 2559 6245
rect 2501 6236 2513 6239
rect 1995 6208 2513 6236
rect 1995 6205 2007 6208
rect 1949 6199 2007 6205
rect 2501 6205 2513 6208
rect 2547 6236 2559 6239
rect 2869 6239 2927 6245
rect 2869 6236 2881 6239
rect 2547 6208 2881 6236
rect 2547 6205 2559 6208
rect 2501 6199 2559 6205
rect 2869 6205 2881 6208
rect 2915 6236 2927 6239
rect 3602 6236 3608 6248
rect 2915 6208 3608 6236
rect 2915 6205 2927 6208
rect 2869 6199 2927 6205
rect 3602 6196 3608 6208
rect 3660 6196 3666 6248
rect 3970 6236 3976 6248
rect 3931 6208 3976 6236
rect 3970 6196 3976 6208
rect 4028 6196 4034 6248
rect 4249 6239 4307 6245
rect 4249 6205 4261 6239
rect 4295 6236 4307 6239
rect 4295 6208 4384 6236
rect 4295 6205 4307 6208
rect 4249 6199 4307 6205
rect 3620 6168 3648 6196
rect 4356 6168 4384 6208
rect 3620 6140 4384 6168
rect 106 6060 112 6112
rect 164 6100 170 6112
rect 1489 6103 1547 6109
rect 1489 6100 1501 6103
rect 164 6072 1501 6100
rect 164 6060 170 6072
rect 1489 6069 1501 6072
rect 1535 6069 1547 6103
rect 4706 6100 4712 6112
rect 4667 6072 4712 6100
rect 1489 6063 1547 6069
rect 4706 6060 4712 6072
rect 4764 6060 4770 6112
rect 1104 6010 22816 6032
rect 1104 5958 8982 6010
rect 9034 5958 9046 6010
rect 9098 5958 9110 6010
rect 9162 5958 9174 6010
rect 9226 5958 16982 6010
rect 17034 5958 17046 6010
rect 17098 5958 17110 6010
rect 17162 5958 17174 6010
rect 17226 5958 22816 6010
rect 1104 5936 22816 5958
rect 106 5856 112 5908
rect 164 5896 170 5908
rect 1673 5899 1731 5905
rect 1673 5896 1685 5899
rect 164 5868 1685 5896
rect 164 5856 170 5868
rect 1673 5865 1685 5868
rect 1719 5865 1731 5899
rect 1673 5859 1731 5865
rect 1854 5856 1860 5908
rect 1912 5896 1918 5908
rect 2685 5899 2743 5905
rect 2685 5896 2697 5899
rect 1912 5868 2697 5896
rect 1912 5856 1918 5868
rect 2685 5865 2697 5868
rect 2731 5896 2743 5899
rect 2866 5896 2872 5908
rect 2731 5868 2872 5896
rect 2731 5865 2743 5868
rect 2685 5859 2743 5865
rect 2866 5856 2872 5868
rect 2924 5856 2930 5908
rect 3050 5896 3056 5908
rect 3011 5868 3056 5896
rect 3050 5856 3056 5868
rect 3108 5856 3114 5908
rect 3881 5899 3939 5905
rect 3881 5865 3893 5899
rect 3927 5896 3939 5899
rect 3970 5896 3976 5908
rect 3927 5868 3976 5896
rect 3927 5865 3939 5868
rect 3881 5859 3939 5865
rect 3970 5856 3976 5868
rect 4028 5856 4034 5908
rect 4157 5899 4215 5905
rect 4157 5865 4169 5899
rect 4203 5865 4215 5899
rect 4157 5859 4215 5865
rect 198 5788 204 5840
rect 256 5828 262 5840
rect 4172 5828 4200 5859
rect 256 5800 4200 5828
rect 256 5788 262 5800
rect 1486 5720 1492 5772
rect 1544 5760 1550 5772
rect 1854 5760 1860 5772
rect 1544 5732 1860 5760
rect 1544 5720 1550 5732
rect 1854 5720 1860 5732
rect 1912 5720 1918 5772
rect 2038 5760 2044 5772
rect 1999 5732 2044 5760
rect 2038 5720 2044 5732
rect 2096 5720 2102 5772
rect 3234 5720 3240 5772
rect 3292 5760 3298 5772
rect 4065 5763 4123 5769
rect 4065 5760 4077 5763
rect 3292 5732 4077 5760
rect 3292 5720 3298 5732
rect 4065 5729 4077 5732
rect 4111 5760 4123 5763
rect 4430 5760 4436 5772
rect 4111 5732 4436 5760
rect 4111 5729 4123 5732
rect 4065 5723 4123 5729
rect 4430 5720 4436 5732
rect 4488 5720 4494 5772
rect 4525 5763 4583 5769
rect 4525 5729 4537 5763
rect 4571 5760 4583 5763
rect 4706 5760 4712 5772
rect 4571 5732 4712 5760
rect 4571 5729 4583 5732
rect 4525 5723 4583 5729
rect 1670 5652 1676 5704
rect 1728 5692 1734 5704
rect 3421 5695 3479 5701
rect 3421 5692 3433 5695
rect 1728 5664 3433 5692
rect 1728 5652 1734 5664
rect 3421 5661 3433 5664
rect 3467 5692 3479 5695
rect 3510 5692 3516 5704
rect 3467 5664 3516 5692
rect 3467 5661 3479 5664
rect 3421 5655 3479 5661
rect 3510 5652 3516 5664
rect 3568 5652 3574 5704
rect 4540 5692 4568 5723
rect 4706 5720 4712 5732
rect 4764 5720 4770 5772
rect 4080 5664 4568 5692
rect 4080 5636 4108 5664
rect 4062 5584 4068 5636
rect 4120 5584 4126 5636
rect 1104 5466 22816 5488
rect 1104 5414 4982 5466
rect 5034 5414 5046 5466
rect 5098 5414 5110 5466
rect 5162 5414 5174 5466
rect 5226 5414 12982 5466
rect 13034 5414 13046 5466
rect 13098 5414 13110 5466
rect 13162 5414 13174 5466
rect 13226 5414 20982 5466
rect 21034 5414 21046 5466
rect 21098 5414 21110 5466
rect 21162 5414 21174 5466
rect 21226 5414 22816 5466
rect 1104 5392 22816 5414
rect 4430 5352 4436 5364
rect 4391 5324 4436 5352
rect 4430 5312 4436 5324
rect 4488 5312 4494 5364
rect 5169 5355 5227 5361
rect 5169 5321 5181 5355
rect 5215 5352 5227 5355
rect 5442 5352 5448 5364
rect 5215 5324 5448 5352
rect 5215 5321 5227 5324
rect 5169 5315 5227 5321
rect 4522 5284 4528 5296
rect 4126 5256 4528 5284
rect 2884 5188 3556 5216
rect 2884 5160 2912 5188
rect 1670 5148 1676 5160
rect 1631 5120 1676 5148
rect 1670 5108 1676 5120
rect 1728 5108 1734 5160
rect 2038 5148 2044 5160
rect 1999 5120 2044 5148
rect 2038 5108 2044 5120
rect 2096 5148 2102 5160
rect 2501 5151 2559 5157
rect 2501 5148 2513 5151
rect 2096 5120 2513 5148
rect 2096 5108 2102 5120
rect 2501 5117 2513 5120
rect 2547 5148 2559 5151
rect 2866 5148 2872 5160
rect 2547 5120 2872 5148
rect 2547 5117 2559 5120
rect 2501 5111 2559 5117
rect 2866 5108 2872 5120
rect 2924 5108 2930 5160
rect 3050 5148 3056 5160
rect 3011 5120 3056 5148
rect 3050 5108 3056 5120
rect 3108 5108 3114 5160
rect 3528 5157 3556 5188
rect 3513 5151 3571 5157
rect 3513 5117 3525 5151
rect 3559 5148 3571 5151
rect 4126 5148 4154 5256
rect 4522 5244 4528 5256
rect 4580 5284 4586 5296
rect 4801 5287 4859 5293
rect 4801 5284 4813 5287
rect 4580 5256 4813 5284
rect 4580 5244 4586 5256
rect 4801 5253 4813 5256
rect 4847 5253 4859 5287
rect 4801 5247 4859 5253
rect 3559 5120 4154 5148
rect 4617 5151 4675 5157
rect 3559 5117 3571 5120
rect 3513 5111 3571 5117
rect 4617 5117 4629 5151
rect 4663 5148 4675 5151
rect 5184 5148 5212 5315
rect 5442 5312 5448 5324
rect 5500 5312 5506 5364
rect 4663 5120 5212 5148
rect 4663 5117 4675 5120
rect 4617 5111 4675 5117
rect 14 5040 20 5092
rect 72 5080 78 5092
rect 72 5052 3004 5080
rect 72 5040 78 5052
rect 106 4972 112 5024
rect 164 5012 170 5024
rect 1581 5015 1639 5021
rect 1581 5012 1593 5015
rect 164 4984 1593 5012
rect 164 4972 170 4984
rect 1581 4981 1593 4984
rect 1627 4981 1639 5015
rect 2976 5012 3004 5052
rect 3145 5015 3203 5021
rect 3145 5012 3157 5015
rect 2976 4984 3157 5012
rect 1581 4975 1639 4981
rect 3145 4981 3157 4984
rect 3191 4981 3203 5015
rect 4062 5012 4068 5024
rect 4023 4984 4068 5012
rect 3145 4975 3203 4981
rect 4062 4972 4068 4984
rect 4120 4972 4126 5024
rect 1104 4922 22816 4944
rect 1104 4870 8982 4922
rect 9034 4870 9046 4922
rect 9098 4870 9110 4922
rect 9162 4870 9174 4922
rect 9226 4870 16982 4922
rect 17034 4870 17046 4922
rect 17098 4870 17110 4922
rect 17162 4870 17174 4922
rect 17226 4870 22816 4922
rect 1104 4848 22816 4870
rect 14 4768 20 4820
rect 72 4808 78 4820
rect 1673 4811 1731 4817
rect 1673 4808 1685 4811
rect 72 4780 1685 4808
rect 72 4768 78 4780
rect 1673 4777 1685 4780
rect 1719 4777 1731 4811
rect 1673 4771 1731 4777
rect 2866 4768 2872 4820
rect 2924 4808 2930 4820
rect 3053 4811 3111 4817
rect 3053 4808 3065 4811
rect 2924 4780 3065 4808
rect 2924 4768 2930 4780
rect 3053 4777 3065 4780
rect 3099 4777 3111 4811
rect 3510 4808 3516 4820
rect 3471 4780 3516 4808
rect 3053 4771 3111 4777
rect 3510 4768 3516 4780
rect 3568 4768 3574 4820
rect 3881 4811 3939 4817
rect 3881 4777 3893 4811
rect 3927 4808 3939 4811
rect 3970 4808 3976 4820
rect 3927 4780 3976 4808
rect 3927 4777 3939 4780
rect 3881 4771 3939 4777
rect 3970 4768 3976 4780
rect 4028 4768 4034 4820
rect 4154 4808 4160 4820
rect 4115 4780 4160 4808
rect 4154 4768 4160 4780
rect 4212 4768 4218 4820
rect 1857 4675 1915 4681
rect 1857 4641 1869 4675
rect 1903 4641 1915 4675
rect 2130 4672 2136 4684
rect 2091 4644 2136 4672
rect 1857 4635 1915 4641
rect 1872 4604 1900 4635
rect 2130 4632 2136 4644
rect 2188 4632 2194 4684
rect 2685 4675 2743 4681
rect 2685 4641 2697 4675
rect 2731 4672 2743 4675
rect 2774 4672 2780 4684
rect 2731 4644 2780 4672
rect 2731 4641 2743 4644
rect 2685 4635 2743 4641
rect 2700 4604 2728 4635
rect 2774 4632 2780 4644
rect 2832 4672 2838 4684
rect 3050 4672 3056 4684
rect 2832 4644 3056 4672
rect 2832 4632 2838 4644
rect 3050 4632 3056 4644
rect 3108 4632 3114 4684
rect 3988 4672 4016 4768
rect 4065 4675 4123 4681
rect 4065 4672 4077 4675
rect 3988 4644 4077 4672
rect 4065 4641 4077 4644
rect 4111 4672 4123 4675
rect 4338 4672 4344 4684
rect 4111 4644 4344 4672
rect 4111 4641 4123 4644
rect 4065 4635 4123 4641
rect 4338 4632 4344 4644
rect 4396 4632 4402 4684
rect 4522 4672 4528 4684
rect 4483 4644 4528 4672
rect 4522 4632 4528 4644
rect 4580 4632 4586 4684
rect 1872 4576 2728 4604
rect 1104 4378 22816 4400
rect 1104 4326 4982 4378
rect 5034 4326 5046 4378
rect 5098 4326 5110 4378
rect 5162 4326 5174 4378
rect 5226 4326 12982 4378
rect 13034 4326 13046 4378
rect 13098 4326 13110 4378
rect 13162 4326 13174 4378
rect 13226 4326 20982 4378
rect 21034 4326 21046 4378
rect 21098 4326 21110 4378
rect 21162 4326 21174 4378
rect 21226 4326 22816 4378
rect 1104 4304 22816 4326
rect 5353 4267 5411 4273
rect 5353 4264 5365 4267
rect 4264 4236 5365 4264
rect 2409 4199 2467 4205
rect 2409 4165 2421 4199
rect 2455 4196 2467 4199
rect 2685 4199 2743 4205
rect 2685 4196 2697 4199
rect 2455 4168 2697 4196
rect 2455 4165 2467 4168
rect 2409 4159 2467 4165
rect 2685 4165 2697 4168
rect 2731 4196 2743 4199
rect 3053 4199 3111 4205
rect 3053 4196 3065 4199
rect 2731 4168 3065 4196
rect 2731 4165 2743 4168
rect 2685 4159 2743 4165
rect 3053 4165 3065 4168
rect 3099 4196 3111 4199
rect 3513 4199 3571 4205
rect 3513 4196 3525 4199
rect 3099 4168 3525 4196
rect 3099 4165 3111 4168
rect 3053 4159 3111 4165
rect 3513 4165 3525 4168
rect 3559 4196 3571 4199
rect 4264 4196 4292 4236
rect 5353 4233 5365 4236
rect 5399 4233 5411 4267
rect 5353 4227 5411 4233
rect 3559 4168 4292 4196
rect 3559 4165 3571 4168
rect 3513 4159 3571 4165
rect 106 4088 112 4140
rect 164 4128 170 4140
rect 4157 4131 4215 4137
rect 4157 4128 4169 4131
rect 164 4100 4169 4128
rect 164 4088 170 4100
rect 4157 4097 4169 4100
rect 4203 4097 4215 4131
rect 4157 4091 4215 4097
rect 1486 4020 1492 4072
rect 1544 4060 1550 4072
rect 1581 4063 1639 4069
rect 1581 4060 1593 4063
rect 1544 4032 1593 4060
rect 1544 4020 1550 4032
rect 1581 4029 1593 4032
rect 1627 4029 1639 4063
rect 2130 4060 2136 4072
rect 2091 4032 2136 4060
rect 1581 4023 1639 4029
rect 2130 4020 2136 4032
rect 2188 4060 2194 4072
rect 2409 4063 2467 4069
rect 2409 4060 2421 4063
rect 2188 4032 2421 4060
rect 2188 4020 2194 4032
rect 2409 4029 2421 4032
rect 2455 4029 2467 4063
rect 2409 4023 2467 4029
rect 3789 4063 3847 4069
rect 3789 4029 3801 4063
rect 3835 4060 3847 4063
rect 3878 4060 3884 4072
rect 3835 4032 3884 4060
rect 3835 4029 3847 4032
rect 3789 4023 3847 4029
rect 3878 4020 3884 4032
rect 3936 4020 3942 4072
rect 4065 4063 4123 4069
rect 4065 4029 4077 4063
rect 4111 4060 4123 4063
rect 4264 4060 4292 4168
rect 4522 4156 4528 4208
rect 4580 4196 4586 4208
rect 4617 4199 4675 4205
rect 4617 4196 4629 4199
rect 4580 4168 4629 4196
rect 4580 4156 4586 4168
rect 4617 4165 4629 4168
rect 4663 4165 4675 4199
rect 4617 4159 4675 4165
rect 4338 4088 4344 4140
rect 4396 4128 4402 4140
rect 4985 4131 5043 4137
rect 4985 4128 4997 4131
rect 4396 4100 4997 4128
rect 4396 4088 4402 4100
rect 4985 4097 4997 4100
rect 5031 4097 5043 4131
rect 4985 4091 5043 4097
rect 4111 4032 4292 4060
rect 4111 4029 4123 4032
rect 4065 4023 4123 4029
rect 4430 4020 4436 4072
rect 4488 4060 4494 4072
rect 5169 4063 5227 4069
rect 5169 4060 5181 4063
rect 4488 4032 5181 4060
rect 4488 4020 4494 4032
rect 5169 4029 5181 4032
rect 5215 4060 5227 4063
rect 5629 4063 5687 4069
rect 5629 4060 5641 4063
rect 5215 4032 5641 4060
rect 5215 4029 5227 4032
rect 5169 4023 5227 4029
rect 5629 4029 5641 4032
rect 5675 4029 5687 4063
rect 5629 4023 5687 4029
rect 106 3884 112 3936
rect 164 3924 170 3936
rect 1673 3927 1731 3933
rect 1673 3924 1685 3927
rect 164 3896 1685 3924
rect 164 3884 170 3896
rect 1673 3893 1685 3896
rect 1719 3893 1731 3927
rect 1673 3887 1731 3893
rect 1104 3834 22816 3856
rect 1104 3782 8982 3834
rect 9034 3782 9046 3834
rect 9098 3782 9110 3834
rect 9162 3782 9174 3834
rect 9226 3782 16982 3834
rect 17034 3782 17046 3834
rect 17098 3782 17110 3834
rect 17162 3782 17174 3834
rect 17226 3782 22816 3834
rect 1104 3760 22816 3782
rect 14 3680 20 3732
rect 72 3720 78 3732
rect 1765 3723 1823 3729
rect 1765 3720 1777 3723
rect 72 3692 1777 3720
rect 72 3680 78 3692
rect 1765 3689 1777 3692
rect 1811 3689 1823 3723
rect 3510 3720 3516 3732
rect 3471 3692 3516 3720
rect 1765 3683 1823 3689
rect 3510 3680 3516 3692
rect 3568 3680 3574 3732
rect 3878 3720 3884 3732
rect 3839 3692 3884 3720
rect 3878 3680 3884 3692
rect 3936 3680 3942 3732
rect 2685 3655 2743 3661
rect 2685 3652 2697 3655
rect 1688 3624 2697 3652
rect 1486 3544 1492 3596
rect 1544 3584 1550 3596
rect 1688 3593 1716 3624
rect 2685 3621 2697 3624
rect 2731 3652 2743 3655
rect 3053 3655 3111 3661
rect 3053 3652 3065 3655
rect 2731 3624 3065 3652
rect 2731 3621 2743 3624
rect 2685 3615 2743 3621
rect 3053 3621 3065 3624
rect 3099 3621 3111 3655
rect 3053 3615 3111 3621
rect 1673 3587 1731 3593
rect 1673 3584 1685 3587
rect 1544 3556 1685 3584
rect 1544 3544 1550 3556
rect 1673 3553 1685 3556
rect 1719 3553 1731 3587
rect 2222 3584 2228 3596
rect 2183 3556 2228 3584
rect 1673 3547 1731 3553
rect 2222 3544 2228 3556
rect 2280 3544 2286 3596
rect 3896 3584 3924 3680
rect 4065 3587 4123 3593
rect 4065 3584 4077 3587
rect 3896 3556 4077 3584
rect 4065 3553 4077 3556
rect 4111 3553 4123 3587
rect 4614 3584 4620 3596
rect 4575 3556 4620 3584
rect 4065 3547 4123 3553
rect 4614 3544 4620 3556
rect 4672 3544 4678 3596
rect 382 3476 388 3528
rect 440 3516 446 3528
rect 4525 3519 4583 3525
rect 4525 3516 4537 3519
rect 440 3488 4537 3516
rect 440 3476 446 3488
rect 4525 3485 4537 3488
rect 4571 3485 4583 3519
rect 4525 3479 4583 3485
rect 1104 3290 22816 3312
rect 1104 3238 4982 3290
rect 5034 3238 5046 3290
rect 5098 3238 5110 3290
rect 5162 3238 5174 3290
rect 5226 3238 12982 3290
rect 13034 3238 13046 3290
rect 13098 3238 13110 3290
rect 13162 3238 13174 3290
rect 13226 3238 20982 3290
rect 21034 3238 21046 3290
rect 21098 3238 21110 3290
rect 21162 3238 21174 3290
rect 21226 3238 22816 3290
rect 1104 3216 22816 3238
rect 4338 3136 4344 3188
rect 4396 3176 4402 3188
rect 5077 3179 5135 3185
rect 5077 3176 5089 3179
rect 4396 3148 5089 3176
rect 4396 3136 4402 3148
rect 5077 3145 5089 3148
rect 5123 3145 5135 3179
rect 5077 3139 5135 3145
rect 5813 3179 5871 3185
rect 5813 3145 5825 3179
rect 5859 3176 5871 3179
rect 5902 3176 5908 3188
rect 5859 3148 5908 3176
rect 5859 3145 5871 3148
rect 5813 3139 5871 3145
rect 4614 3068 4620 3120
rect 4672 3108 4678 3120
rect 4801 3111 4859 3117
rect 4801 3108 4813 3111
rect 4672 3080 4813 3108
rect 4672 3068 4678 3080
rect 4801 3077 4813 3080
rect 4847 3108 4859 3111
rect 5445 3111 5503 3117
rect 5445 3108 5457 3111
rect 4847 3080 5457 3108
rect 4847 3077 4859 3080
rect 4801 3071 4859 3077
rect 5445 3077 5457 3080
rect 5491 3077 5503 3111
rect 5445 3071 5503 3077
rect 3605 3043 3663 3049
rect 3605 3009 3617 3043
rect 3651 3040 3663 3043
rect 4062 3040 4068 3052
rect 3651 3012 4068 3040
rect 3651 3009 3663 3012
rect 3605 3003 3663 3009
rect 4062 3000 4068 3012
rect 4120 3040 4126 3052
rect 4120 3012 4292 3040
rect 4120 3000 4126 3012
rect 1762 2972 1768 2984
rect 1723 2944 1768 2972
rect 1762 2932 1768 2944
rect 1820 2932 1826 2984
rect 2130 2972 2136 2984
rect 2043 2944 2136 2972
rect 2130 2932 2136 2944
rect 2188 2972 2194 2984
rect 2593 2975 2651 2981
rect 2593 2972 2605 2975
rect 2188 2944 2605 2972
rect 2188 2932 2194 2944
rect 2593 2941 2605 2944
rect 2639 2941 2651 2975
rect 3878 2972 3884 2984
rect 3839 2944 3884 2972
rect 2593 2935 2651 2941
rect 3878 2932 3884 2944
rect 3936 2932 3942 2984
rect 4264 2981 4292 3012
rect 4249 2975 4307 2981
rect 4249 2941 4261 2975
rect 4295 2941 4307 2975
rect 4249 2935 4307 2941
rect 5261 2975 5319 2981
rect 5261 2941 5273 2975
rect 5307 2972 5319 2975
rect 5828 2972 5856 3139
rect 5902 3136 5908 3148
rect 5960 3136 5966 3188
rect 5307 2944 5856 2972
rect 5307 2941 5319 2944
rect 5261 2935 5319 2941
rect 106 2796 112 2848
rect 164 2836 170 2848
rect 1673 2839 1731 2845
rect 1673 2836 1685 2839
rect 164 2808 1685 2836
rect 164 2796 170 2808
rect 1673 2805 1685 2808
rect 1719 2805 1731 2839
rect 1673 2799 1731 2805
rect 2222 2796 2228 2848
rect 2280 2836 2286 2848
rect 2961 2839 3019 2845
rect 2961 2836 2973 2839
rect 2280 2808 2973 2836
rect 2280 2796 2286 2808
rect 2961 2805 2973 2808
rect 3007 2805 3019 2839
rect 3786 2836 3792 2848
rect 3747 2808 3792 2836
rect 2961 2799 3019 2805
rect 3786 2796 3792 2808
rect 3844 2796 3850 2848
rect 1104 2746 22816 2768
rect 1104 2694 8982 2746
rect 9034 2694 9046 2746
rect 9098 2694 9110 2746
rect 9162 2694 9174 2746
rect 9226 2694 16982 2746
rect 17034 2694 17046 2746
rect 17098 2694 17110 2746
rect 17162 2694 17174 2746
rect 17226 2694 22816 2746
rect 1104 2672 22816 2694
rect 106 2592 112 2644
rect 164 2632 170 2644
rect 1765 2635 1823 2641
rect 1765 2632 1777 2635
rect 164 2604 1777 2632
rect 164 2592 170 2604
rect 1765 2601 1777 2604
rect 1811 2601 1823 2635
rect 1765 2595 1823 2601
rect 3145 2635 3203 2641
rect 3145 2601 3157 2635
rect 3191 2632 3203 2635
rect 3510 2632 3516 2644
rect 3191 2604 3516 2632
rect 3191 2601 3203 2604
rect 3145 2595 3203 2601
rect 3510 2592 3516 2604
rect 3568 2592 3574 2644
rect 2774 2524 2780 2576
rect 2832 2564 2838 2576
rect 3421 2567 3479 2573
rect 3421 2564 3433 2567
rect 2832 2536 3433 2564
rect 2832 2524 2838 2536
rect 3421 2533 3433 2536
rect 3467 2533 3479 2567
rect 3421 2527 3479 2533
rect 3697 2567 3755 2573
rect 3697 2533 3709 2567
rect 3743 2564 3755 2567
rect 3743 2536 4660 2564
rect 3743 2533 3755 2536
rect 3697 2527 3755 2533
rect 1762 2496 1768 2508
rect 1723 2468 1768 2496
rect 1762 2456 1768 2468
rect 1820 2456 1826 2508
rect 2222 2496 2228 2508
rect 2183 2468 2228 2496
rect 2222 2456 2228 2468
rect 2280 2496 2286 2508
rect 2685 2499 2743 2505
rect 2685 2496 2697 2499
rect 2280 2468 2697 2496
rect 2280 2456 2286 2468
rect 2685 2465 2697 2468
rect 2731 2465 2743 2499
rect 3436 2496 3464 2527
rect 4632 2508 4660 2536
rect 4065 2499 4123 2505
rect 4065 2496 4077 2499
rect 3436 2468 4077 2496
rect 2685 2459 2743 2465
rect 4065 2465 4077 2468
rect 4111 2465 4123 2499
rect 4614 2496 4620 2508
rect 4575 2468 4620 2496
rect 4065 2459 4123 2465
rect 2700 2428 2728 2459
rect 4614 2456 4620 2468
rect 4672 2456 4678 2508
rect 3697 2431 3755 2437
rect 3697 2428 3709 2431
rect 2700 2400 3709 2428
rect 3697 2397 3709 2400
rect 3743 2428 3755 2431
rect 3789 2431 3847 2437
rect 3789 2428 3801 2431
rect 3743 2400 3801 2428
rect 3743 2397 3755 2400
rect 3697 2391 3755 2397
rect 3789 2397 3801 2400
rect 3835 2397 3847 2431
rect 4525 2431 4583 2437
rect 4525 2428 4537 2431
rect 3789 2391 3847 2397
rect 4080 2400 4537 2428
rect 382 2320 388 2372
rect 440 2360 446 2372
rect 4080 2360 4108 2400
rect 4525 2397 4537 2400
rect 4571 2397 4583 2431
rect 4525 2391 4583 2397
rect 440 2332 4108 2360
rect 440 2320 446 2332
rect 1104 2202 22816 2224
rect 1104 2150 4982 2202
rect 5034 2150 5046 2202
rect 5098 2150 5110 2202
rect 5162 2150 5174 2202
rect 5226 2150 12982 2202
rect 13034 2150 13046 2202
rect 13098 2150 13110 2202
rect 13162 2150 13174 2202
rect 13226 2150 20982 2202
rect 21034 2150 21046 2202
rect 21098 2150 21110 2202
rect 21162 2150 21174 2202
rect 21226 2150 22816 2202
rect 1104 2128 22816 2150
rect 106 1300 112 1352
rect 164 1340 170 1352
rect 3786 1340 3792 1352
rect 164 1312 3792 1340
rect 164 1300 170 1312
rect 3786 1300 3792 1312
rect 3844 1300 3850 1352
<< via1 >>
rect 1952 23536 2004 23588
rect 2596 23536 2648 23588
rect 112 21836 164 21888
rect 4160 21836 4212 21888
rect 4982 21734 5034 21786
rect 5046 21734 5098 21786
rect 5110 21734 5162 21786
rect 5174 21734 5226 21786
rect 12982 21734 13034 21786
rect 13046 21734 13098 21786
rect 13110 21734 13162 21786
rect 13174 21734 13226 21786
rect 20982 21734 21034 21786
rect 21046 21734 21098 21786
rect 21110 21734 21162 21786
rect 21174 21734 21226 21786
rect 112 21360 164 21412
rect 2136 21292 2188 21344
rect 8982 21190 9034 21242
rect 9046 21190 9098 21242
rect 9110 21190 9162 21242
rect 9174 21190 9226 21242
rect 16982 21190 17034 21242
rect 17046 21190 17098 21242
rect 17110 21190 17162 21242
rect 17174 21190 17226 21242
rect 4160 21131 4212 21140
rect 4160 21097 4169 21131
rect 4169 21097 4203 21131
rect 4203 21097 4212 21131
rect 4160 21088 4212 21097
rect 2136 20952 2188 21004
rect 4068 20995 4120 21004
rect 4068 20961 4077 20995
rect 4077 20961 4111 20995
rect 4111 20961 4120 20995
rect 4068 20952 4120 20961
rect 2504 20884 2556 20936
rect 2136 20748 2188 20800
rect 3516 20748 3568 20800
rect 5356 20748 5408 20800
rect 4982 20646 5034 20698
rect 5046 20646 5098 20698
rect 5110 20646 5162 20698
rect 5174 20646 5226 20698
rect 12982 20646 13034 20698
rect 13046 20646 13098 20698
rect 13110 20646 13162 20698
rect 13174 20646 13226 20698
rect 20982 20646 21034 20698
rect 21046 20646 21098 20698
rect 21110 20646 21162 20698
rect 21174 20646 21226 20698
rect 20 20408 72 20460
rect 112 20204 164 20256
rect 2136 20340 2188 20392
rect 3516 20383 3568 20392
rect 2412 20247 2464 20256
rect 2412 20213 2421 20247
rect 2421 20213 2455 20247
rect 2455 20213 2464 20247
rect 2412 20204 2464 20213
rect 2504 20204 2556 20256
rect 3516 20349 3525 20383
rect 3525 20349 3559 20383
rect 3559 20349 3568 20383
rect 3516 20340 3568 20349
rect 4528 20383 4580 20392
rect 4528 20349 4537 20383
rect 4537 20349 4571 20383
rect 4571 20349 4580 20383
rect 4528 20340 4580 20349
rect 5356 20340 5408 20392
rect 7012 20340 7064 20392
rect 4068 20247 4120 20256
rect 4068 20213 4077 20247
rect 4077 20213 4111 20247
rect 4111 20213 4120 20247
rect 4068 20204 4120 20213
rect 4712 20247 4764 20256
rect 4712 20213 4721 20247
rect 4721 20213 4755 20247
rect 4755 20213 4764 20247
rect 4712 20204 4764 20213
rect 8982 20102 9034 20154
rect 9046 20102 9098 20154
rect 9110 20102 9162 20154
rect 9174 20102 9226 20154
rect 16982 20102 17034 20154
rect 17046 20102 17098 20154
rect 17110 20102 17162 20154
rect 17174 20102 17226 20154
rect 388 20000 440 20052
rect 4620 20043 4672 20052
rect 4620 20009 4629 20043
rect 4629 20009 4663 20043
rect 4663 20009 4672 20043
rect 4620 20000 4672 20009
rect 4344 19975 4396 19984
rect 4344 19941 4353 19975
rect 4353 19941 4387 19975
rect 4387 19941 4396 19975
rect 4344 19932 4396 19941
rect 5356 19932 5408 19984
rect 1676 19907 1728 19916
rect 1676 19873 1685 19907
rect 1685 19873 1719 19907
rect 1719 19873 1728 19907
rect 1676 19864 1728 19873
rect 2136 19864 2188 19916
rect 4528 19907 4580 19916
rect 4528 19873 4537 19907
rect 4537 19873 4571 19907
rect 4571 19873 4580 19907
rect 4528 19864 4580 19873
rect 4160 19796 4212 19848
rect 6276 19864 6328 19916
rect 2504 19660 2556 19712
rect 4982 19558 5034 19610
rect 5046 19558 5098 19610
rect 5110 19558 5162 19610
rect 5174 19558 5226 19610
rect 12982 19558 13034 19610
rect 13046 19558 13098 19610
rect 13110 19558 13162 19610
rect 13174 19558 13226 19610
rect 20982 19558 21034 19610
rect 21046 19558 21098 19610
rect 21110 19558 21162 19610
rect 21174 19558 21226 19610
rect 2136 19456 2188 19508
rect 4528 19499 4580 19508
rect 4528 19465 4537 19499
rect 4537 19465 4571 19499
rect 4571 19465 4580 19499
rect 4528 19456 4580 19465
rect 7012 19499 7064 19508
rect 7012 19465 7021 19499
rect 7021 19465 7055 19499
rect 7055 19465 7064 19499
rect 7012 19456 7064 19465
rect 204 19320 256 19372
rect 1676 19295 1728 19304
rect 1676 19261 1685 19295
rect 1685 19261 1719 19295
rect 1719 19261 1728 19295
rect 1676 19252 1728 19261
rect 2688 19252 2740 19304
rect 3608 19295 3660 19304
rect 3608 19261 3617 19295
rect 3617 19261 3651 19295
rect 3651 19261 3660 19295
rect 3608 19252 3660 19261
rect 4344 19252 4396 19304
rect 4528 19252 4580 19304
rect 4804 19252 4856 19304
rect 6828 19295 6880 19304
rect 296 19184 348 19236
rect 1860 19116 1912 19168
rect 2412 19116 2464 19168
rect 6828 19261 6837 19295
rect 6837 19261 6871 19295
rect 6871 19261 6880 19295
rect 6828 19252 6880 19261
rect 5908 19159 5960 19168
rect 5908 19125 5917 19159
rect 5917 19125 5951 19159
rect 5951 19125 5960 19159
rect 5908 19116 5960 19125
rect 6276 19159 6328 19168
rect 6276 19125 6285 19159
rect 6285 19125 6319 19159
rect 6319 19125 6328 19159
rect 6276 19116 6328 19125
rect 8982 19014 9034 19066
rect 9046 19014 9098 19066
rect 9110 19014 9162 19066
rect 9174 19014 9226 19066
rect 16982 19014 17034 19066
rect 17046 19014 17098 19066
rect 17110 19014 17162 19066
rect 17174 19014 17226 19066
rect 1768 18955 1820 18964
rect 1768 18921 1777 18955
rect 1777 18921 1811 18955
rect 1811 18921 1820 18955
rect 1768 18912 1820 18921
rect 3608 18912 3660 18964
rect 4160 18912 4212 18964
rect 4252 18912 4304 18964
rect 2228 18819 2280 18828
rect 2228 18785 2237 18819
rect 2237 18785 2271 18819
rect 2271 18785 2280 18819
rect 2228 18776 2280 18785
rect 4068 18819 4120 18828
rect 4068 18785 4077 18819
rect 4077 18785 4111 18819
rect 4111 18785 4120 18819
rect 4068 18776 4120 18785
rect 4620 18819 4672 18828
rect 4620 18785 4629 18819
rect 4629 18785 4663 18819
rect 4663 18785 4672 18819
rect 5632 18819 5684 18828
rect 4620 18776 4672 18785
rect 5632 18785 5641 18819
rect 5641 18785 5675 18819
rect 5675 18785 5684 18819
rect 5632 18776 5684 18785
rect 2412 18708 2464 18760
rect 5448 18572 5500 18624
rect 6184 18615 6236 18624
rect 6184 18581 6193 18615
rect 6193 18581 6227 18615
rect 6227 18581 6236 18615
rect 6184 18572 6236 18581
rect 4982 18470 5034 18522
rect 5046 18470 5098 18522
rect 5110 18470 5162 18522
rect 5174 18470 5226 18522
rect 12982 18470 13034 18522
rect 13046 18470 13098 18522
rect 13110 18470 13162 18522
rect 13174 18470 13226 18522
rect 20982 18470 21034 18522
rect 21046 18470 21098 18522
rect 21110 18470 21162 18522
rect 21174 18470 21226 18522
rect 5448 18411 5500 18420
rect 5448 18377 5457 18411
rect 5457 18377 5491 18411
rect 5491 18377 5500 18411
rect 5448 18368 5500 18377
rect 6276 18368 6328 18420
rect 112 18232 164 18284
rect 2688 18232 2740 18284
rect 4068 18232 4120 18284
rect 5540 18275 5592 18284
rect 5540 18241 5549 18275
rect 5549 18241 5583 18275
rect 5583 18241 5592 18275
rect 5540 18232 5592 18241
rect 2228 18207 2280 18216
rect 2228 18173 2237 18207
rect 2237 18173 2271 18207
rect 2271 18173 2280 18207
rect 2228 18164 2280 18173
rect 3792 18207 3844 18216
rect 3792 18173 3801 18207
rect 3801 18173 3835 18207
rect 3835 18173 3844 18207
rect 3792 18164 3844 18173
rect 4620 18164 4672 18216
rect 6184 18164 6236 18216
rect 6920 18164 6972 18216
rect 4804 18096 4856 18148
rect 5172 18139 5224 18148
rect 5172 18105 5181 18139
rect 5181 18105 5215 18139
rect 5215 18105 5224 18139
rect 5172 18096 5224 18105
rect 1768 18028 1820 18080
rect 2412 18028 2464 18080
rect 3240 18071 3292 18080
rect 3240 18037 3249 18071
rect 3249 18037 3283 18071
rect 3283 18037 3292 18071
rect 3240 18028 3292 18037
rect 3424 18071 3476 18080
rect 3424 18037 3433 18071
rect 3433 18037 3467 18071
rect 3467 18037 3476 18071
rect 3424 18028 3476 18037
rect 6552 18071 6604 18080
rect 6552 18037 6561 18071
rect 6561 18037 6595 18071
rect 6595 18037 6604 18071
rect 6552 18028 6604 18037
rect 7012 18071 7064 18080
rect 7012 18037 7021 18071
rect 7021 18037 7055 18071
rect 7055 18037 7064 18071
rect 7012 18028 7064 18037
rect 8982 17926 9034 17978
rect 9046 17926 9098 17978
rect 9110 17926 9162 17978
rect 9174 17926 9226 17978
rect 16982 17926 17034 17978
rect 17046 17926 17098 17978
rect 17110 17926 17162 17978
rect 17174 17926 17226 17978
rect 20 17824 72 17876
rect 2228 17824 2280 17876
rect 3792 17867 3844 17876
rect 3792 17833 3801 17867
rect 3801 17833 3835 17867
rect 3835 17833 3844 17867
rect 3792 17824 3844 17833
rect 6184 17867 6236 17876
rect 6184 17833 6193 17867
rect 6193 17833 6227 17867
rect 6227 17833 6236 17867
rect 6920 17867 6972 17876
rect 6184 17824 6236 17833
rect 6920 17833 6929 17867
rect 6929 17833 6963 17867
rect 6963 17833 6972 17867
rect 6920 17824 6972 17833
rect 5632 17756 5684 17808
rect 6552 17756 6604 17808
rect 1952 17731 2004 17740
rect 1952 17697 1961 17731
rect 1961 17697 1995 17731
rect 1995 17697 2004 17731
rect 1952 17688 2004 17697
rect 4436 17688 4488 17740
rect 2412 17620 2464 17672
rect 4252 17527 4304 17536
rect 4252 17493 4261 17527
rect 4261 17493 4295 17527
rect 4295 17493 4304 17527
rect 4252 17484 4304 17493
rect 4528 17527 4580 17536
rect 4528 17493 4537 17527
rect 4537 17493 4571 17527
rect 4571 17493 4580 17527
rect 5172 17688 5224 17740
rect 6644 17688 6696 17740
rect 5632 17620 5684 17672
rect 5724 17620 5776 17672
rect 7012 17620 7064 17672
rect 6184 17552 6236 17604
rect 4528 17484 4580 17493
rect 5448 17484 5500 17536
rect 6092 17484 6144 17536
rect 20 17459 72 17468
rect 20 17425 29 17459
rect 29 17425 63 17459
rect 63 17425 72 17459
rect 20 17416 72 17425
rect 4982 17382 5034 17434
rect 5046 17382 5098 17434
rect 5110 17382 5162 17434
rect 5174 17382 5226 17434
rect 12982 17382 13034 17434
rect 13046 17382 13098 17434
rect 13110 17382 13162 17434
rect 13174 17382 13226 17434
rect 20982 17382 21034 17434
rect 21046 17382 21098 17434
rect 21110 17382 21162 17434
rect 21174 17382 21226 17434
rect 5724 17280 5776 17332
rect 6828 17280 6880 17332
rect 20 17144 72 17196
rect 5356 17144 5408 17196
rect 6092 17212 6144 17264
rect 1768 17076 1820 17128
rect 1952 17119 2004 17128
rect 1952 17085 1961 17119
rect 1961 17085 1995 17119
rect 1995 17085 2004 17119
rect 1952 17076 2004 17085
rect 3516 17119 3568 17128
rect 3240 17008 3292 17060
rect 3516 17085 3525 17119
rect 3525 17085 3559 17119
rect 3559 17085 3568 17119
rect 3516 17076 3568 17085
rect 5632 17144 5684 17196
rect 6920 17144 6972 17196
rect 3700 17008 3752 17060
rect 112 16940 164 16992
rect 2412 16983 2464 16992
rect 2412 16949 2421 16983
rect 2421 16949 2455 16983
rect 2455 16949 2464 16983
rect 2412 16940 2464 16949
rect 4344 16983 4396 16992
rect 4344 16949 4353 16983
rect 4353 16949 4387 16983
rect 4387 16949 4396 16983
rect 7380 17076 7432 17128
rect 5172 17051 5224 17060
rect 5172 17017 5181 17051
rect 5181 17017 5215 17051
rect 5215 17017 5224 17051
rect 5172 17008 5224 17017
rect 4344 16940 4396 16949
rect 5356 16940 5408 16992
rect 6644 16983 6696 16992
rect 6644 16949 6653 16983
rect 6653 16949 6687 16983
rect 6687 16949 6696 16983
rect 6644 16940 6696 16949
rect 7380 16983 7432 16992
rect 7380 16949 7389 16983
rect 7389 16949 7423 16983
rect 7423 16949 7432 16983
rect 7380 16940 7432 16949
rect 8982 16838 9034 16890
rect 9046 16838 9098 16890
rect 9110 16838 9162 16890
rect 9174 16838 9226 16890
rect 16982 16838 17034 16890
rect 17046 16838 17098 16890
rect 17110 16838 17162 16890
rect 17174 16838 17226 16890
rect 1952 16668 2004 16720
rect 2872 16668 2924 16720
rect 3516 16668 3568 16720
rect 6920 16779 6972 16788
rect 6920 16745 6929 16779
rect 6929 16745 6963 16779
rect 6963 16745 6972 16779
rect 6920 16736 6972 16745
rect 5632 16668 5684 16720
rect 5908 16711 5960 16720
rect 5908 16677 5917 16711
rect 5917 16677 5951 16711
rect 5951 16677 5960 16711
rect 5908 16668 5960 16677
rect 3976 16600 4028 16652
rect 4528 16600 4580 16652
rect 5172 16643 5224 16652
rect 5172 16609 5181 16643
rect 5181 16609 5215 16643
rect 5215 16609 5224 16643
rect 5172 16600 5224 16609
rect 6368 16600 6420 16652
rect 6736 16643 6788 16652
rect 6736 16609 6745 16643
rect 6745 16609 6779 16643
rect 6779 16609 6788 16643
rect 6736 16600 6788 16609
rect 2688 16532 2740 16584
rect 4436 16532 4488 16584
rect 5540 16575 5592 16584
rect 5540 16541 5549 16575
rect 5549 16541 5583 16575
rect 5583 16541 5592 16575
rect 5540 16532 5592 16541
rect 1768 16396 1820 16448
rect 5724 16464 5776 16516
rect 5448 16439 5500 16448
rect 5448 16405 5457 16439
rect 5457 16405 5491 16439
rect 5491 16405 5500 16439
rect 5448 16396 5500 16405
rect 4982 16294 5034 16346
rect 5046 16294 5098 16346
rect 5110 16294 5162 16346
rect 5174 16294 5226 16346
rect 12982 16294 13034 16346
rect 13046 16294 13098 16346
rect 13110 16294 13162 16346
rect 13174 16294 13226 16346
rect 20982 16294 21034 16346
rect 21046 16294 21098 16346
rect 21110 16294 21162 16346
rect 21174 16294 21226 16346
rect 4436 16192 4488 16244
rect 5540 16192 5592 16244
rect 6368 16192 6420 16244
rect 7748 16235 7800 16244
rect 7748 16201 7757 16235
rect 7757 16201 7791 16235
rect 7791 16201 7800 16235
rect 7748 16192 7800 16201
rect 5356 16124 5408 16176
rect 5632 16124 5684 16176
rect 2412 16056 2464 16108
rect 1584 16031 1636 16040
rect 1584 15997 1593 16031
rect 1593 15997 1627 16031
rect 1627 15997 1636 16031
rect 1584 15988 1636 15997
rect 2136 16031 2188 16040
rect 2136 15997 2145 16031
rect 2145 15997 2179 16031
rect 2179 15997 2188 16031
rect 2136 15988 2188 15997
rect 4344 16056 4396 16108
rect 4068 15988 4120 16040
rect 4859 16031 4911 16040
rect 4859 15997 4868 16031
rect 4868 15997 4902 16031
rect 4902 15997 4911 16031
rect 4859 15988 4911 15997
rect 6644 16056 6696 16108
rect 5448 15988 5500 16040
rect 7840 16031 7892 16040
rect 7840 15997 7849 16031
rect 7849 15997 7883 16031
rect 7883 15997 7892 16031
rect 7840 15988 7892 15997
rect 20 15920 72 15972
rect 4528 15920 4580 15972
rect 6736 15920 6788 15972
rect 7564 15920 7616 15972
rect 9588 15920 9640 15972
rect 2688 15895 2740 15904
rect 2688 15861 2697 15895
rect 2697 15861 2731 15895
rect 2731 15861 2740 15895
rect 2688 15852 2740 15861
rect 3240 15895 3292 15904
rect 3240 15861 3249 15895
rect 3249 15861 3283 15895
rect 3283 15861 3292 15895
rect 3240 15852 3292 15861
rect 6368 15852 6420 15904
rect 8982 15750 9034 15802
rect 9046 15750 9098 15802
rect 9110 15750 9162 15802
rect 9174 15750 9226 15802
rect 16982 15750 17034 15802
rect 17046 15750 17098 15802
rect 17110 15750 17162 15802
rect 17174 15750 17226 15802
rect 204 15648 256 15700
rect 2872 15691 2924 15700
rect 2872 15657 2881 15691
rect 2881 15657 2915 15691
rect 2915 15657 2924 15691
rect 2872 15648 2924 15657
rect 3976 15648 4028 15700
rect 4712 15648 4764 15700
rect 5632 15648 5684 15700
rect 5724 15648 5776 15700
rect 6460 15691 6512 15700
rect 6460 15657 6469 15691
rect 6469 15657 6503 15691
rect 6503 15657 6512 15691
rect 6460 15648 6512 15657
rect 2136 15580 2188 15632
rect 1860 15555 1912 15564
rect 1860 15521 1869 15555
rect 1869 15521 1903 15555
rect 1903 15521 1912 15555
rect 1860 15512 1912 15521
rect 3332 15580 3384 15632
rect 4252 15580 4304 15632
rect 7840 15580 7892 15632
rect 3792 15512 3844 15564
rect 4528 15512 4580 15564
rect 6276 15512 6328 15564
rect 4804 15444 4856 15496
rect 5540 15444 5592 15496
rect 7656 15444 7708 15496
rect 3976 15376 4028 15428
rect 1584 15351 1636 15360
rect 1584 15317 1593 15351
rect 1593 15317 1627 15351
rect 1627 15317 1636 15351
rect 1584 15308 1636 15317
rect 4712 15308 4764 15360
rect 5356 15308 5408 15360
rect 5448 15308 5500 15360
rect 4982 15206 5034 15258
rect 5046 15206 5098 15258
rect 5110 15206 5162 15258
rect 5174 15206 5226 15258
rect 12982 15206 13034 15258
rect 13046 15206 13098 15258
rect 13110 15206 13162 15258
rect 13174 15206 13226 15258
rect 20982 15206 21034 15258
rect 21046 15206 21098 15258
rect 21110 15206 21162 15258
rect 21174 15206 21226 15258
rect 112 15104 164 15156
rect 3332 15147 3384 15156
rect 3332 15113 3341 15147
rect 3341 15113 3375 15147
rect 3375 15113 3384 15147
rect 3332 15104 3384 15113
rect 3792 15147 3844 15156
rect 3792 15113 3801 15147
rect 3801 15113 3835 15147
rect 3835 15113 3844 15147
rect 3792 15104 3844 15113
rect 4068 15147 4120 15156
rect 4068 15113 4077 15147
rect 4077 15113 4111 15147
rect 4111 15113 4120 15147
rect 4068 15104 4120 15113
rect 4804 15104 4856 15156
rect 6644 15147 6696 15156
rect 6644 15113 6653 15147
rect 6653 15113 6687 15147
rect 6687 15113 6696 15147
rect 6644 15104 6696 15113
rect 5264 14968 5316 15020
rect 6092 15036 6144 15088
rect 6276 15079 6328 15088
rect 6276 15045 6285 15079
rect 6285 15045 6319 15079
rect 6319 15045 6328 15079
rect 6276 15036 6328 15045
rect 2780 14943 2832 14952
rect 2780 14909 2789 14943
rect 2789 14909 2823 14943
rect 2823 14909 2832 14943
rect 2780 14900 2832 14909
rect 3332 14900 3384 14952
rect 4252 14900 4304 14952
rect 5448 14900 5500 14952
rect 7196 15011 7248 15020
rect 7196 14977 7205 15011
rect 7205 14977 7239 15011
rect 7239 14977 7248 15011
rect 7196 14968 7248 14977
rect 7288 15011 7340 15020
rect 7288 14977 7297 15011
rect 7297 14977 7331 15011
rect 7331 14977 7340 15011
rect 7288 14968 7340 14977
rect 2688 14832 2740 14884
rect 3608 14832 3660 14884
rect 6828 14875 6880 14884
rect 6828 14841 6837 14875
rect 6837 14841 6871 14875
rect 6871 14841 6880 14875
rect 6828 14832 6880 14841
rect 1860 14807 1912 14816
rect 1860 14773 1869 14807
rect 1869 14773 1903 14807
rect 1903 14773 1912 14807
rect 1860 14764 1912 14773
rect 4068 14764 4120 14816
rect 4436 14764 4488 14816
rect 4528 14764 4580 14816
rect 8982 14662 9034 14714
rect 9046 14662 9098 14714
rect 9110 14662 9162 14714
rect 9174 14662 9226 14714
rect 16982 14662 17034 14714
rect 17046 14662 17098 14714
rect 17110 14662 17162 14714
rect 17174 14662 17226 14714
rect 20 14560 72 14612
rect 4252 14560 4304 14612
rect 4804 14492 4856 14544
rect 6276 14560 6328 14612
rect 6828 14560 6880 14612
rect 7840 14560 7892 14612
rect 5540 14492 5592 14544
rect 7196 14492 7248 14544
rect 1676 14424 1728 14476
rect 2780 14467 2832 14476
rect 2780 14433 2789 14467
rect 2789 14433 2823 14467
rect 2823 14433 2832 14467
rect 2780 14424 2832 14433
rect 3884 14424 3936 14476
rect 4528 14424 4580 14476
rect 4712 14424 4764 14476
rect 6092 14467 6144 14476
rect 6092 14433 6101 14467
rect 6101 14433 6135 14467
rect 6135 14433 6144 14467
rect 6092 14424 6144 14433
rect 6276 14424 6328 14476
rect 5448 14399 5500 14408
rect 5448 14365 5457 14399
rect 5457 14365 5491 14399
rect 5491 14365 5500 14399
rect 5448 14356 5500 14365
rect 1952 14288 2004 14340
rect 4436 14288 4488 14340
rect 4252 14263 4304 14272
rect 4252 14229 4261 14263
rect 4261 14229 4295 14263
rect 4295 14229 4304 14263
rect 4252 14220 4304 14229
rect 4344 14220 4396 14272
rect 5264 14288 5316 14340
rect 4712 14263 4764 14272
rect 4712 14229 4721 14263
rect 4721 14229 4755 14263
rect 4755 14229 4764 14263
rect 4712 14220 4764 14229
rect 5724 14263 5776 14272
rect 5724 14229 5733 14263
rect 5733 14229 5767 14263
rect 5767 14229 5776 14263
rect 5724 14220 5776 14229
rect 6368 14220 6420 14272
rect 4982 14118 5034 14170
rect 5046 14118 5098 14170
rect 5110 14118 5162 14170
rect 5174 14118 5226 14170
rect 12982 14118 13034 14170
rect 13046 14118 13098 14170
rect 13110 14118 13162 14170
rect 13174 14118 13226 14170
rect 20982 14118 21034 14170
rect 21046 14118 21098 14170
rect 21110 14118 21162 14170
rect 21174 14118 21226 14170
rect 2780 14016 2832 14068
rect 4804 14016 4856 14068
rect 2136 13948 2188 14000
rect 1676 13855 1728 13864
rect 1676 13821 1685 13855
rect 1685 13821 1719 13855
rect 1719 13821 1728 13855
rect 1676 13812 1728 13821
rect 1952 13855 2004 13864
rect 1952 13821 1961 13855
rect 1961 13821 1995 13855
rect 1995 13821 2004 13855
rect 1952 13812 2004 13821
rect 4252 13880 4304 13932
rect 5632 14016 5684 14068
rect 6276 14016 6328 14068
rect 5264 13855 5316 13864
rect 5264 13821 5270 13855
rect 5270 13821 5316 13855
rect 2872 13787 2924 13796
rect 2872 13753 2881 13787
rect 2881 13753 2915 13787
rect 2915 13753 2924 13787
rect 5264 13812 5316 13821
rect 2872 13744 2924 13753
rect 4804 13744 4856 13796
rect 5540 13880 5592 13932
rect 6092 13880 6144 13932
rect 7472 13880 7524 13932
rect 7288 13855 7340 13864
rect 7288 13821 7297 13855
rect 7297 13821 7331 13855
rect 7331 13821 7340 13855
rect 7288 13812 7340 13821
rect 112 13676 164 13728
rect 3056 13719 3108 13728
rect 3056 13685 3065 13719
rect 3065 13685 3099 13719
rect 3099 13685 3108 13719
rect 3056 13676 3108 13685
rect 5908 13676 5960 13728
rect 6920 13719 6972 13728
rect 6920 13685 6929 13719
rect 6929 13685 6963 13719
rect 6963 13685 6972 13719
rect 6920 13676 6972 13685
rect 8982 13574 9034 13626
rect 9046 13574 9098 13626
rect 9110 13574 9162 13626
rect 9174 13574 9226 13626
rect 16982 13574 17034 13626
rect 17046 13574 17098 13626
rect 17110 13574 17162 13626
rect 17174 13574 17226 13626
rect 1584 13515 1636 13524
rect 1584 13481 1593 13515
rect 1593 13481 1627 13515
rect 1627 13481 1636 13515
rect 1584 13472 1636 13481
rect 1952 13515 2004 13524
rect 1952 13481 1961 13515
rect 1961 13481 1995 13515
rect 1995 13481 2004 13515
rect 1952 13472 2004 13481
rect 3884 13515 3936 13524
rect 112 13404 164 13456
rect 3884 13481 3893 13515
rect 3893 13481 3927 13515
rect 3927 13481 3936 13515
rect 3884 13472 3936 13481
rect 4344 13515 4396 13524
rect 4344 13481 4353 13515
rect 4353 13481 4387 13515
rect 4387 13481 4396 13515
rect 4344 13472 4396 13481
rect 4436 13472 4488 13524
rect 5540 13472 5592 13524
rect 7288 13472 7340 13524
rect 5632 13404 5684 13456
rect 6092 13404 6144 13456
rect 2136 13336 2188 13388
rect 2228 13336 2280 13388
rect 2872 13379 2924 13388
rect 2872 13345 2881 13379
rect 2881 13345 2915 13379
rect 2915 13345 2924 13379
rect 2872 13336 2924 13345
rect 4620 13336 4672 13388
rect 5264 13336 5316 13388
rect 7564 13379 7616 13388
rect 7564 13345 7573 13379
rect 7573 13345 7607 13379
rect 7607 13345 7616 13379
rect 7564 13336 7616 13345
rect 5448 13268 5500 13320
rect 7288 13311 7340 13320
rect 7288 13277 7297 13311
rect 7297 13277 7331 13311
rect 7331 13277 7340 13311
rect 7288 13268 7340 13277
rect 2780 13200 2832 13252
rect 7472 13200 7524 13252
rect 3424 13175 3476 13184
rect 3424 13141 3433 13175
rect 3433 13141 3467 13175
rect 3467 13141 3476 13175
rect 3424 13132 3476 13141
rect 5356 13132 5408 13184
rect 4982 13030 5034 13082
rect 5046 13030 5098 13082
rect 5110 13030 5162 13082
rect 5174 13030 5226 13082
rect 12982 13030 13034 13082
rect 13046 13030 13098 13082
rect 13110 13030 13162 13082
rect 13174 13030 13226 13082
rect 20982 13030 21034 13082
rect 21046 13030 21098 13082
rect 21110 13030 21162 13082
rect 21174 13030 21226 13082
rect 1860 12928 1912 12980
rect 3240 12928 3292 12980
rect 4804 12971 4856 12980
rect 4804 12937 4813 12971
rect 4813 12937 4847 12971
rect 4847 12937 4856 12971
rect 4804 12928 4856 12937
rect 2228 12724 2280 12776
rect 2780 12767 2832 12776
rect 2780 12733 2789 12767
rect 2789 12733 2823 12767
rect 2823 12733 2832 12767
rect 2780 12724 2832 12733
rect 2872 12724 2924 12776
rect 4252 12724 4304 12776
rect 4712 12792 4764 12844
rect 5632 12928 5684 12980
rect 7564 12928 7616 12980
rect 4620 12656 4672 12708
rect 5356 12724 5408 12776
rect 7380 12767 7432 12776
rect 7380 12733 7389 12767
rect 7389 12733 7423 12767
rect 7423 12733 7432 12767
rect 7380 12724 7432 12733
rect 5632 12656 5684 12708
rect 6092 12656 6144 12708
rect 20 12588 72 12640
rect 5540 12631 5592 12640
rect 5540 12597 5549 12631
rect 5549 12597 5583 12631
rect 5583 12597 5592 12631
rect 5540 12588 5592 12597
rect 6368 12631 6420 12640
rect 6368 12597 6377 12631
rect 6377 12597 6411 12631
rect 6411 12597 6420 12631
rect 6368 12588 6420 12597
rect 8982 12486 9034 12538
rect 9046 12486 9098 12538
rect 9110 12486 9162 12538
rect 9174 12486 9226 12538
rect 16982 12486 17034 12538
rect 17046 12486 17098 12538
rect 17110 12486 17162 12538
rect 17174 12486 17226 12538
rect 112 12384 164 12436
rect 204 12316 256 12368
rect 5448 12427 5500 12436
rect 5448 12393 5457 12427
rect 5457 12393 5491 12427
rect 5491 12393 5500 12427
rect 5448 12384 5500 12393
rect 6644 12384 6696 12436
rect 7380 12384 7432 12436
rect 3700 12316 3752 12368
rect 4804 12316 4856 12368
rect 6092 12359 6144 12368
rect 6092 12325 6101 12359
rect 6101 12325 6135 12359
rect 6135 12325 6144 12359
rect 6092 12316 6144 12325
rect 1676 12248 1728 12300
rect 2872 12291 2924 12300
rect 2872 12257 2881 12291
rect 2881 12257 2915 12291
rect 2915 12257 2924 12291
rect 2872 12248 2924 12257
rect 4252 12291 4304 12300
rect 4252 12257 4261 12291
rect 4261 12257 4295 12291
rect 4295 12257 4304 12291
rect 4252 12248 4304 12257
rect 4528 12291 4580 12300
rect 4528 12257 4537 12291
rect 4537 12257 4571 12291
rect 4571 12257 4580 12291
rect 4528 12248 4580 12257
rect 6184 12248 6236 12300
rect 7564 12248 7616 12300
rect 2688 12180 2740 12232
rect 3424 12223 3476 12232
rect 3424 12189 3433 12223
rect 3433 12189 3467 12223
rect 3467 12189 3476 12223
rect 3424 12180 3476 12189
rect 6460 12223 6512 12232
rect 6460 12189 6469 12223
rect 6469 12189 6503 12223
rect 6503 12189 6512 12223
rect 6460 12180 6512 12189
rect 2136 12112 2188 12164
rect 3516 12112 3568 12164
rect 4620 12112 4672 12164
rect 6368 12155 6420 12164
rect 6368 12121 6377 12155
rect 6377 12121 6411 12155
rect 6411 12121 6420 12155
rect 6368 12112 6420 12121
rect 7104 12112 7156 12164
rect 7932 12155 7984 12164
rect 7932 12121 7941 12155
rect 7941 12121 7975 12155
rect 7975 12121 7984 12155
rect 7932 12112 7984 12121
rect 1584 12087 1636 12096
rect 1584 12053 1593 12087
rect 1593 12053 1627 12087
rect 1627 12053 1636 12087
rect 1584 12044 1636 12053
rect 1952 12087 2004 12096
rect 1952 12053 1961 12087
rect 1961 12053 1995 12087
rect 1995 12053 2004 12087
rect 1952 12044 2004 12053
rect 2320 12087 2372 12096
rect 2320 12053 2329 12087
rect 2329 12053 2363 12087
rect 2363 12053 2372 12087
rect 2320 12044 2372 12053
rect 5356 12044 5408 12096
rect 6736 12087 6788 12096
rect 6736 12053 6745 12087
rect 6745 12053 6779 12087
rect 6779 12053 6788 12087
rect 6736 12044 6788 12053
rect 8024 12044 8076 12096
rect 4982 11942 5034 11994
rect 5046 11942 5098 11994
rect 5110 11942 5162 11994
rect 5174 11942 5226 11994
rect 12982 11942 13034 11994
rect 13046 11942 13098 11994
rect 13110 11942 13162 11994
rect 13174 11942 13226 11994
rect 20982 11942 21034 11994
rect 21046 11942 21098 11994
rect 21110 11942 21162 11994
rect 21174 11942 21226 11994
rect 2872 11840 2924 11892
rect 4528 11840 4580 11892
rect 4620 11840 4672 11892
rect 5356 11840 5408 11892
rect 6184 11883 6236 11892
rect 6184 11849 6193 11883
rect 6193 11849 6227 11883
rect 6227 11849 6236 11883
rect 6184 11840 6236 11849
rect 6644 11883 6696 11892
rect 6644 11849 6653 11883
rect 6653 11849 6687 11883
rect 6687 11849 6696 11883
rect 6644 11840 6696 11849
rect 7288 11840 7340 11892
rect 7380 11840 7432 11892
rect 1952 11704 2004 11756
rect 6460 11772 6512 11824
rect 7104 11815 7156 11824
rect 7104 11781 7113 11815
rect 7113 11781 7147 11815
rect 7147 11781 7156 11815
rect 7104 11772 7156 11781
rect 7564 11772 7616 11824
rect 1676 11679 1728 11688
rect 1676 11645 1685 11679
rect 1685 11645 1719 11679
rect 1719 11645 1728 11679
rect 1676 11636 1728 11645
rect 2320 11636 2372 11688
rect 2780 11636 2832 11688
rect 3516 11679 3568 11688
rect 3516 11645 3525 11679
rect 3525 11645 3559 11679
rect 3559 11645 3568 11679
rect 3516 11636 3568 11645
rect 20 11568 72 11620
rect 112 11500 164 11552
rect 5724 11636 5776 11688
rect 6092 11636 6144 11688
rect 6644 11636 6696 11688
rect 7012 11636 7064 11688
rect 4804 11568 4856 11620
rect 4528 11543 4580 11552
rect 4528 11509 4537 11543
rect 4537 11509 4571 11543
rect 4571 11509 4580 11543
rect 4528 11500 4580 11509
rect 6920 11500 6972 11552
rect 8982 11398 9034 11450
rect 9046 11398 9098 11450
rect 9110 11398 9162 11450
rect 9174 11398 9226 11450
rect 16982 11398 17034 11450
rect 17046 11398 17098 11450
rect 17110 11398 17162 11450
rect 17174 11398 17226 11450
rect 112 11296 164 11348
rect 2688 11296 2740 11348
rect 4528 11296 4580 11348
rect 6460 11296 6512 11348
rect 7932 11296 7984 11348
rect 1676 11203 1728 11212
rect 1676 11169 1685 11203
rect 1685 11169 1719 11203
rect 1719 11169 1728 11203
rect 1676 11160 1728 11169
rect 3516 11228 3568 11280
rect 5724 11271 5776 11280
rect 5724 11237 5733 11271
rect 5733 11237 5767 11271
rect 5767 11237 5776 11271
rect 5724 11228 5776 11237
rect 2780 11160 2832 11212
rect 4252 11160 4304 11212
rect 4620 11203 4672 11212
rect 4620 11169 4629 11203
rect 4629 11169 4663 11203
rect 4663 11169 4672 11203
rect 4620 11160 4672 11169
rect 6184 11160 6236 11212
rect 7196 11160 7248 11212
rect 7472 11160 7524 11212
rect 6092 11135 6144 11144
rect 6092 11101 6101 11135
rect 6101 11101 6135 11135
rect 6135 11101 6144 11135
rect 6092 11092 6144 11101
rect 6460 11092 6512 11144
rect 4160 11024 4212 11076
rect 7012 11024 7064 11076
rect 3148 10999 3200 11008
rect 3148 10965 3157 10999
rect 3157 10965 3191 10999
rect 3191 10965 3200 10999
rect 3148 10956 3200 10965
rect 4252 10999 4304 11008
rect 4252 10965 4261 10999
rect 4261 10965 4295 10999
rect 4295 10965 4304 10999
rect 4252 10956 4304 10965
rect 6368 10956 6420 11008
rect 7472 10999 7524 11008
rect 7472 10965 7481 10999
rect 7481 10965 7515 10999
rect 7515 10965 7524 10999
rect 7472 10956 7524 10965
rect 4982 10854 5034 10906
rect 5046 10854 5098 10906
rect 5110 10854 5162 10906
rect 5174 10854 5226 10906
rect 12982 10854 13034 10906
rect 13046 10854 13098 10906
rect 13110 10854 13162 10906
rect 13174 10854 13226 10906
rect 20982 10854 21034 10906
rect 21046 10854 21098 10906
rect 21110 10854 21162 10906
rect 21174 10854 21226 10906
rect 1676 10752 1728 10804
rect 2780 10795 2832 10804
rect 2780 10761 2789 10795
rect 2789 10761 2823 10795
rect 2823 10761 2832 10795
rect 2780 10752 2832 10761
rect 4160 10752 4212 10804
rect 6092 10795 6144 10804
rect 6092 10761 6101 10795
rect 6101 10761 6135 10795
rect 6135 10761 6144 10795
rect 6092 10752 6144 10761
rect 6368 10795 6420 10804
rect 6368 10761 6377 10795
rect 6377 10761 6411 10795
rect 6411 10761 6420 10795
rect 6368 10752 6420 10761
rect 7288 10795 7340 10804
rect 7288 10761 7297 10795
rect 7297 10761 7331 10795
rect 7331 10761 7340 10795
rect 7288 10752 7340 10761
rect 7564 10752 7616 10804
rect 2596 10684 2648 10736
rect 204 10616 256 10668
rect 2504 10616 2556 10668
rect 1676 10591 1728 10600
rect 1676 10557 1685 10591
rect 1685 10557 1719 10591
rect 1719 10557 1728 10591
rect 1676 10548 1728 10557
rect 2320 10548 2372 10600
rect 2872 10548 2924 10600
rect 3884 10616 3936 10668
rect 4528 10616 4580 10668
rect 3792 10548 3844 10600
rect 20 10480 72 10532
rect 112 10480 164 10532
rect 4988 10523 5040 10532
rect 4988 10489 4997 10523
rect 4997 10489 5031 10523
rect 5031 10489 5040 10523
rect 4988 10480 5040 10489
rect 6736 10548 6788 10600
rect 4620 10412 4672 10464
rect 5356 10412 5408 10464
rect 8982 10310 9034 10362
rect 9046 10310 9098 10362
rect 9110 10310 9162 10362
rect 9174 10310 9226 10362
rect 16982 10310 17034 10362
rect 17046 10310 17098 10362
rect 17110 10310 17162 10362
rect 17174 10310 17226 10362
rect 1676 10208 1728 10260
rect 2320 10251 2372 10260
rect 2320 10217 2329 10251
rect 2329 10217 2363 10251
rect 2363 10217 2372 10251
rect 2320 10208 2372 10217
rect 2504 10251 2556 10260
rect 2504 10217 2513 10251
rect 2513 10217 2547 10251
rect 2547 10217 2556 10251
rect 2504 10208 2556 10217
rect 3516 10208 3568 10260
rect 4252 10251 4304 10260
rect 4252 10217 4261 10251
rect 4261 10217 4295 10251
rect 4295 10217 4304 10251
rect 4252 10208 4304 10217
rect 4528 10251 4580 10260
rect 4528 10217 4537 10251
rect 4537 10217 4571 10251
rect 4571 10217 4580 10251
rect 4528 10208 4580 10217
rect 4988 10251 5040 10260
rect 4988 10217 4997 10251
rect 4997 10217 5031 10251
rect 5031 10217 5040 10251
rect 4988 10208 5040 10217
rect 5724 10208 5776 10260
rect 1400 10115 1452 10124
rect 1400 10081 1409 10115
rect 1409 10081 1443 10115
rect 1443 10081 1452 10115
rect 1400 10072 1452 10081
rect 4160 10140 4212 10192
rect 3792 10004 3844 10056
rect 4712 10072 4764 10124
rect 6000 10140 6052 10192
rect 6184 10183 6236 10192
rect 6184 10149 6193 10183
rect 6193 10149 6227 10183
rect 6227 10149 6236 10183
rect 6184 10140 6236 10149
rect 5724 10072 5776 10124
rect 6644 10115 6696 10124
rect 6644 10081 6653 10115
rect 6653 10081 6687 10115
rect 6687 10081 6696 10115
rect 6644 10072 6696 10081
rect 7288 10072 7340 10124
rect 4620 10004 4672 10056
rect 4528 9936 4580 9988
rect 4804 9936 4856 9988
rect 5356 9936 5408 9988
rect 4252 9868 4304 9920
rect 6736 9979 6788 9988
rect 6736 9945 6745 9979
rect 6745 9945 6779 9979
rect 6779 9945 6788 9979
rect 6736 9936 6788 9945
rect 4982 9766 5034 9818
rect 5046 9766 5098 9818
rect 5110 9766 5162 9818
rect 5174 9766 5226 9818
rect 12982 9766 13034 9818
rect 13046 9766 13098 9818
rect 13110 9766 13162 9818
rect 13174 9766 13226 9818
rect 20982 9766 21034 9818
rect 21046 9766 21098 9818
rect 21110 9766 21162 9818
rect 21174 9766 21226 9818
rect 1400 9664 1452 9716
rect 2688 9707 2740 9716
rect 2688 9673 2697 9707
rect 2697 9673 2731 9707
rect 2731 9673 2740 9707
rect 2688 9664 2740 9673
rect 4712 9664 4764 9716
rect 5356 9664 5408 9716
rect 6736 9664 6788 9716
rect 1584 9596 1636 9648
rect 4068 9596 4120 9648
rect 5172 9596 5224 9648
rect 3056 9528 3108 9580
rect 6644 9528 6696 9580
rect 3792 9503 3844 9512
rect 1860 9392 1912 9444
rect 3792 9469 3801 9503
rect 3801 9469 3835 9503
rect 3835 9469 3844 9503
rect 3792 9460 3844 9469
rect 5080 9503 5132 9512
rect 5080 9469 5089 9503
rect 5089 9469 5123 9503
rect 5123 9469 5132 9503
rect 5080 9460 5132 9469
rect 5172 9503 5224 9512
rect 5172 9469 5181 9503
rect 5181 9469 5215 9503
rect 5215 9469 5224 9503
rect 5172 9460 5224 9469
rect 5724 9460 5776 9512
rect 3148 9392 3200 9444
rect 112 9324 164 9376
rect 3332 9367 3384 9376
rect 3332 9333 3341 9367
rect 3341 9333 3375 9367
rect 3375 9333 3384 9367
rect 3332 9324 3384 9333
rect 4988 9324 5040 9376
rect 7288 9324 7340 9376
rect 8982 9222 9034 9274
rect 9046 9222 9098 9274
rect 9110 9222 9162 9274
rect 9174 9222 9226 9274
rect 16982 9222 17034 9274
rect 17046 9222 17098 9274
rect 17110 9222 17162 9274
rect 17174 9222 17226 9274
rect 112 9120 164 9172
rect 3056 9163 3108 9172
rect 3056 9129 3065 9163
rect 3065 9129 3099 9163
rect 3099 9129 3108 9163
rect 3056 9120 3108 9129
rect 3148 9120 3200 9172
rect 4712 9120 4764 9172
rect 2688 9052 2740 9104
rect 6644 9163 6696 9172
rect 6644 9129 6653 9163
rect 6653 9129 6687 9163
rect 6687 9129 6696 9163
rect 6644 9120 6696 9129
rect 5080 9095 5132 9104
rect 5080 9061 5089 9095
rect 5089 9061 5123 9095
rect 5123 9061 5132 9095
rect 5080 9052 5132 9061
rect 5356 9052 5408 9104
rect 1860 9027 1912 9036
rect 1860 8993 1869 9027
rect 1869 8993 1903 9027
rect 1903 8993 1912 9027
rect 1860 8984 1912 8993
rect 2044 9027 2096 9036
rect 2044 8993 2053 9027
rect 2053 8993 2087 9027
rect 2087 8993 2096 9027
rect 2044 8984 2096 8993
rect 3516 8984 3568 9036
rect 4620 8984 4672 9036
rect 4988 8984 5040 9036
rect 4252 8916 4304 8968
rect 4804 8916 4856 8968
rect 5724 8984 5776 9036
rect 5172 8848 5224 8900
rect 5540 8848 5592 8900
rect 4982 8678 5034 8730
rect 5046 8678 5098 8730
rect 5110 8678 5162 8730
rect 5174 8678 5226 8730
rect 12982 8678 13034 8730
rect 13046 8678 13098 8730
rect 13110 8678 13162 8730
rect 13174 8678 13226 8730
rect 20982 8678 21034 8730
rect 21046 8678 21098 8730
rect 21110 8678 21162 8730
rect 21174 8678 21226 8730
rect 4804 8619 4856 8628
rect 4804 8585 4813 8619
rect 4813 8585 4847 8619
rect 4847 8585 4856 8619
rect 4804 8576 4856 8585
rect 5356 8619 5408 8628
rect 5356 8585 5365 8619
rect 5365 8585 5399 8619
rect 5399 8585 5408 8619
rect 5356 8576 5408 8585
rect 5724 8508 5776 8560
rect 2872 8440 2924 8492
rect 4804 8440 4856 8492
rect 2044 8415 2096 8424
rect 2044 8381 2053 8415
rect 2053 8381 2087 8415
rect 2087 8381 2096 8415
rect 2044 8372 2096 8381
rect 3608 8415 3660 8424
rect 20 8304 72 8356
rect 3608 8381 3617 8415
rect 3617 8381 3651 8415
rect 3651 8381 3660 8415
rect 3608 8372 3660 8381
rect 112 8236 164 8288
rect 3516 8304 3568 8356
rect 6184 8304 6236 8356
rect 3608 8236 3660 8288
rect 3976 8236 4028 8288
rect 5264 8236 5316 8288
rect 8982 8134 9034 8186
rect 9046 8134 9098 8186
rect 9110 8134 9162 8186
rect 9174 8134 9226 8186
rect 16982 8134 17034 8186
rect 17046 8134 17098 8186
rect 17110 8134 17162 8186
rect 17174 8134 17226 8186
rect 112 8032 164 8084
rect 1860 8032 1912 8084
rect 3516 8032 3568 8084
rect 5264 8075 5316 8084
rect 5264 8041 5273 8075
rect 5273 8041 5307 8075
rect 5307 8041 5316 8075
rect 5264 8032 5316 8041
rect 5540 8007 5592 8016
rect 5540 7973 5549 8007
rect 5549 7973 5583 8007
rect 5583 7973 5592 8007
rect 5540 7964 5592 7973
rect 1584 7939 1636 7948
rect 1584 7905 1593 7939
rect 1593 7905 1627 7939
rect 1627 7905 1636 7939
rect 1584 7896 1636 7905
rect 2044 7939 2096 7948
rect 2044 7905 2053 7939
rect 2053 7905 2087 7939
rect 2087 7905 2096 7939
rect 2044 7896 2096 7905
rect 2320 7896 2372 7948
rect 4344 7896 4396 7948
rect 4620 7939 4672 7948
rect 4620 7905 4629 7939
rect 4629 7905 4663 7939
rect 4663 7905 4672 7939
rect 4620 7896 4672 7905
rect 4712 7896 4764 7948
rect 6092 7939 6144 7948
rect 6092 7905 6101 7939
rect 6101 7905 6135 7939
rect 6135 7905 6144 7939
rect 6092 7896 6144 7905
rect 6920 7896 6972 7948
rect 2872 7760 2924 7812
rect 3884 7760 3936 7812
rect 6184 7760 6236 7812
rect 4982 7590 5034 7642
rect 5046 7590 5098 7642
rect 5110 7590 5162 7642
rect 5174 7590 5226 7642
rect 12982 7590 13034 7642
rect 13046 7590 13098 7642
rect 13110 7590 13162 7642
rect 13174 7590 13226 7642
rect 20982 7590 21034 7642
rect 21046 7590 21098 7642
rect 21110 7590 21162 7642
rect 21174 7590 21226 7642
rect 2044 7488 2096 7540
rect 4344 7531 4396 7540
rect 4344 7497 4353 7531
rect 4353 7497 4387 7531
rect 4387 7497 4396 7531
rect 4344 7488 4396 7497
rect 4712 7488 4764 7540
rect 6092 7531 6144 7540
rect 6092 7497 6101 7531
rect 6101 7497 6135 7531
rect 6135 7497 6144 7531
rect 6092 7488 6144 7497
rect 7288 7531 7340 7540
rect 7288 7497 7297 7531
rect 7297 7497 7331 7531
rect 7331 7497 7340 7531
rect 7288 7488 7340 7497
rect 1860 7284 1912 7336
rect 1952 7284 2004 7336
rect 3700 7284 3752 7336
rect 3884 7327 3936 7336
rect 3884 7293 3893 7327
rect 3893 7293 3927 7327
rect 3927 7293 3936 7327
rect 3884 7284 3936 7293
rect 8024 7420 8076 7472
rect 12072 7284 12124 7336
rect 1584 7191 1636 7200
rect 1584 7157 1593 7191
rect 1593 7157 1627 7191
rect 1627 7157 1636 7191
rect 1584 7148 1636 7157
rect 3424 7191 3476 7200
rect 3424 7157 3433 7191
rect 3433 7157 3467 7191
rect 3467 7157 3476 7191
rect 3424 7148 3476 7157
rect 3608 7148 3660 7200
rect 8982 7046 9034 7098
rect 9046 7046 9098 7098
rect 9110 7046 9162 7098
rect 9174 7046 9226 7098
rect 16982 7046 17034 7098
rect 17046 7046 17098 7098
rect 17110 7046 17162 7098
rect 17174 7046 17226 7098
rect 112 6944 164 6996
rect 1860 6944 1912 6996
rect 3056 6944 3108 6996
rect 3700 6987 3752 6996
rect 3700 6953 3709 6987
rect 3709 6953 3743 6987
rect 3743 6953 3752 6987
rect 3700 6944 3752 6953
rect 296 6876 348 6928
rect 1952 6851 2004 6860
rect 1952 6817 1961 6851
rect 1961 6817 1995 6851
rect 1995 6817 2004 6851
rect 1952 6808 2004 6817
rect 2872 6851 2924 6860
rect 2872 6817 2881 6851
rect 2881 6817 2915 6851
rect 2915 6817 2924 6851
rect 2872 6808 2924 6817
rect 4528 6808 4580 6860
rect 5632 6851 5684 6860
rect 3884 6604 3936 6656
rect 5632 6817 5641 6851
rect 5641 6817 5675 6851
rect 5675 6817 5684 6851
rect 5632 6808 5684 6817
rect 4712 6604 4764 6656
rect 4982 6502 5034 6554
rect 5046 6502 5098 6554
rect 5110 6502 5162 6554
rect 5174 6502 5226 6554
rect 12982 6502 13034 6554
rect 13046 6502 13098 6554
rect 13110 6502 13162 6554
rect 13174 6502 13226 6554
rect 20982 6502 21034 6554
rect 21046 6502 21098 6554
rect 21110 6502 21162 6554
rect 21174 6502 21226 6554
rect 4528 6400 4580 6452
rect 5632 6443 5684 6452
rect 5632 6409 5641 6443
rect 5641 6409 5675 6443
rect 5675 6409 5684 6443
rect 5632 6400 5684 6409
rect 20 6264 72 6316
rect 1676 6239 1728 6248
rect 1676 6205 1685 6239
rect 1685 6205 1719 6239
rect 1719 6205 1728 6239
rect 1676 6196 1728 6205
rect 3608 6239 3660 6248
rect 3608 6205 3617 6239
rect 3617 6205 3651 6239
rect 3651 6205 3660 6239
rect 3608 6196 3660 6205
rect 3976 6239 4028 6248
rect 3976 6205 3985 6239
rect 3985 6205 4019 6239
rect 4019 6205 4028 6239
rect 3976 6196 4028 6205
rect 112 6060 164 6112
rect 4712 6103 4764 6112
rect 4712 6069 4721 6103
rect 4721 6069 4755 6103
rect 4755 6069 4764 6103
rect 4712 6060 4764 6069
rect 8982 5958 9034 6010
rect 9046 5958 9098 6010
rect 9110 5958 9162 6010
rect 9174 5958 9226 6010
rect 16982 5958 17034 6010
rect 17046 5958 17098 6010
rect 17110 5958 17162 6010
rect 17174 5958 17226 6010
rect 112 5856 164 5908
rect 1860 5856 1912 5908
rect 2872 5856 2924 5908
rect 3056 5899 3108 5908
rect 3056 5865 3065 5899
rect 3065 5865 3099 5899
rect 3099 5865 3108 5899
rect 3056 5856 3108 5865
rect 3976 5856 4028 5908
rect 204 5788 256 5840
rect 1492 5720 1544 5772
rect 1860 5763 1912 5772
rect 1860 5729 1869 5763
rect 1869 5729 1903 5763
rect 1903 5729 1912 5763
rect 1860 5720 1912 5729
rect 2044 5763 2096 5772
rect 2044 5729 2053 5763
rect 2053 5729 2087 5763
rect 2087 5729 2096 5763
rect 2044 5720 2096 5729
rect 3240 5720 3292 5772
rect 4436 5720 4488 5772
rect 1676 5652 1728 5704
rect 3516 5652 3568 5704
rect 4712 5720 4764 5772
rect 4068 5584 4120 5636
rect 4982 5414 5034 5466
rect 5046 5414 5098 5466
rect 5110 5414 5162 5466
rect 5174 5414 5226 5466
rect 12982 5414 13034 5466
rect 13046 5414 13098 5466
rect 13110 5414 13162 5466
rect 13174 5414 13226 5466
rect 20982 5414 21034 5466
rect 21046 5414 21098 5466
rect 21110 5414 21162 5466
rect 21174 5414 21226 5466
rect 4436 5355 4488 5364
rect 4436 5321 4445 5355
rect 4445 5321 4479 5355
rect 4479 5321 4488 5355
rect 4436 5312 4488 5321
rect 1676 5151 1728 5160
rect 1676 5117 1685 5151
rect 1685 5117 1719 5151
rect 1719 5117 1728 5151
rect 1676 5108 1728 5117
rect 2044 5151 2096 5160
rect 2044 5117 2053 5151
rect 2053 5117 2087 5151
rect 2087 5117 2096 5151
rect 2044 5108 2096 5117
rect 2872 5151 2924 5160
rect 2872 5117 2881 5151
rect 2881 5117 2915 5151
rect 2915 5117 2924 5151
rect 2872 5108 2924 5117
rect 3056 5151 3108 5160
rect 3056 5117 3065 5151
rect 3065 5117 3099 5151
rect 3099 5117 3108 5151
rect 3056 5108 3108 5117
rect 4528 5244 4580 5296
rect 5448 5312 5500 5364
rect 20 5040 72 5092
rect 112 4972 164 5024
rect 4068 5015 4120 5024
rect 4068 4981 4077 5015
rect 4077 4981 4111 5015
rect 4111 4981 4120 5015
rect 4068 4972 4120 4981
rect 8982 4870 9034 4922
rect 9046 4870 9098 4922
rect 9110 4870 9162 4922
rect 9174 4870 9226 4922
rect 16982 4870 17034 4922
rect 17046 4870 17098 4922
rect 17110 4870 17162 4922
rect 17174 4870 17226 4922
rect 20 4768 72 4820
rect 2872 4768 2924 4820
rect 3516 4811 3568 4820
rect 3516 4777 3525 4811
rect 3525 4777 3559 4811
rect 3559 4777 3568 4811
rect 3516 4768 3568 4777
rect 3976 4768 4028 4820
rect 4160 4811 4212 4820
rect 4160 4777 4169 4811
rect 4169 4777 4203 4811
rect 4203 4777 4212 4811
rect 4160 4768 4212 4777
rect 2136 4675 2188 4684
rect 2136 4641 2145 4675
rect 2145 4641 2179 4675
rect 2179 4641 2188 4675
rect 2136 4632 2188 4641
rect 2780 4632 2832 4684
rect 3056 4632 3108 4684
rect 4344 4632 4396 4684
rect 4528 4675 4580 4684
rect 4528 4641 4537 4675
rect 4537 4641 4571 4675
rect 4571 4641 4580 4675
rect 4528 4632 4580 4641
rect 4982 4326 5034 4378
rect 5046 4326 5098 4378
rect 5110 4326 5162 4378
rect 5174 4326 5226 4378
rect 12982 4326 13034 4378
rect 13046 4326 13098 4378
rect 13110 4326 13162 4378
rect 13174 4326 13226 4378
rect 20982 4326 21034 4378
rect 21046 4326 21098 4378
rect 21110 4326 21162 4378
rect 21174 4326 21226 4378
rect 112 4088 164 4140
rect 1492 4020 1544 4072
rect 2136 4063 2188 4072
rect 2136 4029 2145 4063
rect 2145 4029 2179 4063
rect 2179 4029 2188 4063
rect 2136 4020 2188 4029
rect 3884 4020 3936 4072
rect 4528 4156 4580 4208
rect 4344 4088 4396 4140
rect 4436 4020 4488 4072
rect 112 3884 164 3936
rect 8982 3782 9034 3834
rect 9046 3782 9098 3834
rect 9110 3782 9162 3834
rect 9174 3782 9226 3834
rect 16982 3782 17034 3834
rect 17046 3782 17098 3834
rect 17110 3782 17162 3834
rect 17174 3782 17226 3834
rect 20 3680 72 3732
rect 3516 3723 3568 3732
rect 3516 3689 3525 3723
rect 3525 3689 3559 3723
rect 3559 3689 3568 3723
rect 3516 3680 3568 3689
rect 3884 3723 3936 3732
rect 3884 3689 3893 3723
rect 3893 3689 3927 3723
rect 3927 3689 3936 3723
rect 3884 3680 3936 3689
rect 1492 3544 1544 3596
rect 2228 3587 2280 3596
rect 2228 3553 2237 3587
rect 2237 3553 2271 3587
rect 2271 3553 2280 3587
rect 2228 3544 2280 3553
rect 4620 3587 4672 3596
rect 4620 3553 4629 3587
rect 4629 3553 4663 3587
rect 4663 3553 4672 3587
rect 4620 3544 4672 3553
rect 388 3476 440 3528
rect 4982 3238 5034 3290
rect 5046 3238 5098 3290
rect 5110 3238 5162 3290
rect 5174 3238 5226 3290
rect 12982 3238 13034 3290
rect 13046 3238 13098 3290
rect 13110 3238 13162 3290
rect 13174 3238 13226 3290
rect 20982 3238 21034 3290
rect 21046 3238 21098 3290
rect 21110 3238 21162 3290
rect 21174 3238 21226 3290
rect 4344 3136 4396 3188
rect 4620 3068 4672 3120
rect 4068 3000 4120 3052
rect 1768 2975 1820 2984
rect 1768 2941 1777 2975
rect 1777 2941 1811 2975
rect 1811 2941 1820 2975
rect 1768 2932 1820 2941
rect 2136 2975 2188 2984
rect 2136 2941 2145 2975
rect 2145 2941 2179 2975
rect 2179 2941 2188 2975
rect 2136 2932 2188 2941
rect 3884 2975 3936 2984
rect 3884 2941 3893 2975
rect 3893 2941 3927 2975
rect 3927 2941 3936 2975
rect 3884 2932 3936 2941
rect 5908 3136 5960 3188
rect 112 2796 164 2848
rect 2228 2796 2280 2848
rect 3792 2839 3844 2848
rect 3792 2805 3801 2839
rect 3801 2805 3835 2839
rect 3835 2805 3844 2839
rect 3792 2796 3844 2805
rect 8982 2694 9034 2746
rect 9046 2694 9098 2746
rect 9110 2694 9162 2746
rect 9174 2694 9226 2746
rect 16982 2694 17034 2746
rect 17046 2694 17098 2746
rect 17110 2694 17162 2746
rect 17174 2694 17226 2746
rect 112 2592 164 2644
rect 3516 2592 3568 2644
rect 2780 2524 2832 2576
rect 1768 2499 1820 2508
rect 1768 2465 1777 2499
rect 1777 2465 1811 2499
rect 1811 2465 1820 2499
rect 1768 2456 1820 2465
rect 2228 2499 2280 2508
rect 2228 2465 2237 2499
rect 2237 2465 2271 2499
rect 2271 2465 2280 2499
rect 2228 2456 2280 2465
rect 4620 2499 4672 2508
rect 4620 2465 4629 2499
rect 4629 2465 4663 2499
rect 4663 2465 4672 2499
rect 4620 2456 4672 2465
rect 388 2320 440 2372
rect 4982 2150 5034 2202
rect 5046 2150 5098 2202
rect 5110 2150 5162 2202
rect 5174 2150 5226 2202
rect 12982 2150 13034 2202
rect 13046 2150 13098 2202
rect 13110 2150 13162 2202
rect 13174 2150 13226 2202
rect 20982 2150 21034 2202
rect 21046 2150 21098 2202
rect 21110 2150 21162 2202
rect 21174 2150 21226 2202
rect 112 1300 164 1352
rect 3792 1300 3844 1352
<< metal2 >>
rect 110 23760 166 23769
rect 166 23718 336 23746
rect 110 23695 166 23704
rect 18 23352 74 23361
rect 18 23287 74 23296
rect 32 20466 60 23287
rect 110 22944 166 22953
rect 166 22902 244 22930
rect 110 22879 166 22888
rect 110 22536 166 22545
rect 110 22471 166 22480
rect 124 21894 152 22471
rect 112 21888 164 21894
rect 112 21830 164 21836
rect 110 21720 166 21729
rect 110 21655 166 21664
rect 124 21418 152 21655
rect 112 21412 164 21418
rect 112 21354 164 21360
rect 110 21312 166 21321
rect 110 21247 166 21256
rect 20 20460 72 20466
rect 20 20402 72 20408
rect 124 20262 152 21247
rect 112 20256 164 20262
rect 112 20198 164 20204
rect 110 19816 166 19825
rect 110 19751 166 19760
rect 18 18592 74 18601
rect 18 18527 74 18536
rect 32 17882 60 18527
rect 124 18290 152 19751
rect 216 19378 244 22902
rect 204 19372 256 19378
rect 204 19314 256 19320
rect 308 19242 336 23718
rect 1950 23588 2006 24000
rect 5906 23610 5962 24000
rect 9954 23610 10010 24000
rect 13910 23610 13966 24000
rect 17958 23610 18014 24000
rect 1950 23536 1952 23588
rect 2004 23536 2006 23588
rect 1950 23520 2006 23536
rect 2596 23588 2648 23594
rect 2596 23530 2648 23536
rect 5906 23582 6040 23610
rect 1964 23499 1992 23520
rect 2136 21344 2188 21350
rect 2136 21286 2188 21292
rect 2148 21010 2176 21286
rect 2136 21004 2188 21010
rect 2136 20946 2188 20952
rect 386 20904 442 20913
rect 386 20839 442 20848
rect 400 20058 428 20839
rect 2148 20806 2176 20946
rect 2504 20936 2556 20942
rect 2504 20878 2556 20884
rect 2136 20800 2188 20806
rect 2136 20742 2188 20748
rect 2148 20398 2176 20742
rect 2136 20392 2188 20398
rect 2136 20334 2188 20340
rect 1766 20088 1822 20097
rect 388 20052 440 20058
rect 1766 20023 1822 20032
rect 388 19994 440 20000
rect 1676 19916 1728 19922
rect 1676 19858 1728 19864
rect 1688 19310 1716 19858
rect 1676 19304 1728 19310
rect 1676 19246 1728 19252
rect 296 19236 348 19242
rect 296 19178 348 19184
rect 1780 18970 1808 20023
rect 2148 19922 2176 20334
rect 2516 20262 2544 20878
rect 2412 20256 2464 20262
rect 2412 20198 2464 20204
rect 2504 20256 2556 20262
rect 2504 20198 2556 20204
rect 2136 19916 2188 19922
rect 2136 19858 2188 19864
rect 2148 19514 2176 19858
rect 2136 19508 2188 19514
rect 2136 19450 2188 19456
rect 2424 19174 2452 20198
rect 2516 19718 2544 20198
rect 2504 19712 2556 19718
rect 2504 19654 2556 19660
rect 1860 19168 1912 19174
rect 1860 19110 1912 19116
rect 2412 19168 2464 19174
rect 2412 19110 2464 19116
rect 1768 18964 1820 18970
rect 1768 18906 1820 18912
rect 112 18284 164 18290
rect 112 18226 164 18232
rect 110 18184 166 18193
rect 110 18119 166 18128
rect 20 17876 72 17882
rect 20 17818 72 17824
rect 18 17776 74 17785
rect 18 17711 74 17720
rect 32 17474 60 17711
rect 20 17468 72 17474
rect 20 17410 72 17416
rect 18 17368 74 17377
rect 18 17303 74 17312
rect 32 17202 60 17303
rect 20 17196 72 17202
rect 20 17138 72 17144
rect 18 17096 74 17105
rect 18 17031 74 17040
rect 32 15978 60 17031
rect 124 16998 152 18119
rect 1768 18080 1820 18086
rect 1872 18068 1900 19110
rect 2228 18828 2280 18834
rect 2228 18770 2280 18776
rect 2240 18222 2268 18770
rect 2412 18760 2464 18766
rect 2516 18748 2544 19654
rect 2464 18720 2544 18748
rect 2412 18702 2464 18708
rect 2228 18216 2280 18222
rect 2228 18158 2280 18164
rect 1820 18040 1900 18068
rect 1768 18022 1820 18028
rect 1780 17134 1808 18022
rect 2240 17882 2268 18158
rect 2424 18086 2452 18702
rect 2412 18080 2464 18086
rect 2412 18022 2464 18028
rect 2228 17876 2280 17882
rect 2228 17818 2280 17824
rect 1952 17740 2004 17746
rect 1952 17682 2004 17688
rect 1964 17134 1992 17682
rect 2424 17678 2452 18022
rect 2412 17672 2464 17678
rect 2412 17614 2464 17620
rect 1768 17128 1820 17134
rect 1768 17070 1820 17076
rect 1952 17128 2004 17134
rect 1952 17070 2004 17076
rect 112 16992 164 16998
rect 112 16934 164 16940
rect 110 16688 166 16697
rect 166 16646 244 16674
rect 110 16623 166 16632
rect 110 16280 166 16289
rect 110 16215 166 16224
rect 20 15972 72 15978
rect 20 15914 72 15920
rect 18 15872 74 15881
rect 18 15807 74 15816
rect 32 14618 60 15807
rect 124 15162 152 16215
rect 216 15706 244 16646
rect 1780 16454 1808 17070
rect 1964 16726 1992 17070
rect 2424 16998 2452 17614
rect 2412 16992 2464 16998
rect 2412 16934 2464 16940
rect 1952 16720 2004 16726
rect 1952 16662 2004 16668
rect 1768 16448 1820 16454
rect 1768 16390 1820 16396
rect 1584 16040 1636 16046
rect 1584 15982 1636 15988
rect 204 15700 256 15706
rect 204 15642 256 15648
rect 1596 15366 1624 15982
rect 1780 15552 1808 16390
rect 2424 16114 2452 16934
rect 2412 16108 2464 16114
rect 2412 16050 2464 16056
rect 2136 16040 2188 16046
rect 2136 15982 2188 15988
rect 2148 15638 2176 15982
rect 2136 15632 2188 15638
rect 2136 15574 2188 15580
rect 1860 15564 1912 15570
rect 1780 15524 1860 15552
rect 1860 15506 1912 15512
rect 1584 15360 1636 15366
rect 1584 15302 1636 15308
rect 112 15156 164 15162
rect 112 15098 164 15104
rect 110 15056 166 15065
rect 166 15014 244 15042
rect 110 14991 166 15000
rect 20 14612 72 14618
rect 20 14554 72 14560
rect 110 14240 166 14249
rect 110 14175 166 14184
rect 124 13734 152 14175
rect 112 13728 164 13734
rect 112 13670 164 13676
rect 110 13560 166 13569
rect 110 13495 166 13504
rect 124 13462 152 13495
rect 112 13456 164 13462
rect 112 13398 164 13404
rect 18 13152 74 13161
rect 18 13087 74 13096
rect 32 12646 60 13087
rect 110 12744 166 12753
rect 110 12679 166 12688
rect 20 12640 72 12646
rect 20 12582 72 12588
rect 124 12442 152 12679
rect 112 12436 164 12442
rect 112 12378 164 12384
rect 216 12374 244 15014
rect 1596 13530 1624 15302
rect 1872 14822 1900 15506
rect 1860 14816 1912 14822
rect 1860 14758 1912 14764
rect 1676 14476 1728 14482
rect 1676 14418 1728 14424
rect 1688 13870 1716 14418
rect 1676 13864 1728 13870
rect 1676 13806 1728 13812
rect 1584 13524 1636 13530
rect 1584 13466 1636 13472
rect 204 12368 256 12374
rect 18 12336 74 12345
rect 204 12310 256 12316
rect 1688 12306 1716 13806
rect 1872 12986 1900 14758
rect 1952 14340 2004 14346
rect 1952 14282 2004 14288
rect 1964 13870 1992 14282
rect 2136 14000 2188 14006
rect 2136 13942 2188 13948
rect 1952 13864 2004 13870
rect 1952 13806 2004 13812
rect 1964 13530 1992 13806
rect 1952 13524 2004 13530
rect 1952 13466 2004 13472
rect 2148 13394 2176 13942
rect 2136 13388 2188 13394
rect 2136 13330 2188 13336
rect 2228 13388 2280 13394
rect 2228 13330 2280 13336
rect 1860 12980 1912 12986
rect 1860 12922 1912 12928
rect 18 12271 74 12280
rect 1676 12300 1728 12306
rect 32 11626 60 12271
rect 1676 12242 1728 12248
rect 2148 12170 2176 13330
rect 2240 12782 2268 13330
rect 2228 12776 2280 12782
rect 2228 12718 2280 12724
rect 2136 12164 2188 12170
rect 2136 12106 2188 12112
rect 1584 12096 1636 12102
rect 1584 12038 1636 12044
rect 1952 12096 2004 12102
rect 2240 12084 2268 12718
rect 2320 12096 2372 12102
rect 2240 12056 2320 12084
rect 1952 12038 2004 12044
rect 2320 12038 2372 12044
rect 110 11928 166 11937
rect 110 11863 166 11872
rect 20 11620 72 11626
rect 20 11562 72 11568
rect 124 11558 152 11863
rect 112 11552 164 11558
rect 18 11520 74 11529
rect 112 11494 164 11500
rect 18 11455 74 11464
rect 32 10538 60 11455
rect 112 11348 164 11354
rect 112 11290 164 11296
rect 124 11121 152 11290
rect 110 11112 166 11121
rect 110 11047 166 11056
rect 110 10704 166 10713
rect 166 10674 244 10690
rect 166 10668 256 10674
rect 166 10662 204 10668
rect 110 10639 166 10648
rect 204 10610 256 10616
rect 20 10532 72 10538
rect 20 10474 72 10480
rect 112 10532 164 10538
rect 112 10474 164 10480
rect 18 10432 74 10441
rect 18 10367 74 10376
rect 32 9674 60 10367
rect 124 10033 152 10474
rect 1400 10124 1452 10130
rect 1400 10066 1452 10072
rect 110 10024 166 10033
rect 110 9959 166 9968
rect 1412 9722 1440 10066
rect 1400 9716 1452 9722
rect 32 9646 152 9674
rect 1400 9658 1452 9664
rect 1596 9654 1624 12038
rect 1964 11762 1992 12038
rect 1952 11756 2004 11762
rect 1952 11698 2004 11704
rect 2332 11694 2360 12038
rect 1676 11688 1728 11694
rect 1676 11630 1728 11636
rect 2320 11688 2372 11694
rect 2320 11630 2372 11636
rect 1688 11218 1716 11630
rect 1676 11212 1728 11218
rect 1676 11154 1728 11160
rect 1688 10810 1716 11154
rect 1676 10804 1728 10810
rect 1676 10746 1728 10752
rect 1688 10606 1716 10746
rect 2608 10742 2636 23530
rect 5906 23520 5962 23582
rect 4160 21888 4212 21894
rect 4160 21830 4212 21836
rect 4172 21146 4200 21830
rect 4956 21788 5252 21808
rect 5012 21786 5036 21788
rect 5092 21786 5116 21788
rect 5172 21786 5196 21788
rect 5034 21734 5036 21786
rect 5098 21734 5110 21786
rect 5172 21734 5174 21786
rect 5012 21732 5036 21734
rect 5092 21732 5116 21734
rect 5172 21732 5196 21734
rect 4956 21712 5252 21732
rect 4710 21448 4766 21457
rect 4710 21383 4766 21392
rect 4160 21140 4212 21146
rect 4160 21082 4212 21088
rect 4068 21004 4120 21010
rect 4068 20946 4120 20952
rect 3516 20800 3568 20806
rect 3516 20742 3568 20748
rect 3528 20398 3556 20742
rect 3516 20392 3568 20398
rect 3516 20334 3568 20340
rect 4080 20262 4108 20946
rect 4528 20392 4580 20398
rect 4528 20334 4580 20340
rect 4068 20256 4120 20262
rect 4068 20198 4120 20204
rect 2688 19304 2740 19310
rect 2688 19246 2740 19252
rect 3608 19304 3660 19310
rect 3608 19246 3660 19252
rect 2700 18290 2728 19246
rect 3620 18970 3648 19246
rect 3608 18964 3660 18970
rect 3608 18906 3660 18912
rect 4080 18834 4108 20198
rect 4344 19984 4396 19990
rect 4344 19926 4396 19932
rect 4160 19848 4212 19854
rect 4160 19790 4212 19796
rect 4172 18970 4200 19790
rect 4356 19310 4384 19926
rect 4540 19922 4568 20334
rect 4724 20262 4752 21383
rect 5356 20800 5408 20806
rect 5356 20742 5408 20748
rect 4956 20700 5252 20720
rect 5012 20698 5036 20700
rect 5092 20698 5116 20700
rect 5172 20698 5196 20700
rect 5034 20646 5036 20698
rect 5098 20646 5110 20698
rect 5172 20646 5174 20698
rect 5012 20644 5036 20646
rect 5092 20644 5116 20646
rect 5172 20644 5196 20646
rect 4956 20624 5252 20644
rect 5368 20398 5396 20742
rect 5356 20392 5408 20398
rect 5356 20334 5408 20340
rect 4712 20256 4764 20262
rect 4618 20224 4674 20233
rect 4712 20198 4764 20204
rect 4618 20159 4674 20168
rect 4632 20058 4660 20159
rect 4620 20052 4672 20058
rect 4620 19994 4672 20000
rect 5368 19990 5396 20334
rect 5356 19984 5408 19990
rect 5356 19926 5408 19932
rect 4528 19916 4580 19922
rect 4528 19858 4580 19864
rect 4540 19514 4568 19858
rect 4956 19612 5252 19632
rect 5012 19610 5036 19612
rect 5092 19610 5116 19612
rect 5172 19610 5196 19612
rect 5034 19558 5036 19610
rect 5098 19558 5110 19610
rect 5172 19558 5174 19610
rect 5012 19556 5036 19558
rect 5092 19556 5116 19558
rect 5172 19556 5196 19558
rect 4956 19536 5252 19556
rect 4528 19508 4580 19514
rect 4528 19450 4580 19456
rect 4540 19310 4568 19450
rect 4344 19304 4396 19310
rect 4250 19272 4306 19281
rect 4344 19246 4396 19252
rect 4528 19304 4580 19310
rect 4528 19246 4580 19252
rect 4804 19304 4856 19310
rect 4804 19246 4856 19252
rect 4250 19207 4306 19216
rect 4264 18970 4292 19207
rect 4160 18964 4212 18970
rect 4160 18906 4212 18912
rect 4252 18964 4304 18970
rect 4252 18906 4304 18912
rect 4068 18828 4120 18834
rect 4068 18770 4120 18776
rect 4620 18828 4672 18834
rect 4620 18770 4672 18776
rect 3422 18728 3478 18737
rect 3422 18663 3478 18672
rect 2688 18284 2740 18290
rect 2688 18226 2740 18232
rect 2700 16590 2728 18226
rect 3436 18086 3464 18663
rect 4080 18290 4108 18770
rect 4068 18284 4120 18290
rect 4068 18226 4120 18232
rect 4632 18222 4660 18770
rect 3792 18216 3844 18222
rect 3792 18158 3844 18164
rect 4620 18216 4672 18222
rect 4620 18158 4672 18164
rect 3240 18080 3292 18086
rect 3240 18022 3292 18028
rect 3424 18080 3476 18086
rect 3424 18022 3476 18028
rect 3252 17066 3280 18022
rect 3804 17882 3832 18158
rect 4816 18154 4844 19246
rect 5908 19168 5960 19174
rect 5908 19110 5960 19116
rect 5632 18828 5684 18834
rect 5632 18770 5684 18776
rect 5448 18624 5500 18630
rect 5448 18566 5500 18572
rect 4956 18524 5252 18544
rect 5012 18522 5036 18524
rect 5092 18522 5116 18524
rect 5172 18522 5196 18524
rect 5034 18470 5036 18522
rect 5098 18470 5110 18522
rect 5172 18470 5174 18522
rect 5012 18468 5036 18470
rect 5092 18468 5116 18470
rect 5172 18468 5196 18470
rect 4956 18448 5252 18468
rect 5460 18426 5488 18566
rect 5448 18420 5500 18426
rect 5448 18362 5500 18368
rect 4804 18148 4856 18154
rect 4804 18090 4856 18096
rect 5172 18148 5224 18154
rect 5172 18090 5224 18096
rect 3792 17876 3844 17882
rect 3792 17818 3844 17824
rect 5184 17746 5212 18090
rect 4436 17740 4488 17746
rect 4436 17682 4488 17688
rect 5172 17740 5224 17746
rect 5172 17682 5224 17688
rect 4252 17536 4304 17542
rect 4252 17478 4304 17484
rect 3516 17128 3568 17134
rect 3516 17070 3568 17076
rect 3240 17060 3292 17066
rect 3240 17002 3292 17008
rect 3528 16726 3556 17070
rect 3700 17060 3752 17066
rect 3700 17002 3752 17008
rect 2872 16720 2924 16726
rect 2872 16662 2924 16668
rect 3516 16720 3568 16726
rect 3516 16662 3568 16668
rect 2688 16584 2740 16590
rect 2688 16526 2740 16532
rect 2700 15910 2728 16526
rect 2688 15904 2740 15910
rect 2688 15846 2740 15852
rect 2700 14890 2728 15846
rect 2884 15706 2912 16662
rect 3238 16008 3294 16017
rect 3238 15943 3294 15952
rect 3252 15910 3280 15943
rect 3240 15904 3292 15910
rect 3240 15846 3292 15852
rect 2872 15700 2924 15706
rect 2872 15642 2924 15648
rect 3332 15632 3384 15638
rect 3332 15574 3384 15580
rect 3344 15162 3372 15574
rect 3332 15156 3384 15162
rect 3332 15098 3384 15104
rect 3344 14958 3372 15098
rect 2780 14952 2832 14958
rect 2780 14894 2832 14900
rect 3332 14952 3384 14958
rect 3332 14894 3384 14900
rect 2688 14884 2740 14890
rect 2688 14826 2740 14832
rect 2792 14482 2820 14894
rect 3608 14884 3660 14890
rect 3608 14826 3660 14832
rect 2780 14476 2832 14482
rect 2780 14418 2832 14424
rect 2792 14074 2820 14418
rect 2780 14068 2832 14074
rect 2780 14010 2832 14016
rect 3054 13832 3110 13841
rect 2872 13796 2924 13802
rect 3054 13767 3110 13776
rect 2872 13738 2924 13744
rect 2884 13394 2912 13738
rect 3068 13734 3096 13767
rect 3056 13728 3108 13734
rect 3056 13670 3108 13676
rect 2872 13388 2924 13394
rect 2872 13330 2924 13336
rect 2780 13252 2832 13258
rect 2780 13194 2832 13200
rect 2792 12782 2820 13194
rect 2884 12782 2912 13330
rect 3424 13184 3476 13190
rect 3424 13126 3476 13132
rect 3240 12980 3292 12986
rect 3240 12922 3292 12928
rect 2780 12776 2832 12782
rect 2780 12718 2832 12724
rect 2872 12776 2924 12782
rect 2872 12718 2924 12724
rect 2688 12232 2740 12238
rect 2688 12174 2740 12180
rect 2700 11354 2728 12174
rect 2792 11778 2820 12718
rect 2884 12306 2912 12718
rect 2872 12300 2924 12306
rect 2872 12242 2924 12248
rect 2884 11898 2912 12242
rect 2872 11892 2924 11898
rect 2872 11834 2924 11840
rect 2792 11750 2912 11778
rect 2780 11688 2832 11694
rect 2780 11630 2832 11636
rect 2688 11348 2740 11354
rect 2688 11290 2740 11296
rect 2792 11218 2820 11630
rect 2780 11212 2832 11218
rect 2780 11154 2832 11160
rect 2792 10810 2820 11154
rect 2780 10804 2832 10810
rect 2780 10746 2832 10752
rect 2596 10736 2648 10742
rect 2596 10678 2648 10684
rect 2504 10668 2556 10674
rect 2504 10610 2556 10616
rect 1676 10600 1728 10606
rect 1676 10542 1728 10548
rect 2320 10600 2372 10606
rect 2320 10542 2372 10548
rect 1688 10266 1716 10542
rect 2332 10266 2360 10542
rect 2516 10266 2544 10610
rect 2884 10606 2912 11750
rect 3148 11008 3200 11014
rect 3148 10950 3200 10956
rect 2872 10600 2924 10606
rect 2872 10542 2924 10548
rect 1676 10260 1728 10266
rect 1676 10202 1728 10208
rect 2320 10260 2372 10266
rect 2320 10202 2372 10208
rect 2504 10260 2556 10266
rect 2504 10202 2556 10208
rect 124 9382 152 9646
rect 1584 9648 1636 9654
rect 1584 9590 1636 9596
rect 112 9376 164 9382
rect 112 9318 164 9324
rect 18 9208 74 9217
rect 18 9143 74 9152
rect 112 9172 164 9178
rect 32 8362 60 9143
rect 112 9114 164 9120
rect 124 8809 152 9114
rect 110 8800 166 8809
rect 110 8735 166 8744
rect 110 8392 166 8401
rect 20 8356 72 8362
rect 110 8327 166 8336
rect 20 8298 72 8304
rect 124 8294 152 8327
rect 112 8288 164 8294
rect 112 8230 164 8236
rect 112 8084 164 8090
rect 112 8026 164 8032
rect 124 7993 152 8026
rect 110 7984 166 7993
rect 1596 7954 1624 9590
rect 1860 9444 1912 9450
rect 1860 9386 1912 9392
rect 1872 9042 1900 9386
rect 1860 9036 1912 9042
rect 1860 8978 1912 8984
rect 2044 9036 2096 9042
rect 2044 8978 2096 8984
rect 1872 8090 1900 8978
rect 2056 8430 2084 8978
rect 2044 8424 2096 8430
rect 2044 8366 2096 8372
rect 1860 8084 1912 8090
rect 1860 8026 1912 8032
rect 110 7919 166 7928
rect 1584 7948 1636 7954
rect 1636 7908 1716 7936
rect 1584 7890 1636 7896
rect 18 7576 74 7585
rect 18 7511 74 7520
rect 32 6322 60 7511
rect 1582 7304 1638 7313
rect 1582 7239 1638 7248
rect 1596 7206 1624 7239
rect 1584 7200 1636 7206
rect 1584 7142 1636 7148
rect 112 6996 164 7002
rect 112 6938 164 6944
rect 124 6905 152 6938
rect 296 6928 348 6934
rect 110 6896 166 6905
rect 296 6870 348 6876
rect 110 6831 166 6840
rect 110 6488 166 6497
rect 110 6423 166 6432
rect 20 6316 72 6322
rect 20 6258 72 6264
rect 124 6118 152 6423
rect 112 6112 164 6118
rect 112 6054 164 6060
rect 112 5908 164 5914
rect 112 5850 164 5856
rect 18 5672 74 5681
rect 18 5607 74 5616
rect 32 5098 60 5607
rect 124 5273 152 5850
rect 204 5840 256 5846
rect 204 5782 256 5788
rect 110 5264 166 5273
rect 110 5199 166 5208
rect 20 5092 72 5098
rect 20 5034 72 5040
rect 112 5024 164 5030
rect 112 4966 164 4972
rect 124 4865 152 4966
rect 110 4856 166 4865
rect 20 4820 72 4826
rect 110 4791 166 4800
rect 20 4762 72 4768
rect 32 4049 60 4762
rect 110 4448 166 4457
rect 110 4383 166 4392
rect 124 4146 152 4383
rect 112 4140 164 4146
rect 112 4082 164 4088
rect 18 4040 74 4049
rect 18 3975 74 3984
rect 112 3936 164 3942
rect 112 3878 164 3884
rect 20 3732 72 3738
rect 20 3674 72 3680
rect 32 2145 60 3674
rect 124 3641 152 3878
rect 110 3632 166 3641
rect 110 3567 166 3576
rect 110 3360 166 3369
rect 110 3295 166 3304
rect 124 2854 152 3295
rect 112 2848 164 2854
rect 112 2790 164 2796
rect 112 2644 164 2650
rect 112 2586 164 2592
rect 18 2136 74 2145
rect 18 2071 74 2080
rect 124 1737 152 2586
rect 110 1728 166 1737
rect 110 1663 166 1672
rect 112 1352 164 1358
rect 18 1320 74 1329
rect 74 1300 112 1306
rect 74 1294 164 1300
rect 74 1278 152 1294
rect 18 1255 74 1264
rect 110 912 166 921
rect 216 898 244 5782
rect 166 870 244 898
rect 110 847 166 856
rect 110 232 166 241
rect 308 218 336 6870
rect 1688 6254 1716 7908
rect 1872 7342 1900 8026
rect 2056 7954 2084 8366
rect 2332 7954 2360 10202
rect 2688 9716 2740 9722
rect 2688 9658 2740 9664
rect 2700 9110 2728 9658
rect 3056 9580 3108 9586
rect 3056 9522 3108 9528
rect 3068 9178 3096 9522
rect 3160 9450 3188 10950
rect 3148 9444 3200 9450
rect 3148 9386 3200 9392
rect 3160 9178 3188 9386
rect 3056 9172 3108 9178
rect 3056 9114 3108 9120
rect 3148 9172 3200 9178
rect 3148 9114 3200 9120
rect 2688 9104 2740 9110
rect 2688 9046 2740 9052
rect 2872 8492 2924 8498
rect 2872 8434 2924 8440
rect 2044 7948 2096 7954
rect 2044 7890 2096 7896
rect 2320 7948 2372 7954
rect 2320 7890 2372 7896
rect 2056 7546 2084 7890
rect 2884 7818 2912 8434
rect 2872 7812 2924 7818
rect 2872 7754 2924 7760
rect 2044 7540 2096 7546
rect 2044 7482 2096 7488
rect 1860 7336 1912 7342
rect 1860 7278 1912 7284
rect 1952 7336 2004 7342
rect 1952 7278 2004 7284
rect 1872 7002 1900 7278
rect 1860 6996 1912 7002
rect 1860 6938 1912 6944
rect 1964 6866 1992 7278
rect 2884 6866 2912 7754
rect 3056 6996 3108 7002
rect 3056 6938 3108 6944
rect 1952 6860 2004 6866
rect 1952 6802 2004 6808
rect 2872 6860 2924 6866
rect 2872 6802 2924 6808
rect 1676 6248 1728 6254
rect 1676 6190 1728 6196
rect 1492 5772 1544 5778
rect 1492 5714 1544 5720
rect 1504 4078 1532 5714
rect 1688 5710 1716 6190
rect 2884 5914 2912 6802
rect 3068 5914 3096 6938
rect 1860 5908 1912 5914
rect 1860 5850 1912 5856
rect 2872 5908 2924 5914
rect 2872 5850 2924 5856
rect 3056 5908 3108 5914
rect 3056 5850 3108 5856
rect 1872 5778 1900 5850
rect 1860 5772 1912 5778
rect 1860 5714 1912 5720
rect 2044 5772 2096 5778
rect 2044 5714 2096 5720
rect 1676 5704 1728 5710
rect 1676 5646 1728 5652
rect 1688 5166 1716 5646
rect 2056 5166 2084 5714
rect 3068 5166 3096 5850
rect 3252 5778 3280 12922
rect 3436 12238 3464 13126
rect 3424 12232 3476 12238
rect 3424 12174 3476 12180
rect 3516 12164 3568 12170
rect 3516 12106 3568 12112
rect 3528 11694 3556 12106
rect 3516 11688 3568 11694
rect 3516 11630 3568 11636
rect 3528 11286 3556 11630
rect 3516 11280 3568 11286
rect 3516 11222 3568 11228
rect 3528 10266 3556 11222
rect 3620 10713 3648 14826
rect 3712 12374 3740 17002
rect 3976 16652 4028 16658
rect 3976 16594 4028 16600
rect 3988 15706 4016 16594
rect 4068 16040 4120 16046
rect 4068 15982 4120 15988
rect 3976 15700 4028 15706
rect 3976 15642 4028 15648
rect 3792 15564 3844 15570
rect 3792 15506 3844 15512
rect 3804 15162 3832 15506
rect 3988 15434 4016 15642
rect 3976 15428 4028 15434
rect 3976 15370 4028 15376
rect 4080 15162 4108 15982
rect 4264 15638 4292 17478
rect 4344 16992 4396 16998
rect 4344 16934 4396 16940
rect 4356 16114 4384 16934
rect 4448 16590 4476 17682
rect 5460 17542 5488 18362
rect 5540 18284 5592 18290
rect 5540 18226 5592 18232
rect 4528 17536 4580 17542
rect 4528 17478 4580 17484
rect 5448 17536 5500 17542
rect 5448 17478 5500 17484
rect 4540 16658 4568 17478
rect 4956 17436 5252 17456
rect 5012 17434 5036 17436
rect 5092 17434 5116 17436
rect 5172 17434 5196 17436
rect 5034 17382 5036 17434
rect 5098 17382 5110 17434
rect 5172 17382 5174 17434
rect 5012 17380 5036 17382
rect 5092 17380 5116 17382
rect 5172 17380 5196 17382
rect 4956 17360 5252 17380
rect 5356 17196 5408 17202
rect 5356 17138 5408 17144
rect 5172 17060 5224 17066
rect 5172 17002 5224 17008
rect 5184 16658 5212 17002
rect 5368 16998 5396 17138
rect 5356 16992 5408 16998
rect 5356 16934 5408 16940
rect 4528 16652 4580 16658
rect 4528 16594 4580 16600
rect 5172 16652 5224 16658
rect 5172 16594 5224 16600
rect 4436 16584 4488 16590
rect 4436 16526 4488 16532
rect 4448 16250 4476 16526
rect 4436 16244 4488 16250
rect 4436 16186 4488 16192
rect 4344 16108 4396 16114
rect 4344 16050 4396 16056
rect 4540 15978 4568 16594
rect 5368 16436 5396 16934
rect 5552 16590 5580 18226
rect 5644 17814 5672 18770
rect 5632 17808 5684 17814
rect 5632 17750 5684 17756
rect 5632 17672 5684 17678
rect 5632 17614 5684 17620
rect 5724 17672 5776 17678
rect 5724 17614 5776 17620
rect 5644 17202 5672 17614
rect 5736 17338 5764 17614
rect 5724 17332 5776 17338
rect 5724 17274 5776 17280
rect 5632 17196 5684 17202
rect 5632 17138 5684 17144
rect 5632 16720 5684 16726
rect 5632 16662 5684 16668
rect 5540 16584 5592 16590
rect 5540 16526 5592 16532
rect 5448 16448 5500 16454
rect 5368 16408 5448 16436
rect 4956 16348 5252 16368
rect 5012 16346 5036 16348
rect 5092 16346 5116 16348
rect 5172 16346 5196 16348
rect 5034 16294 5036 16346
rect 5098 16294 5110 16346
rect 5172 16294 5174 16346
rect 5012 16292 5036 16294
rect 5092 16292 5116 16294
rect 5172 16292 5196 16294
rect 4956 16272 5252 16292
rect 5368 16182 5396 16408
rect 5448 16390 5500 16396
rect 5552 16250 5580 16526
rect 5540 16244 5592 16250
rect 5540 16186 5592 16192
rect 5356 16176 5408 16182
rect 5356 16118 5408 16124
rect 4859 16040 4911 16046
rect 4724 16000 4859 16028
rect 4528 15972 4580 15978
rect 4528 15914 4580 15920
rect 4252 15632 4304 15638
rect 4252 15574 4304 15580
rect 4540 15570 4568 15914
rect 4724 15706 4752 16000
rect 4859 15982 4911 15988
rect 4712 15700 4764 15706
rect 4712 15642 4764 15648
rect 4528 15564 4580 15570
rect 4528 15506 4580 15512
rect 4724 15366 4752 15642
rect 4804 15496 4856 15502
rect 4804 15438 4856 15444
rect 4712 15360 4764 15366
rect 4712 15302 4764 15308
rect 3792 15156 3844 15162
rect 3792 15098 3844 15104
rect 4068 15156 4120 15162
rect 4068 15098 4120 15104
rect 4080 14822 4108 15098
rect 4252 14952 4304 14958
rect 4342 14920 4398 14929
rect 4304 14900 4342 14906
rect 4252 14894 4342 14900
rect 4264 14878 4342 14894
rect 4068 14816 4120 14822
rect 4068 14758 4120 14764
rect 4264 14618 4292 14878
rect 4342 14855 4398 14864
rect 4436 14816 4488 14822
rect 4436 14758 4488 14764
rect 4528 14816 4580 14822
rect 4528 14758 4580 14764
rect 4252 14612 4304 14618
rect 4252 14554 4304 14560
rect 3884 14476 3936 14482
rect 3884 14418 3936 14424
rect 3896 13530 3924 14418
rect 4448 14346 4476 14758
rect 4540 14482 4568 14758
rect 4724 14482 4752 15302
rect 4816 15162 4844 15438
rect 5368 15366 5396 16118
rect 5448 16040 5500 16046
rect 5448 15982 5500 15988
rect 5460 15366 5488 15982
rect 5552 15502 5580 16186
rect 5644 16182 5672 16662
rect 5736 16522 5764 17274
rect 5920 16726 5948 19110
rect 5908 16720 5960 16726
rect 5908 16662 5960 16668
rect 5724 16516 5776 16522
rect 5724 16458 5776 16464
rect 5632 16176 5684 16182
rect 5632 16118 5684 16124
rect 5644 15706 5672 16118
rect 5736 15706 5764 16458
rect 5632 15700 5684 15706
rect 5632 15642 5684 15648
rect 5724 15700 5776 15706
rect 5724 15642 5776 15648
rect 5540 15496 5592 15502
rect 5540 15438 5592 15444
rect 5356 15360 5408 15366
rect 5356 15302 5408 15308
rect 5448 15360 5500 15366
rect 5448 15302 5500 15308
rect 4956 15260 5252 15280
rect 5012 15258 5036 15260
rect 5092 15258 5116 15260
rect 5172 15258 5196 15260
rect 5034 15206 5036 15258
rect 5098 15206 5110 15258
rect 5172 15206 5174 15258
rect 5012 15204 5036 15206
rect 5092 15204 5116 15206
rect 5172 15204 5196 15206
rect 4956 15184 5252 15204
rect 4804 15156 4856 15162
rect 4804 15098 4856 15104
rect 5264 15020 5316 15026
rect 5264 14962 5316 14968
rect 4804 14544 4856 14550
rect 4804 14486 4856 14492
rect 4528 14476 4580 14482
rect 4528 14418 4580 14424
rect 4712 14476 4764 14482
rect 4712 14418 4764 14424
rect 4436 14340 4488 14346
rect 4436 14282 4488 14288
rect 4252 14272 4304 14278
rect 4252 14214 4304 14220
rect 4344 14272 4396 14278
rect 4344 14214 4396 14220
rect 4264 13938 4292 14214
rect 4252 13932 4304 13938
rect 4252 13874 4304 13880
rect 4356 13530 4384 14214
rect 4448 13705 4476 14282
rect 4712 14272 4764 14278
rect 4712 14214 4764 14220
rect 4434 13696 4490 13705
rect 4490 13654 4568 13682
rect 4434 13631 4490 13640
rect 3884 13524 3936 13530
rect 3884 13466 3936 13472
rect 4344 13524 4396 13530
rect 4344 13466 4396 13472
rect 4436 13524 4488 13530
rect 4436 13466 4488 13472
rect 4252 12776 4304 12782
rect 4252 12718 4304 12724
rect 3700 12368 3752 12374
rect 3700 12310 3752 12316
rect 4264 12306 4292 12718
rect 4252 12300 4304 12306
rect 4252 12242 4304 12248
rect 4264 11218 4292 12242
rect 4252 11212 4304 11218
rect 4252 11154 4304 11160
rect 4160 11076 4212 11082
rect 4160 11018 4212 11024
rect 4172 10810 4200 11018
rect 4264 11014 4292 11154
rect 4252 11008 4304 11014
rect 4252 10950 4304 10956
rect 4160 10804 4212 10810
rect 4160 10746 4212 10752
rect 3606 10704 3662 10713
rect 3662 10662 3740 10690
rect 3606 10639 3662 10648
rect 3516 10260 3568 10266
rect 3516 10202 3568 10208
rect 3330 9480 3386 9489
rect 3330 9415 3386 9424
rect 3344 9382 3372 9415
rect 3332 9376 3384 9382
rect 3332 9318 3384 9324
rect 3528 9042 3556 10202
rect 3516 9036 3568 9042
rect 3516 8978 3568 8984
rect 3608 8424 3660 8430
rect 3608 8366 3660 8372
rect 3516 8356 3568 8362
rect 3516 8298 3568 8304
rect 3528 8090 3556 8298
rect 3620 8294 3648 8366
rect 3608 8288 3660 8294
rect 3608 8230 3660 8236
rect 3516 8084 3568 8090
rect 3516 8026 3568 8032
rect 3712 7342 3740 10662
rect 3884 10668 3936 10674
rect 3884 10610 3936 10616
rect 3792 10600 3844 10606
rect 3792 10542 3844 10548
rect 3804 10062 3832 10542
rect 3792 10056 3844 10062
rect 3792 9998 3844 10004
rect 3804 9518 3832 9998
rect 3792 9512 3844 9518
rect 3792 9454 3844 9460
rect 3896 7818 3924 10610
rect 4264 10266 4292 10950
rect 4252 10260 4304 10266
rect 4252 10202 4304 10208
rect 4160 10192 4212 10198
rect 4160 10134 4212 10140
rect 4172 9674 4200 10134
rect 4252 9920 4304 9926
rect 4252 9862 4304 9868
rect 4080 9654 4200 9674
rect 4068 9648 4200 9654
rect 4120 9646 4200 9648
rect 4068 9590 4120 9596
rect 4264 8974 4292 9862
rect 4252 8968 4304 8974
rect 4252 8910 4304 8916
rect 3976 8288 4028 8294
rect 3976 8230 4028 8236
rect 3884 7812 3936 7818
rect 3884 7754 3936 7760
rect 3700 7336 3752 7342
rect 3700 7278 3752 7284
rect 3884 7336 3936 7342
rect 3884 7278 3936 7284
rect 3424 7200 3476 7206
rect 3424 7142 3476 7148
rect 3608 7200 3660 7206
rect 3608 7142 3660 7148
rect 3240 5772 3292 5778
rect 3240 5714 3292 5720
rect 1676 5160 1728 5166
rect 2044 5160 2096 5166
rect 1728 5120 1808 5148
rect 1676 5102 1728 5108
rect 1492 4072 1544 4078
rect 1492 4014 1544 4020
rect 1504 3602 1532 4014
rect 1492 3596 1544 3602
rect 1492 3538 1544 3544
rect 388 3528 440 3534
rect 388 3470 440 3476
rect 400 2961 428 3470
rect 1780 2990 1808 5120
rect 2044 5102 2096 5108
rect 2872 5160 2924 5166
rect 2872 5102 2924 5108
rect 3056 5160 3108 5166
rect 3056 5102 3108 5108
rect 2884 4826 2912 5102
rect 2872 4820 2924 4826
rect 2872 4762 2924 4768
rect 3068 4690 3096 5102
rect 2136 4684 2188 4690
rect 2136 4626 2188 4632
rect 2780 4684 2832 4690
rect 2780 4626 2832 4632
rect 3056 4684 3108 4690
rect 3056 4626 3108 4632
rect 2148 4078 2176 4626
rect 2136 4072 2188 4078
rect 2136 4014 2188 4020
rect 2148 2990 2176 4014
rect 2228 3596 2280 3602
rect 2228 3538 2280 3544
rect 1768 2984 1820 2990
rect 386 2952 442 2961
rect 1768 2926 1820 2932
rect 2136 2984 2188 2990
rect 2136 2926 2188 2932
rect 386 2887 442 2896
rect 386 2544 442 2553
rect 1780 2514 1808 2926
rect 2240 2854 2268 3538
rect 2228 2848 2280 2854
rect 2228 2790 2280 2796
rect 2240 2514 2268 2790
rect 2792 2582 2820 4626
rect 2780 2576 2832 2582
rect 2780 2518 2832 2524
rect 386 2479 442 2488
rect 1768 2508 1820 2514
rect 400 2378 428 2479
rect 1768 2450 1820 2456
rect 2228 2508 2280 2514
rect 2228 2450 2280 2456
rect 388 2372 440 2378
rect 388 2314 440 2320
rect 3436 649 3464 7142
rect 3620 6254 3648 7142
rect 3712 7002 3740 7278
rect 3700 6996 3752 7002
rect 3700 6938 3752 6944
rect 3896 6662 3924 7278
rect 3884 6656 3936 6662
rect 3884 6598 3936 6604
rect 3988 6254 4016 8230
rect 4344 7948 4396 7954
rect 4344 7890 4396 7896
rect 4356 7546 4384 7890
rect 4344 7540 4396 7546
rect 4344 7482 4396 7488
rect 3608 6248 3660 6254
rect 3608 6190 3660 6196
rect 3976 6248 4028 6254
rect 3976 6190 4028 6196
rect 3988 5914 4016 6190
rect 3976 5908 4028 5914
rect 4448 5896 4476 13466
rect 4540 12306 4568 13654
rect 4620 13388 4672 13394
rect 4620 13330 4672 13336
rect 4632 12714 4660 13330
rect 4724 12850 4752 14214
rect 4816 14074 4844 14486
rect 5276 14346 5304 14962
rect 5264 14340 5316 14346
rect 5264 14282 5316 14288
rect 4956 14172 5252 14192
rect 5012 14170 5036 14172
rect 5092 14170 5116 14172
rect 5172 14170 5196 14172
rect 5034 14118 5036 14170
rect 5098 14118 5110 14170
rect 5172 14118 5174 14170
rect 5012 14116 5036 14118
rect 5092 14116 5116 14118
rect 5172 14116 5196 14118
rect 4956 14096 5252 14116
rect 4804 14068 4856 14074
rect 4804 14010 4856 14016
rect 5264 13864 5316 13870
rect 5264 13806 5316 13812
rect 4804 13796 4856 13802
rect 4804 13738 4856 13744
rect 4816 12986 4844 13738
rect 5276 13394 5304 13806
rect 5264 13388 5316 13394
rect 5264 13330 5316 13336
rect 5368 13190 5396 15302
rect 5460 14958 5488 15302
rect 5448 14952 5500 14958
rect 5448 14894 5500 14900
rect 5460 14414 5488 14894
rect 5552 14550 5580 15438
rect 5540 14544 5592 14550
rect 5540 14486 5592 14492
rect 5448 14408 5500 14414
rect 5448 14350 5500 14356
rect 5460 13326 5488 14350
rect 5552 13938 5580 14486
rect 5644 14074 5672 15642
rect 5724 14272 5776 14278
rect 5724 14214 5776 14220
rect 5632 14068 5684 14074
rect 5632 14010 5684 14016
rect 5540 13932 5592 13938
rect 5540 13874 5592 13880
rect 5552 13530 5580 13874
rect 5540 13524 5592 13530
rect 5540 13466 5592 13472
rect 5644 13462 5672 14010
rect 5632 13456 5684 13462
rect 5632 13398 5684 13404
rect 5448 13320 5500 13326
rect 5448 13262 5500 13268
rect 5356 13184 5408 13190
rect 5356 13126 5408 13132
rect 4956 13084 5252 13104
rect 5012 13082 5036 13084
rect 5092 13082 5116 13084
rect 5172 13082 5196 13084
rect 5034 13030 5036 13082
rect 5098 13030 5110 13082
rect 5172 13030 5174 13082
rect 5012 13028 5036 13030
rect 5092 13028 5116 13030
rect 5172 13028 5196 13030
rect 4956 13008 5252 13028
rect 4804 12980 4856 12986
rect 4804 12922 4856 12928
rect 4712 12844 4764 12850
rect 4712 12786 4764 12792
rect 5368 12782 5396 13126
rect 5356 12776 5408 12782
rect 5356 12718 5408 12724
rect 4620 12708 4672 12714
rect 4620 12650 4672 12656
rect 4528 12300 4580 12306
rect 4528 12242 4580 12248
rect 4540 11898 4568 12242
rect 4632 12170 4660 12650
rect 4804 12368 4856 12374
rect 4804 12310 4856 12316
rect 4620 12164 4672 12170
rect 4620 12106 4672 12112
rect 4632 11898 4660 12106
rect 4528 11892 4580 11898
rect 4528 11834 4580 11840
rect 4620 11892 4672 11898
rect 4620 11834 4672 11840
rect 4816 11626 4844 12310
rect 5368 12102 5396 12718
rect 5460 12442 5488 13262
rect 5644 12986 5672 13398
rect 5632 12980 5684 12986
rect 5632 12922 5684 12928
rect 5644 12714 5672 12922
rect 5632 12708 5684 12714
rect 5632 12650 5684 12656
rect 5540 12640 5592 12646
rect 5540 12582 5592 12588
rect 5448 12436 5500 12442
rect 5448 12378 5500 12384
rect 5356 12096 5408 12102
rect 5356 12038 5408 12044
rect 4956 11996 5252 12016
rect 5012 11994 5036 11996
rect 5092 11994 5116 11996
rect 5172 11994 5196 11996
rect 5034 11942 5036 11994
rect 5098 11942 5110 11994
rect 5172 11942 5174 11994
rect 5012 11940 5036 11942
rect 5092 11940 5116 11942
rect 5172 11940 5196 11942
rect 4956 11920 5252 11940
rect 5368 11898 5396 12038
rect 5356 11892 5408 11898
rect 5356 11834 5408 11840
rect 4804 11620 4856 11626
rect 4804 11562 4856 11568
rect 4528 11552 4580 11558
rect 4528 11494 4580 11500
rect 4540 11354 4568 11494
rect 4528 11348 4580 11354
rect 4528 11290 4580 11296
rect 4620 11212 4672 11218
rect 4620 11154 4672 11160
rect 4528 10668 4580 10674
rect 4528 10610 4580 10616
rect 4540 10266 4568 10610
rect 4632 10470 4660 11154
rect 4620 10464 4672 10470
rect 4620 10406 4672 10412
rect 4528 10260 4580 10266
rect 4528 10202 4580 10208
rect 4632 10062 4660 10406
rect 4712 10124 4764 10130
rect 4712 10066 4764 10072
rect 4620 10056 4672 10062
rect 4620 9998 4672 10004
rect 4528 9988 4580 9994
rect 4528 9930 4580 9936
rect 4540 6866 4568 9930
rect 4724 9722 4752 10066
rect 4816 9994 4844 11562
rect 4956 10908 5252 10928
rect 5012 10906 5036 10908
rect 5092 10906 5116 10908
rect 5172 10906 5196 10908
rect 5034 10854 5036 10906
rect 5098 10854 5110 10906
rect 5172 10854 5174 10906
rect 5012 10852 5036 10854
rect 5092 10852 5116 10854
rect 5172 10852 5196 10854
rect 4956 10832 5252 10852
rect 4988 10532 5040 10538
rect 4988 10474 5040 10480
rect 5000 10266 5028 10474
rect 5356 10464 5408 10470
rect 5356 10406 5408 10412
rect 4988 10260 5040 10266
rect 4988 10202 5040 10208
rect 5368 9994 5396 10406
rect 4804 9988 4856 9994
rect 4804 9930 4856 9936
rect 5356 9988 5408 9994
rect 5356 9930 5408 9936
rect 4956 9820 5252 9840
rect 5012 9818 5036 9820
rect 5092 9818 5116 9820
rect 5172 9818 5196 9820
rect 5034 9766 5036 9818
rect 5098 9766 5110 9818
rect 5172 9766 5174 9818
rect 5012 9764 5036 9766
rect 5092 9764 5116 9766
rect 5172 9764 5196 9766
rect 4956 9744 5252 9764
rect 5368 9722 5396 9930
rect 4712 9716 4764 9722
rect 5356 9716 5408 9722
rect 4764 9676 4844 9704
rect 4712 9658 4764 9664
rect 4712 9172 4764 9178
rect 4712 9114 4764 9120
rect 4620 9036 4672 9042
rect 4620 8978 4672 8984
rect 4632 7954 4660 8978
rect 4724 7954 4752 9114
rect 4816 8974 4844 9676
rect 5356 9658 5408 9664
rect 5172 9648 5224 9654
rect 5172 9590 5224 9596
rect 5184 9518 5212 9590
rect 5080 9512 5132 9518
rect 5080 9454 5132 9460
rect 5172 9512 5224 9518
rect 5172 9454 5224 9460
rect 4988 9376 5040 9382
rect 4988 9318 5040 9324
rect 5000 9042 5028 9318
rect 5092 9110 5120 9454
rect 5080 9104 5132 9110
rect 5080 9046 5132 9052
rect 4988 9036 5040 9042
rect 4988 8978 5040 8984
rect 4804 8968 4856 8974
rect 4804 8910 4856 8916
rect 4816 8634 4844 8910
rect 5184 8906 5212 9454
rect 5356 9104 5408 9110
rect 5356 9046 5408 9052
rect 5172 8900 5224 8906
rect 5172 8842 5224 8848
rect 4956 8732 5252 8752
rect 5012 8730 5036 8732
rect 5092 8730 5116 8732
rect 5172 8730 5196 8732
rect 5034 8678 5036 8730
rect 5098 8678 5110 8730
rect 5172 8678 5174 8730
rect 5012 8676 5036 8678
rect 5092 8676 5116 8678
rect 5172 8676 5196 8678
rect 4956 8656 5252 8676
rect 5368 8634 5396 9046
rect 5552 9024 5580 12582
rect 5736 11914 5764 14214
rect 5908 13728 5960 13734
rect 5908 13670 5960 13676
rect 5460 8996 5580 9024
rect 5644 11886 5764 11914
rect 4804 8628 4856 8634
rect 4804 8570 4856 8576
rect 5356 8628 5408 8634
rect 5356 8570 5408 8576
rect 4816 8498 4844 8570
rect 4804 8492 4856 8498
rect 4804 8434 4856 8440
rect 5264 8288 5316 8294
rect 5264 8230 5316 8236
rect 5276 8090 5304 8230
rect 5264 8084 5316 8090
rect 5264 8026 5316 8032
rect 4620 7948 4672 7954
rect 4620 7890 4672 7896
rect 4712 7948 4764 7954
rect 4712 7890 4764 7896
rect 4724 7546 4752 7890
rect 4956 7644 5252 7664
rect 5012 7642 5036 7644
rect 5092 7642 5116 7644
rect 5172 7642 5196 7644
rect 5034 7590 5036 7642
rect 5098 7590 5110 7642
rect 5172 7590 5174 7642
rect 5012 7588 5036 7590
rect 5092 7588 5116 7590
rect 5172 7588 5196 7590
rect 4956 7568 5252 7588
rect 4712 7540 4764 7546
rect 4712 7482 4764 7488
rect 4528 6860 4580 6866
rect 4528 6802 4580 6808
rect 4540 6458 4568 6802
rect 4712 6656 4764 6662
rect 4712 6598 4764 6604
rect 4528 6452 4580 6458
rect 4528 6394 4580 6400
rect 4724 6118 4752 6598
rect 4956 6556 5252 6576
rect 5012 6554 5036 6556
rect 5092 6554 5116 6556
rect 5172 6554 5196 6556
rect 5034 6502 5036 6554
rect 5098 6502 5110 6554
rect 5172 6502 5174 6554
rect 5012 6500 5036 6502
rect 5092 6500 5116 6502
rect 5172 6500 5196 6502
rect 4956 6480 5252 6500
rect 4712 6112 4764 6118
rect 4712 6054 4764 6060
rect 3976 5850 4028 5856
rect 4356 5868 4476 5896
rect 3516 5704 3568 5710
rect 3516 5646 3568 5652
rect 3528 4826 3556 5646
rect 3988 4826 4016 5850
rect 4068 5636 4120 5642
rect 4068 5578 4120 5584
rect 4080 5030 4108 5578
rect 4356 5250 4384 5868
rect 4724 5778 4752 6054
rect 4436 5772 4488 5778
rect 4436 5714 4488 5720
rect 4712 5772 4764 5778
rect 4712 5714 4764 5720
rect 4448 5370 4476 5714
rect 4956 5468 5252 5488
rect 5012 5466 5036 5468
rect 5092 5466 5116 5468
rect 5172 5466 5196 5468
rect 5034 5414 5036 5466
rect 5098 5414 5110 5466
rect 5172 5414 5174 5466
rect 5012 5412 5036 5414
rect 5092 5412 5116 5414
rect 5172 5412 5196 5414
rect 4956 5392 5252 5412
rect 5460 5370 5488 8996
rect 5540 8900 5592 8906
rect 5540 8842 5592 8848
rect 5552 8022 5580 8842
rect 5540 8016 5592 8022
rect 5540 7958 5592 7964
rect 5644 6866 5672 11886
rect 5724 11688 5776 11694
rect 5724 11630 5776 11636
rect 5736 11286 5764 11630
rect 5724 11280 5776 11286
rect 5724 11222 5776 11228
rect 5736 10266 5764 11222
rect 5724 10260 5776 10266
rect 5724 10202 5776 10208
rect 5724 10124 5776 10130
rect 5724 10066 5776 10072
rect 5736 9518 5764 10066
rect 5724 9512 5776 9518
rect 5724 9454 5776 9460
rect 5736 9042 5764 9454
rect 5724 9036 5776 9042
rect 5724 8978 5776 8984
rect 5736 8566 5764 8978
rect 5724 8560 5776 8566
rect 5724 8502 5776 8508
rect 5632 6860 5684 6866
rect 5632 6802 5684 6808
rect 5644 6458 5672 6802
rect 5632 6452 5684 6458
rect 5632 6394 5684 6400
rect 4436 5364 4488 5370
rect 4436 5306 4488 5312
rect 5448 5364 5500 5370
rect 5448 5306 5500 5312
rect 4528 5296 4580 5302
rect 4356 5222 4476 5250
rect 4528 5238 4580 5244
rect 4068 5024 4120 5030
rect 4068 4966 4120 4972
rect 4158 4992 4214 5001
rect 3516 4820 3568 4826
rect 3976 4820 4028 4826
rect 3516 4762 3568 4768
rect 3896 4780 3976 4808
rect 3528 3738 3556 4762
rect 3896 4078 3924 4780
rect 3976 4762 4028 4768
rect 3884 4072 3936 4078
rect 3884 4014 3936 4020
rect 3896 3738 3924 4014
rect 3516 3732 3568 3738
rect 3516 3674 3568 3680
rect 3884 3732 3936 3738
rect 3884 3674 3936 3680
rect 3528 2650 3556 3674
rect 3896 2990 3924 3674
rect 4080 3058 4108 4966
rect 4158 4927 4214 4936
rect 4172 4826 4200 4927
rect 4160 4820 4212 4826
rect 4160 4762 4212 4768
rect 4344 4684 4396 4690
rect 4344 4626 4396 4632
rect 4356 4146 4384 4626
rect 4344 4140 4396 4146
rect 4344 4082 4396 4088
rect 4356 3194 4384 4082
rect 4448 4078 4476 5222
rect 4540 4690 4568 5238
rect 4528 4684 4580 4690
rect 4528 4626 4580 4632
rect 4540 4214 4568 4626
rect 4956 4380 5252 4400
rect 5012 4378 5036 4380
rect 5092 4378 5116 4380
rect 5172 4378 5196 4380
rect 5034 4326 5036 4378
rect 5098 4326 5110 4378
rect 5172 4326 5174 4378
rect 5012 4324 5036 4326
rect 5092 4324 5116 4326
rect 5172 4324 5196 4326
rect 4956 4304 5252 4324
rect 4528 4208 4580 4214
rect 4528 4150 4580 4156
rect 4436 4072 4488 4078
rect 4436 4014 4488 4020
rect 4620 3596 4672 3602
rect 4620 3538 4672 3544
rect 4344 3188 4396 3194
rect 4344 3130 4396 3136
rect 4632 3126 4660 3538
rect 4956 3292 5252 3312
rect 5012 3290 5036 3292
rect 5092 3290 5116 3292
rect 5172 3290 5196 3292
rect 5034 3238 5036 3290
rect 5098 3238 5110 3290
rect 5172 3238 5174 3290
rect 5012 3236 5036 3238
rect 5092 3236 5116 3238
rect 5172 3236 5196 3238
rect 4956 3216 5252 3236
rect 5920 3194 5948 13670
rect 6012 10198 6040 23582
rect 9600 23582 10010 23610
rect 8956 21244 9252 21264
rect 9012 21242 9036 21244
rect 9092 21242 9116 21244
rect 9172 21242 9196 21244
rect 9034 21190 9036 21242
rect 9098 21190 9110 21242
rect 9172 21190 9174 21242
rect 9012 21188 9036 21190
rect 9092 21188 9116 21190
rect 9172 21188 9196 21190
rect 8956 21168 9252 21188
rect 7012 20392 7064 20398
rect 7012 20334 7064 20340
rect 6276 19916 6328 19922
rect 6276 19858 6328 19864
rect 6288 19174 6316 19858
rect 7024 19514 7052 20334
rect 8956 20156 9252 20176
rect 9012 20154 9036 20156
rect 9092 20154 9116 20156
rect 9172 20154 9196 20156
rect 9034 20102 9036 20154
rect 9098 20102 9110 20154
rect 9172 20102 9174 20154
rect 9012 20100 9036 20102
rect 9092 20100 9116 20102
rect 9172 20100 9196 20102
rect 8956 20080 9252 20100
rect 7012 19508 7064 19514
rect 7012 19450 7064 19456
rect 6828 19304 6880 19310
rect 6828 19246 6880 19252
rect 6276 19168 6328 19174
rect 6276 19110 6328 19116
rect 6184 18624 6236 18630
rect 6184 18566 6236 18572
rect 6196 18222 6224 18566
rect 6288 18426 6316 19110
rect 6276 18420 6328 18426
rect 6276 18362 6328 18368
rect 6184 18216 6236 18222
rect 6184 18158 6236 18164
rect 6196 17882 6224 18158
rect 6552 18080 6604 18086
rect 6552 18022 6604 18028
rect 6184 17876 6236 17882
rect 6184 17818 6236 17824
rect 6196 17610 6224 17818
rect 6564 17814 6592 18022
rect 6552 17808 6604 17814
rect 6552 17750 6604 17756
rect 6644 17740 6696 17746
rect 6644 17682 6696 17688
rect 6184 17604 6236 17610
rect 6184 17546 6236 17552
rect 6092 17536 6144 17542
rect 6092 17478 6144 17484
rect 6104 17270 6132 17478
rect 6092 17264 6144 17270
rect 6092 17206 6144 17212
rect 6104 15094 6132 17206
rect 6656 16998 6684 17682
rect 6840 17338 6868 19246
rect 8956 19068 9252 19088
rect 9012 19066 9036 19068
rect 9092 19066 9116 19068
rect 9172 19066 9196 19068
rect 9034 19014 9036 19066
rect 9098 19014 9110 19066
rect 9172 19014 9174 19066
rect 9012 19012 9036 19014
rect 9092 19012 9116 19014
rect 9172 19012 9196 19014
rect 8956 18992 9252 19012
rect 6920 18216 6972 18222
rect 6920 18158 6972 18164
rect 6932 17882 6960 18158
rect 7012 18080 7064 18086
rect 7012 18022 7064 18028
rect 6920 17876 6972 17882
rect 6920 17818 6972 17824
rect 7024 17678 7052 18022
rect 8956 17980 9252 18000
rect 9012 17978 9036 17980
rect 9092 17978 9116 17980
rect 9172 17978 9196 17980
rect 9034 17926 9036 17978
rect 9098 17926 9110 17978
rect 9172 17926 9174 17978
rect 9012 17924 9036 17926
rect 9092 17924 9116 17926
rect 9172 17924 9196 17926
rect 8956 17904 9252 17924
rect 7012 17672 7064 17678
rect 7012 17614 7064 17620
rect 6828 17332 6880 17338
rect 6828 17274 6880 17280
rect 6920 17196 6972 17202
rect 6920 17138 6972 17144
rect 6644 16992 6696 16998
rect 6644 16934 6696 16940
rect 6368 16652 6420 16658
rect 6368 16594 6420 16600
rect 6380 16250 6408 16594
rect 6368 16244 6420 16250
rect 6368 16186 6420 16192
rect 6380 15910 6408 16186
rect 6656 16114 6684 16934
rect 6932 16794 6960 17138
rect 7380 17128 7432 17134
rect 7378 17096 7380 17105
rect 7432 17096 7434 17105
rect 7378 17031 7434 17040
rect 7392 16998 7420 17031
rect 7380 16992 7432 16998
rect 7380 16934 7432 16940
rect 6920 16788 6972 16794
rect 6920 16730 6972 16736
rect 6736 16652 6788 16658
rect 6736 16594 6788 16600
rect 6644 16108 6696 16114
rect 6644 16050 6696 16056
rect 6368 15904 6420 15910
rect 6368 15846 6420 15852
rect 6460 15700 6512 15706
rect 6460 15642 6512 15648
rect 6276 15564 6328 15570
rect 6276 15506 6328 15512
rect 6288 15094 6316 15506
rect 6092 15088 6144 15094
rect 6092 15030 6144 15036
rect 6276 15088 6328 15094
rect 6276 15030 6328 15036
rect 6104 14482 6132 15030
rect 6288 14618 6316 15030
rect 6276 14612 6328 14618
rect 6276 14554 6328 14560
rect 6288 14482 6316 14554
rect 6092 14476 6144 14482
rect 6092 14418 6144 14424
rect 6276 14476 6328 14482
rect 6276 14418 6328 14424
rect 6104 13938 6132 14418
rect 6288 14074 6316 14418
rect 6368 14272 6420 14278
rect 6368 14214 6420 14220
rect 6276 14068 6328 14074
rect 6276 14010 6328 14016
rect 6092 13932 6144 13938
rect 6092 13874 6144 13880
rect 6104 13462 6132 13874
rect 6092 13456 6144 13462
rect 6092 13398 6144 13404
rect 6092 12708 6144 12714
rect 6092 12650 6144 12656
rect 6104 12374 6132 12650
rect 6380 12646 6408 14214
rect 6368 12640 6420 12646
rect 6368 12582 6420 12588
rect 6092 12368 6144 12374
rect 6092 12310 6144 12316
rect 6104 11694 6132 12310
rect 6184 12300 6236 12306
rect 6184 12242 6236 12248
rect 6196 11898 6224 12242
rect 6380 12170 6408 12582
rect 6472 12238 6500 15642
rect 6656 15162 6684 16050
rect 6748 15978 6776 16594
rect 6736 15972 6788 15978
rect 6736 15914 6788 15920
rect 6644 15156 6696 15162
rect 6644 15098 6696 15104
rect 7196 15020 7248 15026
rect 7196 14962 7248 14968
rect 7288 15020 7340 15026
rect 7288 14962 7340 14968
rect 6828 14884 6880 14890
rect 6828 14826 6880 14832
rect 6840 14618 6868 14826
rect 6828 14612 6880 14618
rect 6828 14554 6880 14560
rect 7208 14550 7236 14962
rect 7300 14929 7328 14962
rect 7286 14920 7342 14929
rect 7286 14855 7342 14864
rect 7196 14544 7248 14550
rect 7196 14486 7248 14492
rect 6918 13968 6974 13977
rect 6918 13903 6974 13912
rect 6932 13734 6960 13903
rect 7288 13864 7340 13870
rect 7288 13806 7340 13812
rect 6920 13728 6972 13734
rect 7300 13705 7328 13806
rect 6920 13670 6972 13676
rect 7286 13696 7342 13705
rect 7286 13631 7342 13640
rect 7300 13530 7328 13631
rect 7288 13524 7340 13530
rect 7288 13466 7340 13472
rect 7288 13320 7340 13326
rect 7288 13262 7340 13268
rect 6644 12436 6696 12442
rect 6644 12378 6696 12384
rect 6460 12232 6512 12238
rect 6460 12174 6512 12180
rect 6368 12164 6420 12170
rect 6368 12106 6420 12112
rect 6184 11892 6236 11898
rect 6184 11834 6236 11840
rect 6092 11688 6144 11694
rect 6092 11630 6144 11636
rect 6184 11212 6236 11218
rect 6184 11154 6236 11160
rect 6092 11144 6144 11150
rect 6092 11086 6144 11092
rect 6104 10810 6132 11086
rect 6092 10804 6144 10810
rect 6092 10746 6144 10752
rect 6196 10198 6224 11154
rect 6380 11014 6408 12106
rect 6472 11830 6500 12174
rect 6656 11898 6684 12378
rect 7104 12164 7156 12170
rect 7104 12106 7156 12112
rect 6736 12096 6788 12102
rect 6736 12038 6788 12044
rect 6644 11892 6696 11898
rect 6644 11834 6696 11840
rect 6460 11824 6512 11830
rect 6460 11766 6512 11772
rect 6472 11354 6500 11766
rect 6656 11694 6684 11834
rect 6644 11688 6696 11694
rect 6644 11630 6696 11636
rect 6460 11348 6512 11354
rect 6460 11290 6512 11296
rect 6472 11150 6500 11290
rect 6460 11144 6512 11150
rect 6460 11086 6512 11092
rect 6368 11008 6420 11014
rect 6368 10950 6420 10956
rect 6380 10810 6408 10950
rect 6368 10804 6420 10810
rect 6368 10746 6420 10752
rect 6748 10606 6776 12038
rect 7116 11830 7144 12106
rect 7300 11898 7328 13262
rect 7392 12782 7420 16934
rect 8956 16892 9252 16912
rect 9012 16890 9036 16892
rect 9092 16890 9116 16892
rect 9172 16890 9196 16892
rect 9034 16838 9036 16890
rect 9098 16838 9110 16890
rect 9172 16838 9174 16890
rect 9012 16836 9036 16838
rect 9092 16836 9116 16838
rect 9172 16836 9196 16838
rect 8956 16816 9252 16836
rect 7746 16688 7802 16697
rect 7746 16623 7802 16632
rect 7760 16250 7788 16623
rect 7748 16244 7800 16250
rect 7748 16186 7800 16192
rect 7840 16040 7892 16046
rect 7840 15982 7892 15988
rect 7564 15972 7616 15978
rect 7564 15914 7616 15920
rect 7472 13932 7524 13938
rect 7472 13874 7524 13880
rect 7484 13258 7512 13874
rect 7576 13394 7604 15914
rect 7852 15638 7880 15982
rect 9600 15978 9628 23582
rect 9954 23520 10010 23582
rect 13832 23582 13966 23610
rect 12956 21788 13252 21808
rect 13012 21786 13036 21788
rect 13092 21786 13116 21788
rect 13172 21786 13196 21788
rect 13034 21734 13036 21786
rect 13098 21734 13110 21786
rect 13172 21734 13174 21786
rect 13012 21732 13036 21734
rect 13092 21732 13116 21734
rect 13172 21732 13196 21734
rect 12956 21712 13252 21732
rect 12956 20700 13252 20720
rect 13012 20698 13036 20700
rect 13092 20698 13116 20700
rect 13172 20698 13196 20700
rect 13034 20646 13036 20698
rect 13098 20646 13110 20698
rect 13172 20646 13174 20698
rect 13012 20644 13036 20646
rect 13092 20644 13116 20646
rect 13172 20644 13196 20646
rect 12956 20624 13252 20644
rect 12956 19612 13252 19632
rect 13012 19610 13036 19612
rect 13092 19610 13116 19612
rect 13172 19610 13196 19612
rect 13034 19558 13036 19610
rect 13098 19558 13110 19610
rect 13172 19558 13174 19610
rect 13012 19556 13036 19558
rect 13092 19556 13116 19558
rect 13172 19556 13196 19558
rect 12956 19536 13252 19556
rect 12956 18524 13252 18544
rect 13012 18522 13036 18524
rect 13092 18522 13116 18524
rect 13172 18522 13196 18524
rect 13034 18470 13036 18522
rect 13098 18470 13110 18522
rect 13172 18470 13174 18522
rect 13012 18468 13036 18470
rect 13092 18468 13116 18470
rect 13172 18468 13196 18470
rect 12956 18448 13252 18468
rect 12956 17436 13252 17456
rect 13012 17434 13036 17436
rect 13092 17434 13116 17436
rect 13172 17434 13196 17436
rect 13034 17382 13036 17434
rect 13098 17382 13110 17434
rect 13172 17382 13174 17434
rect 13012 17380 13036 17382
rect 13092 17380 13116 17382
rect 13172 17380 13196 17382
rect 12956 17360 13252 17380
rect 13832 17105 13860 23582
rect 13910 23520 13966 23582
rect 17696 23582 18014 23610
rect 16956 21244 17252 21264
rect 17012 21242 17036 21244
rect 17092 21242 17116 21244
rect 17172 21242 17196 21244
rect 17034 21190 17036 21242
rect 17098 21190 17110 21242
rect 17172 21190 17174 21242
rect 17012 21188 17036 21190
rect 17092 21188 17116 21190
rect 17172 21188 17196 21190
rect 16956 21168 17252 21188
rect 16956 20156 17252 20176
rect 17012 20154 17036 20156
rect 17092 20154 17116 20156
rect 17172 20154 17196 20156
rect 17034 20102 17036 20154
rect 17098 20102 17110 20154
rect 17172 20102 17174 20154
rect 17012 20100 17036 20102
rect 17092 20100 17116 20102
rect 17172 20100 17196 20102
rect 16956 20080 17252 20100
rect 16956 19068 17252 19088
rect 17012 19066 17036 19068
rect 17092 19066 17116 19068
rect 17172 19066 17196 19068
rect 17034 19014 17036 19066
rect 17098 19014 17110 19066
rect 17172 19014 17174 19066
rect 17012 19012 17036 19014
rect 17092 19012 17116 19014
rect 17172 19012 17196 19014
rect 16956 18992 17252 19012
rect 16956 17980 17252 18000
rect 17012 17978 17036 17980
rect 17092 17978 17116 17980
rect 17172 17978 17196 17980
rect 17034 17926 17036 17978
rect 17098 17926 17110 17978
rect 17172 17926 17174 17978
rect 17012 17924 17036 17926
rect 17092 17924 17116 17926
rect 17172 17924 17196 17926
rect 16956 17904 17252 17924
rect 13818 17096 13874 17105
rect 13818 17031 13874 17040
rect 16956 16892 17252 16912
rect 17012 16890 17036 16892
rect 17092 16890 17116 16892
rect 17172 16890 17196 16892
rect 17034 16838 17036 16890
rect 17098 16838 17110 16890
rect 17172 16838 17174 16890
rect 17012 16836 17036 16838
rect 17092 16836 17116 16838
rect 17172 16836 17196 16838
rect 16956 16816 17252 16836
rect 17696 16697 17724 23582
rect 17958 23520 18014 23582
rect 21914 23610 21970 24000
rect 21914 23582 22048 23610
rect 21914 23520 21970 23582
rect 20956 21788 21252 21808
rect 21012 21786 21036 21788
rect 21092 21786 21116 21788
rect 21172 21786 21196 21788
rect 21034 21734 21036 21786
rect 21098 21734 21110 21786
rect 21172 21734 21174 21786
rect 21012 21732 21036 21734
rect 21092 21732 21116 21734
rect 21172 21732 21196 21734
rect 20956 21712 21252 21732
rect 20956 20700 21252 20720
rect 21012 20698 21036 20700
rect 21092 20698 21116 20700
rect 21172 20698 21196 20700
rect 21034 20646 21036 20698
rect 21098 20646 21110 20698
rect 21172 20646 21174 20698
rect 21012 20644 21036 20646
rect 21092 20644 21116 20646
rect 21172 20644 21196 20646
rect 20956 20624 21252 20644
rect 20956 19612 21252 19632
rect 21012 19610 21036 19612
rect 21092 19610 21116 19612
rect 21172 19610 21196 19612
rect 21034 19558 21036 19610
rect 21098 19558 21110 19610
rect 21172 19558 21174 19610
rect 21012 19556 21036 19558
rect 21092 19556 21116 19558
rect 21172 19556 21196 19558
rect 20956 19536 21252 19556
rect 20956 18524 21252 18544
rect 21012 18522 21036 18524
rect 21092 18522 21116 18524
rect 21172 18522 21196 18524
rect 21034 18470 21036 18522
rect 21098 18470 21110 18522
rect 21172 18470 21174 18522
rect 21012 18468 21036 18470
rect 21092 18468 21116 18470
rect 21172 18468 21196 18470
rect 20956 18448 21252 18468
rect 20956 17436 21252 17456
rect 21012 17434 21036 17436
rect 21092 17434 21116 17436
rect 21172 17434 21196 17436
rect 21034 17382 21036 17434
rect 21098 17382 21110 17434
rect 21172 17382 21174 17434
rect 21012 17380 21036 17382
rect 21092 17380 21116 17382
rect 21172 17380 21196 17382
rect 20956 17360 21252 17380
rect 17682 16688 17738 16697
rect 17682 16623 17738 16632
rect 12956 16348 13252 16368
rect 13012 16346 13036 16348
rect 13092 16346 13116 16348
rect 13172 16346 13196 16348
rect 13034 16294 13036 16346
rect 13098 16294 13110 16346
rect 13172 16294 13174 16346
rect 13012 16292 13036 16294
rect 13092 16292 13116 16294
rect 13172 16292 13196 16294
rect 12956 16272 13252 16292
rect 20956 16348 21252 16368
rect 21012 16346 21036 16348
rect 21092 16346 21116 16348
rect 21172 16346 21196 16348
rect 21034 16294 21036 16346
rect 21098 16294 21110 16346
rect 21172 16294 21174 16346
rect 21012 16292 21036 16294
rect 21092 16292 21116 16294
rect 21172 16292 21196 16294
rect 20956 16272 21252 16292
rect 9588 15972 9640 15978
rect 9588 15914 9640 15920
rect 8956 15804 9252 15824
rect 9012 15802 9036 15804
rect 9092 15802 9116 15804
rect 9172 15802 9196 15804
rect 9034 15750 9036 15802
rect 9098 15750 9110 15802
rect 9172 15750 9174 15802
rect 9012 15748 9036 15750
rect 9092 15748 9116 15750
rect 9172 15748 9196 15750
rect 8956 15728 9252 15748
rect 16956 15804 17252 15824
rect 17012 15802 17036 15804
rect 17092 15802 17116 15804
rect 17172 15802 17196 15804
rect 17034 15750 17036 15802
rect 17098 15750 17110 15802
rect 17172 15750 17174 15802
rect 17012 15748 17036 15750
rect 17092 15748 17116 15750
rect 17172 15748 17196 15750
rect 16956 15728 17252 15748
rect 7840 15632 7892 15638
rect 7654 15600 7710 15609
rect 22020 15609 22048 23582
rect 7840 15574 7892 15580
rect 22006 15600 22062 15609
rect 7654 15535 7710 15544
rect 7668 15502 7696 15535
rect 7656 15496 7708 15502
rect 7656 15438 7708 15444
rect 7852 14618 7880 15574
rect 22006 15535 22062 15544
rect 12956 15260 13252 15280
rect 13012 15258 13036 15260
rect 13092 15258 13116 15260
rect 13172 15258 13196 15260
rect 13034 15206 13036 15258
rect 13098 15206 13110 15258
rect 13172 15206 13174 15258
rect 13012 15204 13036 15206
rect 13092 15204 13116 15206
rect 13172 15204 13196 15206
rect 12956 15184 13252 15204
rect 20956 15260 21252 15280
rect 21012 15258 21036 15260
rect 21092 15258 21116 15260
rect 21172 15258 21196 15260
rect 21034 15206 21036 15258
rect 21098 15206 21110 15258
rect 21172 15206 21174 15258
rect 21012 15204 21036 15206
rect 21092 15204 21116 15206
rect 21172 15204 21196 15206
rect 20956 15184 21252 15204
rect 8956 14716 9252 14736
rect 9012 14714 9036 14716
rect 9092 14714 9116 14716
rect 9172 14714 9196 14716
rect 9034 14662 9036 14714
rect 9098 14662 9110 14714
rect 9172 14662 9174 14714
rect 9012 14660 9036 14662
rect 9092 14660 9116 14662
rect 9172 14660 9196 14662
rect 8956 14640 9252 14660
rect 16956 14716 17252 14736
rect 17012 14714 17036 14716
rect 17092 14714 17116 14716
rect 17172 14714 17196 14716
rect 17034 14662 17036 14714
rect 17098 14662 17110 14714
rect 17172 14662 17174 14714
rect 17012 14660 17036 14662
rect 17092 14660 17116 14662
rect 17172 14660 17196 14662
rect 16956 14640 17252 14660
rect 7840 14612 7892 14618
rect 7840 14554 7892 14560
rect 12956 14172 13252 14192
rect 13012 14170 13036 14172
rect 13092 14170 13116 14172
rect 13172 14170 13196 14172
rect 13034 14118 13036 14170
rect 13098 14118 13110 14170
rect 13172 14118 13174 14170
rect 13012 14116 13036 14118
rect 13092 14116 13116 14118
rect 13172 14116 13196 14118
rect 12956 14096 13252 14116
rect 20956 14172 21252 14192
rect 21012 14170 21036 14172
rect 21092 14170 21116 14172
rect 21172 14170 21196 14172
rect 21034 14118 21036 14170
rect 21098 14118 21110 14170
rect 21172 14118 21174 14170
rect 21012 14116 21036 14118
rect 21092 14116 21116 14118
rect 21172 14116 21196 14118
rect 20956 14096 21252 14116
rect 8956 13628 9252 13648
rect 9012 13626 9036 13628
rect 9092 13626 9116 13628
rect 9172 13626 9196 13628
rect 9034 13574 9036 13626
rect 9098 13574 9110 13626
rect 9172 13574 9174 13626
rect 9012 13572 9036 13574
rect 9092 13572 9116 13574
rect 9172 13572 9196 13574
rect 8956 13552 9252 13572
rect 16956 13628 17252 13648
rect 17012 13626 17036 13628
rect 17092 13626 17116 13628
rect 17172 13626 17196 13628
rect 17034 13574 17036 13626
rect 17098 13574 17110 13626
rect 17172 13574 17174 13626
rect 17012 13572 17036 13574
rect 17092 13572 17116 13574
rect 17172 13572 17196 13574
rect 16956 13552 17252 13572
rect 7564 13388 7616 13394
rect 7564 13330 7616 13336
rect 7472 13252 7524 13258
rect 7472 13194 7524 13200
rect 7380 12776 7432 12782
rect 7380 12718 7432 12724
rect 7392 12442 7420 12718
rect 7380 12436 7432 12442
rect 7380 12378 7432 12384
rect 7392 11898 7420 12378
rect 7288 11892 7340 11898
rect 7288 11834 7340 11840
rect 7380 11892 7432 11898
rect 7380 11834 7432 11840
rect 7104 11824 7156 11830
rect 7104 11766 7156 11772
rect 7012 11688 7064 11694
rect 7012 11630 7064 11636
rect 6920 11552 6972 11558
rect 6920 11494 6972 11500
rect 6736 10600 6788 10606
rect 6736 10542 6788 10548
rect 6000 10192 6052 10198
rect 6000 10134 6052 10140
rect 6184 10192 6236 10198
rect 6184 10134 6236 10140
rect 6644 10124 6696 10130
rect 6644 10066 6696 10072
rect 6656 9586 6684 10066
rect 6736 9988 6788 9994
rect 6736 9930 6788 9936
rect 6748 9722 6776 9930
rect 6736 9716 6788 9722
rect 6736 9658 6788 9664
rect 6644 9580 6696 9586
rect 6644 9522 6696 9528
rect 6656 9178 6684 9522
rect 6644 9172 6696 9178
rect 6644 9114 6696 9120
rect 6184 8356 6236 8362
rect 6184 8298 6236 8304
rect 6092 7948 6144 7954
rect 6092 7890 6144 7896
rect 6104 7546 6132 7890
rect 6196 7818 6224 8298
rect 6932 7954 6960 11494
rect 7024 11082 7052 11630
rect 7196 11212 7248 11218
rect 7300 11200 7328 11834
rect 7484 11218 7512 13194
rect 7576 12986 7604 13330
rect 12956 13084 13252 13104
rect 13012 13082 13036 13084
rect 13092 13082 13116 13084
rect 13172 13082 13196 13084
rect 13034 13030 13036 13082
rect 13098 13030 13110 13082
rect 13172 13030 13174 13082
rect 13012 13028 13036 13030
rect 13092 13028 13116 13030
rect 13172 13028 13196 13030
rect 12956 13008 13252 13028
rect 20956 13084 21252 13104
rect 21012 13082 21036 13084
rect 21092 13082 21116 13084
rect 21172 13082 21196 13084
rect 21034 13030 21036 13082
rect 21098 13030 21110 13082
rect 21172 13030 21174 13082
rect 21012 13028 21036 13030
rect 21092 13028 21116 13030
rect 21172 13028 21196 13030
rect 20956 13008 21252 13028
rect 7564 12980 7616 12986
rect 7564 12922 7616 12928
rect 7576 12306 7604 12922
rect 8956 12540 9252 12560
rect 9012 12538 9036 12540
rect 9092 12538 9116 12540
rect 9172 12538 9196 12540
rect 9034 12486 9036 12538
rect 9098 12486 9110 12538
rect 9172 12486 9174 12538
rect 9012 12484 9036 12486
rect 9092 12484 9116 12486
rect 9172 12484 9196 12486
rect 8956 12464 9252 12484
rect 16956 12540 17252 12560
rect 17012 12538 17036 12540
rect 17092 12538 17116 12540
rect 17172 12538 17196 12540
rect 17034 12486 17036 12538
rect 17098 12486 17110 12538
rect 17172 12486 17174 12538
rect 17012 12484 17036 12486
rect 17092 12484 17116 12486
rect 17172 12484 17196 12486
rect 16956 12464 17252 12484
rect 7564 12300 7616 12306
rect 7564 12242 7616 12248
rect 7576 11830 7604 12242
rect 7932 12164 7984 12170
rect 7932 12106 7984 12112
rect 7564 11824 7616 11830
rect 7564 11766 7616 11772
rect 7944 11354 7972 12106
rect 8024 12096 8076 12102
rect 8024 12038 8076 12044
rect 7932 11348 7984 11354
rect 7932 11290 7984 11296
rect 7248 11172 7328 11200
rect 7196 11154 7248 11160
rect 7012 11076 7064 11082
rect 7012 11018 7064 11024
rect 7300 10810 7328 11172
rect 7472 11212 7524 11218
rect 7524 11172 7604 11200
rect 7472 11154 7524 11160
rect 7472 11008 7524 11014
rect 7472 10950 7524 10956
rect 7288 10804 7340 10810
rect 7288 10746 7340 10752
rect 7484 10713 7512 10950
rect 7576 10810 7604 11172
rect 7564 10804 7616 10810
rect 7564 10746 7616 10752
rect 7470 10704 7526 10713
rect 7470 10639 7526 10648
rect 7288 10124 7340 10130
rect 7288 10066 7340 10072
rect 7300 9382 7328 10066
rect 7288 9376 7340 9382
rect 7288 9318 7340 9324
rect 6920 7948 6972 7954
rect 6920 7890 6972 7896
rect 6184 7812 6236 7818
rect 6184 7754 6236 7760
rect 7300 7546 7328 9318
rect 6092 7540 6144 7546
rect 6092 7482 6144 7488
rect 7288 7540 7340 7546
rect 7288 7482 7340 7488
rect 8036 7478 8064 12038
rect 12956 11996 13252 12016
rect 13012 11994 13036 11996
rect 13092 11994 13116 11996
rect 13172 11994 13196 11996
rect 13034 11942 13036 11994
rect 13098 11942 13110 11994
rect 13172 11942 13174 11994
rect 13012 11940 13036 11942
rect 13092 11940 13116 11942
rect 13172 11940 13196 11942
rect 12956 11920 13252 11940
rect 20956 11996 21252 12016
rect 21012 11994 21036 11996
rect 21092 11994 21116 11996
rect 21172 11994 21196 11996
rect 21034 11942 21036 11994
rect 21098 11942 21110 11994
rect 21172 11942 21174 11994
rect 21012 11940 21036 11942
rect 21092 11940 21116 11942
rect 21172 11940 21196 11942
rect 20956 11920 21252 11940
rect 8956 11452 9252 11472
rect 9012 11450 9036 11452
rect 9092 11450 9116 11452
rect 9172 11450 9196 11452
rect 9034 11398 9036 11450
rect 9098 11398 9110 11450
rect 9172 11398 9174 11450
rect 9012 11396 9036 11398
rect 9092 11396 9116 11398
rect 9172 11396 9196 11398
rect 8956 11376 9252 11396
rect 16956 11452 17252 11472
rect 17012 11450 17036 11452
rect 17092 11450 17116 11452
rect 17172 11450 17196 11452
rect 17034 11398 17036 11450
rect 17098 11398 17110 11450
rect 17172 11398 17174 11450
rect 17012 11396 17036 11398
rect 17092 11396 17116 11398
rect 17172 11396 17196 11398
rect 16956 11376 17252 11396
rect 12956 10908 13252 10928
rect 13012 10906 13036 10908
rect 13092 10906 13116 10908
rect 13172 10906 13196 10908
rect 13034 10854 13036 10906
rect 13098 10854 13110 10906
rect 13172 10854 13174 10906
rect 13012 10852 13036 10854
rect 13092 10852 13116 10854
rect 13172 10852 13196 10854
rect 12956 10832 13252 10852
rect 20956 10908 21252 10928
rect 21012 10906 21036 10908
rect 21092 10906 21116 10908
rect 21172 10906 21196 10908
rect 21034 10854 21036 10906
rect 21098 10854 21110 10906
rect 21172 10854 21174 10906
rect 21012 10852 21036 10854
rect 21092 10852 21116 10854
rect 21172 10852 21196 10854
rect 20956 10832 21252 10852
rect 8956 10364 9252 10384
rect 9012 10362 9036 10364
rect 9092 10362 9116 10364
rect 9172 10362 9196 10364
rect 9034 10310 9036 10362
rect 9098 10310 9110 10362
rect 9172 10310 9174 10362
rect 9012 10308 9036 10310
rect 9092 10308 9116 10310
rect 9172 10308 9196 10310
rect 8956 10288 9252 10308
rect 16956 10364 17252 10384
rect 17012 10362 17036 10364
rect 17092 10362 17116 10364
rect 17172 10362 17196 10364
rect 17034 10310 17036 10362
rect 17098 10310 17110 10362
rect 17172 10310 17174 10362
rect 17012 10308 17036 10310
rect 17092 10308 17116 10310
rect 17172 10308 17196 10310
rect 16956 10288 17252 10308
rect 12956 9820 13252 9840
rect 13012 9818 13036 9820
rect 13092 9818 13116 9820
rect 13172 9818 13196 9820
rect 13034 9766 13036 9818
rect 13098 9766 13110 9818
rect 13172 9766 13174 9818
rect 13012 9764 13036 9766
rect 13092 9764 13116 9766
rect 13172 9764 13196 9766
rect 12956 9744 13252 9764
rect 20956 9820 21252 9840
rect 21012 9818 21036 9820
rect 21092 9818 21116 9820
rect 21172 9818 21196 9820
rect 21034 9766 21036 9818
rect 21098 9766 21110 9818
rect 21172 9766 21174 9818
rect 21012 9764 21036 9766
rect 21092 9764 21116 9766
rect 21172 9764 21196 9766
rect 20956 9744 21252 9764
rect 8956 9276 9252 9296
rect 9012 9274 9036 9276
rect 9092 9274 9116 9276
rect 9172 9274 9196 9276
rect 9034 9222 9036 9274
rect 9098 9222 9110 9274
rect 9172 9222 9174 9274
rect 9012 9220 9036 9222
rect 9092 9220 9116 9222
rect 9172 9220 9196 9222
rect 8956 9200 9252 9220
rect 16956 9276 17252 9296
rect 17012 9274 17036 9276
rect 17092 9274 17116 9276
rect 17172 9274 17196 9276
rect 17034 9222 17036 9274
rect 17098 9222 17110 9274
rect 17172 9222 17174 9274
rect 17012 9220 17036 9222
rect 17092 9220 17116 9222
rect 17172 9220 17196 9222
rect 16956 9200 17252 9220
rect 12956 8732 13252 8752
rect 13012 8730 13036 8732
rect 13092 8730 13116 8732
rect 13172 8730 13196 8732
rect 13034 8678 13036 8730
rect 13098 8678 13110 8730
rect 13172 8678 13174 8730
rect 13012 8676 13036 8678
rect 13092 8676 13116 8678
rect 13172 8676 13196 8678
rect 12956 8656 13252 8676
rect 20956 8732 21252 8752
rect 21012 8730 21036 8732
rect 21092 8730 21116 8732
rect 21172 8730 21196 8732
rect 21034 8678 21036 8730
rect 21098 8678 21110 8730
rect 21172 8678 21174 8730
rect 21012 8676 21036 8678
rect 21092 8676 21116 8678
rect 21172 8676 21196 8678
rect 20956 8656 21252 8676
rect 8956 8188 9252 8208
rect 9012 8186 9036 8188
rect 9092 8186 9116 8188
rect 9172 8186 9196 8188
rect 9034 8134 9036 8186
rect 9098 8134 9110 8186
rect 9172 8134 9174 8186
rect 9012 8132 9036 8134
rect 9092 8132 9116 8134
rect 9172 8132 9196 8134
rect 8956 8112 9252 8132
rect 16956 8188 17252 8208
rect 17012 8186 17036 8188
rect 17092 8186 17116 8188
rect 17172 8186 17196 8188
rect 17034 8134 17036 8186
rect 17098 8134 17110 8186
rect 17172 8134 17174 8186
rect 17012 8132 17036 8134
rect 17092 8132 17116 8134
rect 17172 8132 17196 8134
rect 16956 8112 17252 8132
rect 12956 7644 13252 7664
rect 13012 7642 13036 7644
rect 13092 7642 13116 7644
rect 13172 7642 13196 7644
rect 13034 7590 13036 7642
rect 13098 7590 13110 7642
rect 13172 7590 13174 7642
rect 13012 7588 13036 7590
rect 13092 7588 13116 7590
rect 13172 7588 13196 7590
rect 12956 7568 13252 7588
rect 20956 7644 21252 7664
rect 21012 7642 21036 7644
rect 21092 7642 21116 7644
rect 21172 7642 21196 7644
rect 21034 7590 21036 7642
rect 21098 7590 21110 7642
rect 21172 7590 21174 7642
rect 21012 7588 21036 7590
rect 21092 7588 21116 7590
rect 21172 7588 21196 7590
rect 20956 7568 21252 7588
rect 8024 7472 8076 7478
rect 8024 7414 8076 7420
rect 12072 7336 12124 7342
rect 12072 7278 12124 7284
rect 8956 7100 9252 7120
rect 9012 7098 9036 7100
rect 9092 7098 9116 7100
rect 9172 7098 9196 7100
rect 9034 7046 9036 7098
rect 9098 7046 9110 7098
rect 9172 7046 9174 7098
rect 9012 7044 9036 7046
rect 9092 7044 9116 7046
rect 9172 7044 9196 7046
rect 8956 7024 9252 7044
rect 8956 6012 9252 6032
rect 9012 6010 9036 6012
rect 9092 6010 9116 6012
rect 9172 6010 9196 6012
rect 9034 5958 9036 6010
rect 9098 5958 9110 6010
rect 9172 5958 9174 6010
rect 9012 5956 9036 5958
rect 9092 5956 9116 5958
rect 9172 5956 9196 5958
rect 8956 5936 9252 5956
rect 8956 4924 9252 4944
rect 9012 4922 9036 4924
rect 9092 4922 9116 4924
rect 9172 4922 9196 4924
rect 9034 4870 9036 4922
rect 9098 4870 9110 4922
rect 9172 4870 9174 4922
rect 9012 4868 9036 4870
rect 9092 4868 9116 4870
rect 9172 4868 9196 4870
rect 8956 4848 9252 4868
rect 8956 3836 9252 3856
rect 9012 3834 9036 3836
rect 9092 3834 9116 3836
rect 9172 3834 9196 3836
rect 9034 3782 9036 3834
rect 9098 3782 9110 3834
rect 9172 3782 9174 3834
rect 9012 3780 9036 3782
rect 9092 3780 9116 3782
rect 9172 3780 9196 3782
rect 8956 3760 9252 3780
rect 5908 3188 5960 3194
rect 5908 3130 5960 3136
rect 4620 3120 4672 3126
rect 4620 3062 4672 3068
rect 4068 3052 4120 3058
rect 4068 2994 4120 3000
rect 3884 2984 3936 2990
rect 3884 2926 3936 2932
rect 3792 2848 3844 2854
rect 3792 2790 3844 2796
rect 3516 2644 3568 2650
rect 3516 2586 3568 2592
rect 3804 1358 3832 2790
rect 4632 2514 4660 3062
rect 8956 2748 9252 2768
rect 9012 2746 9036 2748
rect 9092 2746 9116 2748
rect 9172 2746 9196 2748
rect 9034 2694 9036 2746
rect 9098 2694 9110 2746
rect 9172 2694 9174 2746
rect 9012 2692 9036 2694
rect 9092 2692 9116 2694
rect 9172 2692 9196 2694
rect 8956 2672 9252 2692
rect 4620 2508 4672 2514
rect 4620 2450 4672 2456
rect 4956 2204 5252 2224
rect 5012 2202 5036 2204
rect 5092 2202 5116 2204
rect 5172 2202 5196 2204
rect 5034 2150 5036 2202
rect 5098 2150 5110 2202
rect 5172 2150 5174 2202
rect 5012 2148 5036 2150
rect 5092 2148 5116 2150
rect 5172 2148 5196 2150
rect 4956 2128 5252 2148
rect 3792 1352 3844 1358
rect 3792 1294 3844 1300
rect 3422 640 3478 649
rect 3422 575 3478 584
rect 166 190 336 218
rect 110 167 166 176
rect 11978 82 12034 480
rect 12084 82 12112 7278
rect 16956 7100 17252 7120
rect 17012 7098 17036 7100
rect 17092 7098 17116 7100
rect 17172 7098 17196 7100
rect 17034 7046 17036 7098
rect 17098 7046 17110 7098
rect 17172 7046 17174 7098
rect 17012 7044 17036 7046
rect 17092 7044 17116 7046
rect 17172 7044 17196 7046
rect 16956 7024 17252 7044
rect 12956 6556 13252 6576
rect 13012 6554 13036 6556
rect 13092 6554 13116 6556
rect 13172 6554 13196 6556
rect 13034 6502 13036 6554
rect 13098 6502 13110 6554
rect 13172 6502 13174 6554
rect 13012 6500 13036 6502
rect 13092 6500 13116 6502
rect 13172 6500 13196 6502
rect 12956 6480 13252 6500
rect 20956 6556 21252 6576
rect 21012 6554 21036 6556
rect 21092 6554 21116 6556
rect 21172 6554 21196 6556
rect 21034 6502 21036 6554
rect 21098 6502 21110 6554
rect 21172 6502 21174 6554
rect 21012 6500 21036 6502
rect 21092 6500 21116 6502
rect 21172 6500 21196 6502
rect 20956 6480 21252 6500
rect 16956 6012 17252 6032
rect 17012 6010 17036 6012
rect 17092 6010 17116 6012
rect 17172 6010 17196 6012
rect 17034 5958 17036 6010
rect 17098 5958 17110 6010
rect 17172 5958 17174 6010
rect 17012 5956 17036 5958
rect 17092 5956 17116 5958
rect 17172 5956 17196 5958
rect 16956 5936 17252 5956
rect 12956 5468 13252 5488
rect 13012 5466 13036 5468
rect 13092 5466 13116 5468
rect 13172 5466 13196 5468
rect 13034 5414 13036 5466
rect 13098 5414 13110 5466
rect 13172 5414 13174 5466
rect 13012 5412 13036 5414
rect 13092 5412 13116 5414
rect 13172 5412 13196 5414
rect 12956 5392 13252 5412
rect 20956 5468 21252 5488
rect 21012 5466 21036 5468
rect 21092 5466 21116 5468
rect 21172 5466 21196 5468
rect 21034 5414 21036 5466
rect 21098 5414 21110 5466
rect 21172 5414 21174 5466
rect 21012 5412 21036 5414
rect 21092 5412 21116 5414
rect 21172 5412 21196 5414
rect 20956 5392 21252 5412
rect 16956 4924 17252 4944
rect 17012 4922 17036 4924
rect 17092 4922 17116 4924
rect 17172 4922 17196 4924
rect 17034 4870 17036 4922
rect 17098 4870 17110 4922
rect 17172 4870 17174 4922
rect 17012 4868 17036 4870
rect 17092 4868 17116 4870
rect 17172 4868 17196 4870
rect 16956 4848 17252 4868
rect 12956 4380 13252 4400
rect 13012 4378 13036 4380
rect 13092 4378 13116 4380
rect 13172 4378 13196 4380
rect 13034 4326 13036 4378
rect 13098 4326 13110 4378
rect 13172 4326 13174 4378
rect 13012 4324 13036 4326
rect 13092 4324 13116 4326
rect 13172 4324 13196 4326
rect 12956 4304 13252 4324
rect 20956 4380 21252 4400
rect 21012 4378 21036 4380
rect 21092 4378 21116 4380
rect 21172 4378 21196 4380
rect 21034 4326 21036 4378
rect 21098 4326 21110 4378
rect 21172 4326 21174 4378
rect 21012 4324 21036 4326
rect 21092 4324 21116 4326
rect 21172 4324 21196 4326
rect 20956 4304 21252 4324
rect 16956 3836 17252 3856
rect 17012 3834 17036 3836
rect 17092 3834 17116 3836
rect 17172 3834 17196 3836
rect 17034 3782 17036 3834
rect 17098 3782 17110 3834
rect 17172 3782 17174 3834
rect 17012 3780 17036 3782
rect 17092 3780 17116 3782
rect 17172 3780 17196 3782
rect 16956 3760 17252 3780
rect 12956 3292 13252 3312
rect 13012 3290 13036 3292
rect 13092 3290 13116 3292
rect 13172 3290 13196 3292
rect 13034 3238 13036 3290
rect 13098 3238 13110 3290
rect 13172 3238 13174 3290
rect 13012 3236 13036 3238
rect 13092 3236 13116 3238
rect 13172 3236 13196 3238
rect 12956 3216 13252 3236
rect 20956 3292 21252 3312
rect 21012 3290 21036 3292
rect 21092 3290 21116 3292
rect 21172 3290 21196 3292
rect 21034 3238 21036 3290
rect 21098 3238 21110 3290
rect 21172 3238 21174 3290
rect 21012 3236 21036 3238
rect 21092 3236 21116 3238
rect 21172 3236 21196 3238
rect 20956 3216 21252 3236
rect 16956 2748 17252 2768
rect 17012 2746 17036 2748
rect 17092 2746 17116 2748
rect 17172 2746 17196 2748
rect 17034 2694 17036 2746
rect 17098 2694 17110 2746
rect 17172 2694 17174 2746
rect 17012 2692 17036 2694
rect 17092 2692 17116 2694
rect 17172 2692 17196 2694
rect 16956 2672 17252 2692
rect 12956 2204 13252 2224
rect 13012 2202 13036 2204
rect 13092 2202 13116 2204
rect 13172 2202 13196 2204
rect 13034 2150 13036 2202
rect 13098 2150 13110 2202
rect 13172 2150 13174 2202
rect 13012 2148 13036 2150
rect 13092 2148 13116 2150
rect 13172 2148 13196 2150
rect 12956 2128 13252 2148
rect 20956 2204 21252 2224
rect 21012 2202 21036 2204
rect 21092 2202 21116 2204
rect 21172 2202 21196 2204
rect 21034 2150 21036 2202
rect 21098 2150 21110 2202
rect 21172 2150 21174 2202
rect 21012 2148 21036 2150
rect 21092 2148 21116 2150
rect 21172 2148 21196 2150
rect 20956 2128 21252 2148
rect 11978 54 12112 82
rect 11978 0 12034 54
<< via2 >>
rect 110 23704 166 23760
rect 18 23296 74 23352
rect 110 22888 166 22944
rect 110 22480 166 22536
rect 110 21664 166 21720
rect 110 21256 166 21312
rect 110 19760 166 19816
rect 18 18536 74 18592
rect 386 20848 442 20904
rect 1766 20032 1822 20088
rect 110 18128 166 18184
rect 18 17720 74 17776
rect 18 17312 74 17368
rect 18 17040 74 17096
rect 110 16632 166 16688
rect 110 16224 166 16280
rect 18 15816 74 15872
rect 110 15000 166 15056
rect 110 14184 166 14240
rect 110 13504 166 13560
rect 18 13096 74 13152
rect 110 12688 166 12744
rect 18 12280 74 12336
rect 110 11872 166 11928
rect 18 11464 74 11520
rect 110 11056 166 11112
rect 110 10648 166 10704
rect 18 10376 74 10432
rect 110 9968 166 10024
rect 4956 21786 5012 21788
rect 5036 21786 5092 21788
rect 5116 21786 5172 21788
rect 5196 21786 5252 21788
rect 4956 21734 4982 21786
rect 4982 21734 5012 21786
rect 5036 21734 5046 21786
rect 5046 21734 5092 21786
rect 5116 21734 5162 21786
rect 5162 21734 5172 21786
rect 5196 21734 5226 21786
rect 5226 21734 5252 21786
rect 4956 21732 5012 21734
rect 5036 21732 5092 21734
rect 5116 21732 5172 21734
rect 5196 21732 5252 21734
rect 4710 21392 4766 21448
rect 4956 20698 5012 20700
rect 5036 20698 5092 20700
rect 5116 20698 5172 20700
rect 5196 20698 5252 20700
rect 4956 20646 4982 20698
rect 4982 20646 5012 20698
rect 5036 20646 5046 20698
rect 5046 20646 5092 20698
rect 5116 20646 5162 20698
rect 5162 20646 5172 20698
rect 5196 20646 5226 20698
rect 5226 20646 5252 20698
rect 4956 20644 5012 20646
rect 5036 20644 5092 20646
rect 5116 20644 5172 20646
rect 5196 20644 5252 20646
rect 4618 20168 4674 20224
rect 4956 19610 5012 19612
rect 5036 19610 5092 19612
rect 5116 19610 5172 19612
rect 5196 19610 5252 19612
rect 4956 19558 4982 19610
rect 4982 19558 5012 19610
rect 5036 19558 5046 19610
rect 5046 19558 5092 19610
rect 5116 19558 5162 19610
rect 5162 19558 5172 19610
rect 5196 19558 5226 19610
rect 5226 19558 5252 19610
rect 4956 19556 5012 19558
rect 5036 19556 5092 19558
rect 5116 19556 5172 19558
rect 5196 19556 5252 19558
rect 4250 19216 4306 19272
rect 3422 18672 3478 18728
rect 4956 18522 5012 18524
rect 5036 18522 5092 18524
rect 5116 18522 5172 18524
rect 5196 18522 5252 18524
rect 4956 18470 4982 18522
rect 4982 18470 5012 18522
rect 5036 18470 5046 18522
rect 5046 18470 5092 18522
rect 5116 18470 5162 18522
rect 5162 18470 5172 18522
rect 5196 18470 5226 18522
rect 5226 18470 5252 18522
rect 4956 18468 5012 18470
rect 5036 18468 5092 18470
rect 5116 18468 5172 18470
rect 5196 18468 5252 18470
rect 3238 15952 3294 16008
rect 3054 13776 3110 13832
rect 18 9152 74 9208
rect 110 8744 166 8800
rect 110 8336 166 8392
rect 110 7928 166 7984
rect 18 7520 74 7576
rect 1582 7248 1638 7304
rect 110 6840 166 6896
rect 110 6432 166 6488
rect 18 5616 74 5672
rect 110 5208 166 5264
rect 110 4800 166 4856
rect 110 4392 166 4448
rect 18 3984 74 4040
rect 110 3576 166 3632
rect 110 3304 166 3360
rect 18 2080 74 2136
rect 110 1672 166 1728
rect 18 1264 74 1320
rect 110 856 166 912
rect 110 176 166 232
rect 4956 17434 5012 17436
rect 5036 17434 5092 17436
rect 5116 17434 5172 17436
rect 5196 17434 5252 17436
rect 4956 17382 4982 17434
rect 4982 17382 5012 17434
rect 5036 17382 5046 17434
rect 5046 17382 5092 17434
rect 5116 17382 5162 17434
rect 5162 17382 5172 17434
rect 5196 17382 5226 17434
rect 5226 17382 5252 17434
rect 4956 17380 5012 17382
rect 5036 17380 5092 17382
rect 5116 17380 5172 17382
rect 5196 17380 5252 17382
rect 4956 16346 5012 16348
rect 5036 16346 5092 16348
rect 5116 16346 5172 16348
rect 5196 16346 5252 16348
rect 4956 16294 4982 16346
rect 4982 16294 5012 16346
rect 5036 16294 5046 16346
rect 5046 16294 5092 16346
rect 5116 16294 5162 16346
rect 5162 16294 5172 16346
rect 5196 16294 5226 16346
rect 5226 16294 5252 16346
rect 4956 16292 5012 16294
rect 5036 16292 5092 16294
rect 5116 16292 5172 16294
rect 5196 16292 5252 16294
rect 4342 14864 4398 14920
rect 4956 15258 5012 15260
rect 5036 15258 5092 15260
rect 5116 15258 5172 15260
rect 5196 15258 5252 15260
rect 4956 15206 4982 15258
rect 4982 15206 5012 15258
rect 5036 15206 5046 15258
rect 5046 15206 5092 15258
rect 5116 15206 5162 15258
rect 5162 15206 5172 15258
rect 5196 15206 5226 15258
rect 5226 15206 5252 15258
rect 4956 15204 5012 15206
rect 5036 15204 5092 15206
rect 5116 15204 5172 15206
rect 5196 15204 5252 15206
rect 4434 13640 4490 13696
rect 3606 10648 3662 10704
rect 3330 9424 3386 9480
rect 386 2896 442 2952
rect 386 2488 442 2544
rect 4956 14170 5012 14172
rect 5036 14170 5092 14172
rect 5116 14170 5172 14172
rect 5196 14170 5252 14172
rect 4956 14118 4982 14170
rect 4982 14118 5012 14170
rect 5036 14118 5046 14170
rect 5046 14118 5092 14170
rect 5116 14118 5162 14170
rect 5162 14118 5172 14170
rect 5196 14118 5226 14170
rect 5226 14118 5252 14170
rect 4956 14116 5012 14118
rect 5036 14116 5092 14118
rect 5116 14116 5172 14118
rect 5196 14116 5252 14118
rect 4956 13082 5012 13084
rect 5036 13082 5092 13084
rect 5116 13082 5172 13084
rect 5196 13082 5252 13084
rect 4956 13030 4982 13082
rect 4982 13030 5012 13082
rect 5036 13030 5046 13082
rect 5046 13030 5092 13082
rect 5116 13030 5162 13082
rect 5162 13030 5172 13082
rect 5196 13030 5226 13082
rect 5226 13030 5252 13082
rect 4956 13028 5012 13030
rect 5036 13028 5092 13030
rect 5116 13028 5172 13030
rect 5196 13028 5252 13030
rect 4956 11994 5012 11996
rect 5036 11994 5092 11996
rect 5116 11994 5172 11996
rect 5196 11994 5252 11996
rect 4956 11942 4982 11994
rect 4982 11942 5012 11994
rect 5036 11942 5046 11994
rect 5046 11942 5092 11994
rect 5116 11942 5162 11994
rect 5162 11942 5172 11994
rect 5196 11942 5226 11994
rect 5226 11942 5252 11994
rect 4956 11940 5012 11942
rect 5036 11940 5092 11942
rect 5116 11940 5172 11942
rect 5196 11940 5252 11942
rect 4956 10906 5012 10908
rect 5036 10906 5092 10908
rect 5116 10906 5172 10908
rect 5196 10906 5252 10908
rect 4956 10854 4982 10906
rect 4982 10854 5012 10906
rect 5036 10854 5046 10906
rect 5046 10854 5092 10906
rect 5116 10854 5162 10906
rect 5162 10854 5172 10906
rect 5196 10854 5226 10906
rect 5226 10854 5252 10906
rect 4956 10852 5012 10854
rect 5036 10852 5092 10854
rect 5116 10852 5172 10854
rect 5196 10852 5252 10854
rect 4956 9818 5012 9820
rect 5036 9818 5092 9820
rect 5116 9818 5172 9820
rect 5196 9818 5252 9820
rect 4956 9766 4982 9818
rect 4982 9766 5012 9818
rect 5036 9766 5046 9818
rect 5046 9766 5092 9818
rect 5116 9766 5162 9818
rect 5162 9766 5172 9818
rect 5196 9766 5226 9818
rect 5226 9766 5252 9818
rect 4956 9764 5012 9766
rect 5036 9764 5092 9766
rect 5116 9764 5172 9766
rect 5196 9764 5252 9766
rect 4956 8730 5012 8732
rect 5036 8730 5092 8732
rect 5116 8730 5172 8732
rect 5196 8730 5252 8732
rect 4956 8678 4982 8730
rect 4982 8678 5012 8730
rect 5036 8678 5046 8730
rect 5046 8678 5092 8730
rect 5116 8678 5162 8730
rect 5162 8678 5172 8730
rect 5196 8678 5226 8730
rect 5226 8678 5252 8730
rect 4956 8676 5012 8678
rect 5036 8676 5092 8678
rect 5116 8676 5172 8678
rect 5196 8676 5252 8678
rect 4956 7642 5012 7644
rect 5036 7642 5092 7644
rect 5116 7642 5172 7644
rect 5196 7642 5252 7644
rect 4956 7590 4982 7642
rect 4982 7590 5012 7642
rect 5036 7590 5046 7642
rect 5046 7590 5092 7642
rect 5116 7590 5162 7642
rect 5162 7590 5172 7642
rect 5196 7590 5226 7642
rect 5226 7590 5252 7642
rect 4956 7588 5012 7590
rect 5036 7588 5092 7590
rect 5116 7588 5172 7590
rect 5196 7588 5252 7590
rect 4956 6554 5012 6556
rect 5036 6554 5092 6556
rect 5116 6554 5172 6556
rect 5196 6554 5252 6556
rect 4956 6502 4982 6554
rect 4982 6502 5012 6554
rect 5036 6502 5046 6554
rect 5046 6502 5092 6554
rect 5116 6502 5162 6554
rect 5162 6502 5172 6554
rect 5196 6502 5226 6554
rect 5226 6502 5252 6554
rect 4956 6500 5012 6502
rect 5036 6500 5092 6502
rect 5116 6500 5172 6502
rect 5196 6500 5252 6502
rect 4956 5466 5012 5468
rect 5036 5466 5092 5468
rect 5116 5466 5172 5468
rect 5196 5466 5252 5468
rect 4956 5414 4982 5466
rect 4982 5414 5012 5466
rect 5036 5414 5046 5466
rect 5046 5414 5092 5466
rect 5116 5414 5162 5466
rect 5162 5414 5172 5466
rect 5196 5414 5226 5466
rect 5226 5414 5252 5466
rect 4956 5412 5012 5414
rect 5036 5412 5092 5414
rect 5116 5412 5172 5414
rect 5196 5412 5252 5414
rect 4158 4936 4214 4992
rect 4956 4378 5012 4380
rect 5036 4378 5092 4380
rect 5116 4378 5172 4380
rect 5196 4378 5252 4380
rect 4956 4326 4982 4378
rect 4982 4326 5012 4378
rect 5036 4326 5046 4378
rect 5046 4326 5092 4378
rect 5116 4326 5162 4378
rect 5162 4326 5172 4378
rect 5196 4326 5226 4378
rect 5226 4326 5252 4378
rect 4956 4324 5012 4326
rect 5036 4324 5092 4326
rect 5116 4324 5172 4326
rect 5196 4324 5252 4326
rect 4956 3290 5012 3292
rect 5036 3290 5092 3292
rect 5116 3290 5172 3292
rect 5196 3290 5252 3292
rect 4956 3238 4982 3290
rect 4982 3238 5012 3290
rect 5036 3238 5046 3290
rect 5046 3238 5092 3290
rect 5116 3238 5162 3290
rect 5162 3238 5172 3290
rect 5196 3238 5226 3290
rect 5226 3238 5252 3290
rect 4956 3236 5012 3238
rect 5036 3236 5092 3238
rect 5116 3236 5172 3238
rect 5196 3236 5252 3238
rect 8956 21242 9012 21244
rect 9036 21242 9092 21244
rect 9116 21242 9172 21244
rect 9196 21242 9252 21244
rect 8956 21190 8982 21242
rect 8982 21190 9012 21242
rect 9036 21190 9046 21242
rect 9046 21190 9092 21242
rect 9116 21190 9162 21242
rect 9162 21190 9172 21242
rect 9196 21190 9226 21242
rect 9226 21190 9252 21242
rect 8956 21188 9012 21190
rect 9036 21188 9092 21190
rect 9116 21188 9172 21190
rect 9196 21188 9252 21190
rect 8956 20154 9012 20156
rect 9036 20154 9092 20156
rect 9116 20154 9172 20156
rect 9196 20154 9252 20156
rect 8956 20102 8982 20154
rect 8982 20102 9012 20154
rect 9036 20102 9046 20154
rect 9046 20102 9092 20154
rect 9116 20102 9162 20154
rect 9162 20102 9172 20154
rect 9196 20102 9226 20154
rect 9226 20102 9252 20154
rect 8956 20100 9012 20102
rect 9036 20100 9092 20102
rect 9116 20100 9172 20102
rect 9196 20100 9252 20102
rect 8956 19066 9012 19068
rect 9036 19066 9092 19068
rect 9116 19066 9172 19068
rect 9196 19066 9252 19068
rect 8956 19014 8982 19066
rect 8982 19014 9012 19066
rect 9036 19014 9046 19066
rect 9046 19014 9092 19066
rect 9116 19014 9162 19066
rect 9162 19014 9172 19066
rect 9196 19014 9226 19066
rect 9226 19014 9252 19066
rect 8956 19012 9012 19014
rect 9036 19012 9092 19014
rect 9116 19012 9172 19014
rect 9196 19012 9252 19014
rect 8956 17978 9012 17980
rect 9036 17978 9092 17980
rect 9116 17978 9172 17980
rect 9196 17978 9252 17980
rect 8956 17926 8982 17978
rect 8982 17926 9012 17978
rect 9036 17926 9046 17978
rect 9046 17926 9092 17978
rect 9116 17926 9162 17978
rect 9162 17926 9172 17978
rect 9196 17926 9226 17978
rect 9226 17926 9252 17978
rect 8956 17924 9012 17926
rect 9036 17924 9092 17926
rect 9116 17924 9172 17926
rect 9196 17924 9252 17926
rect 7378 17076 7380 17096
rect 7380 17076 7432 17096
rect 7432 17076 7434 17096
rect 7378 17040 7434 17076
rect 7286 14864 7342 14920
rect 6918 13912 6974 13968
rect 7286 13640 7342 13696
rect 8956 16890 9012 16892
rect 9036 16890 9092 16892
rect 9116 16890 9172 16892
rect 9196 16890 9252 16892
rect 8956 16838 8982 16890
rect 8982 16838 9012 16890
rect 9036 16838 9046 16890
rect 9046 16838 9092 16890
rect 9116 16838 9162 16890
rect 9162 16838 9172 16890
rect 9196 16838 9226 16890
rect 9226 16838 9252 16890
rect 8956 16836 9012 16838
rect 9036 16836 9092 16838
rect 9116 16836 9172 16838
rect 9196 16836 9252 16838
rect 7746 16632 7802 16688
rect 12956 21786 13012 21788
rect 13036 21786 13092 21788
rect 13116 21786 13172 21788
rect 13196 21786 13252 21788
rect 12956 21734 12982 21786
rect 12982 21734 13012 21786
rect 13036 21734 13046 21786
rect 13046 21734 13092 21786
rect 13116 21734 13162 21786
rect 13162 21734 13172 21786
rect 13196 21734 13226 21786
rect 13226 21734 13252 21786
rect 12956 21732 13012 21734
rect 13036 21732 13092 21734
rect 13116 21732 13172 21734
rect 13196 21732 13252 21734
rect 12956 20698 13012 20700
rect 13036 20698 13092 20700
rect 13116 20698 13172 20700
rect 13196 20698 13252 20700
rect 12956 20646 12982 20698
rect 12982 20646 13012 20698
rect 13036 20646 13046 20698
rect 13046 20646 13092 20698
rect 13116 20646 13162 20698
rect 13162 20646 13172 20698
rect 13196 20646 13226 20698
rect 13226 20646 13252 20698
rect 12956 20644 13012 20646
rect 13036 20644 13092 20646
rect 13116 20644 13172 20646
rect 13196 20644 13252 20646
rect 12956 19610 13012 19612
rect 13036 19610 13092 19612
rect 13116 19610 13172 19612
rect 13196 19610 13252 19612
rect 12956 19558 12982 19610
rect 12982 19558 13012 19610
rect 13036 19558 13046 19610
rect 13046 19558 13092 19610
rect 13116 19558 13162 19610
rect 13162 19558 13172 19610
rect 13196 19558 13226 19610
rect 13226 19558 13252 19610
rect 12956 19556 13012 19558
rect 13036 19556 13092 19558
rect 13116 19556 13172 19558
rect 13196 19556 13252 19558
rect 12956 18522 13012 18524
rect 13036 18522 13092 18524
rect 13116 18522 13172 18524
rect 13196 18522 13252 18524
rect 12956 18470 12982 18522
rect 12982 18470 13012 18522
rect 13036 18470 13046 18522
rect 13046 18470 13092 18522
rect 13116 18470 13162 18522
rect 13162 18470 13172 18522
rect 13196 18470 13226 18522
rect 13226 18470 13252 18522
rect 12956 18468 13012 18470
rect 13036 18468 13092 18470
rect 13116 18468 13172 18470
rect 13196 18468 13252 18470
rect 12956 17434 13012 17436
rect 13036 17434 13092 17436
rect 13116 17434 13172 17436
rect 13196 17434 13252 17436
rect 12956 17382 12982 17434
rect 12982 17382 13012 17434
rect 13036 17382 13046 17434
rect 13046 17382 13092 17434
rect 13116 17382 13162 17434
rect 13162 17382 13172 17434
rect 13196 17382 13226 17434
rect 13226 17382 13252 17434
rect 12956 17380 13012 17382
rect 13036 17380 13092 17382
rect 13116 17380 13172 17382
rect 13196 17380 13252 17382
rect 16956 21242 17012 21244
rect 17036 21242 17092 21244
rect 17116 21242 17172 21244
rect 17196 21242 17252 21244
rect 16956 21190 16982 21242
rect 16982 21190 17012 21242
rect 17036 21190 17046 21242
rect 17046 21190 17092 21242
rect 17116 21190 17162 21242
rect 17162 21190 17172 21242
rect 17196 21190 17226 21242
rect 17226 21190 17252 21242
rect 16956 21188 17012 21190
rect 17036 21188 17092 21190
rect 17116 21188 17172 21190
rect 17196 21188 17252 21190
rect 16956 20154 17012 20156
rect 17036 20154 17092 20156
rect 17116 20154 17172 20156
rect 17196 20154 17252 20156
rect 16956 20102 16982 20154
rect 16982 20102 17012 20154
rect 17036 20102 17046 20154
rect 17046 20102 17092 20154
rect 17116 20102 17162 20154
rect 17162 20102 17172 20154
rect 17196 20102 17226 20154
rect 17226 20102 17252 20154
rect 16956 20100 17012 20102
rect 17036 20100 17092 20102
rect 17116 20100 17172 20102
rect 17196 20100 17252 20102
rect 16956 19066 17012 19068
rect 17036 19066 17092 19068
rect 17116 19066 17172 19068
rect 17196 19066 17252 19068
rect 16956 19014 16982 19066
rect 16982 19014 17012 19066
rect 17036 19014 17046 19066
rect 17046 19014 17092 19066
rect 17116 19014 17162 19066
rect 17162 19014 17172 19066
rect 17196 19014 17226 19066
rect 17226 19014 17252 19066
rect 16956 19012 17012 19014
rect 17036 19012 17092 19014
rect 17116 19012 17172 19014
rect 17196 19012 17252 19014
rect 16956 17978 17012 17980
rect 17036 17978 17092 17980
rect 17116 17978 17172 17980
rect 17196 17978 17252 17980
rect 16956 17926 16982 17978
rect 16982 17926 17012 17978
rect 17036 17926 17046 17978
rect 17046 17926 17092 17978
rect 17116 17926 17162 17978
rect 17162 17926 17172 17978
rect 17196 17926 17226 17978
rect 17226 17926 17252 17978
rect 16956 17924 17012 17926
rect 17036 17924 17092 17926
rect 17116 17924 17172 17926
rect 17196 17924 17252 17926
rect 13818 17040 13874 17096
rect 16956 16890 17012 16892
rect 17036 16890 17092 16892
rect 17116 16890 17172 16892
rect 17196 16890 17252 16892
rect 16956 16838 16982 16890
rect 16982 16838 17012 16890
rect 17036 16838 17046 16890
rect 17046 16838 17092 16890
rect 17116 16838 17162 16890
rect 17162 16838 17172 16890
rect 17196 16838 17226 16890
rect 17226 16838 17252 16890
rect 16956 16836 17012 16838
rect 17036 16836 17092 16838
rect 17116 16836 17172 16838
rect 17196 16836 17252 16838
rect 20956 21786 21012 21788
rect 21036 21786 21092 21788
rect 21116 21786 21172 21788
rect 21196 21786 21252 21788
rect 20956 21734 20982 21786
rect 20982 21734 21012 21786
rect 21036 21734 21046 21786
rect 21046 21734 21092 21786
rect 21116 21734 21162 21786
rect 21162 21734 21172 21786
rect 21196 21734 21226 21786
rect 21226 21734 21252 21786
rect 20956 21732 21012 21734
rect 21036 21732 21092 21734
rect 21116 21732 21172 21734
rect 21196 21732 21252 21734
rect 20956 20698 21012 20700
rect 21036 20698 21092 20700
rect 21116 20698 21172 20700
rect 21196 20698 21252 20700
rect 20956 20646 20982 20698
rect 20982 20646 21012 20698
rect 21036 20646 21046 20698
rect 21046 20646 21092 20698
rect 21116 20646 21162 20698
rect 21162 20646 21172 20698
rect 21196 20646 21226 20698
rect 21226 20646 21252 20698
rect 20956 20644 21012 20646
rect 21036 20644 21092 20646
rect 21116 20644 21172 20646
rect 21196 20644 21252 20646
rect 20956 19610 21012 19612
rect 21036 19610 21092 19612
rect 21116 19610 21172 19612
rect 21196 19610 21252 19612
rect 20956 19558 20982 19610
rect 20982 19558 21012 19610
rect 21036 19558 21046 19610
rect 21046 19558 21092 19610
rect 21116 19558 21162 19610
rect 21162 19558 21172 19610
rect 21196 19558 21226 19610
rect 21226 19558 21252 19610
rect 20956 19556 21012 19558
rect 21036 19556 21092 19558
rect 21116 19556 21172 19558
rect 21196 19556 21252 19558
rect 20956 18522 21012 18524
rect 21036 18522 21092 18524
rect 21116 18522 21172 18524
rect 21196 18522 21252 18524
rect 20956 18470 20982 18522
rect 20982 18470 21012 18522
rect 21036 18470 21046 18522
rect 21046 18470 21092 18522
rect 21116 18470 21162 18522
rect 21162 18470 21172 18522
rect 21196 18470 21226 18522
rect 21226 18470 21252 18522
rect 20956 18468 21012 18470
rect 21036 18468 21092 18470
rect 21116 18468 21172 18470
rect 21196 18468 21252 18470
rect 20956 17434 21012 17436
rect 21036 17434 21092 17436
rect 21116 17434 21172 17436
rect 21196 17434 21252 17436
rect 20956 17382 20982 17434
rect 20982 17382 21012 17434
rect 21036 17382 21046 17434
rect 21046 17382 21092 17434
rect 21116 17382 21162 17434
rect 21162 17382 21172 17434
rect 21196 17382 21226 17434
rect 21226 17382 21252 17434
rect 20956 17380 21012 17382
rect 21036 17380 21092 17382
rect 21116 17380 21172 17382
rect 21196 17380 21252 17382
rect 17682 16632 17738 16688
rect 12956 16346 13012 16348
rect 13036 16346 13092 16348
rect 13116 16346 13172 16348
rect 13196 16346 13252 16348
rect 12956 16294 12982 16346
rect 12982 16294 13012 16346
rect 13036 16294 13046 16346
rect 13046 16294 13092 16346
rect 13116 16294 13162 16346
rect 13162 16294 13172 16346
rect 13196 16294 13226 16346
rect 13226 16294 13252 16346
rect 12956 16292 13012 16294
rect 13036 16292 13092 16294
rect 13116 16292 13172 16294
rect 13196 16292 13252 16294
rect 20956 16346 21012 16348
rect 21036 16346 21092 16348
rect 21116 16346 21172 16348
rect 21196 16346 21252 16348
rect 20956 16294 20982 16346
rect 20982 16294 21012 16346
rect 21036 16294 21046 16346
rect 21046 16294 21092 16346
rect 21116 16294 21162 16346
rect 21162 16294 21172 16346
rect 21196 16294 21226 16346
rect 21226 16294 21252 16346
rect 20956 16292 21012 16294
rect 21036 16292 21092 16294
rect 21116 16292 21172 16294
rect 21196 16292 21252 16294
rect 8956 15802 9012 15804
rect 9036 15802 9092 15804
rect 9116 15802 9172 15804
rect 9196 15802 9252 15804
rect 8956 15750 8982 15802
rect 8982 15750 9012 15802
rect 9036 15750 9046 15802
rect 9046 15750 9092 15802
rect 9116 15750 9162 15802
rect 9162 15750 9172 15802
rect 9196 15750 9226 15802
rect 9226 15750 9252 15802
rect 8956 15748 9012 15750
rect 9036 15748 9092 15750
rect 9116 15748 9172 15750
rect 9196 15748 9252 15750
rect 16956 15802 17012 15804
rect 17036 15802 17092 15804
rect 17116 15802 17172 15804
rect 17196 15802 17252 15804
rect 16956 15750 16982 15802
rect 16982 15750 17012 15802
rect 17036 15750 17046 15802
rect 17046 15750 17092 15802
rect 17116 15750 17162 15802
rect 17162 15750 17172 15802
rect 17196 15750 17226 15802
rect 17226 15750 17252 15802
rect 16956 15748 17012 15750
rect 17036 15748 17092 15750
rect 17116 15748 17172 15750
rect 17196 15748 17252 15750
rect 7654 15544 7710 15600
rect 22006 15544 22062 15600
rect 12956 15258 13012 15260
rect 13036 15258 13092 15260
rect 13116 15258 13172 15260
rect 13196 15258 13252 15260
rect 12956 15206 12982 15258
rect 12982 15206 13012 15258
rect 13036 15206 13046 15258
rect 13046 15206 13092 15258
rect 13116 15206 13162 15258
rect 13162 15206 13172 15258
rect 13196 15206 13226 15258
rect 13226 15206 13252 15258
rect 12956 15204 13012 15206
rect 13036 15204 13092 15206
rect 13116 15204 13172 15206
rect 13196 15204 13252 15206
rect 20956 15258 21012 15260
rect 21036 15258 21092 15260
rect 21116 15258 21172 15260
rect 21196 15258 21252 15260
rect 20956 15206 20982 15258
rect 20982 15206 21012 15258
rect 21036 15206 21046 15258
rect 21046 15206 21092 15258
rect 21116 15206 21162 15258
rect 21162 15206 21172 15258
rect 21196 15206 21226 15258
rect 21226 15206 21252 15258
rect 20956 15204 21012 15206
rect 21036 15204 21092 15206
rect 21116 15204 21172 15206
rect 21196 15204 21252 15206
rect 8956 14714 9012 14716
rect 9036 14714 9092 14716
rect 9116 14714 9172 14716
rect 9196 14714 9252 14716
rect 8956 14662 8982 14714
rect 8982 14662 9012 14714
rect 9036 14662 9046 14714
rect 9046 14662 9092 14714
rect 9116 14662 9162 14714
rect 9162 14662 9172 14714
rect 9196 14662 9226 14714
rect 9226 14662 9252 14714
rect 8956 14660 9012 14662
rect 9036 14660 9092 14662
rect 9116 14660 9172 14662
rect 9196 14660 9252 14662
rect 16956 14714 17012 14716
rect 17036 14714 17092 14716
rect 17116 14714 17172 14716
rect 17196 14714 17252 14716
rect 16956 14662 16982 14714
rect 16982 14662 17012 14714
rect 17036 14662 17046 14714
rect 17046 14662 17092 14714
rect 17116 14662 17162 14714
rect 17162 14662 17172 14714
rect 17196 14662 17226 14714
rect 17226 14662 17252 14714
rect 16956 14660 17012 14662
rect 17036 14660 17092 14662
rect 17116 14660 17172 14662
rect 17196 14660 17252 14662
rect 12956 14170 13012 14172
rect 13036 14170 13092 14172
rect 13116 14170 13172 14172
rect 13196 14170 13252 14172
rect 12956 14118 12982 14170
rect 12982 14118 13012 14170
rect 13036 14118 13046 14170
rect 13046 14118 13092 14170
rect 13116 14118 13162 14170
rect 13162 14118 13172 14170
rect 13196 14118 13226 14170
rect 13226 14118 13252 14170
rect 12956 14116 13012 14118
rect 13036 14116 13092 14118
rect 13116 14116 13172 14118
rect 13196 14116 13252 14118
rect 20956 14170 21012 14172
rect 21036 14170 21092 14172
rect 21116 14170 21172 14172
rect 21196 14170 21252 14172
rect 20956 14118 20982 14170
rect 20982 14118 21012 14170
rect 21036 14118 21046 14170
rect 21046 14118 21092 14170
rect 21116 14118 21162 14170
rect 21162 14118 21172 14170
rect 21196 14118 21226 14170
rect 21226 14118 21252 14170
rect 20956 14116 21012 14118
rect 21036 14116 21092 14118
rect 21116 14116 21172 14118
rect 21196 14116 21252 14118
rect 8956 13626 9012 13628
rect 9036 13626 9092 13628
rect 9116 13626 9172 13628
rect 9196 13626 9252 13628
rect 8956 13574 8982 13626
rect 8982 13574 9012 13626
rect 9036 13574 9046 13626
rect 9046 13574 9092 13626
rect 9116 13574 9162 13626
rect 9162 13574 9172 13626
rect 9196 13574 9226 13626
rect 9226 13574 9252 13626
rect 8956 13572 9012 13574
rect 9036 13572 9092 13574
rect 9116 13572 9172 13574
rect 9196 13572 9252 13574
rect 16956 13626 17012 13628
rect 17036 13626 17092 13628
rect 17116 13626 17172 13628
rect 17196 13626 17252 13628
rect 16956 13574 16982 13626
rect 16982 13574 17012 13626
rect 17036 13574 17046 13626
rect 17046 13574 17092 13626
rect 17116 13574 17162 13626
rect 17162 13574 17172 13626
rect 17196 13574 17226 13626
rect 17226 13574 17252 13626
rect 16956 13572 17012 13574
rect 17036 13572 17092 13574
rect 17116 13572 17172 13574
rect 17196 13572 17252 13574
rect 12956 13082 13012 13084
rect 13036 13082 13092 13084
rect 13116 13082 13172 13084
rect 13196 13082 13252 13084
rect 12956 13030 12982 13082
rect 12982 13030 13012 13082
rect 13036 13030 13046 13082
rect 13046 13030 13092 13082
rect 13116 13030 13162 13082
rect 13162 13030 13172 13082
rect 13196 13030 13226 13082
rect 13226 13030 13252 13082
rect 12956 13028 13012 13030
rect 13036 13028 13092 13030
rect 13116 13028 13172 13030
rect 13196 13028 13252 13030
rect 20956 13082 21012 13084
rect 21036 13082 21092 13084
rect 21116 13082 21172 13084
rect 21196 13082 21252 13084
rect 20956 13030 20982 13082
rect 20982 13030 21012 13082
rect 21036 13030 21046 13082
rect 21046 13030 21092 13082
rect 21116 13030 21162 13082
rect 21162 13030 21172 13082
rect 21196 13030 21226 13082
rect 21226 13030 21252 13082
rect 20956 13028 21012 13030
rect 21036 13028 21092 13030
rect 21116 13028 21172 13030
rect 21196 13028 21252 13030
rect 8956 12538 9012 12540
rect 9036 12538 9092 12540
rect 9116 12538 9172 12540
rect 9196 12538 9252 12540
rect 8956 12486 8982 12538
rect 8982 12486 9012 12538
rect 9036 12486 9046 12538
rect 9046 12486 9092 12538
rect 9116 12486 9162 12538
rect 9162 12486 9172 12538
rect 9196 12486 9226 12538
rect 9226 12486 9252 12538
rect 8956 12484 9012 12486
rect 9036 12484 9092 12486
rect 9116 12484 9172 12486
rect 9196 12484 9252 12486
rect 16956 12538 17012 12540
rect 17036 12538 17092 12540
rect 17116 12538 17172 12540
rect 17196 12538 17252 12540
rect 16956 12486 16982 12538
rect 16982 12486 17012 12538
rect 17036 12486 17046 12538
rect 17046 12486 17092 12538
rect 17116 12486 17162 12538
rect 17162 12486 17172 12538
rect 17196 12486 17226 12538
rect 17226 12486 17252 12538
rect 16956 12484 17012 12486
rect 17036 12484 17092 12486
rect 17116 12484 17172 12486
rect 17196 12484 17252 12486
rect 7470 10648 7526 10704
rect 12956 11994 13012 11996
rect 13036 11994 13092 11996
rect 13116 11994 13172 11996
rect 13196 11994 13252 11996
rect 12956 11942 12982 11994
rect 12982 11942 13012 11994
rect 13036 11942 13046 11994
rect 13046 11942 13092 11994
rect 13116 11942 13162 11994
rect 13162 11942 13172 11994
rect 13196 11942 13226 11994
rect 13226 11942 13252 11994
rect 12956 11940 13012 11942
rect 13036 11940 13092 11942
rect 13116 11940 13172 11942
rect 13196 11940 13252 11942
rect 20956 11994 21012 11996
rect 21036 11994 21092 11996
rect 21116 11994 21172 11996
rect 21196 11994 21252 11996
rect 20956 11942 20982 11994
rect 20982 11942 21012 11994
rect 21036 11942 21046 11994
rect 21046 11942 21092 11994
rect 21116 11942 21162 11994
rect 21162 11942 21172 11994
rect 21196 11942 21226 11994
rect 21226 11942 21252 11994
rect 20956 11940 21012 11942
rect 21036 11940 21092 11942
rect 21116 11940 21172 11942
rect 21196 11940 21252 11942
rect 8956 11450 9012 11452
rect 9036 11450 9092 11452
rect 9116 11450 9172 11452
rect 9196 11450 9252 11452
rect 8956 11398 8982 11450
rect 8982 11398 9012 11450
rect 9036 11398 9046 11450
rect 9046 11398 9092 11450
rect 9116 11398 9162 11450
rect 9162 11398 9172 11450
rect 9196 11398 9226 11450
rect 9226 11398 9252 11450
rect 8956 11396 9012 11398
rect 9036 11396 9092 11398
rect 9116 11396 9172 11398
rect 9196 11396 9252 11398
rect 16956 11450 17012 11452
rect 17036 11450 17092 11452
rect 17116 11450 17172 11452
rect 17196 11450 17252 11452
rect 16956 11398 16982 11450
rect 16982 11398 17012 11450
rect 17036 11398 17046 11450
rect 17046 11398 17092 11450
rect 17116 11398 17162 11450
rect 17162 11398 17172 11450
rect 17196 11398 17226 11450
rect 17226 11398 17252 11450
rect 16956 11396 17012 11398
rect 17036 11396 17092 11398
rect 17116 11396 17172 11398
rect 17196 11396 17252 11398
rect 12956 10906 13012 10908
rect 13036 10906 13092 10908
rect 13116 10906 13172 10908
rect 13196 10906 13252 10908
rect 12956 10854 12982 10906
rect 12982 10854 13012 10906
rect 13036 10854 13046 10906
rect 13046 10854 13092 10906
rect 13116 10854 13162 10906
rect 13162 10854 13172 10906
rect 13196 10854 13226 10906
rect 13226 10854 13252 10906
rect 12956 10852 13012 10854
rect 13036 10852 13092 10854
rect 13116 10852 13172 10854
rect 13196 10852 13252 10854
rect 20956 10906 21012 10908
rect 21036 10906 21092 10908
rect 21116 10906 21172 10908
rect 21196 10906 21252 10908
rect 20956 10854 20982 10906
rect 20982 10854 21012 10906
rect 21036 10854 21046 10906
rect 21046 10854 21092 10906
rect 21116 10854 21162 10906
rect 21162 10854 21172 10906
rect 21196 10854 21226 10906
rect 21226 10854 21252 10906
rect 20956 10852 21012 10854
rect 21036 10852 21092 10854
rect 21116 10852 21172 10854
rect 21196 10852 21252 10854
rect 8956 10362 9012 10364
rect 9036 10362 9092 10364
rect 9116 10362 9172 10364
rect 9196 10362 9252 10364
rect 8956 10310 8982 10362
rect 8982 10310 9012 10362
rect 9036 10310 9046 10362
rect 9046 10310 9092 10362
rect 9116 10310 9162 10362
rect 9162 10310 9172 10362
rect 9196 10310 9226 10362
rect 9226 10310 9252 10362
rect 8956 10308 9012 10310
rect 9036 10308 9092 10310
rect 9116 10308 9172 10310
rect 9196 10308 9252 10310
rect 16956 10362 17012 10364
rect 17036 10362 17092 10364
rect 17116 10362 17172 10364
rect 17196 10362 17252 10364
rect 16956 10310 16982 10362
rect 16982 10310 17012 10362
rect 17036 10310 17046 10362
rect 17046 10310 17092 10362
rect 17116 10310 17162 10362
rect 17162 10310 17172 10362
rect 17196 10310 17226 10362
rect 17226 10310 17252 10362
rect 16956 10308 17012 10310
rect 17036 10308 17092 10310
rect 17116 10308 17172 10310
rect 17196 10308 17252 10310
rect 12956 9818 13012 9820
rect 13036 9818 13092 9820
rect 13116 9818 13172 9820
rect 13196 9818 13252 9820
rect 12956 9766 12982 9818
rect 12982 9766 13012 9818
rect 13036 9766 13046 9818
rect 13046 9766 13092 9818
rect 13116 9766 13162 9818
rect 13162 9766 13172 9818
rect 13196 9766 13226 9818
rect 13226 9766 13252 9818
rect 12956 9764 13012 9766
rect 13036 9764 13092 9766
rect 13116 9764 13172 9766
rect 13196 9764 13252 9766
rect 20956 9818 21012 9820
rect 21036 9818 21092 9820
rect 21116 9818 21172 9820
rect 21196 9818 21252 9820
rect 20956 9766 20982 9818
rect 20982 9766 21012 9818
rect 21036 9766 21046 9818
rect 21046 9766 21092 9818
rect 21116 9766 21162 9818
rect 21162 9766 21172 9818
rect 21196 9766 21226 9818
rect 21226 9766 21252 9818
rect 20956 9764 21012 9766
rect 21036 9764 21092 9766
rect 21116 9764 21172 9766
rect 21196 9764 21252 9766
rect 8956 9274 9012 9276
rect 9036 9274 9092 9276
rect 9116 9274 9172 9276
rect 9196 9274 9252 9276
rect 8956 9222 8982 9274
rect 8982 9222 9012 9274
rect 9036 9222 9046 9274
rect 9046 9222 9092 9274
rect 9116 9222 9162 9274
rect 9162 9222 9172 9274
rect 9196 9222 9226 9274
rect 9226 9222 9252 9274
rect 8956 9220 9012 9222
rect 9036 9220 9092 9222
rect 9116 9220 9172 9222
rect 9196 9220 9252 9222
rect 16956 9274 17012 9276
rect 17036 9274 17092 9276
rect 17116 9274 17172 9276
rect 17196 9274 17252 9276
rect 16956 9222 16982 9274
rect 16982 9222 17012 9274
rect 17036 9222 17046 9274
rect 17046 9222 17092 9274
rect 17116 9222 17162 9274
rect 17162 9222 17172 9274
rect 17196 9222 17226 9274
rect 17226 9222 17252 9274
rect 16956 9220 17012 9222
rect 17036 9220 17092 9222
rect 17116 9220 17172 9222
rect 17196 9220 17252 9222
rect 12956 8730 13012 8732
rect 13036 8730 13092 8732
rect 13116 8730 13172 8732
rect 13196 8730 13252 8732
rect 12956 8678 12982 8730
rect 12982 8678 13012 8730
rect 13036 8678 13046 8730
rect 13046 8678 13092 8730
rect 13116 8678 13162 8730
rect 13162 8678 13172 8730
rect 13196 8678 13226 8730
rect 13226 8678 13252 8730
rect 12956 8676 13012 8678
rect 13036 8676 13092 8678
rect 13116 8676 13172 8678
rect 13196 8676 13252 8678
rect 20956 8730 21012 8732
rect 21036 8730 21092 8732
rect 21116 8730 21172 8732
rect 21196 8730 21252 8732
rect 20956 8678 20982 8730
rect 20982 8678 21012 8730
rect 21036 8678 21046 8730
rect 21046 8678 21092 8730
rect 21116 8678 21162 8730
rect 21162 8678 21172 8730
rect 21196 8678 21226 8730
rect 21226 8678 21252 8730
rect 20956 8676 21012 8678
rect 21036 8676 21092 8678
rect 21116 8676 21172 8678
rect 21196 8676 21252 8678
rect 8956 8186 9012 8188
rect 9036 8186 9092 8188
rect 9116 8186 9172 8188
rect 9196 8186 9252 8188
rect 8956 8134 8982 8186
rect 8982 8134 9012 8186
rect 9036 8134 9046 8186
rect 9046 8134 9092 8186
rect 9116 8134 9162 8186
rect 9162 8134 9172 8186
rect 9196 8134 9226 8186
rect 9226 8134 9252 8186
rect 8956 8132 9012 8134
rect 9036 8132 9092 8134
rect 9116 8132 9172 8134
rect 9196 8132 9252 8134
rect 16956 8186 17012 8188
rect 17036 8186 17092 8188
rect 17116 8186 17172 8188
rect 17196 8186 17252 8188
rect 16956 8134 16982 8186
rect 16982 8134 17012 8186
rect 17036 8134 17046 8186
rect 17046 8134 17092 8186
rect 17116 8134 17162 8186
rect 17162 8134 17172 8186
rect 17196 8134 17226 8186
rect 17226 8134 17252 8186
rect 16956 8132 17012 8134
rect 17036 8132 17092 8134
rect 17116 8132 17172 8134
rect 17196 8132 17252 8134
rect 12956 7642 13012 7644
rect 13036 7642 13092 7644
rect 13116 7642 13172 7644
rect 13196 7642 13252 7644
rect 12956 7590 12982 7642
rect 12982 7590 13012 7642
rect 13036 7590 13046 7642
rect 13046 7590 13092 7642
rect 13116 7590 13162 7642
rect 13162 7590 13172 7642
rect 13196 7590 13226 7642
rect 13226 7590 13252 7642
rect 12956 7588 13012 7590
rect 13036 7588 13092 7590
rect 13116 7588 13172 7590
rect 13196 7588 13252 7590
rect 20956 7642 21012 7644
rect 21036 7642 21092 7644
rect 21116 7642 21172 7644
rect 21196 7642 21252 7644
rect 20956 7590 20982 7642
rect 20982 7590 21012 7642
rect 21036 7590 21046 7642
rect 21046 7590 21092 7642
rect 21116 7590 21162 7642
rect 21162 7590 21172 7642
rect 21196 7590 21226 7642
rect 21226 7590 21252 7642
rect 20956 7588 21012 7590
rect 21036 7588 21092 7590
rect 21116 7588 21172 7590
rect 21196 7588 21252 7590
rect 8956 7098 9012 7100
rect 9036 7098 9092 7100
rect 9116 7098 9172 7100
rect 9196 7098 9252 7100
rect 8956 7046 8982 7098
rect 8982 7046 9012 7098
rect 9036 7046 9046 7098
rect 9046 7046 9092 7098
rect 9116 7046 9162 7098
rect 9162 7046 9172 7098
rect 9196 7046 9226 7098
rect 9226 7046 9252 7098
rect 8956 7044 9012 7046
rect 9036 7044 9092 7046
rect 9116 7044 9172 7046
rect 9196 7044 9252 7046
rect 8956 6010 9012 6012
rect 9036 6010 9092 6012
rect 9116 6010 9172 6012
rect 9196 6010 9252 6012
rect 8956 5958 8982 6010
rect 8982 5958 9012 6010
rect 9036 5958 9046 6010
rect 9046 5958 9092 6010
rect 9116 5958 9162 6010
rect 9162 5958 9172 6010
rect 9196 5958 9226 6010
rect 9226 5958 9252 6010
rect 8956 5956 9012 5958
rect 9036 5956 9092 5958
rect 9116 5956 9172 5958
rect 9196 5956 9252 5958
rect 8956 4922 9012 4924
rect 9036 4922 9092 4924
rect 9116 4922 9172 4924
rect 9196 4922 9252 4924
rect 8956 4870 8982 4922
rect 8982 4870 9012 4922
rect 9036 4870 9046 4922
rect 9046 4870 9092 4922
rect 9116 4870 9162 4922
rect 9162 4870 9172 4922
rect 9196 4870 9226 4922
rect 9226 4870 9252 4922
rect 8956 4868 9012 4870
rect 9036 4868 9092 4870
rect 9116 4868 9172 4870
rect 9196 4868 9252 4870
rect 8956 3834 9012 3836
rect 9036 3834 9092 3836
rect 9116 3834 9172 3836
rect 9196 3834 9252 3836
rect 8956 3782 8982 3834
rect 8982 3782 9012 3834
rect 9036 3782 9046 3834
rect 9046 3782 9092 3834
rect 9116 3782 9162 3834
rect 9162 3782 9172 3834
rect 9196 3782 9226 3834
rect 9226 3782 9252 3834
rect 8956 3780 9012 3782
rect 9036 3780 9092 3782
rect 9116 3780 9172 3782
rect 9196 3780 9252 3782
rect 8956 2746 9012 2748
rect 9036 2746 9092 2748
rect 9116 2746 9172 2748
rect 9196 2746 9252 2748
rect 8956 2694 8982 2746
rect 8982 2694 9012 2746
rect 9036 2694 9046 2746
rect 9046 2694 9092 2746
rect 9116 2694 9162 2746
rect 9162 2694 9172 2746
rect 9196 2694 9226 2746
rect 9226 2694 9252 2746
rect 8956 2692 9012 2694
rect 9036 2692 9092 2694
rect 9116 2692 9172 2694
rect 9196 2692 9252 2694
rect 4956 2202 5012 2204
rect 5036 2202 5092 2204
rect 5116 2202 5172 2204
rect 5196 2202 5252 2204
rect 4956 2150 4982 2202
rect 4982 2150 5012 2202
rect 5036 2150 5046 2202
rect 5046 2150 5092 2202
rect 5116 2150 5162 2202
rect 5162 2150 5172 2202
rect 5196 2150 5226 2202
rect 5226 2150 5252 2202
rect 4956 2148 5012 2150
rect 5036 2148 5092 2150
rect 5116 2148 5172 2150
rect 5196 2148 5252 2150
rect 3422 584 3478 640
rect 16956 7098 17012 7100
rect 17036 7098 17092 7100
rect 17116 7098 17172 7100
rect 17196 7098 17252 7100
rect 16956 7046 16982 7098
rect 16982 7046 17012 7098
rect 17036 7046 17046 7098
rect 17046 7046 17092 7098
rect 17116 7046 17162 7098
rect 17162 7046 17172 7098
rect 17196 7046 17226 7098
rect 17226 7046 17252 7098
rect 16956 7044 17012 7046
rect 17036 7044 17092 7046
rect 17116 7044 17172 7046
rect 17196 7044 17252 7046
rect 12956 6554 13012 6556
rect 13036 6554 13092 6556
rect 13116 6554 13172 6556
rect 13196 6554 13252 6556
rect 12956 6502 12982 6554
rect 12982 6502 13012 6554
rect 13036 6502 13046 6554
rect 13046 6502 13092 6554
rect 13116 6502 13162 6554
rect 13162 6502 13172 6554
rect 13196 6502 13226 6554
rect 13226 6502 13252 6554
rect 12956 6500 13012 6502
rect 13036 6500 13092 6502
rect 13116 6500 13172 6502
rect 13196 6500 13252 6502
rect 20956 6554 21012 6556
rect 21036 6554 21092 6556
rect 21116 6554 21172 6556
rect 21196 6554 21252 6556
rect 20956 6502 20982 6554
rect 20982 6502 21012 6554
rect 21036 6502 21046 6554
rect 21046 6502 21092 6554
rect 21116 6502 21162 6554
rect 21162 6502 21172 6554
rect 21196 6502 21226 6554
rect 21226 6502 21252 6554
rect 20956 6500 21012 6502
rect 21036 6500 21092 6502
rect 21116 6500 21172 6502
rect 21196 6500 21252 6502
rect 16956 6010 17012 6012
rect 17036 6010 17092 6012
rect 17116 6010 17172 6012
rect 17196 6010 17252 6012
rect 16956 5958 16982 6010
rect 16982 5958 17012 6010
rect 17036 5958 17046 6010
rect 17046 5958 17092 6010
rect 17116 5958 17162 6010
rect 17162 5958 17172 6010
rect 17196 5958 17226 6010
rect 17226 5958 17252 6010
rect 16956 5956 17012 5958
rect 17036 5956 17092 5958
rect 17116 5956 17172 5958
rect 17196 5956 17252 5958
rect 12956 5466 13012 5468
rect 13036 5466 13092 5468
rect 13116 5466 13172 5468
rect 13196 5466 13252 5468
rect 12956 5414 12982 5466
rect 12982 5414 13012 5466
rect 13036 5414 13046 5466
rect 13046 5414 13092 5466
rect 13116 5414 13162 5466
rect 13162 5414 13172 5466
rect 13196 5414 13226 5466
rect 13226 5414 13252 5466
rect 12956 5412 13012 5414
rect 13036 5412 13092 5414
rect 13116 5412 13172 5414
rect 13196 5412 13252 5414
rect 20956 5466 21012 5468
rect 21036 5466 21092 5468
rect 21116 5466 21172 5468
rect 21196 5466 21252 5468
rect 20956 5414 20982 5466
rect 20982 5414 21012 5466
rect 21036 5414 21046 5466
rect 21046 5414 21092 5466
rect 21116 5414 21162 5466
rect 21162 5414 21172 5466
rect 21196 5414 21226 5466
rect 21226 5414 21252 5466
rect 20956 5412 21012 5414
rect 21036 5412 21092 5414
rect 21116 5412 21172 5414
rect 21196 5412 21252 5414
rect 16956 4922 17012 4924
rect 17036 4922 17092 4924
rect 17116 4922 17172 4924
rect 17196 4922 17252 4924
rect 16956 4870 16982 4922
rect 16982 4870 17012 4922
rect 17036 4870 17046 4922
rect 17046 4870 17092 4922
rect 17116 4870 17162 4922
rect 17162 4870 17172 4922
rect 17196 4870 17226 4922
rect 17226 4870 17252 4922
rect 16956 4868 17012 4870
rect 17036 4868 17092 4870
rect 17116 4868 17172 4870
rect 17196 4868 17252 4870
rect 12956 4378 13012 4380
rect 13036 4378 13092 4380
rect 13116 4378 13172 4380
rect 13196 4378 13252 4380
rect 12956 4326 12982 4378
rect 12982 4326 13012 4378
rect 13036 4326 13046 4378
rect 13046 4326 13092 4378
rect 13116 4326 13162 4378
rect 13162 4326 13172 4378
rect 13196 4326 13226 4378
rect 13226 4326 13252 4378
rect 12956 4324 13012 4326
rect 13036 4324 13092 4326
rect 13116 4324 13172 4326
rect 13196 4324 13252 4326
rect 20956 4378 21012 4380
rect 21036 4378 21092 4380
rect 21116 4378 21172 4380
rect 21196 4378 21252 4380
rect 20956 4326 20982 4378
rect 20982 4326 21012 4378
rect 21036 4326 21046 4378
rect 21046 4326 21092 4378
rect 21116 4326 21162 4378
rect 21162 4326 21172 4378
rect 21196 4326 21226 4378
rect 21226 4326 21252 4378
rect 20956 4324 21012 4326
rect 21036 4324 21092 4326
rect 21116 4324 21172 4326
rect 21196 4324 21252 4326
rect 16956 3834 17012 3836
rect 17036 3834 17092 3836
rect 17116 3834 17172 3836
rect 17196 3834 17252 3836
rect 16956 3782 16982 3834
rect 16982 3782 17012 3834
rect 17036 3782 17046 3834
rect 17046 3782 17092 3834
rect 17116 3782 17162 3834
rect 17162 3782 17172 3834
rect 17196 3782 17226 3834
rect 17226 3782 17252 3834
rect 16956 3780 17012 3782
rect 17036 3780 17092 3782
rect 17116 3780 17172 3782
rect 17196 3780 17252 3782
rect 12956 3290 13012 3292
rect 13036 3290 13092 3292
rect 13116 3290 13172 3292
rect 13196 3290 13252 3292
rect 12956 3238 12982 3290
rect 12982 3238 13012 3290
rect 13036 3238 13046 3290
rect 13046 3238 13092 3290
rect 13116 3238 13162 3290
rect 13162 3238 13172 3290
rect 13196 3238 13226 3290
rect 13226 3238 13252 3290
rect 12956 3236 13012 3238
rect 13036 3236 13092 3238
rect 13116 3236 13172 3238
rect 13196 3236 13252 3238
rect 20956 3290 21012 3292
rect 21036 3290 21092 3292
rect 21116 3290 21172 3292
rect 21196 3290 21252 3292
rect 20956 3238 20982 3290
rect 20982 3238 21012 3290
rect 21036 3238 21046 3290
rect 21046 3238 21092 3290
rect 21116 3238 21162 3290
rect 21162 3238 21172 3290
rect 21196 3238 21226 3290
rect 21226 3238 21252 3290
rect 20956 3236 21012 3238
rect 21036 3236 21092 3238
rect 21116 3236 21172 3238
rect 21196 3236 21252 3238
rect 16956 2746 17012 2748
rect 17036 2746 17092 2748
rect 17116 2746 17172 2748
rect 17196 2746 17252 2748
rect 16956 2694 16982 2746
rect 16982 2694 17012 2746
rect 17036 2694 17046 2746
rect 17046 2694 17092 2746
rect 17116 2694 17162 2746
rect 17162 2694 17172 2746
rect 17196 2694 17226 2746
rect 17226 2694 17252 2746
rect 16956 2692 17012 2694
rect 17036 2692 17092 2694
rect 17116 2692 17172 2694
rect 17196 2692 17252 2694
rect 12956 2202 13012 2204
rect 13036 2202 13092 2204
rect 13116 2202 13172 2204
rect 13196 2202 13252 2204
rect 12956 2150 12982 2202
rect 12982 2150 13012 2202
rect 13036 2150 13046 2202
rect 13046 2150 13092 2202
rect 13116 2150 13162 2202
rect 13162 2150 13172 2202
rect 13196 2150 13226 2202
rect 13226 2150 13252 2202
rect 12956 2148 13012 2150
rect 13036 2148 13092 2150
rect 13116 2148 13172 2150
rect 13196 2148 13252 2150
rect 20956 2202 21012 2204
rect 21036 2202 21092 2204
rect 21116 2202 21172 2204
rect 21196 2202 21252 2204
rect 20956 2150 20982 2202
rect 20982 2150 21012 2202
rect 21036 2150 21046 2202
rect 21046 2150 21092 2202
rect 21116 2150 21162 2202
rect 21162 2150 21172 2202
rect 21196 2150 21226 2202
rect 21226 2150 21252 2202
rect 20956 2148 21012 2150
rect 21036 2148 21092 2150
rect 21116 2148 21172 2150
rect 21196 2148 21252 2150
<< metal3 >>
rect 0 23760 480 23792
rect 0 23704 110 23760
rect 166 23704 480 23760
rect 0 23672 480 23704
rect 0 23352 480 23384
rect 0 23296 18 23352
rect 74 23296 480 23352
rect 0 23264 480 23296
rect 0 22944 480 22976
rect 0 22888 110 22944
rect 166 22888 480 22944
rect 0 22856 480 22888
rect 0 22536 480 22568
rect 0 22480 110 22536
rect 166 22480 480 22536
rect 0 22448 480 22480
rect 0 22132 480 22160
rect 0 22068 60 22132
rect 124 22068 480 22132
rect 0 22040 480 22068
rect 4944 21792 5264 21793
rect 0 21720 480 21752
rect 4944 21728 4952 21792
rect 5016 21728 5032 21792
rect 5096 21728 5112 21792
rect 5176 21728 5192 21792
rect 5256 21728 5264 21792
rect 4944 21727 5264 21728
rect 12944 21792 13264 21793
rect 12944 21728 12952 21792
rect 13016 21728 13032 21792
rect 13096 21728 13112 21792
rect 13176 21728 13192 21792
rect 13256 21728 13264 21792
rect 12944 21727 13264 21728
rect 20944 21792 21264 21793
rect 20944 21728 20952 21792
rect 21016 21728 21032 21792
rect 21096 21728 21112 21792
rect 21176 21728 21192 21792
rect 21256 21728 21264 21792
rect 20944 21727 21264 21728
rect 0 21664 110 21720
rect 166 21664 480 21720
rect 0 21632 480 21664
rect 606 21388 612 21452
rect 676 21450 682 21452
rect 4705 21450 4771 21453
rect 676 21448 4771 21450
rect 676 21392 4710 21448
rect 4766 21392 4771 21448
rect 676 21390 4771 21392
rect 676 21388 682 21390
rect 4705 21387 4771 21390
rect 0 21312 480 21344
rect 0 21256 110 21312
rect 166 21256 480 21312
rect 0 21224 480 21256
rect 8944 21248 9264 21249
rect 8944 21184 8952 21248
rect 9016 21184 9032 21248
rect 9096 21184 9112 21248
rect 9176 21184 9192 21248
rect 9256 21184 9264 21248
rect 8944 21183 9264 21184
rect 16944 21248 17264 21249
rect 16944 21184 16952 21248
rect 17016 21184 17032 21248
rect 17096 21184 17112 21248
rect 17176 21184 17192 21248
rect 17256 21184 17264 21248
rect 16944 21183 17264 21184
rect 0 20904 480 20936
rect 0 20848 386 20904
rect 442 20848 480 20904
rect 0 20816 480 20848
rect 4944 20704 5264 20705
rect 0 20636 480 20664
rect 4944 20640 4952 20704
rect 5016 20640 5032 20704
rect 5096 20640 5112 20704
rect 5176 20640 5192 20704
rect 5256 20640 5264 20704
rect 4944 20639 5264 20640
rect 12944 20704 13264 20705
rect 12944 20640 12952 20704
rect 13016 20640 13032 20704
rect 13096 20640 13112 20704
rect 13176 20640 13192 20704
rect 13256 20640 13264 20704
rect 12944 20639 13264 20640
rect 20944 20704 21264 20705
rect 20944 20640 20952 20704
rect 21016 20640 21032 20704
rect 21096 20640 21112 20704
rect 21176 20640 21192 20704
rect 21256 20640 21264 20704
rect 20944 20639 21264 20640
rect 0 20572 60 20636
rect 124 20572 480 20636
rect 0 20544 480 20572
rect 54 20334 60 20398
rect 124 20396 130 20398
rect 124 20336 674 20396
rect 124 20334 130 20336
rect 0 20228 480 20256
rect 0 20164 60 20228
rect 124 20164 480 20228
rect 614 20226 674 20336
rect 4613 20226 4679 20229
rect 614 20224 4679 20226
rect 614 20168 4618 20224
rect 4674 20168 4679 20224
rect 614 20166 4679 20168
rect 0 20136 480 20164
rect 4613 20163 4679 20166
rect 8944 20160 9264 20161
rect 8944 20096 8952 20160
rect 9016 20096 9032 20160
rect 9096 20096 9112 20160
rect 9176 20096 9192 20160
rect 9256 20096 9264 20160
rect 8944 20095 9264 20096
rect 16944 20160 17264 20161
rect 16944 20096 16952 20160
rect 17016 20096 17032 20160
rect 17096 20096 17112 20160
rect 17176 20096 17192 20160
rect 17256 20096 17264 20160
rect 16944 20095 17264 20096
rect 606 20028 612 20092
rect 676 20090 682 20092
rect 1761 20090 1827 20093
rect 676 20088 1827 20090
rect 676 20032 1766 20088
rect 1822 20032 1827 20088
rect 676 20030 1827 20032
rect 676 20028 682 20030
rect 1761 20027 1827 20030
rect 0 19816 480 19848
rect 0 19760 110 19816
rect 166 19760 480 19816
rect 0 19728 480 19760
rect 4944 19616 5264 19617
rect 4944 19552 4952 19616
rect 5016 19552 5032 19616
rect 5096 19552 5112 19616
rect 5176 19552 5192 19616
rect 5256 19552 5264 19616
rect 4944 19551 5264 19552
rect 12944 19616 13264 19617
rect 12944 19552 12952 19616
rect 13016 19552 13032 19616
rect 13096 19552 13112 19616
rect 13176 19552 13192 19616
rect 13256 19552 13264 19616
rect 12944 19551 13264 19552
rect 20944 19616 21264 19617
rect 20944 19552 20952 19616
rect 21016 19552 21032 19616
rect 21096 19552 21112 19616
rect 21176 19552 21192 19616
rect 21256 19552 21264 19616
rect 20944 19551 21264 19552
rect 0 19350 480 19440
rect 0 19320 674 19350
rect 62 19290 674 19320
rect 614 19274 674 19290
rect 4245 19274 4311 19277
rect 614 19272 4311 19274
rect 614 19216 4250 19272
rect 4306 19216 4311 19272
rect 614 19214 4311 19216
rect 4245 19211 4311 19214
rect 8944 19072 9264 19073
rect 0 19004 480 19032
rect 8944 19008 8952 19072
rect 9016 19008 9032 19072
rect 9096 19008 9112 19072
rect 9176 19008 9192 19072
rect 9256 19008 9264 19072
rect 8944 19007 9264 19008
rect 16944 19072 17264 19073
rect 16944 19008 16952 19072
rect 17016 19008 17032 19072
rect 17096 19008 17112 19072
rect 17176 19008 17192 19072
rect 17256 19008 17264 19072
rect 16944 19007 17264 19008
rect 0 18940 60 19004
rect 124 18940 480 19004
rect 0 18912 480 18940
rect 606 18668 612 18732
rect 676 18730 682 18732
rect 3417 18730 3483 18733
rect 676 18728 3483 18730
rect 676 18672 3422 18728
rect 3478 18672 3483 18728
rect 676 18670 3483 18672
rect 676 18668 682 18670
rect 3417 18667 3483 18670
rect 0 18592 480 18624
rect 0 18536 18 18592
rect 74 18536 480 18592
rect 0 18504 480 18536
rect 4944 18528 5264 18529
rect 4944 18464 4952 18528
rect 5016 18464 5032 18528
rect 5096 18464 5112 18528
rect 5176 18464 5192 18528
rect 5256 18464 5264 18528
rect 4944 18463 5264 18464
rect 12944 18528 13264 18529
rect 12944 18464 12952 18528
rect 13016 18464 13032 18528
rect 13096 18464 13112 18528
rect 13176 18464 13192 18528
rect 13256 18464 13264 18528
rect 12944 18463 13264 18464
rect 20944 18528 21264 18529
rect 20944 18464 20952 18528
rect 21016 18464 21032 18528
rect 21096 18464 21112 18528
rect 21176 18464 21192 18528
rect 21256 18464 21264 18528
rect 20944 18463 21264 18464
rect 0 18184 480 18216
rect 0 18128 110 18184
rect 166 18128 480 18184
rect 0 18096 480 18128
rect 8944 17984 9264 17985
rect 8944 17920 8952 17984
rect 9016 17920 9032 17984
rect 9096 17920 9112 17984
rect 9176 17920 9192 17984
rect 9256 17920 9264 17984
rect 8944 17919 9264 17920
rect 16944 17984 17264 17985
rect 16944 17920 16952 17984
rect 17016 17920 17032 17984
rect 17096 17920 17112 17984
rect 17176 17920 17192 17984
rect 17256 17920 17264 17984
rect 16944 17919 17264 17920
rect 0 17776 480 17808
rect 0 17720 18 17776
rect 74 17720 480 17776
rect 0 17688 480 17720
rect 4944 17440 5264 17441
rect 0 17368 480 17400
rect 4944 17376 4952 17440
rect 5016 17376 5032 17440
rect 5096 17376 5112 17440
rect 5176 17376 5192 17440
rect 5256 17376 5264 17440
rect 4944 17375 5264 17376
rect 12944 17440 13264 17441
rect 12944 17376 12952 17440
rect 13016 17376 13032 17440
rect 13096 17376 13112 17440
rect 13176 17376 13192 17440
rect 13256 17376 13264 17440
rect 12944 17375 13264 17376
rect 20944 17440 21264 17441
rect 20944 17376 20952 17440
rect 21016 17376 21032 17440
rect 21096 17376 21112 17440
rect 21176 17376 21192 17440
rect 21256 17376 21264 17440
rect 20944 17375 21264 17376
rect 0 17312 18 17368
rect 74 17312 480 17368
rect 0 17280 480 17312
rect 0 17096 480 17128
rect 0 17040 18 17096
rect 74 17040 480 17096
rect 0 17008 480 17040
rect 7373 17098 7439 17101
rect 13813 17098 13879 17101
rect 7373 17096 13879 17098
rect 7373 17040 7378 17096
rect 7434 17040 13818 17096
rect 13874 17040 13879 17096
rect 7373 17038 13879 17040
rect 7373 17035 7439 17038
rect 13813 17035 13879 17038
rect 8944 16896 9264 16897
rect 8944 16832 8952 16896
rect 9016 16832 9032 16896
rect 9096 16832 9112 16896
rect 9176 16832 9192 16896
rect 9256 16832 9264 16896
rect 8944 16831 9264 16832
rect 16944 16896 17264 16897
rect 16944 16832 16952 16896
rect 17016 16832 17032 16896
rect 17096 16832 17112 16896
rect 17176 16832 17192 16896
rect 17256 16832 17264 16896
rect 16944 16831 17264 16832
rect 0 16688 480 16720
rect 0 16632 110 16688
rect 166 16632 480 16688
rect 0 16600 480 16632
rect 7741 16690 7807 16693
rect 17677 16690 17743 16693
rect 7741 16688 17743 16690
rect 7741 16632 7746 16688
rect 7802 16632 17682 16688
rect 17738 16632 17743 16688
rect 7741 16630 17743 16632
rect 7741 16627 7807 16630
rect 17677 16627 17743 16630
rect 4944 16352 5264 16353
rect 0 16280 480 16312
rect 4944 16288 4952 16352
rect 5016 16288 5032 16352
rect 5096 16288 5112 16352
rect 5176 16288 5192 16352
rect 5256 16288 5264 16352
rect 4944 16287 5264 16288
rect 12944 16352 13264 16353
rect 12944 16288 12952 16352
rect 13016 16288 13032 16352
rect 13096 16288 13112 16352
rect 13176 16288 13192 16352
rect 13256 16288 13264 16352
rect 12944 16287 13264 16288
rect 20944 16352 21264 16353
rect 20944 16288 20952 16352
rect 21016 16288 21032 16352
rect 21096 16288 21112 16352
rect 21176 16288 21192 16352
rect 21256 16288 21264 16352
rect 20944 16287 21264 16288
rect 0 16224 110 16280
rect 166 16224 480 16280
rect 0 16192 480 16224
rect 606 15948 612 16012
rect 676 16010 682 16012
rect 3233 16010 3299 16013
rect 676 16008 3299 16010
rect 676 15952 3238 16008
rect 3294 15952 3299 16008
rect 676 15950 3299 15952
rect 676 15948 682 15950
rect 3233 15947 3299 15950
rect 0 15872 480 15904
rect 0 15816 18 15872
rect 74 15816 480 15872
rect 0 15784 480 15816
rect 8944 15808 9264 15809
rect 8944 15744 8952 15808
rect 9016 15744 9032 15808
rect 9096 15744 9112 15808
rect 9176 15744 9192 15808
rect 9256 15744 9264 15808
rect 8944 15743 9264 15744
rect 16944 15808 17264 15809
rect 16944 15744 16952 15808
rect 17016 15744 17032 15808
rect 17096 15744 17112 15808
rect 17176 15744 17192 15808
rect 17256 15744 17264 15808
rect 16944 15743 17264 15744
rect 7649 15602 7715 15605
rect 22001 15602 22067 15605
rect 7649 15600 22067 15602
rect 7649 15544 7654 15600
rect 7710 15544 22006 15600
rect 22062 15544 22067 15600
rect 7649 15542 22067 15544
rect 7649 15539 7715 15542
rect 22001 15539 22067 15542
rect 0 15468 480 15496
rect 0 15404 60 15468
rect 124 15404 480 15468
rect 0 15376 480 15404
rect 4944 15264 5264 15265
rect 4944 15200 4952 15264
rect 5016 15200 5032 15264
rect 5096 15200 5112 15264
rect 5176 15200 5192 15264
rect 5256 15200 5264 15264
rect 4944 15199 5264 15200
rect 12944 15264 13264 15265
rect 12944 15200 12952 15264
rect 13016 15200 13032 15264
rect 13096 15200 13112 15264
rect 13176 15200 13192 15264
rect 13256 15200 13264 15264
rect 12944 15199 13264 15200
rect 20944 15264 21264 15265
rect 20944 15200 20952 15264
rect 21016 15200 21032 15264
rect 21096 15200 21112 15264
rect 21176 15200 21192 15264
rect 21256 15200 21264 15264
rect 20944 15199 21264 15200
rect 0 15056 480 15088
rect 0 15000 110 15056
rect 166 15000 480 15056
rect 0 14968 480 15000
rect 4337 14922 4403 14925
rect 7281 14922 7347 14925
rect 4337 14920 7347 14922
rect 4337 14864 4342 14920
rect 4398 14864 7286 14920
rect 7342 14864 7347 14920
rect 4337 14862 7347 14864
rect 4337 14859 4403 14862
rect 7281 14859 7347 14862
rect 8944 14720 9264 14721
rect 0 14652 480 14680
rect 8944 14656 8952 14720
rect 9016 14656 9032 14720
rect 9096 14656 9112 14720
rect 9176 14656 9192 14720
rect 9256 14656 9264 14720
rect 8944 14655 9264 14656
rect 16944 14720 17264 14721
rect 16944 14656 16952 14720
rect 17016 14656 17032 14720
rect 17096 14656 17112 14720
rect 17176 14656 17192 14720
rect 17256 14656 17264 14720
rect 16944 14655 17264 14656
rect 0 14588 60 14652
rect 124 14588 480 14652
rect 0 14560 480 14588
rect 0 14240 480 14272
rect 0 14184 110 14240
rect 166 14184 480 14240
rect 0 14152 480 14184
rect 4944 14176 5264 14177
rect 4944 14112 4952 14176
rect 5016 14112 5032 14176
rect 5096 14112 5112 14176
rect 5176 14112 5192 14176
rect 5256 14112 5264 14176
rect 4944 14111 5264 14112
rect 12944 14176 13264 14177
rect 12944 14112 12952 14176
rect 13016 14112 13032 14176
rect 13096 14112 13112 14176
rect 13176 14112 13192 14176
rect 13256 14112 13264 14176
rect 12944 14111 13264 14112
rect 20944 14176 21264 14177
rect 20944 14112 20952 14176
rect 21016 14112 21032 14176
rect 21096 14112 21112 14176
rect 21176 14112 21192 14176
rect 21256 14112 21264 14176
rect 20944 14111 21264 14112
rect 606 13908 612 13972
rect 676 13970 682 13972
rect 6913 13970 6979 13973
rect 676 13968 6979 13970
rect 676 13912 6918 13968
rect 6974 13912 6979 13968
rect 676 13910 6979 13912
rect 676 13908 682 13910
rect 6913 13907 6979 13910
rect 0 13836 480 13864
rect 0 13772 60 13836
rect 124 13772 480 13836
rect 606 13772 612 13836
rect 676 13834 682 13836
rect 3049 13834 3115 13837
rect 676 13832 3115 13834
rect 676 13776 3054 13832
rect 3110 13776 3115 13832
rect 676 13774 3115 13776
rect 676 13772 682 13774
rect 0 13744 480 13772
rect 3049 13771 3115 13774
rect 4429 13698 4495 13701
rect 7281 13698 7347 13701
rect 4429 13696 7347 13698
rect 4429 13640 4434 13696
rect 4490 13640 7286 13696
rect 7342 13640 7347 13696
rect 4429 13638 7347 13640
rect 4429 13635 4495 13638
rect 7281 13635 7347 13638
rect 8944 13632 9264 13633
rect 0 13560 480 13592
rect 8944 13568 8952 13632
rect 9016 13568 9032 13632
rect 9096 13568 9112 13632
rect 9176 13568 9192 13632
rect 9256 13568 9264 13632
rect 8944 13567 9264 13568
rect 16944 13632 17264 13633
rect 16944 13568 16952 13632
rect 17016 13568 17032 13632
rect 17096 13568 17112 13632
rect 17176 13568 17192 13632
rect 17256 13568 17264 13632
rect 16944 13567 17264 13568
rect 0 13504 110 13560
rect 166 13504 480 13560
rect 0 13472 480 13504
rect 0 13152 480 13184
rect 0 13096 18 13152
rect 74 13096 480 13152
rect 0 13064 480 13096
rect 4944 13088 5264 13089
rect 4944 13024 4952 13088
rect 5016 13024 5032 13088
rect 5096 13024 5112 13088
rect 5176 13024 5192 13088
rect 5256 13024 5264 13088
rect 4944 13023 5264 13024
rect 12944 13088 13264 13089
rect 12944 13024 12952 13088
rect 13016 13024 13032 13088
rect 13096 13024 13112 13088
rect 13176 13024 13192 13088
rect 13256 13024 13264 13088
rect 12944 13023 13264 13024
rect 20944 13088 21264 13089
rect 20944 13024 20952 13088
rect 21016 13024 21032 13088
rect 21096 13024 21112 13088
rect 21176 13024 21192 13088
rect 21256 13024 21264 13088
rect 20944 13023 21264 13024
rect 0 12744 480 12776
rect 0 12688 110 12744
rect 166 12688 480 12744
rect 0 12656 480 12688
rect 8944 12544 9264 12545
rect 8944 12480 8952 12544
rect 9016 12480 9032 12544
rect 9096 12480 9112 12544
rect 9176 12480 9192 12544
rect 9256 12480 9264 12544
rect 8944 12479 9264 12480
rect 16944 12544 17264 12545
rect 16944 12480 16952 12544
rect 17016 12480 17032 12544
rect 17096 12480 17112 12544
rect 17176 12480 17192 12544
rect 17256 12480 17264 12544
rect 16944 12479 17264 12480
rect 0 12336 480 12368
rect 0 12280 18 12336
rect 74 12280 480 12336
rect 0 12248 480 12280
rect 4944 12000 5264 12001
rect 0 11928 480 11960
rect 4944 11936 4952 12000
rect 5016 11936 5032 12000
rect 5096 11936 5112 12000
rect 5176 11936 5192 12000
rect 5256 11936 5264 12000
rect 4944 11935 5264 11936
rect 12944 12000 13264 12001
rect 12944 11936 12952 12000
rect 13016 11936 13032 12000
rect 13096 11936 13112 12000
rect 13176 11936 13192 12000
rect 13256 11936 13264 12000
rect 12944 11935 13264 11936
rect 20944 12000 21264 12001
rect 20944 11936 20952 12000
rect 21016 11936 21032 12000
rect 21096 11936 21112 12000
rect 21176 11936 21192 12000
rect 21256 11936 21264 12000
rect 20944 11935 21264 11936
rect 0 11872 110 11928
rect 166 11872 480 11928
rect 0 11840 480 11872
rect 0 11520 480 11552
rect 0 11464 18 11520
rect 74 11464 480 11520
rect 0 11432 480 11464
rect 8944 11456 9264 11457
rect 8944 11392 8952 11456
rect 9016 11392 9032 11456
rect 9096 11392 9112 11456
rect 9176 11392 9192 11456
rect 9256 11392 9264 11456
rect 8944 11391 9264 11392
rect 16944 11456 17264 11457
rect 16944 11392 16952 11456
rect 17016 11392 17032 11456
rect 17096 11392 17112 11456
rect 17176 11392 17192 11456
rect 17256 11392 17264 11456
rect 16944 11391 17264 11392
rect 0 11112 480 11144
rect 0 11056 110 11112
rect 166 11056 480 11112
rect 0 11024 480 11056
rect 4944 10912 5264 10913
rect 4944 10848 4952 10912
rect 5016 10848 5032 10912
rect 5096 10848 5112 10912
rect 5176 10848 5192 10912
rect 5256 10848 5264 10912
rect 4944 10847 5264 10848
rect 12944 10912 13264 10913
rect 12944 10848 12952 10912
rect 13016 10848 13032 10912
rect 13096 10848 13112 10912
rect 13176 10848 13192 10912
rect 13256 10848 13264 10912
rect 12944 10847 13264 10848
rect 20944 10912 21264 10913
rect 20944 10848 20952 10912
rect 21016 10848 21032 10912
rect 21096 10848 21112 10912
rect 21176 10848 21192 10912
rect 21256 10848 21264 10912
rect 20944 10847 21264 10848
rect 0 10704 480 10736
rect 0 10648 110 10704
rect 166 10648 480 10704
rect 0 10616 480 10648
rect 3601 10706 3667 10709
rect 7465 10706 7531 10709
rect 3601 10704 7531 10706
rect 3601 10648 3606 10704
rect 3662 10648 7470 10704
rect 7526 10648 7531 10704
rect 3601 10646 7531 10648
rect 3601 10643 3667 10646
rect 7465 10643 7531 10646
rect 0 10432 480 10464
rect 0 10376 18 10432
rect 74 10376 480 10432
rect 0 10344 480 10376
rect 8944 10368 9264 10369
rect 8944 10304 8952 10368
rect 9016 10304 9032 10368
rect 9096 10304 9112 10368
rect 9176 10304 9192 10368
rect 9256 10304 9264 10368
rect 8944 10303 9264 10304
rect 16944 10368 17264 10369
rect 16944 10304 16952 10368
rect 17016 10304 17032 10368
rect 17096 10304 17112 10368
rect 17176 10304 17192 10368
rect 17256 10304 17264 10368
rect 16944 10303 17264 10304
rect 0 10024 480 10056
rect 0 9968 110 10024
rect 166 9968 480 10024
rect 0 9936 480 9968
rect 4944 9824 5264 9825
rect 4944 9760 4952 9824
rect 5016 9760 5032 9824
rect 5096 9760 5112 9824
rect 5176 9760 5192 9824
rect 5256 9760 5264 9824
rect 4944 9759 5264 9760
rect 12944 9824 13264 9825
rect 12944 9760 12952 9824
rect 13016 9760 13032 9824
rect 13096 9760 13112 9824
rect 13176 9760 13192 9824
rect 13256 9760 13264 9824
rect 12944 9759 13264 9760
rect 20944 9824 21264 9825
rect 20944 9760 20952 9824
rect 21016 9760 21032 9824
rect 21096 9760 21112 9824
rect 21176 9760 21192 9824
rect 21256 9760 21264 9824
rect 20944 9759 21264 9760
rect 0 9528 480 9648
rect 62 9482 122 9528
rect 3325 9482 3391 9485
rect 62 9480 3391 9482
rect 62 9424 3330 9480
rect 3386 9424 3391 9480
rect 62 9422 3391 9424
rect 3325 9419 3391 9422
rect 8944 9280 9264 9281
rect 0 9208 480 9240
rect 8944 9216 8952 9280
rect 9016 9216 9032 9280
rect 9096 9216 9112 9280
rect 9176 9216 9192 9280
rect 9256 9216 9264 9280
rect 8944 9215 9264 9216
rect 16944 9280 17264 9281
rect 16944 9216 16952 9280
rect 17016 9216 17032 9280
rect 17096 9216 17112 9280
rect 17176 9216 17192 9280
rect 17256 9216 17264 9280
rect 16944 9215 17264 9216
rect 0 9152 18 9208
rect 74 9152 480 9208
rect 0 9120 480 9152
rect 0 8800 480 8832
rect 0 8744 110 8800
rect 166 8744 480 8800
rect 0 8712 480 8744
rect 4944 8736 5264 8737
rect 4944 8672 4952 8736
rect 5016 8672 5032 8736
rect 5096 8672 5112 8736
rect 5176 8672 5192 8736
rect 5256 8672 5264 8736
rect 4944 8671 5264 8672
rect 12944 8736 13264 8737
rect 12944 8672 12952 8736
rect 13016 8672 13032 8736
rect 13096 8672 13112 8736
rect 13176 8672 13192 8736
rect 13256 8672 13264 8736
rect 12944 8671 13264 8672
rect 20944 8736 21264 8737
rect 20944 8672 20952 8736
rect 21016 8672 21032 8736
rect 21096 8672 21112 8736
rect 21176 8672 21192 8736
rect 21256 8672 21264 8736
rect 20944 8671 21264 8672
rect 0 8392 480 8424
rect 0 8336 110 8392
rect 166 8336 480 8392
rect 0 8304 480 8336
rect 8944 8192 9264 8193
rect 8944 8128 8952 8192
rect 9016 8128 9032 8192
rect 9096 8128 9112 8192
rect 9176 8128 9192 8192
rect 9256 8128 9264 8192
rect 8944 8127 9264 8128
rect 16944 8192 17264 8193
rect 16944 8128 16952 8192
rect 17016 8128 17032 8192
rect 17096 8128 17112 8192
rect 17176 8128 17192 8192
rect 17256 8128 17264 8192
rect 16944 8127 17264 8128
rect 0 7984 480 8016
rect 0 7928 110 7984
rect 166 7928 480 7984
rect 0 7896 480 7928
rect 4944 7648 5264 7649
rect 0 7576 480 7608
rect 4944 7584 4952 7648
rect 5016 7584 5032 7648
rect 5096 7584 5112 7648
rect 5176 7584 5192 7648
rect 5256 7584 5264 7648
rect 4944 7583 5264 7584
rect 12944 7648 13264 7649
rect 12944 7584 12952 7648
rect 13016 7584 13032 7648
rect 13096 7584 13112 7648
rect 13176 7584 13192 7648
rect 13256 7584 13264 7648
rect 12944 7583 13264 7584
rect 20944 7648 21264 7649
rect 20944 7584 20952 7648
rect 21016 7584 21032 7648
rect 21096 7584 21112 7648
rect 21176 7584 21192 7648
rect 21256 7584 21264 7648
rect 20944 7583 21264 7584
rect 0 7520 18 7576
rect 74 7520 480 7576
rect 0 7488 480 7520
rect 1577 7306 1643 7309
rect 62 7304 1643 7306
rect 62 7248 1582 7304
rect 1638 7248 1643 7304
rect 62 7246 1643 7248
rect 62 7200 122 7246
rect 1577 7243 1643 7246
rect 0 7080 480 7200
rect 8944 7104 9264 7105
rect 8944 7040 8952 7104
rect 9016 7040 9032 7104
rect 9096 7040 9112 7104
rect 9176 7040 9192 7104
rect 9256 7040 9264 7104
rect 8944 7039 9264 7040
rect 16944 7104 17264 7105
rect 16944 7040 16952 7104
rect 17016 7040 17032 7104
rect 17096 7040 17112 7104
rect 17176 7040 17192 7104
rect 17256 7040 17264 7104
rect 16944 7039 17264 7040
rect 0 6896 480 6928
rect 0 6840 110 6896
rect 166 6840 480 6896
rect 0 6808 480 6840
rect 4944 6560 5264 6561
rect 0 6488 480 6520
rect 4944 6496 4952 6560
rect 5016 6496 5032 6560
rect 5096 6496 5112 6560
rect 5176 6496 5192 6560
rect 5256 6496 5264 6560
rect 4944 6495 5264 6496
rect 12944 6560 13264 6561
rect 12944 6496 12952 6560
rect 13016 6496 13032 6560
rect 13096 6496 13112 6560
rect 13176 6496 13192 6560
rect 13256 6496 13264 6560
rect 12944 6495 13264 6496
rect 20944 6560 21264 6561
rect 20944 6496 20952 6560
rect 21016 6496 21032 6560
rect 21096 6496 21112 6560
rect 21176 6496 21192 6560
rect 21256 6496 21264 6560
rect 20944 6495 21264 6496
rect 0 6432 110 6488
rect 166 6432 480 6488
rect 0 6400 480 6432
rect 0 6084 480 6112
rect 0 6020 60 6084
rect 124 6020 480 6084
rect 0 5992 480 6020
rect 8944 6016 9264 6017
rect 8944 5952 8952 6016
rect 9016 5952 9032 6016
rect 9096 5952 9112 6016
rect 9176 5952 9192 6016
rect 9256 5952 9264 6016
rect 8944 5951 9264 5952
rect 16944 6016 17264 6017
rect 16944 5952 16952 6016
rect 17016 5952 17032 6016
rect 17096 5952 17112 6016
rect 17176 5952 17192 6016
rect 17256 5952 17264 6016
rect 16944 5951 17264 5952
rect 0 5672 480 5704
rect 0 5616 18 5672
rect 74 5616 480 5672
rect 0 5584 480 5616
rect 4944 5472 5264 5473
rect 4944 5408 4952 5472
rect 5016 5408 5032 5472
rect 5096 5408 5112 5472
rect 5176 5408 5192 5472
rect 5256 5408 5264 5472
rect 4944 5407 5264 5408
rect 12944 5472 13264 5473
rect 12944 5408 12952 5472
rect 13016 5408 13032 5472
rect 13096 5408 13112 5472
rect 13176 5408 13192 5472
rect 13256 5408 13264 5472
rect 12944 5407 13264 5408
rect 20944 5472 21264 5473
rect 20944 5408 20952 5472
rect 21016 5408 21032 5472
rect 21096 5408 21112 5472
rect 21176 5408 21192 5472
rect 21256 5408 21264 5472
rect 20944 5407 21264 5408
rect 0 5264 480 5296
rect 0 5208 110 5264
rect 166 5208 480 5264
rect 0 5176 480 5208
rect 54 5068 60 5132
rect 124 5130 130 5132
rect 124 5070 4170 5130
rect 124 5068 130 5070
rect 4110 4997 4170 5070
rect 4110 4992 4219 4997
rect 4110 4936 4158 4992
rect 4214 4936 4219 4992
rect 4110 4934 4219 4936
rect 4153 4931 4219 4934
rect 8944 4928 9264 4929
rect 0 4856 480 4888
rect 8944 4864 8952 4928
rect 9016 4864 9032 4928
rect 9096 4864 9112 4928
rect 9176 4864 9192 4928
rect 9256 4864 9264 4928
rect 8944 4863 9264 4864
rect 16944 4928 17264 4929
rect 16944 4864 16952 4928
rect 17016 4864 17032 4928
rect 17096 4864 17112 4928
rect 17176 4864 17192 4928
rect 17256 4864 17264 4928
rect 16944 4863 17264 4864
rect 0 4800 110 4856
rect 166 4800 480 4856
rect 0 4768 480 4800
rect 0 4448 480 4480
rect 0 4392 110 4448
rect 166 4392 480 4448
rect 0 4360 480 4392
rect 4944 4384 5264 4385
rect 4944 4320 4952 4384
rect 5016 4320 5032 4384
rect 5096 4320 5112 4384
rect 5176 4320 5192 4384
rect 5256 4320 5264 4384
rect 4944 4319 5264 4320
rect 12944 4384 13264 4385
rect 12944 4320 12952 4384
rect 13016 4320 13032 4384
rect 13096 4320 13112 4384
rect 13176 4320 13192 4384
rect 13256 4320 13264 4384
rect 12944 4319 13264 4320
rect 20944 4384 21264 4385
rect 20944 4320 20952 4384
rect 21016 4320 21032 4384
rect 21096 4320 21112 4384
rect 21176 4320 21192 4384
rect 21256 4320 21264 4384
rect 20944 4319 21264 4320
rect 0 4040 480 4072
rect 0 3984 18 4040
rect 74 3984 480 4040
rect 0 3952 480 3984
rect 8944 3840 9264 3841
rect 8944 3776 8952 3840
rect 9016 3776 9032 3840
rect 9096 3776 9112 3840
rect 9176 3776 9192 3840
rect 9256 3776 9264 3840
rect 8944 3775 9264 3776
rect 16944 3840 17264 3841
rect 16944 3776 16952 3840
rect 17016 3776 17032 3840
rect 17096 3776 17112 3840
rect 17176 3776 17192 3840
rect 17256 3776 17264 3840
rect 16944 3775 17264 3776
rect 0 3632 480 3664
rect 0 3576 110 3632
rect 166 3576 480 3632
rect 0 3544 480 3576
rect 0 3360 480 3392
rect 0 3304 110 3360
rect 166 3304 480 3360
rect 0 3272 480 3304
rect 4944 3296 5264 3297
rect 4944 3232 4952 3296
rect 5016 3232 5032 3296
rect 5096 3232 5112 3296
rect 5176 3232 5192 3296
rect 5256 3232 5264 3296
rect 4944 3231 5264 3232
rect 12944 3296 13264 3297
rect 12944 3232 12952 3296
rect 13016 3232 13032 3296
rect 13096 3232 13112 3296
rect 13176 3232 13192 3296
rect 13256 3232 13264 3296
rect 12944 3231 13264 3232
rect 20944 3296 21264 3297
rect 20944 3232 20952 3296
rect 21016 3232 21032 3296
rect 21096 3232 21112 3296
rect 21176 3232 21192 3296
rect 21256 3232 21264 3296
rect 20944 3231 21264 3232
rect 0 2952 480 2984
rect 0 2896 386 2952
rect 442 2896 480 2952
rect 0 2864 480 2896
rect 8944 2752 9264 2753
rect 8944 2688 8952 2752
rect 9016 2688 9032 2752
rect 9096 2688 9112 2752
rect 9176 2688 9192 2752
rect 9256 2688 9264 2752
rect 8944 2687 9264 2688
rect 16944 2752 17264 2753
rect 16944 2688 16952 2752
rect 17016 2688 17032 2752
rect 17096 2688 17112 2752
rect 17176 2688 17192 2752
rect 17256 2688 17264 2752
rect 16944 2687 17264 2688
rect 0 2544 480 2576
rect 0 2488 386 2544
rect 442 2488 480 2544
rect 0 2456 480 2488
rect 4944 2208 5264 2209
rect 0 2136 480 2168
rect 4944 2144 4952 2208
rect 5016 2144 5032 2208
rect 5096 2144 5112 2208
rect 5176 2144 5192 2208
rect 5256 2144 5264 2208
rect 4944 2143 5264 2144
rect 12944 2208 13264 2209
rect 12944 2144 12952 2208
rect 13016 2144 13032 2208
rect 13096 2144 13112 2208
rect 13176 2144 13192 2208
rect 13256 2144 13264 2208
rect 12944 2143 13264 2144
rect 20944 2208 21264 2209
rect 20944 2144 20952 2208
rect 21016 2144 21032 2208
rect 21096 2144 21112 2208
rect 21176 2144 21192 2208
rect 21256 2144 21264 2208
rect 20944 2143 21264 2144
rect 0 2080 18 2136
rect 74 2080 480 2136
rect 0 2048 480 2080
rect 0 1728 480 1760
rect 0 1672 110 1728
rect 166 1672 480 1728
rect 0 1640 480 1672
rect 0 1320 480 1352
rect 0 1264 18 1320
rect 74 1264 480 1320
rect 0 1232 480 1264
rect 0 912 480 944
rect 0 856 110 912
rect 166 856 480 912
rect 0 824 480 856
rect 3417 642 3483 645
rect 62 640 3483 642
rect 62 584 3422 640
rect 3478 584 3483 640
rect 62 582 3483 584
rect 62 536 122 582
rect 3417 579 3483 582
rect 0 416 480 536
rect 0 232 480 264
rect 0 176 110 232
rect 166 176 480 232
rect 0 144 480 176
<< via3 >>
rect 60 22068 124 22132
rect 4952 21788 5016 21792
rect 4952 21732 4956 21788
rect 4956 21732 5012 21788
rect 5012 21732 5016 21788
rect 4952 21728 5016 21732
rect 5032 21788 5096 21792
rect 5032 21732 5036 21788
rect 5036 21732 5092 21788
rect 5092 21732 5096 21788
rect 5032 21728 5096 21732
rect 5112 21788 5176 21792
rect 5112 21732 5116 21788
rect 5116 21732 5172 21788
rect 5172 21732 5176 21788
rect 5112 21728 5176 21732
rect 5192 21788 5256 21792
rect 5192 21732 5196 21788
rect 5196 21732 5252 21788
rect 5252 21732 5256 21788
rect 5192 21728 5256 21732
rect 12952 21788 13016 21792
rect 12952 21732 12956 21788
rect 12956 21732 13012 21788
rect 13012 21732 13016 21788
rect 12952 21728 13016 21732
rect 13032 21788 13096 21792
rect 13032 21732 13036 21788
rect 13036 21732 13092 21788
rect 13092 21732 13096 21788
rect 13032 21728 13096 21732
rect 13112 21788 13176 21792
rect 13112 21732 13116 21788
rect 13116 21732 13172 21788
rect 13172 21732 13176 21788
rect 13112 21728 13176 21732
rect 13192 21788 13256 21792
rect 13192 21732 13196 21788
rect 13196 21732 13252 21788
rect 13252 21732 13256 21788
rect 13192 21728 13256 21732
rect 20952 21788 21016 21792
rect 20952 21732 20956 21788
rect 20956 21732 21012 21788
rect 21012 21732 21016 21788
rect 20952 21728 21016 21732
rect 21032 21788 21096 21792
rect 21032 21732 21036 21788
rect 21036 21732 21092 21788
rect 21092 21732 21096 21788
rect 21032 21728 21096 21732
rect 21112 21788 21176 21792
rect 21112 21732 21116 21788
rect 21116 21732 21172 21788
rect 21172 21732 21176 21788
rect 21112 21728 21176 21732
rect 21192 21788 21256 21792
rect 21192 21732 21196 21788
rect 21196 21732 21252 21788
rect 21252 21732 21256 21788
rect 21192 21728 21256 21732
rect 612 21388 676 21452
rect 8952 21244 9016 21248
rect 8952 21188 8956 21244
rect 8956 21188 9012 21244
rect 9012 21188 9016 21244
rect 8952 21184 9016 21188
rect 9032 21244 9096 21248
rect 9032 21188 9036 21244
rect 9036 21188 9092 21244
rect 9092 21188 9096 21244
rect 9032 21184 9096 21188
rect 9112 21244 9176 21248
rect 9112 21188 9116 21244
rect 9116 21188 9172 21244
rect 9172 21188 9176 21244
rect 9112 21184 9176 21188
rect 9192 21244 9256 21248
rect 9192 21188 9196 21244
rect 9196 21188 9252 21244
rect 9252 21188 9256 21244
rect 9192 21184 9256 21188
rect 16952 21244 17016 21248
rect 16952 21188 16956 21244
rect 16956 21188 17012 21244
rect 17012 21188 17016 21244
rect 16952 21184 17016 21188
rect 17032 21244 17096 21248
rect 17032 21188 17036 21244
rect 17036 21188 17092 21244
rect 17092 21188 17096 21244
rect 17032 21184 17096 21188
rect 17112 21244 17176 21248
rect 17112 21188 17116 21244
rect 17116 21188 17172 21244
rect 17172 21188 17176 21244
rect 17112 21184 17176 21188
rect 17192 21244 17256 21248
rect 17192 21188 17196 21244
rect 17196 21188 17252 21244
rect 17252 21188 17256 21244
rect 17192 21184 17256 21188
rect 4952 20700 5016 20704
rect 4952 20644 4956 20700
rect 4956 20644 5012 20700
rect 5012 20644 5016 20700
rect 4952 20640 5016 20644
rect 5032 20700 5096 20704
rect 5032 20644 5036 20700
rect 5036 20644 5092 20700
rect 5092 20644 5096 20700
rect 5032 20640 5096 20644
rect 5112 20700 5176 20704
rect 5112 20644 5116 20700
rect 5116 20644 5172 20700
rect 5172 20644 5176 20700
rect 5112 20640 5176 20644
rect 5192 20700 5256 20704
rect 5192 20644 5196 20700
rect 5196 20644 5252 20700
rect 5252 20644 5256 20700
rect 5192 20640 5256 20644
rect 12952 20700 13016 20704
rect 12952 20644 12956 20700
rect 12956 20644 13012 20700
rect 13012 20644 13016 20700
rect 12952 20640 13016 20644
rect 13032 20700 13096 20704
rect 13032 20644 13036 20700
rect 13036 20644 13092 20700
rect 13092 20644 13096 20700
rect 13032 20640 13096 20644
rect 13112 20700 13176 20704
rect 13112 20644 13116 20700
rect 13116 20644 13172 20700
rect 13172 20644 13176 20700
rect 13112 20640 13176 20644
rect 13192 20700 13256 20704
rect 13192 20644 13196 20700
rect 13196 20644 13252 20700
rect 13252 20644 13256 20700
rect 13192 20640 13256 20644
rect 20952 20700 21016 20704
rect 20952 20644 20956 20700
rect 20956 20644 21012 20700
rect 21012 20644 21016 20700
rect 20952 20640 21016 20644
rect 21032 20700 21096 20704
rect 21032 20644 21036 20700
rect 21036 20644 21092 20700
rect 21092 20644 21096 20700
rect 21032 20640 21096 20644
rect 21112 20700 21176 20704
rect 21112 20644 21116 20700
rect 21116 20644 21172 20700
rect 21172 20644 21176 20700
rect 21112 20640 21176 20644
rect 21192 20700 21256 20704
rect 21192 20644 21196 20700
rect 21196 20644 21252 20700
rect 21252 20644 21256 20700
rect 21192 20640 21256 20644
rect 60 20572 124 20636
rect 60 20334 124 20398
rect 60 20164 124 20228
rect 8952 20156 9016 20160
rect 8952 20100 8956 20156
rect 8956 20100 9012 20156
rect 9012 20100 9016 20156
rect 8952 20096 9016 20100
rect 9032 20156 9096 20160
rect 9032 20100 9036 20156
rect 9036 20100 9092 20156
rect 9092 20100 9096 20156
rect 9032 20096 9096 20100
rect 9112 20156 9176 20160
rect 9112 20100 9116 20156
rect 9116 20100 9172 20156
rect 9172 20100 9176 20156
rect 9112 20096 9176 20100
rect 9192 20156 9256 20160
rect 9192 20100 9196 20156
rect 9196 20100 9252 20156
rect 9252 20100 9256 20156
rect 9192 20096 9256 20100
rect 16952 20156 17016 20160
rect 16952 20100 16956 20156
rect 16956 20100 17012 20156
rect 17012 20100 17016 20156
rect 16952 20096 17016 20100
rect 17032 20156 17096 20160
rect 17032 20100 17036 20156
rect 17036 20100 17092 20156
rect 17092 20100 17096 20156
rect 17032 20096 17096 20100
rect 17112 20156 17176 20160
rect 17112 20100 17116 20156
rect 17116 20100 17172 20156
rect 17172 20100 17176 20156
rect 17112 20096 17176 20100
rect 17192 20156 17256 20160
rect 17192 20100 17196 20156
rect 17196 20100 17252 20156
rect 17252 20100 17256 20156
rect 17192 20096 17256 20100
rect 612 20028 676 20092
rect 4952 19612 5016 19616
rect 4952 19556 4956 19612
rect 4956 19556 5012 19612
rect 5012 19556 5016 19612
rect 4952 19552 5016 19556
rect 5032 19612 5096 19616
rect 5032 19556 5036 19612
rect 5036 19556 5092 19612
rect 5092 19556 5096 19612
rect 5032 19552 5096 19556
rect 5112 19612 5176 19616
rect 5112 19556 5116 19612
rect 5116 19556 5172 19612
rect 5172 19556 5176 19612
rect 5112 19552 5176 19556
rect 5192 19612 5256 19616
rect 5192 19556 5196 19612
rect 5196 19556 5252 19612
rect 5252 19556 5256 19612
rect 5192 19552 5256 19556
rect 12952 19612 13016 19616
rect 12952 19556 12956 19612
rect 12956 19556 13012 19612
rect 13012 19556 13016 19612
rect 12952 19552 13016 19556
rect 13032 19612 13096 19616
rect 13032 19556 13036 19612
rect 13036 19556 13092 19612
rect 13092 19556 13096 19612
rect 13032 19552 13096 19556
rect 13112 19612 13176 19616
rect 13112 19556 13116 19612
rect 13116 19556 13172 19612
rect 13172 19556 13176 19612
rect 13112 19552 13176 19556
rect 13192 19612 13256 19616
rect 13192 19556 13196 19612
rect 13196 19556 13252 19612
rect 13252 19556 13256 19612
rect 13192 19552 13256 19556
rect 20952 19612 21016 19616
rect 20952 19556 20956 19612
rect 20956 19556 21012 19612
rect 21012 19556 21016 19612
rect 20952 19552 21016 19556
rect 21032 19612 21096 19616
rect 21032 19556 21036 19612
rect 21036 19556 21092 19612
rect 21092 19556 21096 19612
rect 21032 19552 21096 19556
rect 21112 19612 21176 19616
rect 21112 19556 21116 19612
rect 21116 19556 21172 19612
rect 21172 19556 21176 19612
rect 21112 19552 21176 19556
rect 21192 19612 21256 19616
rect 21192 19556 21196 19612
rect 21196 19556 21252 19612
rect 21252 19556 21256 19612
rect 21192 19552 21256 19556
rect 8952 19068 9016 19072
rect 8952 19012 8956 19068
rect 8956 19012 9012 19068
rect 9012 19012 9016 19068
rect 8952 19008 9016 19012
rect 9032 19068 9096 19072
rect 9032 19012 9036 19068
rect 9036 19012 9092 19068
rect 9092 19012 9096 19068
rect 9032 19008 9096 19012
rect 9112 19068 9176 19072
rect 9112 19012 9116 19068
rect 9116 19012 9172 19068
rect 9172 19012 9176 19068
rect 9112 19008 9176 19012
rect 9192 19068 9256 19072
rect 9192 19012 9196 19068
rect 9196 19012 9252 19068
rect 9252 19012 9256 19068
rect 9192 19008 9256 19012
rect 16952 19068 17016 19072
rect 16952 19012 16956 19068
rect 16956 19012 17012 19068
rect 17012 19012 17016 19068
rect 16952 19008 17016 19012
rect 17032 19068 17096 19072
rect 17032 19012 17036 19068
rect 17036 19012 17092 19068
rect 17092 19012 17096 19068
rect 17032 19008 17096 19012
rect 17112 19068 17176 19072
rect 17112 19012 17116 19068
rect 17116 19012 17172 19068
rect 17172 19012 17176 19068
rect 17112 19008 17176 19012
rect 17192 19068 17256 19072
rect 17192 19012 17196 19068
rect 17196 19012 17252 19068
rect 17252 19012 17256 19068
rect 17192 19008 17256 19012
rect 60 18940 124 19004
rect 612 18668 676 18732
rect 4952 18524 5016 18528
rect 4952 18468 4956 18524
rect 4956 18468 5012 18524
rect 5012 18468 5016 18524
rect 4952 18464 5016 18468
rect 5032 18524 5096 18528
rect 5032 18468 5036 18524
rect 5036 18468 5092 18524
rect 5092 18468 5096 18524
rect 5032 18464 5096 18468
rect 5112 18524 5176 18528
rect 5112 18468 5116 18524
rect 5116 18468 5172 18524
rect 5172 18468 5176 18524
rect 5112 18464 5176 18468
rect 5192 18524 5256 18528
rect 5192 18468 5196 18524
rect 5196 18468 5252 18524
rect 5252 18468 5256 18524
rect 5192 18464 5256 18468
rect 12952 18524 13016 18528
rect 12952 18468 12956 18524
rect 12956 18468 13012 18524
rect 13012 18468 13016 18524
rect 12952 18464 13016 18468
rect 13032 18524 13096 18528
rect 13032 18468 13036 18524
rect 13036 18468 13092 18524
rect 13092 18468 13096 18524
rect 13032 18464 13096 18468
rect 13112 18524 13176 18528
rect 13112 18468 13116 18524
rect 13116 18468 13172 18524
rect 13172 18468 13176 18524
rect 13112 18464 13176 18468
rect 13192 18524 13256 18528
rect 13192 18468 13196 18524
rect 13196 18468 13252 18524
rect 13252 18468 13256 18524
rect 13192 18464 13256 18468
rect 20952 18524 21016 18528
rect 20952 18468 20956 18524
rect 20956 18468 21012 18524
rect 21012 18468 21016 18524
rect 20952 18464 21016 18468
rect 21032 18524 21096 18528
rect 21032 18468 21036 18524
rect 21036 18468 21092 18524
rect 21092 18468 21096 18524
rect 21032 18464 21096 18468
rect 21112 18524 21176 18528
rect 21112 18468 21116 18524
rect 21116 18468 21172 18524
rect 21172 18468 21176 18524
rect 21112 18464 21176 18468
rect 21192 18524 21256 18528
rect 21192 18468 21196 18524
rect 21196 18468 21252 18524
rect 21252 18468 21256 18524
rect 21192 18464 21256 18468
rect 8952 17980 9016 17984
rect 8952 17924 8956 17980
rect 8956 17924 9012 17980
rect 9012 17924 9016 17980
rect 8952 17920 9016 17924
rect 9032 17980 9096 17984
rect 9032 17924 9036 17980
rect 9036 17924 9092 17980
rect 9092 17924 9096 17980
rect 9032 17920 9096 17924
rect 9112 17980 9176 17984
rect 9112 17924 9116 17980
rect 9116 17924 9172 17980
rect 9172 17924 9176 17980
rect 9112 17920 9176 17924
rect 9192 17980 9256 17984
rect 9192 17924 9196 17980
rect 9196 17924 9252 17980
rect 9252 17924 9256 17980
rect 9192 17920 9256 17924
rect 16952 17980 17016 17984
rect 16952 17924 16956 17980
rect 16956 17924 17012 17980
rect 17012 17924 17016 17980
rect 16952 17920 17016 17924
rect 17032 17980 17096 17984
rect 17032 17924 17036 17980
rect 17036 17924 17092 17980
rect 17092 17924 17096 17980
rect 17032 17920 17096 17924
rect 17112 17980 17176 17984
rect 17112 17924 17116 17980
rect 17116 17924 17172 17980
rect 17172 17924 17176 17980
rect 17112 17920 17176 17924
rect 17192 17980 17256 17984
rect 17192 17924 17196 17980
rect 17196 17924 17252 17980
rect 17252 17924 17256 17980
rect 17192 17920 17256 17924
rect 4952 17436 5016 17440
rect 4952 17380 4956 17436
rect 4956 17380 5012 17436
rect 5012 17380 5016 17436
rect 4952 17376 5016 17380
rect 5032 17436 5096 17440
rect 5032 17380 5036 17436
rect 5036 17380 5092 17436
rect 5092 17380 5096 17436
rect 5032 17376 5096 17380
rect 5112 17436 5176 17440
rect 5112 17380 5116 17436
rect 5116 17380 5172 17436
rect 5172 17380 5176 17436
rect 5112 17376 5176 17380
rect 5192 17436 5256 17440
rect 5192 17380 5196 17436
rect 5196 17380 5252 17436
rect 5252 17380 5256 17436
rect 5192 17376 5256 17380
rect 12952 17436 13016 17440
rect 12952 17380 12956 17436
rect 12956 17380 13012 17436
rect 13012 17380 13016 17436
rect 12952 17376 13016 17380
rect 13032 17436 13096 17440
rect 13032 17380 13036 17436
rect 13036 17380 13092 17436
rect 13092 17380 13096 17436
rect 13032 17376 13096 17380
rect 13112 17436 13176 17440
rect 13112 17380 13116 17436
rect 13116 17380 13172 17436
rect 13172 17380 13176 17436
rect 13112 17376 13176 17380
rect 13192 17436 13256 17440
rect 13192 17380 13196 17436
rect 13196 17380 13252 17436
rect 13252 17380 13256 17436
rect 13192 17376 13256 17380
rect 20952 17436 21016 17440
rect 20952 17380 20956 17436
rect 20956 17380 21012 17436
rect 21012 17380 21016 17436
rect 20952 17376 21016 17380
rect 21032 17436 21096 17440
rect 21032 17380 21036 17436
rect 21036 17380 21092 17436
rect 21092 17380 21096 17436
rect 21032 17376 21096 17380
rect 21112 17436 21176 17440
rect 21112 17380 21116 17436
rect 21116 17380 21172 17436
rect 21172 17380 21176 17436
rect 21112 17376 21176 17380
rect 21192 17436 21256 17440
rect 21192 17380 21196 17436
rect 21196 17380 21252 17436
rect 21252 17380 21256 17436
rect 21192 17376 21256 17380
rect 8952 16892 9016 16896
rect 8952 16836 8956 16892
rect 8956 16836 9012 16892
rect 9012 16836 9016 16892
rect 8952 16832 9016 16836
rect 9032 16892 9096 16896
rect 9032 16836 9036 16892
rect 9036 16836 9092 16892
rect 9092 16836 9096 16892
rect 9032 16832 9096 16836
rect 9112 16892 9176 16896
rect 9112 16836 9116 16892
rect 9116 16836 9172 16892
rect 9172 16836 9176 16892
rect 9112 16832 9176 16836
rect 9192 16892 9256 16896
rect 9192 16836 9196 16892
rect 9196 16836 9252 16892
rect 9252 16836 9256 16892
rect 9192 16832 9256 16836
rect 16952 16892 17016 16896
rect 16952 16836 16956 16892
rect 16956 16836 17012 16892
rect 17012 16836 17016 16892
rect 16952 16832 17016 16836
rect 17032 16892 17096 16896
rect 17032 16836 17036 16892
rect 17036 16836 17092 16892
rect 17092 16836 17096 16892
rect 17032 16832 17096 16836
rect 17112 16892 17176 16896
rect 17112 16836 17116 16892
rect 17116 16836 17172 16892
rect 17172 16836 17176 16892
rect 17112 16832 17176 16836
rect 17192 16892 17256 16896
rect 17192 16836 17196 16892
rect 17196 16836 17252 16892
rect 17252 16836 17256 16892
rect 17192 16832 17256 16836
rect 4952 16348 5016 16352
rect 4952 16292 4956 16348
rect 4956 16292 5012 16348
rect 5012 16292 5016 16348
rect 4952 16288 5016 16292
rect 5032 16348 5096 16352
rect 5032 16292 5036 16348
rect 5036 16292 5092 16348
rect 5092 16292 5096 16348
rect 5032 16288 5096 16292
rect 5112 16348 5176 16352
rect 5112 16292 5116 16348
rect 5116 16292 5172 16348
rect 5172 16292 5176 16348
rect 5112 16288 5176 16292
rect 5192 16348 5256 16352
rect 5192 16292 5196 16348
rect 5196 16292 5252 16348
rect 5252 16292 5256 16348
rect 5192 16288 5256 16292
rect 12952 16348 13016 16352
rect 12952 16292 12956 16348
rect 12956 16292 13012 16348
rect 13012 16292 13016 16348
rect 12952 16288 13016 16292
rect 13032 16348 13096 16352
rect 13032 16292 13036 16348
rect 13036 16292 13092 16348
rect 13092 16292 13096 16348
rect 13032 16288 13096 16292
rect 13112 16348 13176 16352
rect 13112 16292 13116 16348
rect 13116 16292 13172 16348
rect 13172 16292 13176 16348
rect 13112 16288 13176 16292
rect 13192 16348 13256 16352
rect 13192 16292 13196 16348
rect 13196 16292 13252 16348
rect 13252 16292 13256 16348
rect 13192 16288 13256 16292
rect 20952 16348 21016 16352
rect 20952 16292 20956 16348
rect 20956 16292 21012 16348
rect 21012 16292 21016 16348
rect 20952 16288 21016 16292
rect 21032 16348 21096 16352
rect 21032 16292 21036 16348
rect 21036 16292 21092 16348
rect 21092 16292 21096 16348
rect 21032 16288 21096 16292
rect 21112 16348 21176 16352
rect 21112 16292 21116 16348
rect 21116 16292 21172 16348
rect 21172 16292 21176 16348
rect 21112 16288 21176 16292
rect 21192 16348 21256 16352
rect 21192 16292 21196 16348
rect 21196 16292 21252 16348
rect 21252 16292 21256 16348
rect 21192 16288 21256 16292
rect 612 15948 676 16012
rect 8952 15804 9016 15808
rect 8952 15748 8956 15804
rect 8956 15748 9012 15804
rect 9012 15748 9016 15804
rect 8952 15744 9016 15748
rect 9032 15804 9096 15808
rect 9032 15748 9036 15804
rect 9036 15748 9092 15804
rect 9092 15748 9096 15804
rect 9032 15744 9096 15748
rect 9112 15804 9176 15808
rect 9112 15748 9116 15804
rect 9116 15748 9172 15804
rect 9172 15748 9176 15804
rect 9112 15744 9176 15748
rect 9192 15804 9256 15808
rect 9192 15748 9196 15804
rect 9196 15748 9252 15804
rect 9252 15748 9256 15804
rect 9192 15744 9256 15748
rect 16952 15804 17016 15808
rect 16952 15748 16956 15804
rect 16956 15748 17012 15804
rect 17012 15748 17016 15804
rect 16952 15744 17016 15748
rect 17032 15804 17096 15808
rect 17032 15748 17036 15804
rect 17036 15748 17092 15804
rect 17092 15748 17096 15804
rect 17032 15744 17096 15748
rect 17112 15804 17176 15808
rect 17112 15748 17116 15804
rect 17116 15748 17172 15804
rect 17172 15748 17176 15804
rect 17112 15744 17176 15748
rect 17192 15804 17256 15808
rect 17192 15748 17196 15804
rect 17196 15748 17252 15804
rect 17252 15748 17256 15804
rect 17192 15744 17256 15748
rect 60 15404 124 15468
rect 4952 15260 5016 15264
rect 4952 15204 4956 15260
rect 4956 15204 5012 15260
rect 5012 15204 5016 15260
rect 4952 15200 5016 15204
rect 5032 15260 5096 15264
rect 5032 15204 5036 15260
rect 5036 15204 5092 15260
rect 5092 15204 5096 15260
rect 5032 15200 5096 15204
rect 5112 15260 5176 15264
rect 5112 15204 5116 15260
rect 5116 15204 5172 15260
rect 5172 15204 5176 15260
rect 5112 15200 5176 15204
rect 5192 15260 5256 15264
rect 5192 15204 5196 15260
rect 5196 15204 5252 15260
rect 5252 15204 5256 15260
rect 5192 15200 5256 15204
rect 12952 15260 13016 15264
rect 12952 15204 12956 15260
rect 12956 15204 13012 15260
rect 13012 15204 13016 15260
rect 12952 15200 13016 15204
rect 13032 15260 13096 15264
rect 13032 15204 13036 15260
rect 13036 15204 13092 15260
rect 13092 15204 13096 15260
rect 13032 15200 13096 15204
rect 13112 15260 13176 15264
rect 13112 15204 13116 15260
rect 13116 15204 13172 15260
rect 13172 15204 13176 15260
rect 13112 15200 13176 15204
rect 13192 15260 13256 15264
rect 13192 15204 13196 15260
rect 13196 15204 13252 15260
rect 13252 15204 13256 15260
rect 13192 15200 13256 15204
rect 20952 15260 21016 15264
rect 20952 15204 20956 15260
rect 20956 15204 21012 15260
rect 21012 15204 21016 15260
rect 20952 15200 21016 15204
rect 21032 15260 21096 15264
rect 21032 15204 21036 15260
rect 21036 15204 21092 15260
rect 21092 15204 21096 15260
rect 21032 15200 21096 15204
rect 21112 15260 21176 15264
rect 21112 15204 21116 15260
rect 21116 15204 21172 15260
rect 21172 15204 21176 15260
rect 21112 15200 21176 15204
rect 21192 15260 21256 15264
rect 21192 15204 21196 15260
rect 21196 15204 21252 15260
rect 21252 15204 21256 15260
rect 21192 15200 21256 15204
rect 8952 14716 9016 14720
rect 8952 14660 8956 14716
rect 8956 14660 9012 14716
rect 9012 14660 9016 14716
rect 8952 14656 9016 14660
rect 9032 14716 9096 14720
rect 9032 14660 9036 14716
rect 9036 14660 9092 14716
rect 9092 14660 9096 14716
rect 9032 14656 9096 14660
rect 9112 14716 9176 14720
rect 9112 14660 9116 14716
rect 9116 14660 9172 14716
rect 9172 14660 9176 14716
rect 9112 14656 9176 14660
rect 9192 14716 9256 14720
rect 9192 14660 9196 14716
rect 9196 14660 9252 14716
rect 9252 14660 9256 14716
rect 9192 14656 9256 14660
rect 16952 14716 17016 14720
rect 16952 14660 16956 14716
rect 16956 14660 17012 14716
rect 17012 14660 17016 14716
rect 16952 14656 17016 14660
rect 17032 14716 17096 14720
rect 17032 14660 17036 14716
rect 17036 14660 17092 14716
rect 17092 14660 17096 14716
rect 17032 14656 17096 14660
rect 17112 14716 17176 14720
rect 17112 14660 17116 14716
rect 17116 14660 17172 14716
rect 17172 14660 17176 14716
rect 17112 14656 17176 14660
rect 17192 14716 17256 14720
rect 17192 14660 17196 14716
rect 17196 14660 17252 14716
rect 17252 14660 17256 14716
rect 17192 14656 17256 14660
rect 60 14588 124 14652
rect 4952 14172 5016 14176
rect 4952 14116 4956 14172
rect 4956 14116 5012 14172
rect 5012 14116 5016 14172
rect 4952 14112 5016 14116
rect 5032 14172 5096 14176
rect 5032 14116 5036 14172
rect 5036 14116 5092 14172
rect 5092 14116 5096 14172
rect 5032 14112 5096 14116
rect 5112 14172 5176 14176
rect 5112 14116 5116 14172
rect 5116 14116 5172 14172
rect 5172 14116 5176 14172
rect 5112 14112 5176 14116
rect 5192 14172 5256 14176
rect 5192 14116 5196 14172
rect 5196 14116 5252 14172
rect 5252 14116 5256 14172
rect 5192 14112 5256 14116
rect 12952 14172 13016 14176
rect 12952 14116 12956 14172
rect 12956 14116 13012 14172
rect 13012 14116 13016 14172
rect 12952 14112 13016 14116
rect 13032 14172 13096 14176
rect 13032 14116 13036 14172
rect 13036 14116 13092 14172
rect 13092 14116 13096 14172
rect 13032 14112 13096 14116
rect 13112 14172 13176 14176
rect 13112 14116 13116 14172
rect 13116 14116 13172 14172
rect 13172 14116 13176 14172
rect 13112 14112 13176 14116
rect 13192 14172 13256 14176
rect 13192 14116 13196 14172
rect 13196 14116 13252 14172
rect 13252 14116 13256 14172
rect 13192 14112 13256 14116
rect 20952 14172 21016 14176
rect 20952 14116 20956 14172
rect 20956 14116 21012 14172
rect 21012 14116 21016 14172
rect 20952 14112 21016 14116
rect 21032 14172 21096 14176
rect 21032 14116 21036 14172
rect 21036 14116 21092 14172
rect 21092 14116 21096 14172
rect 21032 14112 21096 14116
rect 21112 14172 21176 14176
rect 21112 14116 21116 14172
rect 21116 14116 21172 14172
rect 21172 14116 21176 14172
rect 21112 14112 21176 14116
rect 21192 14172 21256 14176
rect 21192 14116 21196 14172
rect 21196 14116 21252 14172
rect 21252 14116 21256 14172
rect 21192 14112 21256 14116
rect 612 13908 676 13972
rect 60 13772 124 13836
rect 612 13772 676 13836
rect 8952 13628 9016 13632
rect 8952 13572 8956 13628
rect 8956 13572 9012 13628
rect 9012 13572 9016 13628
rect 8952 13568 9016 13572
rect 9032 13628 9096 13632
rect 9032 13572 9036 13628
rect 9036 13572 9092 13628
rect 9092 13572 9096 13628
rect 9032 13568 9096 13572
rect 9112 13628 9176 13632
rect 9112 13572 9116 13628
rect 9116 13572 9172 13628
rect 9172 13572 9176 13628
rect 9112 13568 9176 13572
rect 9192 13628 9256 13632
rect 9192 13572 9196 13628
rect 9196 13572 9252 13628
rect 9252 13572 9256 13628
rect 9192 13568 9256 13572
rect 16952 13628 17016 13632
rect 16952 13572 16956 13628
rect 16956 13572 17012 13628
rect 17012 13572 17016 13628
rect 16952 13568 17016 13572
rect 17032 13628 17096 13632
rect 17032 13572 17036 13628
rect 17036 13572 17092 13628
rect 17092 13572 17096 13628
rect 17032 13568 17096 13572
rect 17112 13628 17176 13632
rect 17112 13572 17116 13628
rect 17116 13572 17172 13628
rect 17172 13572 17176 13628
rect 17112 13568 17176 13572
rect 17192 13628 17256 13632
rect 17192 13572 17196 13628
rect 17196 13572 17252 13628
rect 17252 13572 17256 13628
rect 17192 13568 17256 13572
rect 4952 13084 5016 13088
rect 4952 13028 4956 13084
rect 4956 13028 5012 13084
rect 5012 13028 5016 13084
rect 4952 13024 5016 13028
rect 5032 13084 5096 13088
rect 5032 13028 5036 13084
rect 5036 13028 5092 13084
rect 5092 13028 5096 13084
rect 5032 13024 5096 13028
rect 5112 13084 5176 13088
rect 5112 13028 5116 13084
rect 5116 13028 5172 13084
rect 5172 13028 5176 13084
rect 5112 13024 5176 13028
rect 5192 13084 5256 13088
rect 5192 13028 5196 13084
rect 5196 13028 5252 13084
rect 5252 13028 5256 13084
rect 5192 13024 5256 13028
rect 12952 13084 13016 13088
rect 12952 13028 12956 13084
rect 12956 13028 13012 13084
rect 13012 13028 13016 13084
rect 12952 13024 13016 13028
rect 13032 13084 13096 13088
rect 13032 13028 13036 13084
rect 13036 13028 13092 13084
rect 13092 13028 13096 13084
rect 13032 13024 13096 13028
rect 13112 13084 13176 13088
rect 13112 13028 13116 13084
rect 13116 13028 13172 13084
rect 13172 13028 13176 13084
rect 13112 13024 13176 13028
rect 13192 13084 13256 13088
rect 13192 13028 13196 13084
rect 13196 13028 13252 13084
rect 13252 13028 13256 13084
rect 13192 13024 13256 13028
rect 20952 13084 21016 13088
rect 20952 13028 20956 13084
rect 20956 13028 21012 13084
rect 21012 13028 21016 13084
rect 20952 13024 21016 13028
rect 21032 13084 21096 13088
rect 21032 13028 21036 13084
rect 21036 13028 21092 13084
rect 21092 13028 21096 13084
rect 21032 13024 21096 13028
rect 21112 13084 21176 13088
rect 21112 13028 21116 13084
rect 21116 13028 21172 13084
rect 21172 13028 21176 13084
rect 21112 13024 21176 13028
rect 21192 13084 21256 13088
rect 21192 13028 21196 13084
rect 21196 13028 21252 13084
rect 21252 13028 21256 13084
rect 21192 13024 21256 13028
rect 8952 12540 9016 12544
rect 8952 12484 8956 12540
rect 8956 12484 9012 12540
rect 9012 12484 9016 12540
rect 8952 12480 9016 12484
rect 9032 12540 9096 12544
rect 9032 12484 9036 12540
rect 9036 12484 9092 12540
rect 9092 12484 9096 12540
rect 9032 12480 9096 12484
rect 9112 12540 9176 12544
rect 9112 12484 9116 12540
rect 9116 12484 9172 12540
rect 9172 12484 9176 12540
rect 9112 12480 9176 12484
rect 9192 12540 9256 12544
rect 9192 12484 9196 12540
rect 9196 12484 9252 12540
rect 9252 12484 9256 12540
rect 9192 12480 9256 12484
rect 16952 12540 17016 12544
rect 16952 12484 16956 12540
rect 16956 12484 17012 12540
rect 17012 12484 17016 12540
rect 16952 12480 17016 12484
rect 17032 12540 17096 12544
rect 17032 12484 17036 12540
rect 17036 12484 17092 12540
rect 17092 12484 17096 12540
rect 17032 12480 17096 12484
rect 17112 12540 17176 12544
rect 17112 12484 17116 12540
rect 17116 12484 17172 12540
rect 17172 12484 17176 12540
rect 17112 12480 17176 12484
rect 17192 12540 17256 12544
rect 17192 12484 17196 12540
rect 17196 12484 17252 12540
rect 17252 12484 17256 12540
rect 17192 12480 17256 12484
rect 4952 11996 5016 12000
rect 4952 11940 4956 11996
rect 4956 11940 5012 11996
rect 5012 11940 5016 11996
rect 4952 11936 5016 11940
rect 5032 11996 5096 12000
rect 5032 11940 5036 11996
rect 5036 11940 5092 11996
rect 5092 11940 5096 11996
rect 5032 11936 5096 11940
rect 5112 11996 5176 12000
rect 5112 11940 5116 11996
rect 5116 11940 5172 11996
rect 5172 11940 5176 11996
rect 5112 11936 5176 11940
rect 5192 11996 5256 12000
rect 5192 11940 5196 11996
rect 5196 11940 5252 11996
rect 5252 11940 5256 11996
rect 5192 11936 5256 11940
rect 12952 11996 13016 12000
rect 12952 11940 12956 11996
rect 12956 11940 13012 11996
rect 13012 11940 13016 11996
rect 12952 11936 13016 11940
rect 13032 11996 13096 12000
rect 13032 11940 13036 11996
rect 13036 11940 13092 11996
rect 13092 11940 13096 11996
rect 13032 11936 13096 11940
rect 13112 11996 13176 12000
rect 13112 11940 13116 11996
rect 13116 11940 13172 11996
rect 13172 11940 13176 11996
rect 13112 11936 13176 11940
rect 13192 11996 13256 12000
rect 13192 11940 13196 11996
rect 13196 11940 13252 11996
rect 13252 11940 13256 11996
rect 13192 11936 13256 11940
rect 20952 11996 21016 12000
rect 20952 11940 20956 11996
rect 20956 11940 21012 11996
rect 21012 11940 21016 11996
rect 20952 11936 21016 11940
rect 21032 11996 21096 12000
rect 21032 11940 21036 11996
rect 21036 11940 21092 11996
rect 21092 11940 21096 11996
rect 21032 11936 21096 11940
rect 21112 11996 21176 12000
rect 21112 11940 21116 11996
rect 21116 11940 21172 11996
rect 21172 11940 21176 11996
rect 21112 11936 21176 11940
rect 21192 11996 21256 12000
rect 21192 11940 21196 11996
rect 21196 11940 21252 11996
rect 21252 11940 21256 11996
rect 21192 11936 21256 11940
rect 8952 11452 9016 11456
rect 8952 11396 8956 11452
rect 8956 11396 9012 11452
rect 9012 11396 9016 11452
rect 8952 11392 9016 11396
rect 9032 11452 9096 11456
rect 9032 11396 9036 11452
rect 9036 11396 9092 11452
rect 9092 11396 9096 11452
rect 9032 11392 9096 11396
rect 9112 11452 9176 11456
rect 9112 11396 9116 11452
rect 9116 11396 9172 11452
rect 9172 11396 9176 11452
rect 9112 11392 9176 11396
rect 9192 11452 9256 11456
rect 9192 11396 9196 11452
rect 9196 11396 9252 11452
rect 9252 11396 9256 11452
rect 9192 11392 9256 11396
rect 16952 11452 17016 11456
rect 16952 11396 16956 11452
rect 16956 11396 17012 11452
rect 17012 11396 17016 11452
rect 16952 11392 17016 11396
rect 17032 11452 17096 11456
rect 17032 11396 17036 11452
rect 17036 11396 17092 11452
rect 17092 11396 17096 11452
rect 17032 11392 17096 11396
rect 17112 11452 17176 11456
rect 17112 11396 17116 11452
rect 17116 11396 17172 11452
rect 17172 11396 17176 11452
rect 17112 11392 17176 11396
rect 17192 11452 17256 11456
rect 17192 11396 17196 11452
rect 17196 11396 17252 11452
rect 17252 11396 17256 11452
rect 17192 11392 17256 11396
rect 4952 10908 5016 10912
rect 4952 10852 4956 10908
rect 4956 10852 5012 10908
rect 5012 10852 5016 10908
rect 4952 10848 5016 10852
rect 5032 10908 5096 10912
rect 5032 10852 5036 10908
rect 5036 10852 5092 10908
rect 5092 10852 5096 10908
rect 5032 10848 5096 10852
rect 5112 10908 5176 10912
rect 5112 10852 5116 10908
rect 5116 10852 5172 10908
rect 5172 10852 5176 10908
rect 5112 10848 5176 10852
rect 5192 10908 5256 10912
rect 5192 10852 5196 10908
rect 5196 10852 5252 10908
rect 5252 10852 5256 10908
rect 5192 10848 5256 10852
rect 12952 10908 13016 10912
rect 12952 10852 12956 10908
rect 12956 10852 13012 10908
rect 13012 10852 13016 10908
rect 12952 10848 13016 10852
rect 13032 10908 13096 10912
rect 13032 10852 13036 10908
rect 13036 10852 13092 10908
rect 13092 10852 13096 10908
rect 13032 10848 13096 10852
rect 13112 10908 13176 10912
rect 13112 10852 13116 10908
rect 13116 10852 13172 10908
rect 13172 10852 13176 10908
rect 13112 10848 13176 10852
rect 13192 10908 13256 10912
rect 13192 10852 13196 10908
rect 13196 10852 13252 10908
rect 13252 10852 13256 10908
rect 13192 10848 13256 10852
rect 20952 10908 21016 10912
rect 20952 10852 20956 10908
rect 20956 10852 21012 10908
rect 21012 10852 21016 10908
rect 20952 10848 21016 10852
rect 21032 10908 21096 10912
rect 21032 10852 21036 10908
rect 21036 10852 21092 10908
rect 21092 10852 21096 10908
rect 21032 10848 21096 10852
rect 21112 10908 21176 10912
rect 21112 10852 21116 10908
rect 21116 10852 21172 10908
rect 21172 10852 21176 10908
rect 21112 10848 21176 10852
rect 21192 10908 21256 10912
rect 21192 10852 21196 10908
rect 21196 10852 21252 10908
rect 21252 10852 21256 10908
rect 21192 10848 21256 10852
rect 8952 10364 9016 10368
rect 8952 10308 8956 10364
rect 8956 10308 9012 10364
rect 9012 10308 9016 10364
rect 8952 10304 9016 10308
rect 9032 10364 9096 10368
rect 9032 10308 9036 10364
rect 9036 10308 9092 10364
rect 9092 10308 9096 10364
rect 9032 10304 9096 10308
rect 9112 10364 9176 10368
rect 9112 10308 9116 10364
rect 9116 10308 9172 10364
rect 9172 10308 9176 10364
rect 9112 10304 9176 10308
rect 9192 10364 9256 10368
rect 9192 10308 9196 10364
rect 9196 10308 9252 10364
rect 9252 10308 9256 10364
rect 9192 10304 9256 10308
rect 16952 10364 17016 10368
rect 16952 10308 16956 10364
rect 16956 10308 17012 10364
rect 17012 10308 17016 10364
rect 16952 10304 17016 10308
rect 17032 10364 17096 10368
rect 17032 10308 17036 10364
rect 17036 10308 17092 10364
rect 17092 10308 17096 10364
rect 17032 10304 17096 10308
rect 17112 10364 17176 10368
rect 17112 10308 17116 10364
rect 17116 10308 17172 10364
rect 17172 10308 17176 10364
rect 17112 10304 17176 10308
rect 17192 10364 17256 10368
rect 17192 10308 17196 10364
rect 17196 10308 17252 10364
rect 17252 10308 17256 10364
rect 17192 10304 17256 10308
rect 4952 9820 5016 9824
rect 4952 9764 4956 9820
rect 4956 9764 5012 9820
rect 5012 9764 5016 9820
rect 4952 9760 5016 9764
rect 5032 9820 5096 9824
rect 5032 9764 5036 9820
rect 5036 9764 5092 9820
rect 5092 9764 5096 9820
rect 5032 9760 5096 9764
rect 5112 9820 5176 9824
rect 5112 9764 5116 9820
rect 5116 9764 5172 9820
rect 5172 9764 5176 9820
rect 5112 9760 5176 9764
rect 5192 9820 5256 9824
rect 5192 9764 5196 9820
rect 5196 9764 5252 9820
rect 5252 9764 5256 9820
rect 5192 9760 5256 9764
rect 12952 9820 13016 9824
rect 12952 9764 12956 9820
rect 12956 9764 13012 9820
rect 13012 9764 13016 9820
rect 12952 9760 13016 9764
rect 13032 9820 13096 9824
rect 13032 9764 13036 9820
rect 13036 9764 13092 9820
rect 13092 9764 13096 9820
rect 13032 9760 13096 9764
rect 13112 9820 13176 9824
rect 13112 9764 13116 9820
rect 13116 9764 13172 9820
rect 13172 9764 13176 9820
rect 13112 9760 13176 9764
rect 13192 9820 13256 9824
rect 13192 9764 13196 9820
rect 13196 9764 13252 9820
rect 13252 9764 13256 9820
rect 13192 9760 13256 9764
rect 20952 9820 21016 9824
rect 20952 9764 20956 9820
rect 20956 9764 21012 9820
rect 21012 9764 21016 9820
rect 20952 9760 21016 9764
rect 21032 9820 21096 9824
rect 21032 9764 21036 9820
rect 21036 9764 21092 9820
rect 21092 9764 21096 9820
rect 21032 9760 21096 9764
rect 21112 9820 21176 9824
rect 21112 9764 21116 9820
rect 21116 9764 21172 9820
rect 21172 9764 21176 9820
rect 21112 9760 21176 9764
rect 21192 9820 21256 9824
rect 21192 9764 21196 9820
rect 21196 9764 21252 9820
rect 21252 9764 21256 9820
rect 21192 9760 21256 9764
rect 8952 9276 9016 9280
rect 8952 9220 8956 9276
rect 8956 9220 9012 9276
rect 9012 9220 9016 9276
rect 8952 9216 9016 9220
rect 9032 9276 9096 9280
rect 9032 9220 9036 9276
rect 9036 9220 9092 9276
rect 9092 9220 9096 9276
rect 9032 9216 9096 9220
rect 9112 9276 9176 9280
rect 9112 9220 9116 9276
rect 9116 9220 9172 9276
rect 9172 9220 9176 9276
rect 9112 9216 9176 9220
rect 9192 9276 9256 9280
rect 9192 9220 9196 9276
rect 9196 9220 9252 9276
rect 9252 9220 9256 9276
rect 9192 9216 9256 9220
rect 16952 9276 17016 9280
rect 16952 9220 16956 9276
rect 16956 9220 17012 9276
rect 17012 9220 17016 9276
rect 16952 9216 17016 9220
rect 17032 9276 17096 9280
rect 17032 9220 17036 9276
rect 17036 9220 17092 9276
rect 17092 9220 17096 9276
rect 17032 9216 17096 9220
rect 17112 9276 17176 9280
rect 17112 9220 17116 9276
rect 17116 9220 17172 9276
rect 17172 9220 17176 9276
rect 17112 9216 17176 9220
rect 17192 9276 17256 9280
rect 17192 9220 17196 9276
rect 17196 9220 17252 9276
rect 17252 9220 17256 9276
rect 17192 9216 17256 9220
rect 4952 8732 5016 8736
rect 4952 8676 4956 8732
rect 4956 8676 5012 8732
rect 5012 8676 5016 8732
rect 4952 8672 5016 8676
rect 5032 8732 5096 8736
rect 5032 8676 5036 8732
rect 5036 8676 5092 8732
rect 5092 8676 5096 8732
rect 5032 8672 5096 8676
rect 5112 8732 5176 8736
rect 5112 8676 5116 8732
rect 5116 8676 5172 8732
rect 5172 8676 5176 8732
rect 5112 8672 5176 8676
rect 5192 8732 5256 8736
rect 5192 8676 5196 8732
rect 5196 8676 5252 8732
rect 5252 8676 5256 8732
rect 5192 8672 5256 8676
rect 12952 8732 13016 8736
rect 12952 8676 12956 8732
rect 12956 8676 13012 8732
rect 13012 8676 13016 8732
rect 12952 8672 13016 8676
rect 13032 8732 13096 8736
rect 13032 8676 13036 8732
rect 13036 8676 13092 8732
rect 13092 8676 13096 8732
rect 13032 8672 13096 8676
rect 13112 8732 13176 8736
rect 13112 8676 13116 8732
rect 13116 8676 13172 8732
rect 13172 8676 13176 8732
rect 13112 8672 13176 8676
rect 13192 8732 13256 8736
rect 13192 8676 13196 8732
rect 13196 8676 13252 8732
rect 13252 8676 13256 8732
rect 13192 8672 13256 8676
rect 20952 8732 21016 8736
rect 20952 8676 20956 8732
rect 20956 8676 21012 8732
rect 21012 8676 21016 8732
rect 20952 8672 21016 8676
rect 21032 8732 21096 8736
rect 21032 8676 21036 8732
rect 21036 8676 21092 8732
rect 21092 8676 21096 8732
rect 21032 8672 21096 8676
rect 21112 8732 21176 8736
rect 21112 8676 21116 8732
rect 21116 8676 21172 8732
rect 21172 8676 21176 8732
rect 21112 8672 21176 8676
rect 21192 8732 21256 8736
rect 21192 8676 21196 8732
rect 21196 8676 21252 8732
rect 21252 8676 21256 8732
rect 21192 8672 21256 8676
rect 8952 8188 9016 8192
rect 8952 8132 8956 8188
rect 8956 8132 9012 8188
rect 9012 8132 9016 8188
rect 8952 8128 9016 8132
rect 9032 8188 9096 8192
rect 9032 8132 9036 8188
rect 9036 8132 9092 8188
rect 9092 8132 9096 8188
rect 9032 8128 9096 8132
rect 9112 8188 9176 8192
rect 9112 8132 9116 8188
rect 9116 8132 9172 8188
rect 9172 8132 9176 8188
rect 9112 8128 9176 8132
rect 9192 8188 9256 8192
rect 9192 8132 9196 8188
rect 9196 8132 9252 8188
rect 9252 8132 9256 8188
rect 9192 8128 9256 8132
rect 16952 8188 17016 8192
rect 16952 8132 16956 8188
rect 16956 8132 17012 8188
rect 17012 8132 17016 8188
rect 16952 8128 17016 8132
rect 17032 8188 17096 8192
rect 17032 8132 17036 8188
rect 17036 8132 17092 8188
rect 17092 8132 17096 8188
rect 17032 8128 17096 8132
rect 17112 8188 17176 8192
rect 17112 8132 17116 8188
rect 17116 8132 17172 8188
rect 17172 8132 17176 8188
rect 17112 8128 17176 8132
rect 17192 8188 17256 8192
rect 17192 8132 17196 8188
rect 17196 8132 17252 8188
rect 17252 8132 17256 8188
rect 17192 8128 17256 8132
rect 4952 7644 5016 7648
rect 4952 7588 4956 7644
rect 4956 7588 5012 7644
rect 5012 7588 5016 7644
rect 4952 7584 5016 7588
rect 5032 7644 5096 7648
rect 5032 7588 5036 7644
rect 5036 7588 5092 7644
rect 5092 7588 5096 7644
rect 5032 7584 5096 7588
rect 5112 7644 5176 7648
rect 5112 7588 5116 7644
rect 5116 7588 5172 7644
rect 5172 7588 5176 7644
rect 5112 7584 5176 7588
rect 5192 7644 5256 7648
rect 5192 7588 5196 7644
rect 5196 7588 5252 7644
rect 5252 7588 5256 7644
rect 5192 7584 5256 7588
rect 12952 7644 13016 7648
rect 12952 7588 12956 7644
rect 12956 7588 13012 7644
rect 13012 7588 13016 7644
rect 12952 7584 13016 7588
rect 13032 7644 13096 7648
rect 13032 7588 13036 7644
rect 13036 7588 13092 7644
rect 13092 7588 13096 7644
rect 13032 7584 13096 7588
rect 13112 7644 13176 7648
rect 13112 7588 13116 7644
rect 13116 7588 13172 7644
rect 13172 7588 13176 7644
rect 13112 7584 13176 7588
rect 13192 7644 13256 7648
rect 13192 7588 13196 7644
rect 13196 7588 13252 7644
rect 13252 7588 13256 7644
rect 13192 7584 13256 7588
rect 20952 7644 21016 7648
rect 20952 7588 20956 7644
rect 20956 7588 21012 7644
rect 21012 7588 21016 7644
rect 20952 7584 21016 7588
rect 21032 7644 21096 7648
rect 21032 7588 21036 7644
rect 21036 7588 21092 7644
rect 21092 7588 21096 7644
rect 21032 7584 21096 7588
rect 21112 7644 21176 7648
rect 21112 7588 21116 7644
rect 21116 7588 21172 7644
rect 21172 7588 21176 7644
rect 21112 7584 21176 7588
rect 21192 7644 21256 7648
rect 21192 7588 21196 7644
rect 21196 7588 21252 7644
rect 21252 7588 21256 7644
rect 21192 7584 21256 7588
rect 8952 7100 9016 7104
rect 8952 7044 8956 7100
rect 8956 7044 9012 7100
rect 9012 7044 9016 7100
rect 8952 7040 9016 7044
rect 9032 7100 9096 7104
rect 9032 7044 9036 7100
rect 9036 7044 9092 7100
rect 9092 7044 9096 7100
rect 9032 7040 9096 7044
rect 9112 7100 9176 7104
rect 9112 7044 9116 7100
rect 9116 7044 9172 7100
rect 9172 7044 9176 7100
rect 9112 7040 9176 7044
rect 9192 7100 9256 7104
rect 9192 7044 9196 7100
rect 9196 7044 9252 7100
rect 9252 7044 9256 7100
rect 9192 7040 9256 7044
rect 16952 7100 17016 7104
rect 16952 7044 16956 7100
rect 16956 7044 17012 7100
rect 17012 7044 17016 7100
rect 16952 7040 17016 7044
rect 17032 7100 17096 7104
rect 17032 7044 17036 7100
rect 17036 7044 17092 7100
rect 17092 7044 17096 7100
rect 17032 7040 17096 7044
rect 17112 7100 17176 7104
rect 17112 7044 17116 7100
rect 17116 7044 17172 7100
rect 17172 7044 17176 7100
rect 17112 7040 17176 7044
rect 17192 7100 17256 7104
rect 17192 7044 17196 7100
rect 17196 7044 17252 7100
rect 17252 7044 17256 7100
rect 17192 7040 17256 7044
rect 4952 6556 5016 6560
rect 4952 6500 4956 6556
rect 4956 6500 5012 6556
rect 5012 6500 5016 6556
rect 4952 6496 5016 6500
rect 5032 6556 5096 6560
rect 5032 6500 5036 6556
rect 5036 6500 5092 6556
rect 5092 6500 5096 6556
rect 5032 6496 5096 6500
rect 5112 6556 5176 6560
rect 5112 6500 5116 6556
rect 5116 6500 5172 6556
rect 5172 6500 5176 6556
rect 5112 6496 5176 6500
rect 5192 6556 5256 6560
rect 5192 6500 5196 6556
rect 5196 6500 5252 6556
rect 5252 6500 5256 6556
rect 5192 6496 5256 6500
rect 12952 6556 13016 6560
rect 12952 6500 12956 6556
rect 12956 6500 13012 6556
rect 13012 6500 13016 6556
rect 12952 6496 13016 6500
rect 13032 6556 13096 6560
rect 13032 6500 13036 6556
rect 13036 6500 13092 6556
rect 13092 6500 13096 6556
rect 13032 6496 13096 6500
rect 13112 6556 13176 6560
rect 13112 6500 13116 6556
rect 13116 6500 13172 6556
rect 13172 6500 13176 6556
rect 13112 6496 13176 6500
rect 13192 6556 13256 6560
rect 13192 6500 13196 6556
rect 13196 6500 13252 6556
rect 13252 6500 13256 6556
rect 13192 6496 13256 6500
rect 20952 6556 21016 6560
rect 20952 6500 20956 6556
rect 20956 6500 21012 6556
rect 21012 6500 21016 6556
rect 20952 6496 21016 6500
rect 21032 6556 21096 6560
rect 21032 6500 21036 6556
rect 21036 6500 21092 6556
rect 21092 6500 21096 6556
rect 21032 6496 21096 6500
rect 21112 6556 21176 6560
rect 21112 6500 21116 6556
rect 21116 6500 21172 6556
rect 21172 6500 21176 6556
rect 21112 6496 21176 6500
rect 21192 6556 21256 6560
rect 21192 6500 21196 6556
rect 21196 6500 21252 6556
rect 21252 6500 21256 6556
rect 21192 6496 21256 6500
rect 60 6020 124 6084
rect 8952 6012 9016 6016
rect 8952 5956 8956 6012
rect 8956 5956 9012 6012
rect 9012 5956 9016 6012
rect 8952 5952 9016 5956
rect 9032 6012 9096 6016
rect 9032 5956 9036 6012
rect 9036 5956 9092 6012
rect 9092 5956 9096 6012
rect 9032 5952 9096 5956
rect 9112 6012 9176 6016
rect 9112 5956 9116 6012
rect 9116 5956 9172 6012
rect 9172 5956 9176 6012
rect 9112 5952 9176 5956
rect 9192 6012 9256 6016
rect 9192 5956 9196 6012
rect 9196 5956 9252 6012
rect 9252 5956 9256 6012
rect 9192 5952 9256 5956
rect 16952 6012 17016 6016
rect 16952 5956 16956 6012
rect 16956 5956 17012 6012
rect 17012 5956 17016 6012
rect 16952 5952 17016 5956
rect 17032 6012 17096 6016
rect 17032 5956 17036 6012
rect 17036 5956 17092 6012
rect 17092 5956 17096 6012
rect 17032 5952 17096 5956
rect 17112 6012 17176 6016
rect 17112 5956 17116 6012
rect 17116 5956 17172 6012
rect 17172 5956 17176 6012
rect 17112 5952 17176 5956
rect 17192 6012 17256 6016
rect 17192 5956 17196 6012
rect 17196 5956 17252 6012
rect 17252 5956 17256 6012
rect 17192 5952 17256 5956
rect 4952 5468 5016 5472
rect 4952 5412 4956 5468
rect 4956 5412 5012 5468
rect 5012 5412 5016 5468
rect 4952 5408 5016 5412
rect 5032 5468 5096 5472
rect 5032 5412 5036 5468
rect 5036 5412 5092 5468
rect 5092 5412 5096 5468
rect 5032 5408 5096 5412
rect 5112 5468 5176 5472
rect 5112 5412 5116 5468
rect 5116 5412 5172 5468
rect 5172 5412 5176 5468
rect 5112 5408 5176 5412
rect 5192 5468 5256 5472
rect 5192 5412 5196 5468
rect 5196 5412 5252 5468
rect 5252 5412 5256 5468
rect 5192 5408 5256 5412
rect 12952 5468 13016 5472
rect 12952 5412 12956 5468
rect 12956 5412 13012 5468
rect 13012 5412 13016 5468
rect 12952 5408 13016 5412
rect 13032 5468 13096 5472
rect 13032 5412 13036 5468
rect 13036 5412 13092 5468
rect 13092 5412 13096 5468
rect 13032 5408 13096 5412
rect 13112 5468 13176 5472
rect 13112 5412 13116 5468
rect 13116 5412 13172 5468
rect 13172 5412 13176 5468
rect 13112 5408 13176 5412
rect 13192 5468 13256 5472
rect 13192 5412 13196 5468
rect 13196 5412 13252 5468
rect 13252 5412 13256 5468
rect 13192 5408 13256 5412
rect 20952 5468 21016 5472
rect 20952 5412 20956 5468
rect 20956 5412 21012 5468
rect 21012 5412 21016 5468
rect 20952 5408 21016 5412
rect 21032 5468 21096 5472
rect 21032 5412 21036 5468
rect 21036 5412 21092 5468
rect 21092 5412 21096 5468
rect 21032 5408 21096 5412
rect 21112 5468 21176 5472
rect 21112 5412 21116 5468
rect 21116 5412 21172 5468
rect 21172 5412 21176 5468
rect 21112 5408 21176 5412
rect 21192 5468 21256 5472
rect 21192 5412 21196 5468
rect 21196 5412 21252 5468
rect 21252 5412 21256 5468
rect 21192 5408 21256 5412
rect 60 5068 124 5132
rect 8952 4924 9016 4928
rect 8952 4868 8956 4924
rect 8956 4868 9012 4924
rect 9012 4868 9016 4924
rect 8952 4864 9016 4868
rect 9032 4924 9096 4928
rect 9032 4868 9036 4924
rect 9036 4868 9092 4924
rect 9092 4868 9096 4924
rect 9032 4864 9096 4868
rect 9112 4924 9176 4928
rect 9112 4868 9116 4924
rect 9116 4868 9172 4924
rect 9172 4868 9176 4924
rect 9112 4864 9176 4868
rect 9192 4924 9256 4928
rect 9192 4868 9196 4924
rect 9196 4868 9252 4924
rect 9252 4868 9256 4924
rect 9192 4864 9256 4868
rect 16952 4924 17016 4928
rect 16952 4868 16956 4924
rect 16956 4868 17012 4924
rect 17012 4868 17016 4924
rect 16952 4864 17016 4868
rect 17032 4924 17096 4928
rect 17032 4868 17036 4924
rect 17036 4868 17092 4924
rect 17092 4868 17096 4924
rect 17032 4864 17096 4868
rect 17112 4924 17176 4928
rect 17112 4868 17116 4924
rect 17116 4868 17172 4924
rect 17172 4868 17176 4924
rect 17112 4864 17176 4868
rect 17192 4924 17256 4928
rect 17192 4868 17196 4924
rect 17196 4868 17252 4924
rect 17252 4868 17256 4924
rect 17192 4864 17256 4868
rect 4952 4380 5016 4384
rect 4952 4324 4956 4380
rect 4956 4324 5012 4380
rect 5012 4324 5016 4380
rect 4952 4320 5016 4324
rect 5032 4380 5096 4384
rect 5032 4324 5036 4380
rect 5036 4324 5092 4380
rect 5092 4324 5096 4380
rect 5032 4320 5096 4324
rect 5112 4380 5176 4384
rect 5112 4324 5116 4380
rect 5116 4324 5172 4380
rect 5172 4324 5176 4380
rect 5112 4320 5176 4324
rect 5192 4380 5256 4384
rect 5192 4324 5196 4380
rect 5196 4324 5252 4380
rect 5252 4324 5256 4380
rect 5192 4320 5256 4324
rect 12952 4380 13016 4384
rect 12952 4324 12956 4380
rect 12956 4324 13012 4380
rect 13012 4324 13016 4380
rect 12952 4320 13016 4324
rect 13032 4380 13096 4384
rect 13032 4324 13036 4380
rect 13036 4324 13092 4380
rect 13092 4324 13096 4380
rect 13032 4320 13096 4324
rect 13112 4380 13176 4384
rect 13112 4324 13116 4380
rect 13116 4324 13172 4380
rect 13172 4324 13176 4380
rect 13112 4320 13176 4324
rect 13192 4380 13256 4384
rect 13192 4324 13196 4380
rect 13196 4324 13252 4380
rect 13252 4324 13256 4380
rect 13192 4320 13256 4324
rect 20952 4380 21016 4384
rect 20952 4324 20956 4380
rect 20956 4324 21012 4380
rect 21012 4324 21016 4380
rect 20952 4320 21016 4324
rect 21032 4380 21096 4384
rect 21032 4324 21036 4380
rect 21036 4324 21092 4380
rect 21092 4324 21096 4380
rect 21032 4320 21096 4324
rect 21112 4380 21176 4384
rect 21112 4324 21116 4380
rect 21116 4324 21172 4380
rect 21172 4324 21176 4380
rect 21112 4320 21176 4324
rect 21192 4380 21256 4384
rect 21192 4324 21196 4380
rect 21196 4324 21252 4380
rect 21252 4324 21256 4380
rect 21192 4320 21256 4324
rect 8952 3836 9016 3840
rect 8952 3780 8956 3836
rect 8956 3780 9012 3836
rect 9012 3780 9016 3836
rect 8952 3776 9016 3780
rect 9032 3836 9096 3840
rect 9032 3780 9036 3836
rect 9036 3780 9092 3836
rect 9092 3780 9096 3836
rect 9032 3776 9096 3780
rect 9112 3836 9176 3840
rect 9112 3780 9116 3836
rect 9116 3780 9172 3836
rect 9172 3780 9176 3836
rect 9112 3776 9176 3780
rect 9192 3836 9256 3840
rect 9192 3780 9196 3836
rect 9196 3780 9252 3836
rect 9252 3780 9256 3836
rect 9192 3776 9256 3780
rect 16952 3836 17016 3840
rect 16952 3780 16956 3836
rect 16956 3780 17012 3836
rect 17012 3780 17016 3836
rect 16952 3776 17016 3780
rect 17032 3836 17096 3840
rect 17032 3780 17036 3836
rect 17036 3780 17092 3836
rect 17092 3780 17096 3836
rect 17032 3776 17096 3780
rect 17112 3836 17176 3840
rect 17112 3780 17116 3836
rect 17116 3780 17172 3836
rect 17172 3780 17176 3836
rect 17112 3776 17176 3780
rect 17192 3836 17256 3840
rect 17192 3780 17196 3836
rect 17196 3780 17252 3836
rect 17252 3780 17256 3836
rect 17192 3776 17256 3780
rect 4952 3292 5016 3296
rect 4952 3236 4956 3292
rect 4956 3236 5012 3292
rect 5012 3236 5016 3292
rect 4952 3232 5016 3236
rect 5032 3292 5096 3296
rect 5032 3236 5036 3292
rect 5036 3236 5092 3292
rect 5092 3236 5096 3292
rect 5032 3232 5096 3236
rect 5112 3292 5176 3296
rect 5112 3236 5116 3292
rect 5116 3236 5172 3292
rect 5172 3236 5176 3292
rect 5112 3232 5176 3236
rect 5192 3292 5256 3296
rect 5192 3236 5196 3292
rect 5196 3236 5252 3292
rect 5252 3236 5256 3292
rect 5192 3232 5256 3236
rect 12952 3292 13016 3296
rect 12952 3236 12956 3292
rect 12956 3236 13012 3292
rect 13012 3236 13016 3292
rect 12952 3232 13016 3236
rect 13032 3292 13096 3296
rect 13032 3236 13036 3292
rect 13036 3236 13092 3292
rect 13092 3236 13096 3292
rect 13032 3232 13096 3236
rect 13112 3292 13176 3296
rect 13112 3236 13116 3292
rect 13116 3236 13172 3292
rect 13172 3236 13176 3292
rect 13112 3232 13176 3236
rect 13192 3292 13256 3296
rect 13192 3236 13196 3292
rect 13196 3236 13252 3292
rect 13252 3236 13256 3292
rect 13192 3232 13256 3236
rect 20952 3292 21016 3296
rect 20952 3236 20956 3292
rect 20956 3236 21012 3292
rect 21012 3236 21016 3292
rect 20952 3232 21016 3236
rect 21032 3292 21096 3296
rect 21032 3236 21036 3292
rect 21036 3236 21092 3292
rect 21092 3236 21096 3292
rect 21032 3232 21096 3236
rect 21112 3292 21176 3296
rect 21112 3236 21116 3292
rect 21116 3236 21172 3292
rect 21172 3236 21176 3292
rect 21112 3232 21176 3236
rect 21192 3292 21256 3296
rect 21192 3236 21196 3292
rect 21196 3236 21252 3292
rect 21252 3236 21256 3292
rect 21192 3232 21256 3236
rect 8952 2748 9016 2752
rect 8952 2692 8956 2748
rect 8956 2692 9012 2748
rect 9012 2692 9016 2748
rect 8952 2688 9016 2692
rect 9032 2748 9096 2752
rect 9032 2692 9036 2748
rect 9036 2692 9092 2748
rect 9092 2692 9096 2748
rect 9032 2688 9096 2692
rect 9112 2748 9176 2752
rect 9112 2692 9116 2748
rect 9116 2692 9172 2748
rect 9172 2692 9176 2748
rect 9112 2688 9176 2692
rect 9192 2748 9256 2752
rect 9192 2692 9196 2748
rect 9196 2692 9252 2748
rect 9252 2692 9256 2748
rect 9192 2688 9256 2692
rect 16952 2748 17016 2752
rect 16952 2692 16956 2748
rect 16956 2692 17012 2748
rect 17012 2692 17016 2748
rect 16952 2688 17016 2692
rect 17032 2748 17096 2752
rect 17032 2692 17036 2748
rect 17036 2692 17092 2748
rect 17092 2692 17096 2748
rect 17032 2688 17096 2692
rect 17112 2748 17176 2752
rect 17112 2692 17116 2748
rect 17116 2692 17172 2748
rect 17172 2692 17176 2748
rect 17112 2688 17176 2692
rect 17192 2748 17256 2752
rect 17192 2692 17196 2748
rect 17196 2692 17252 2748
rect 17252 2692 17256 2748
rect 17192 2688 17256 2692
rect 4952 2204 5016 2208
rect 4952 2148 4956 2204
rect 4956 2148 5012 2204
rect 5012 2148 5016 2204
rect 4952 2144 5016 2148
rect 5032 2204 5096 2208
rect 5032 2148 5036 2204
rect 5036 2148 5092 2204
rect 5092 2148 5096 2204
rect 5032 2144 5096 2148
rect 5112 2204 5176 2208
rect 5112 2148 5116 2204
rect 5116 2148 5172 2204
rect 5172 2148 5176 2204
rect 5112 2144 5176 2148
rect 5192 2204 5256 2208
rect 5192 2148 5196 2204
rect 5196 2148 5252 2204
rect 5252 2148 5256 2204
rect 5192 2144 5256 2148
rect 12952 2204 13016 2208
rect 12952 2148 12956 2204
rect 12956 2148 13012 2204
rect 13012 2148 13016 2204
rect 12952 2144 13016 2148
rect 13032 2204 13096 2208
rect 13032 2148 13036 2204
rect 13036 2148 13092 2204
rect 13092 2148 13096 2204
rect 13032 2144 13096 2148
rect 13112 2204 13176 2208
rect 13112 2148 13116 2204
rect 13116 2148 13172 2204
rect 13172 2148 13176 2204
rect 13112 2144 13176 2148
rect 13192 2204 13256 2208
rect 13192 2148 13196 2204
rect 13196 2148 13252 2204
rect 13252 2148 13256 2204
rect 13192 2144 13256 2148
rect 20952 2204 21016 2208
rect 20952 2148 20956 2204
rect 20956 2148 21012 2204
rect 21012 2148 21016 2204
rect 20952 2144 21016 2148
rect 21032 2204 21096 2208
rect 21032 2148 21036 2204
rect 21036 2148 21092 2204
rect 21092 2148 21096 2204
rect 21032 2144 21096 2148
rect 21112 2204 21176 2208
rect 21112 2148 21116 2204
rect 21116 2148 21172 2204
rect 21172 2148 21176 2204
rect 21112 2144 21176 2148
rect 21192 2204 21256 2208
rect 21192 2148 21196 2204
rect 21196 2148 21252 2204
rect 21252 2148 21256 2204
rect 21192 2144 21256 2148
<< metal4 >>
rect 59 22132 125 22133
rect 59 22068 60 22132
rect 124 22068 125 22132
rect 59 22067 125 22068
rect 62 21450 122 22067
rect 4944 21792 5264 21808
rect 4944 21728 4952 21792
rect 5016 21728 5032 21792
rect 5096 21728 5112 21792
rect 5176 21728 5192 21792
rect 5256 21728 5264 21792
rect 611 21452 677 21453
rect 611 21450 612 21452
rect 62 21390 612 21450
rect 611 21388 612 21390
rect 676 21388 677 21452
rect 611 21387 677 21388
rect 4944 20704 5264 21728
rect 4944 20640 4952 20704
rect 5016 20640 5032 20704
rect 5096 20640 5112 20704
rect 5176 20640 5192 20704
rect 5256 20640 5264 20704
rect 59 20636 125 20637
rect 59 20572 60 20636
rect 124 20572 125 20636
rect 59 20571 125 20572
rect 62 20399 122 20571
rect 59 20398 125 20399
rect 59 20334 60 20398
rect 124 20334 125 20398
rect 59 20333 125 20334
rect 59 20228 125 20229
rect 59 20164 60 20228
rect 124 20164 125 20228
rect 59 20163 125 20164
rect 62 20090 122 20163
rect 611 20092 677 20093
rect 611 20090 612 20092
rect 62 20030 612 20090
rect 611 20028 612 20030
rect 676 20028 677 20092
rect 611 20027 677 20028
rect 4944 19616 5264 20640
rect 4944 19552 4952 19616
rect 5016 19552 5032 19616
rect 5096 19552 5112 19616
rect 5176 19552 5192 19616
rect 5256 19552 5264 19616
rect 59 19004 125 19005
rect 59 18940 60 19004
rect 124 18940 125 19004
rect 59 18939 125 18940
rect 62 18730 122 18939
rect 611 18732 677 18733
rect 611 18730 612 18732
rect 62 18670 612 18730
rect 611 18668 612 18670
rect 676 18668 677 18732
rect 611 18667 677 18668
rect 4944 18528 5264 19552
rect 4944 18464 4952 18528
rect 5016 18464 5032 18528
rect 5096 18464 5112 18528
rect 5176 18464 5192 18528
rect 5256 18464 5264 18528
rect 4944 17440 5264 18464
rect 4944 17376 4952 17440
rect 5016 17376 5032 17440
rect 5096 17376 5112 17440
rect 5176 17376 5192 17440
rect 5256 17376 5264 17440
rect 4944 16352 5264 17376
rect 4944 16288 4952 16352
rect 5016 16288 5032 16352
rect 5096 16288 5112 16352
rect 5176 16288 5192 16352
rect 5256 16288 5264 16352
rect 611 16012 677 16013
rect 611 16010 612 16012
rect 62 15950 612 16010
rect 62 15469 122 15950
rect 611 15948 612 15950
rect 676 15948 677 16012
rect 611 15947 677 15948
rect 59 15468 125 15469
rect 59 15404 60 15468
rect 124 15404 125 15468
rect 59 15403 125 15404
rect 4944 15264 5264 16288
rect 4944 15200 4952 15264
rect 5016 15200 5032 15264
rect 5096 15200 5112 15264
rect 5176 15200 5192 15264
rect 5256 15200 5264 15264
rect 59 14652 125 14653
rect 59 14588 60 14652
rect 124 14588 125 14652
rect 59 14587 125 14588
rect 62 13970 122 14587
rect 4944 14176 5264 15200
rect 4944 14112 4952 14176
rect 5016 14112 5032 14176
rect 5096 14112 5112 14176
rect 5176 14112 5192 14176
rect 5256 14112 5264 14176
rect 611 13972 677 13973
rect 611 13970 612 13972
rect 62 13910 612 13970
rect 611 13908 612 13910
rect 676 13908 677 13972
rect 611 13907 677 13908
rect 59 13836 125 13837
rect 59 13772 60 13836
rect 124 13834 125 13836
rect 611 13836 677 13837
rect 611 13834 612 13836
rect 124 13774 612 13834
rect 124 13772 125 13774
rect 59 13771 125 13772
rect 611 13772 612 13774
rect 676 13772 677 13836
rect 611 13771 677 13772
rect 4944 13088 5264 14112
rect 4944 13024 4952 13088
rect 5016 13024 5032 13088
rect 5096 13024 5112 13088
rect 5176 13024 5192 13088
rect 5256 13024 5264 13088
rect 4944 12000 5264 13024
rect 4944 11936 4952 12000
rect 5016 11936 5032 12000
rect 5096 11936 5112 12000
rect 5176 11936 5192 12000
rect 5256 11936 5264 12000
rect 4944 10912 5264 11936
rect 4944 10848 4952 10912
rect 5016 10848 5032 10912
rect 5096 10848 5112 10912
rect 5176 10848 5192 10912
rect 5256 10848 5264 10912
rect 4944 9824 5264 10848
rect 4944 9760 4952 9824
rect 5016 9760 5032 9824
rect 5096 9760 5112 9824
rect 5176 9760 5192 9824
rect 5256 9760 5264 9824
rect 4944 8736 5264 9760
rect 4944 8672 4952 8736
rect 5016 8672 5032 8736
rect 5096 8672 5112 8736
rect 5176 8672 5192 8736
rect 5256 8672 5264 8736
rect 4944 7648 5264 8672
rect 4944 7584 4952 7648
rect 5016 7584 5032 7648
rect 5096 7584 5112 7648
rect 5176 7584 5192 7648
rect 5256 7584 5264 7648
rect 4944 6560 5264 7584
rect 4944 6496 4952 6560
rect 5016 6496 5032 6560
rect 5096 6496 5112 6560
rect 5176 6496 5192 6560
rect 5256 6496 5264 6560
rect 59 6084 125 6085
rect 59 6020 60 6084
rect 124 6020 125 6084
rect 59 6019 125 6020
rect 62 5133 122 6019
rect 4944 5472 5264 6496
rect 4944 5408 4952 5472
rect 5016 5408 5032 5472
rect 5096 5408 5112 5472
rect 5176 5408 5192 5472
rect 5256 5408 5264 5472
rect 59 5132 125 5133
rect 59 5068 60 5132
rect 124 5068 125 5132
rect 59 5067 125 5068
rect 4944 4384 5264 5408
rect 4944 4320 4952 4384
rect 5016 4320 5032 4384
rect 5096 4320 5112 4384
rect 5176 4320 5192 4384
rect 5256 4320 5264 4384
rect 4944 3296 5264 4320
rect 4944 3232 4952 3296
rect 5016 3232 5032 3296
rect 5096 3232 5112 3296
rect 5176 3232 5192 3296
rect 5256 3232 5264 3296
rect 4944 2208 5264 3232
rect 4944 2144 4952 2208
rect 5016 2144 5032 2208
rect 5096 2144 5112 2208
rect 5176 2144 5192 2208
rect 5256 2144 5264 2208
rect 4944 2128 5264 2144
rect 8944 21248 9264 21808
rect 8944 21184 8952 21248
rect 9016 21184 9032 21248
rect 9096 21184 9112 21248
rect 9176 21184 9192 21248
rect 9256 21184 9264 21248
rect 8944 20160 9264 21184
rect 8944 20096 8952 20160
rect 9016 20096 9032 20160
rect 9096 20096 9112 20160
rect 9176 20096 9192 20160
rect 9256 20096 9264 20160
rect 8944 19072 9264 20096
rect 8944 19008 8952 19072
rect 9016 19008 9032 19072
rect 9096 19008 9112 19072
rect 9176 19008 9192 19072
rect 9256 19008 9264 19072
rect 8944 17984 9264 19008
rect 8944 17920 8952 17984
rect 9016 17920 9032 17984
rect 9096 17920 9112 17984
rect 9176 17920 9192 17984
rect 9256 17920 9264 17984
rect 8944 16896 9264 17920
rect 8944 16832 8952 16896
rect 9016 16832 9032 16896
rect 9096 16832 9112 16896
rect 9176 16832 9192 16896
rect 9256 16832 9264 16896
rect 8944 15808 9264 16832
rect 8944 15744 8952 15808
rect 9016 15744 9032 15808
rect 9096 15744 9112 15808
rect 9176 15744 9192 15808
rect 9256 15744 9264 15808
rect 8944 14720 9264 15744
rect 8944 14656 8952 14720
rect 9016 14656 9032 14720
rect 9096 14656 9112 14720
rect 9176 14656 9192 14720
rect 9256 14656 9264 14720
rect 8944 13632 9264 14656
rect 8944 13568 8952 13632
rect 9016 13568 9032 13632
rect 9096 13568 9112 13632
rect 9176 13568 9192 13632
rect 9256 13568 9264 13632
rect 8944 12544 9264 13568
rect 8944 12480 8952 12544
rect 9016 12480 9032 12544
rect 9096 12480 9112 12544
rect 9176 12480 9192 12544
rect 9256 12480 9264 12544
rect 8944 11456 9264 12480
rect 8944 11392 8952 11456
rect 9016 11392 9032 11456
rect 9096 11392 9112 11456
rect 9176 11392 9192 11456
rect 9256 11392 9264 11456
rect 8944 10368 9264 11392
rect 8944 10304 8952 10368
rect 9016 10304 9032 10368
rect 9096 10304 9112 10368
rect 9176 10304 9192 10368
rect 9256 10304 9264 10368
rect 8944 9280 9264 10304
rect 8944 9216 8952 9280
rect 9016 9216 9032 9280
rect 9096 9216 9112 9280
rect 9176 9216 9192 9280
rect 9256 9216 9264 9280
rect 8944 8192 9264 9216
rect 8944 8128 8952 8192
rect 9016 8128 9032 8192
rect 9096 8128 9112 8192
rect 9176 8128 9192 8192
rect 9256 8128 9264 8192
rect 8944 7104 9264 8128
rect 8944 7040 8952 7104
rect 9016 7040 9032 7104
rect 9096 7040 9112 7104
rect 9176 7040 9192 7104
rect 9256 7040 9264 7104
rect 8944 6016 9264 7040
rect 8944 5952 8952 6016
rect 9016 5952 9032 6016
rect 9096 5952 9112 6016
rect 9176 5952 9192 6016
rect 9256 5952 9264 6016
rect 8944 4928 9264 5952
rect 8944 4864 8952 4928
rect 9016 4864 9032 4928
rect 9096 4864 9112 4928
rect 9176 4864 9192 4928
rect 9256 4864 9264 4928
rect 8944 3840 9264 4864
rect 8944 3776 8952 3840
rect 9016 3776 9032 3840
rect 9096 3776 9112 3840
rect 9176 3776 9192 3840
rect 9256 3776 9264 3840
rect 8944 2752 9264 3776
rect 8944 2688 8952 2752
rect 9016 2688 9032 2752
rect 9096 2688 9112 2752
rect 9176 2688 9192 2752
rect 9256 2688 9264 2752
rect 8944 2128 9264 2688
rect 12944 21792 13264 21808
rect 12944 21728 12952 21792
rect 13016 21728 13032 21792
rect 13096 21728 13112 21792
rect 13176 21728 13192 21792
rect 13256 21728 13264 21792
rect 12944 20704 13264 21728
rect 12944 20640 12952 20704
rect 13016 20640 13032 20704
rect 13096 20640 13112 20704
rect 13176 20640 13192 20704
rect 13256 20640 13264 20704
rect 12944 19616 13264 20640
rect 12944 19552 12952 19616
rect 13016 19552 13032 19616
rect 13096 19552 13112 19616
rect 13176 19552 13192 19616
rect 13256 19552 13264 19616
rect 12944 18528 13264 19552
rect 12944 18464 12952 18528
rect 13016 18464 13032 18528
rect 13096 18464 13112 18528
rect 13176 18464 13192 18528
rect 13256 18464 13264 18528
rect 12944 17440 13264 18464
rect 12944 17376 12952 17440
rect 13016 17376 13032 17440
rect 13096 17376 13112 17440
rect 13176 17376 13192 17440
rect 13256 17376 13264 17440
rect 12944 16352 13264 17376
rect 12944 16288 12952 16352
rect 13016 16288 13032 16352
rect 13096 16288 13112 16352
rect 13176 16288 13192 16352
rect 13256 16288 13264 16352
rect 12944 15264 13264 16288
rect 12944 15200 12952 15264
rect 13016 15200 13032 15264
rect 13096 15200 13112 15264
rect 13176 15200 13192 15264
rect 13256 15200 13264 15264
rect 12944 14176 13264 15200
rect 12944 14112 12952 14176
rect 13016 14112 13032 14176
rect 13096 14112 13112 14176
rect 13176 14112 13192 14176
rect 13256 14112 13264 14176
rect 12944 13088 13264 14112
rect 12944 13024 12952 13088
rect 13016 13024 13032 13088
rect 13096 13024 13112 13088
rect 13176 13024 13192 13088
rect 13256 13024 13264 13088
rect 12944 12000 13264 13024
rect 12944 11936 12952 12000
rect 13016 11936 13032 12000
rect 13096 11936 13112 12000
rect 13176 11936 13192 12000
rect 13256 11936 13264 12000
rect 12944 10912 13264 11936
rect 12944 10848 12952 10912
rect 13016 10848 13032 10912
rect 13096 10848 13112 10912
rect 13176 10848 13192 10912
rect 13256 10848 13264 10912
rect 12944 9824 13264 10848
rect 12944 9760 12952 9824
rect 13016 9760 13032 9824
rect 13096 9760 13112 9824
rect 13176 9760 13192 9824
rect 13256 9760 13264 9824
rect 12944 8736 13264 9760
rect 12944 8672 12952 8736
rect 13016 8672 13032 8736
rect 13096 8672 13112 8736
rect 13176 8672 13192 8736
rect 13256 8672 13264 8736
rect 12944 7648 13264 8672
rect 12944 7584 12952 7648
rect 13016 7584 13032 7648
rect 13096 7584 13112 7648
rect 13176 7584 13192 7648
rect 13256 7584 13264 7648
rect 12944 6560 13264 7584
rect 12944 6496 12952 6560
rect 13016 6496 13032 6560
rect 13096 6496 13112 6560
rect 13176 6496 13192 6560
rect 13256 6496 13264 6560
rect 12944 5472 13264 6496
rect 12944 5408 12952 5472
rect 13016 5408 13032 5472
rect 13096 5408 13112 5472
rect 13176 5408 13192 5472
rect 13256 5408 13264 5472
rect 12944 4384 13264 5408
rect 12944 4320 12952 4384
rect 13016 4320 13032 4384
rect 13096 4320 13112 4384
rect 13176 4320 13192 4384
rect 13256 4320 13264 4384
rect 12944 3296 13264 4320
rect 12944 3232 12952 3296
rect 13016 3232 13032 3296
rect 13096 3232 13112 3296
rect 13176 3232 13192 3296
rect 13256 3232 13264 3296
rect 12944 2208 13264 3232
rect 12944 2144 12952 2208
rect 13016 2144 13032 2208
rect 13096 2144 13112 2208
rect 13176 2144 13192 2208
rect 13256 2144 13264 2208
rect 12944 2128 13264 2144
rect 16944 21248 17264 21808
rect 16944 21184 16952 21248
rect 17016 21184 17032 21248
rect 17096 21184 17112 21248
rect 17176 21184 17192 21248
rect 17256 21184 17264 21248
rect 16944 20160 17264 21184
rect 16944 20096 16952 20160
rect 17016 20096 17032 20160
rect 17096 20096 17112 20160
rect 17176 20096 17192 20160
rect 17256 20096 17264 20160
rect 16944 19072 17264 20096
rect 16944 19008 16952 19072
rect 17016 19008 17032 19072
rect 17096 19008 17112 19072
rect 17176 19008 17192 19072
rect 17256 19008 17264 19072
rect 16944 17984 17264 19008
rect 16944 17920 16952 17984
rect 17016 17920 17032 17984
rect 17096 17920 17112 17984
rect 17176 17920 17192 17984
rect 17256 17920 17264 17984
rect 16944 16896 17264 17920
rect 16944 16832 16952 16896
rect 17016 16832 17032 16896
rect 17096 16832 17112 16896
rect 17176 16832 17192 16896
rect 17256 16832 17264 16896
rect 16944 15808 17264 16832
rect 16944 15744 16952 15808
rect 17016 15744 17032 15808
rect 17096 15744 17112 15808
rect 17176 15744 17192 15808
rect 17256 15744 17264 15808
rect 16944 14720 17264 15744
rect 16944 14656 16952 14720
rect 17016 14656 17032 14720
rect 17096 14656 17112 14720
rect 17176 14656 17192 14720
rect 17256 14656 17264 14720
rect 16944 13632 17264 14656
rect 16944 13568 16952 13632
rect 17016 13568 17032 13632
rect 17096 13568 17112 13632
rect 17176 13568 17192 13632
rect 17256 13568 17264 13632
rect 16944 12544 17264 13568
rect 16944 12480 16952 12544
rect 17016 12480 17032 12544
rect 17096 12480 17112 12544
rect 17176 12480 17192 12544
rect 17256 12480 17264 12544
rect 16944 11456 17264 12480
rect 16944 11392 16952 11456
rect 17016 11392 17032 11456
rect 17096 11392 17112 11456
rect 17176 11392 17192 11456
rect 17256 11392 17264 11456
rect 16944 10368 17264 11392
rect 16944 10304 16952 10368
rect 17016 10304 17032 10368
rect 17096 10304 17112 10368
rect 17176 10304 17192 10368
rect 17256 10304 17264 10368
rect 16944 9280 17264 10304
rect 16944 9216 16952 9280
rect 17016 9216 17032 9280
rect 17096 9216 17112 9280
rect 17176 9216 17192 9280
rect 17256 9216 17264 9280
rect 16944 8192 17264 9216
rect 16944 8128 16952 8192
rect 17016 8128 17032 8192
rect 17096 8128 17112 8192
rect 17176 8128 17192 8192
rect 17256 8128 17264 8192
rect 16944 7104 17264 8128
rect 16944 7040 16952 7104
rect 17016 7040 17032 7104
rect 17096 7040 17112 7104
rect 17176 7040 17192 7104
rect 17256 7040 17264 7104
rect 16944 6016 17264 7040
rect 16944 5952 16952 6016
rect 17016 5952 17032 6016
rect 17096 5952 17112 6016
rect 17176 5952 17192 6016
rect 17256 5952 17264 6016
rect 16944 4928 17264 5952
rect 16944 4864 16952 4928
rect 17016 4864 17032 4928
rect 17096 4864 17112 4928
rect 17176 4864 17192 4928
rect 17256 4864 17264 4928
rect 16944 3840 17264 4864
rect 16944 3776 16952 3840
rect 17016 3776 17032 3840
rect 17096 3776 17112 3840
rect 17176 3776 17192 3840
rect 17256 3776 17264 3840
rect 16944 2752 17264 3776
rect 16944 2688 16952 2752
rect 17016 2688 17032 2752
rect 17096 2688 17112 2752
rect 17176 2688 17192 2752
rect 17256 2688 17264 2752
rect 16944 2128 17264 2688
rect 20944 21792 21264 21808
rect 20944 21728 20952 21792
rect 21016 21728 21032 21792
rect 21096 21728 21112 21792
rect 21176 21728 21192 21792
rect 21256 21728 21264 21792
rect 20944 20704 21264 21728
rect 20944 20640 20952 20704
rect 21016 20640 21032 20704
rect 21096 20640 21112 20704
rect 21176 20640 21192 20704
rect 21256 20640 21264 20704
rect 20944 19616 21264 20640
rect 20944 19552 20952 19616
rect 21016 19552 21032 19616
rect 21096 19552 21112 19616
rect 21176 19552 21192 19616
rect 21256 19552 21264 19616
rect 20944 18528 21264 19552
rect 20944 18464 20952 18528
rect 21016 18464 21032 18528
rect 21096 18464 21112 18528
rect 21176 18464 21192 18528
rect 21256 18464 21264 18528
rect 20944 17440 21264 18464
rect 20944 17376 20952 17440
rect 21016 17376 21032 17440
rect 21096 17376 21112 17440
rect 21176 17376 21192 17440
rect 21256 17376 21264 17440
rect 20944 16352 21264 17376
rect 20944 16288 20952 16352
rect 21016 16288 21032 16352
rect 21096 16288 21112 16352
rect 21176 16288 21192 16352
rect 21256 16288 21264 16352
rect 20944 15264 21264 16288
rect 20944 15200 20952 15264
rect 21016 15200 21032 15264
rect 21096 15200 21112 15264
rect 21176 15200 21192 15264
rect 21256 15200 21264 15264
rect 20944 14176 21264 15200
rect 20944 14112 20952 14176
rect 21016 14112 21032 14176
rect 21096 14112 21112 14176
rect 21176 14112 21192 14176
rect 21256 14112 21264 14176
rect 20944 13088 21264 14112
rect 20944 13024 20952 13088
rect 21016 13024 21032 13088
rect 21096 13024 21112 13088
rect 21176 13024 21192 13088
rect 21256 13024 21264 13088
rect 20944 12000 21264 13024
rect 20944 11936 20952 12000
rect 21016 11936 21032 12000
rect 21096 11936 21112 12000
rect 21176 11936 21192 12000
rect 21256 11936 21264 12000
rect 20944 10912 21264 11936
rect 20944 10848 20952 10912
rect 21016 10848 21032 10912
rect 21096 10848 21112 10912
rect 21176 10848 21192 10912
rect 21256 10848 21264 10912
rect 20944 9824 21264 10848
rect 20944 9760 20952 9824
rect 21016 9760 21032 9824
rect 21096 9760 21112 9824
rect 21176 9760 21192 9824
rect 21256 9760 21264 9824
rect 20944 8736 21264 9760
rect 20944 8672 20952 8736
rect 21016 8672 21032 8736
rect 21096 8672 21112 8736
rect 21176 8672 21192 8736
rect 21256 8672 21264 8736
rect 20944 7648 21264 8672
rect 20944 7584 20952 7648
rect 21016 7584 21032 7648
rect 21096 7584 21112 7648
rect 21176 7584 21192 7648
rect 21256 7584 21264 7648
rect 20944 6560 21264 7584
rect 20944 6496 20952 6560
rect 21016 6496 21032 6560
rect 21096 6496 21112 6560
rect 21176 6496 21192 6560
rect 21256 6496 21264 6560
rect 20944 5472 21264 6496
rect 20944 5408 20952 5472
rect 21016 5408 21032 5472
rect 21096 5408 21112 5472
rect 21176 5408 21192 5472
rect 21256 5408 21264 5472
rect 20944 4384 21264 5408
rect 20944 4320 20952 4384
rect 21016 4320 21032 4384
rect 21096 4320 21112 4384
rect 21176 4320 21192 4384
rect 21256 4320 21264 4384
rect 20944 3296 21264 4320
rect 20944 3232 20952 3296
rect 21016 3232 21032 3296
rect 21096 3232 21112 3296
rect 21176 3232 21192 3296
rect 21256 3232 21264 3296
rect 20944 2208 21264 3232
rect 20944 2144 20952 2208
rect 21016 2144 21032 2208
rect 21096 2144 21112 2208
rect 21176 2144 21192 2208
rect 21256 2144 21264 2208
rect 20944 2128 21264 2144
use scs8hd_nor2_4  _120_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1564 0 1 2720
box -38 -48 866 592
use scs8hd_nor2_4  _127_
timestamp 1586364061
transform 1 0 1656 0 -1 2720
box -38 -48 866 592
use scs8hd_decap_3  PHY_0 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1104 0 -1 2720
box -38 -48 314 592
use scs8hd_decap_3  PHY_2
timestamp 1586364061
transform 1 0 1104 0 1 2720
box -38 -48 314 592
use scs8hd_decap_3  FILLER_0_3
timestamp 1586364061
transform 1 0 1380 0 -1 2720
box -38 -48 314 592
use scs8hd_fill_2  FILLER_1_3 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1380 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_14
timestamp 1586364061
transform 1 0 2392 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_15
timestamp 1586364061
transform 1 0 2484 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__127__B tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 2668 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__120__B
timestamp 1586364061
transform 1 0 2576 0 1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_1_22 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 3128 0 1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_1_18
timestamp 1586364061
transform 1 0 2760 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_19
timestamp 1586364061
transform 1 0 2852 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__127__A
timestamp 1586364061
transform 1 0 3036 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__126__B
timestamp 1586364061
transform 1 0 2944 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_23
timestamp 1586364061
transform 1 0 3220 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__125__A
timestamp 1586364061
transform 1 0 3404 0 -1 2720
box -38 -48 222 592
use scs8hd_nor2_4  _125_
timestamp 1586364061
transform 1 0 4048 0 -1 2720
box -38 -48 866 592
use scs8hd_nor2_4  _130_
timestamp 1586364061
transform 1 0 3680 0 1 2720
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_72 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 3956 0 -1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__125__B
timestamp 1586364061
transform 1 0 3772 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__130__B
timestamp 1586364061
transform 1 0 3496 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_27
timestamp 1586364061
transform 1 0 3588 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_37
timestamp 1586364061
transform 1 0 4508 0 1 2720
box -38 -48 222 592
use scs8hd_buf_1  _123_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 5244 0 1 2720
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__123__A
timestamp 1586364061
transform 1 0 5704 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__124__B
timestamp 1586364061
transform 1 0 4692 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__124__A
timestamp 1586364061
transform 1 0 5060 0 1 2720
box -38 -48 222 592
use scs8hd_decap_12  FILLER_0_41 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 4876 0 -1 2720
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_1_41
timestamp 1586364061
transform 1 0 4876 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_48
timestamp 1586364061
transform 1 0 5520 0 1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_73
timestamp 1586364061
transform 1 0 6808 0 -1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_79
timestamp 1586364061
transform 1 0 6716 0 1 2720
box -38 -48 130 592
use scs8hd_decap_8  FILLER_0_53 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 5980 0 -1 2720
box -38 -48 774 592
use scs8hd_fill_1  FILLER_0_61 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 6716 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_12  FILLER_0_63
timestamp 1586364061
transform 1 0 6900 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_1_52
timestamp 1586364061
transform 1 0 5888 0 1 2720
box -38 -48 774 592
use scs8hd_fill_1  FILLER_1_60
timestamp 1586364061
transform 1 0 6624 0 1 2720
box -38 -48 130 592
use scs8hd_decap_12  FILLER_1_62
timestamp 1586364061
transform 1 0 6808 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_75
timestamp 1586364061
transform 1 0 8004 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_74
timestamp 1586364061
transform 1 0 7912 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_0_87 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 9108 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_1_86
timestamp 1586364061
transform 1 0 9016 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_74
timestamp 1586364061
transform 1 0 9660 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_12  FILLER_0_94
timestamp 1586364061
transform 1 0 9752 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_98
timestamp 1586364061
transform 1 0 10120 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_106
timestamp 1586364061
transform 1 0 10856 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_110
timestamp 1586364061
transform 1 0 11224 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_75
timestamp 1586364061
transform 1 0 12512 0 -1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_80
timestamp 1586364061
transform 1 0 12328 0 1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_118
timestamp 1586364061
transform 1 0 11960 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_0_125
timestamp 1586364061
transform 1 0 12604 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_123
timestamp 1586364061
transform 1 0 12420 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_137
timestamp 1586364061
transform 1 0 13708 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_135
timestamp 1586364061
transform 1 0 13524 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_0_149
timestamp 1586364061
transform 1 0 14812 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_1_147
timestamp 1586364061
transform 1 0 14628 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_76
timestamp 1586364061
transform 1 0 15364 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_12  FILLER_0_156
timestamp 1586364061
transform 1 0 15456 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_159
timestamp 1586364061
transform 1 0 15732 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_168
timestamp 1586364061
transform 1 0 16560 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_171
timestamp 1586364061
transform 1 0 16836 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_77
timestamp 1586364061
transform 1 0 18216 0 -1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_81
timestamp 1586364061
transform 1 0 17940 0 1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_180
timestamp 1586364061
transform 1 0 17664 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_0_187
timestamp 1586364061
transform 1 0 18308 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_184
timestamp 1586364061
transform 1 0 18032 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_199
timestamp 1586364061
transform 1 0 19412 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_196
timestamp 1586364061
transform 1 0 19136 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_78
timestamp 1586364061
transform 1 0 21068 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_211
timestamp 1586364061
transform 1 0 20516 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_0_218
timestamp 1586364061
transform 1 0 21160 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_208
timestamp 1586364061
transform 1 0 20240 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_0_230
timestamp 1586364061
transform 1 0 22264 0 -1 2720
box -38 -48 314 592
use scs8hd_decap_12  FILLER_1_220
timestamp 1586364061
transform 1 0 21344 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_3  PHY_1
timestamp 1586364061
transform -1 0 22816 0 -1 2720
box -38 -48 314 592
use scs8hd_decap_3  PHY_3
timestamp 1586364061
transform -1 0 22816 0 1 2720
box -38 -48 314 592
use scs8hd_fill_1  FILLER_1_232
timestamp 1586364061
transform 1 0 22448 0 1 2720
box -38 -48 130 592
use scs8hd_nor2_4  _126_
timestamp 1586364061
transform 1 0 1656 0 -1 3808
box -38 -48 866 592
use scs8hd_decap_3  PHY_4
timestamp 1586364061
transform 1 0 1104 0 -1 3808
box -38 -48 314 592
use scs8hd_decap_3  FILLER_2_3
timestamp 1586364061
transform 1 0 1380 0 -1 3808
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__126__A
timestamp 1586364061
transform 1 0 2668 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__119__A
timestamp 1586364061
transform 1 0 3036 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__120__A
timestamp 1586364061
transform 1 0 3404 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_15
timestamp 1586364061
transform 1 0 2484 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_19
timestamp 1586364061
transform 1 0 2852 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_23
timestamp 1586364061
transform 1 0 3220 0 -1 3808
box -38 -48 222 592
use scs8hd_nor2_4  _124_
timestamp 1586364061
transform 1 0 4048 0 -1 3808
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_82
timestamp 1586364061
transform 1 0 3956 0 -1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__130__A
timestamp 1586364061
transform 1 0 3772 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_27
timestamp 1586364061
transform 1 0 3588 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_12  FILLER_2_41
timestamp 1586364061
transform 1 0 4876 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_53
timestamp 1586364061
transform 1 0 5980 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_65
timestamp 1586364061
transform 1 0 7084 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_77
timestamp 1586364061
transform 1 0 8188 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_2_89
timestamp 1586364061
transform 1 0 9292 0 -1 3808
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_83
timestamp 1586364061
transform 1 0 9568 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_2_93
timestamp 1586364061
transform 1 0 9660 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_105
timestamp 1586364061
transform 1 0 10764 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_117
timestamp 1586364061
transform 1 0 11868 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_129
timestamp 1586364061
transform 1 0 12972 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_141
timestamp 1586364061
transform 1 0 14076 0 -1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_84
timestamp 1586364061
transform 1 0 15180 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_2_154
timestamp 1586364061
transform 1 0 15272 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_166
timestamp 1586364061
transform 1 0 16376 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_178
timestamp 1586364061
transform 1 0 17480 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_190
timestamp 1586364061
transform 1 0 18584 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_202
timestamp 1586364061
transform 1 0 19688 0 -1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_85
timestamp 1586364061
transform 1 0 20792 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_2_215
timestamp 1586364061
transform 1 0 20884 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_2_227
timestamp 1586364061
transform 1 0 21988 0 -1 3808
box -38 -48 590 592
use scs8hd_decap_3  PHY_5
timestamp 1586364061
transform -1 0 22816 0 -1 3808
box -38 -48 314 592
use scs8hd_nor2_4  _119_
timestamp 1586364061
transform 1 0 1564 0 1 3808
box -38 -48 866 592
use scs8hd_decap_3  PHY_6
timestamp 1586364061
transform 1 0 1104 0 1 3808
box -38 -48 314 592
use scs8hd_fill_2  FILLER_3_3
timestamp 1586364061
transform 1 0 1380 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__119__B
timestamp 1586364061
transform 1 0 2576 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__118__B
timestamp 1586364061
transform 1 0 2944 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__117__B
timestamp 1586364061
transform 1 0 3404 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_14
timestamp 1586364061
transform 1 0 2392 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_18
timestamp 1586364061
transform 1 0 2760 0 1 3808
box -38 -48 222 592
use scs8hd_decap_3  FILLER_3_22
timestamp 1586364061
transform 1 0 3128 0 1 3808
box -38 -48 314 592
use scs8hd_nor2_4  _117_
timestamp 1586364061
transform 1 0 3588 0 1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__110__B
timestamp 1586364061
transform 1 0 4600 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_36
timestamp 1586364061
transform 1 0 4416 0 1 3808
box -38 -48 222 592
use scs8hd_buf_1  _116_
timestamp 1586364061
transform 1 0 5152 0 1 3808
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__116__A
timestamp 1586364061
transform 1 0 5612 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__110__A
timestamp 1586364061
transform 1 0 4968 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_40
timestamp 1586364061
transform 1 0 4784 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_47
timestamp 1586364061
transform 1 0 5428 0 1 3808
box -38 -48 222 592
use scs8hd_decap_8  FILLER_3_51
timestamp 1586364061
transform 1 0 5796 0 1 3808
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_86
timestamp 1586364061
transform 1 0 6716 0 1 3808
box -38 -48 130 592
use scs8hd_fill_2  FILLER_3_59
timestamp 1586364061
transform 1 0 6532 0 1 3808
box -38 -48 222 592
use scs8hd_decap_12  FILLER_3_62
timestamp 1586364061
transform 1 0 6808 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_74
timestamp 1586364061
transform 1 0 7912 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_86
timestamp 1586364061
transform 1 0 9016 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_98
timestamp 1586364061
transform 1 0 10120 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_110
timestamp 1586364061
transform 1 0 11224 0 1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_87
timestamp 1586364061
transform 1 0 12328 0 1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_3_123
timestamp 1586364061
transform 1 0 12420 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_135
timestamp 1586364061
transform 1 0 13524 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_147
timestamp 1586364061
transform 1 0 14628 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_159
timestamp 1586364061
transform 1 0 15732 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_171
timestamp 1586364061
transform 1 0 16836 0 1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_88
timestamp 1586364061
transform 1 0 17940 0 1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_3_184
timestamp 1586364061
transform 1 0 18032 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_196
timestamp 1586364061
transform 1 0 19136 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_208
timestamp 1586364061
transform 1 0 20240 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_220
timestamp 1586364061
transform 1 0 21344 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_3  PHY_7
timestamp 1586364061
transform -1 0 22816 0 1 3808
box -38 -48 314 592
use scs8hd_fill_1  FILLER_3_232
timestamp 1586364061
transform 1 0 22448 0 1 3808
box -38 -48 130 592
use scs8hd_nor2_4  _118_
timestamp 1586364061
transform 1 0 1564 0 -1 4896
box -38 -48 866 592
use scs8hd_decap_3  PHY_8
timestamp 1586364061
transform 1 0 1104 0 -1 4896
box -38 -48 314 592
use scs8hd_fill_2  FILLER_4_3
timestamp 1586364061
transform 1 0 1380 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__111__B
timestamp 1586364061
transform 1 0 3036 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__118__A
timestamp 1586364061
transform 1 0 2576 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__113__A
timestamp 1586364061
transform 1 0 3404 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_14
timestamp 1586364061
transform 1 0 2392 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_3  FILLER_4_18
timestamp 1586364061
transform 1 0 2760 0 -1 4896
box -38 -48 314 592
use scs8hd_fill_2  FILLER_4_23
timestamp 1586364061
transform 1 0 3220 0 -1 4896
box -38 -48 222 592
use scs8hd_nor2_4  _110_
timestamp 1586364061
transform 1 0 4048 0 -1 4896
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_89
timestamp 1586364061
transform 1 0 3956 0 -1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__117__A
timestamp 1586364061
transform 1 0 3772 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_27
timestamp 1586364061
transform 1 0 3588 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_12  FILLER_4_41
timestamp 1586364061
transform 1 0 4876 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_53
timestamp 1586364061
transform 1 0 5980 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_65
timestamp 1586364061
transform 1 0 7084 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_77
timestamp 1586364061
transform 1 0 8188 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_4_89
timestamp 1586364061
transform 1 0 9292 0 -1 4896
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_90
timestamp 1586364061
transform 1 0 9568 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_4_93
timestamp 1586364061
transform 1 0 9660 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_105
timestamp 1586364061
transform 1 0 10764 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_117
timestamp 1586364061
transform 1 0 11868 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_129
timestamp 1586364061
transform 1 0 12972 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_141
timestamp 1586364061
transform 1 0 14076 0 -1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_91
timestamp 1586364061
transform 1 0 15180 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_4_154
timestamp 1586364061
transform 1 0 15272 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_166
timestamp 1586364061
transform 1 0 16376 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_178
timestamp 1586364061
transform 1 0 17480 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_190
timestamp 1586364061
transform 1 0 18584 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_202
timestamp 1586364061
transform 1 0 19688 0 -1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_92
timestamp 1586364061
transform 1 0 20792 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_4_215
timestamp 1586364061
transform 1 0 20884 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_4_227
timestamp 1586364061
transform 1 0 21988 0 -1 4896
box -38 -48 590 592
use scs8hd_decap_3  PHY_9
timestamp 1586364061
transform -1 0 22816 0 -1 4896
box -38 -48 314 592
use scs8hd_nor2_4  _113_
timestamp 1586364061
transform 1 0 1472 0 1 4896
box -38 -48 866 592
use scs8hd_decap_3  PHY_10
timestamp 1586364061
transform 1 0 1104 0 1 4896
box -38 -48 314 592
use scs8hd_fill_1  FILLER_5_3
timestamp 1586364061
transform 1 0 1380 0 1 4896
box -38 -48 130 592
use scs8hd_nor2_4  _111_
timestamp 1586364061
transform 1 0 3036 0 1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__113__B
timestamp 1586364061
transform 1 0 2484 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__112__B
timestamp 1586364061
transform 1 0 2852 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_13
timestamp 1586364061
transform 1 0 2300 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_17
timestamp 1586364061
transform 1 0 2668 0 1 4896
box -38 -48 222 592
use scs8hd_buf_1  _109_
timestamp 1586364061
transform 1 0 4600 0 1 4896
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__132__B
timestamp 1586364061
transform 1 0 4048 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__132__A
timestamp 1586364061
transform 1 0 4416 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_30
timestamp 1586364061
transform 1 0 3864 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_34
timestamp 1586364061
transform 1 0 4232 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__109__A
timestamp 1586364061
transform 1 0 5060 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_41
timestamp 1586364061
transform 1 0 4876 0 1 4896
box -38 -48 222 592
use scs8hd_decap_12  FILLER_5_45
timestamp 1586364061
transform 1 0 5244 0 1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_93
timestamp 1586364061
transform 1 0 6716 0 1 4896
box -38 -48 130 592
use scs8hd_decap_4  FILLER_5_57
timestamp 1586364061
transform 1 0 6348 0 1 4896
box -38 -48 406 592
use scs8hd_decap_12  FILLER_5_62
timestamp 1586364061
transform 1 0 6808 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_74
timestamp 1586364061
transform 1 0 7912 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_86
timestamp 1586364061
transform 1 0 9016 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_98
timestamp 1586364061
transform 1 0 10120 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_110
timestamp 1586364061
transform 1 0 11224 0 1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_94
timestamp 1586364061
transform 1 0 12328 0 1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_5_123
timestamp 1586364061
transform 1 0 12420 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_135
timestamp 1586364061
transform 1 0 13524 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_147
timestamp 1586364061
transform 1 0 14628 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_159
timestamp 1586364061
transform 1 0 15732 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_171
timestamp 1586364061
transform 1 0 16836 0 1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_95
timestamp 1586364061
transform 1 0 17940 0 1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_5_184
timestamp 1586364061
transform 1 0 18032 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_196
timestamp 1586364061
transform 1 0 19136 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_208
timestamp 1586364061
transform 1 0 20240 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_220
timestamp 1586364061
transform 1 0 21344 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_3  PHY_11
timestamp 1586364061
transform -1 0 22816 0 1 4896
box -38 -48 314 592
use scs8hd_fill_1  FILLER_5_232
timestamp 1586364061
transform 1 0 22448 0 1 4896
box -38 -48 130 592
use scs8hd_nor2_4  _104_
timestamp 1586364061
transform 1 0 1380 0 1 5984
box -38 -48 866 592
use scs8hd_nor2_4  _112_
timestamp 1586364061
transform 1 0 1564 0 -1 5984
box -38 -48 866 592
use scs8hd_decap_3  PHY_12
timestamp 1586364061
transform 1 0 1104 0 -1 5984
box -38 -48 314 592
use scs8hd_decap_3  PHY_14
timestamp 1586364061
transform 1 0 1104 0 1 5984
box -38 -48 314 592
use scs8hd_fill_2  FILLER_6_3
timestamp 1586364061
transform 1 0 1380 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_12
timestamp 1586364061
transform 1 0 2208 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_16
timestamp 1586364061
transform 1 0 2576 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_14
timestamp 1586364061
transform 1 0 2392 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__112__A
timestamp 1586364061
transform 1 0 2576 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__104__B
timestamp 1586364061
transform 1 0 2392 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_20
timestamp 1586364061
transform 1 0 2944 0 1 5984
box -38 -48 222 592
use scs8hd_decap_3  FILLER_6_18
timestamp 1586364061
transform 1 0 2760 0 -1 5984
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__103__B
timestamp 1586364061
transform 1 0 2760 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_24
timestamp 1586364061
transform 1 0 3312 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_23
timestamp 1586364061
transform 1 0 3220 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__111__A
timestamp 1586364061
transform 1 0 3036 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__136__A
timestamp 1586364061
transform 1 0 3128 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__104__A
timestamp 1586364061
transform 1 0 3404 0 -1 5984
box -38 -48 222 592
use scs8hd_nor2_4  _101_
timestamp 1586364061
transform 1 0 3680 0 1 5984
box -38 -48 866 592
use scs8hd_nor2_4  _132_
timestamp 1586364061
transform 1 0 4048 0 -1 5984
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_96
timestamp 1586364061
transform 1 0 3956 0 -1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__101__B
timestamp 1586364061
transform 1 0 3496 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__101__A
timestamp 1586364061
transform 1 0 3772 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_27
timestamp 1586364061
transform 1 0 3588 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_37
timestamp 1586364061
transform 1 0 4508 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__129__A
timestamp 1586364061
transform 1 0 5612 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__136__B
timestamp 1586364061
transform 1 0 4692 0 1 5984
box -38 -48 222 592
use scs8hd_decap_12  FILLER_6_41
timestamp 1586364061
transform 1 0 4876 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_7_41
timestamp 1586364061
transform 1 0 4876 0 1 5984
box -38 -48 774 592
use scs8hd_decap_8  FILLER_7_51
timestamp 1586364061
transform 1 0 5796 0 1 5984
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_100
timestamp 1586364061
transform 1 0 6716 0 1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_53
timestamp 1586364061
transform 1 0 5980 0 -1 5984
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_7_59
timestamp 1586364061
transform 1 0 6532 0 1 5984
box -38 -48 222 592
use scs8hd_decap_12  FILLER_7_62
timestamp 1586364061
transform 1 0 6808 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_65
timestamp 1586364061
transform 1 0 7084 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_77
timestamp 1586364061
transform 1 0 8188 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_74
timestamp 1586364061
transform 1 0 7912 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_6_89
timestamp 1586364061
transform 1 0 9292 0 -1 5984
box -38 -48 314 592
use scs8hd_decap_12  FILLER_7_86
timestamp 1586364061
transform 1 0 9016 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_97
timestamp 1586364061
transform 1 0 9568 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_93
timestamp 1586364061
transform 1 0 9660 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_98
timestamp 1586364061
transform 1 0 10120 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_105
timestamp 1586364061
transform 1 0 10764 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_110
timestamp 1586364061
transform 1 0 11224 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_101
timestamp 1586364061
transform 1 0 12328 0 1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_117
timestamp 1586364061
transform 1 0 11868 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_123
timestamp 1586364061
transform 1 0 12420 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_129
timestamp 1586364061
transform 1 0 12972 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_141
timestamp 1586364061
transform 1 0 14076 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_135
timestamp 1586364061
transform 1 0 13524 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_98
timestamp 1586364061
transform 1 0 15180 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_154
timestamp 1586364061
transform 1 0 15272 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_147
timestamp 1586364061
transform 1 0 14628 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_166
timestamp 1586364061
transform 1 0 16376 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_159
timestamp 1586364061
transform 1 0 15732 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_178
timestamp 1586364061
transform 1 0 17480 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_171
timestamp 1586364061
transform 1 0 16836 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_102
timestamp 1586364061
transform 1 0 17940 0 1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_190
timestamp 1586364061
transform 1 0 18584 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_184
timestamp 1586364061
transform 1 0 18032 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_202
timestamp 1586364061
transform 1 0 19688 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_196
timestamp 1586364061
transform 1 0 19136 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_99
timestamp 1586364061
transform 1 0 20792 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_215
timestamp 1586364061
transform 1 0 20884 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_208
timestamp 1586364061
transform 1 0 20240 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_6_227
timestamp 1586364061
transform 1 0 21988 0 -1 5984
box -38 -48 590 592
use scs8hd_decap_12  FILLER_7_220
timestamp 1586364061
transform 1 0 21344 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_3  PHY_13
timestamp 1586364061
transform -1 0 22816 0 -1 5984
box -38 -48 314 592
use scs8hd_decap_3  PHY_15
timestamp 1586364061
transform -1 0 22816 0 1 5984
box -38 -48 314 592
use scs8hd_fill_1  FILLER_7_232
timestamp 1586364061
transform 1 0 22448 0 1 5984
box -38 -48 130 592
use scs8hd_nor2_4  _103_
timestamp 1586364061
transform 1 0 1380 0 -1 7072
box -38 -48 866 592
use scs8hd_decap_3  PHY_16
timestamp 1586364061
transform 1 0 1104 0 -1 7072
box -38 -48 314 592
use scs8hd_fill_2  FILLER_8_12
timestamp 1586364061
transform 1 0 2208 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__134__B
timestamp 1586364061
transform 1 0 3312 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__102__A
timestamp 1586364061
transform 1 0 2392 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__103__A
timestamp 1586364061
transform 1 0 2760 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_16
timestamp 1586364061
transform 1 0 2576 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_8_20
timestamp 1586364061
transform 1 0 2944 0 -1 7072
box -38 -48 406 592
use scs8hd_nor2_4  _136_
timestamp 1586364061
transform 1 0 4048 0 -1 7072
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_103
timestamp 1586364061
transform 1 0 3956 0 -1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__134__A
timestamp 1586364061
transform 1 0 3680 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_26
timestamp 1586364061
transform 1 0 3496 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_1  FILLER_8_30
timestamp 1586364061
transform 1 0 3864 0 -1 7072
box -38 -48 130 592
use scs8hd_buf_1  _129_
timestamp 1586364061
transform 1 0 5612 0 -1 7072
box -38 -48 314 592
use scs8hd_decap_8  FILLER_8_41
timestamp 1586364061
transform 1 0 4876 0 -1 7072
box -38 -48 774 592
use scs8hd_decap_12  FILLER_8_52
timestamp 1586364061
transform 1 0 5888 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_64
timestamp 1586364061
transform 1 0 6992 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_76
timestamp 1586364061
transform 1 0 8096 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_8_88
timestamp 1586364061
transform 1 0 9200 0 -1 7072
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_104
timestamp 1586364061
transform 1 0 9568 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_8_93
timestamp 1586364061
transform 1 0 9660 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_105
timestamp 1586364061
transform 1 0 10764 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_117
timestamp 1586364061
transform 1 0 11868 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_129
timestamp 1586364061
transform 1 0 12972 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_141
timestamp 1586364061
transform 1 0 14076 0 -1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_105
timestamp 1586364061
transform 1 0 15180 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_8_154
timestamp 1586364061
transform 1 0 15272 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_166
timestamp 1586364061
transform 1 0 16376 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_178
timestamp 1586364061
transform 1 0 17480 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_190
timestamp 1586364061
transform 1 0 18584 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_202
timestamp 1586364061
transform 1 0 19688 0 -1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_106
timestamp 1586364061
transform 1 0 20792 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_8_215
timestamp 1586364061
transform 1 0 20884 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_8_227
timestamp 1586364061
transform 1 0 21988 0 -1 7072
box -38 -48 590 592
use scs8hd_decap_3  PHY_17
timestamp 1586364061
transform -1 0 22816 0 -1 7072
box -38 -48 314 592
use scs8hd_nor2_4  _102_
timestamp 1586364061
transform 1 0 1472 0 1 7072
box -38 -48 866 592
use scs8hd_decap_3  PHY_18
timestamp 1586364061
transform 1 0 1104 0 1 7072
box -38 -48 314 592
use scs8hd_fill_1  FILLER_9_3
timestamp 1586364061
transform 1 0 1380 0 1 7072
box -38 -48 130 592
use scs8hd_nor2_4  _134_
timestamp 1586364061
transform 1 0 3312 0 1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__098__B
timestamp 1586364061
transform 1 0 2484 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__102__B
timestamp 1586364061
transform 1 0 2852 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_13
timestamp 1586364061
transform 1 0 2300 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_17
timestamp 1586364061
transform 1 0 2668 0 1 7072
box -38 -48 222 592
use scs8hd_decap_3  FILLER_9_21
timestamp 1586364061
transform 1 0 3036 0 1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__088__A
timestamp 1586364061
transform 1 0 4324 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_33
timestamp 1586364061
transform 1 0 4140 0 1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_9_37
timestamp 1586364061
transform 1 0 4508 0 1 7072
box -38 -48 406 592
use scs8hd_buf_1  _100_
timestamp 1586364061
transform 1 0 5428 0 1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__100__A
timestamp 1586364061
transform 1 0 5244 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__092__A
timestamp 1586364061
transform 1 0 4876 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_43
timestamp 1586364061
transform 1 0 5060 0 1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_9_50
timestamp 1586364061
transform 1 0 5704 0 1 7072
box -38 -48 406 592
use scs8hd_inv_8  _069_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 6808 0 1 7072
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_107
timestamp 1586364061
transform 1 0 6716 0 1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__069__A
timestamp 1586364061
transform 1 0 6532 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__094__A
timestamp 1586364061
transform 1 0 6072 0 1 7072
box -38 -48 222 592
use scs8hd_decap_3  FILLER_9_56
timestamp 1586364061
transform 1 0 6256 0 1 7072
box -38 -48 314 592
use scs8hd_decap_12  FILLER_9_71
timestamp 1586364061
transform 1 0 7636 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_83
timestamp 1586364061
transform 1 0 8740 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_95
timestamp 1586364061
transform 1 0 9844 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_107
timestamp 1586364061
transform 1 0 10948 0 1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_108
timestamp 1586364061
transform 1 0 12328 0 1 7072
box -38 -48 130 592
use scs8hd_decap_3  FILLER_9_119
timestamp 1586364061
transform 1 0 12052 0 1 7072
box -38 -48 314 592
use scs8hd_decap_12  FILLER_9_123
timestamp 1586364061
transform 1 0 12420 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_135
timestamp 1586364061
transform 1 0 13524 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_147
timestamp 1586364061
transform 1 0 14628 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_159
timestamp 1586364061
transform 1 0 15732 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_171
timestamp 1586364061
transform 1 0 16836 0 1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_109
timestamp 1586364061
transform 1 0 17940 0 1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_9_184
timestamp 1586364061
transform 1 0 18032 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_196
timestamp 1586364061
transform 1 0 19136 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_208
timestamp 1586364061
transform 1 0 20240 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_220
timestamp 1586364061
transform 1 0 21344 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_3  PHY_19
timestamp 1586364061
transform -1 0 22816 0 1 7072
box -38 -48 314 592
use scs8hd_fill_1  FILLER_9_232
timestamp 1586364061
transform 1 0 22448 0 1 7072
box -38 -48 130 592
use scs8hd_nor2_4  _098_
timestamp 1586364061
transform 1 0 1472 0 -1 8160
box -38 -48 866 592
use scs8hd_decap_3  PHY_20
timestamp 1586364061
transform 1 0 1104 0 -1 8160
box -38 -48 314 592
use scs8hd_fill_1  FILLER_10_3
timestamp 1586364061
transform 1 0 1380 0 -1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__095__B
timestamp 1586364061
transform 1 0 3312 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__096__A
timestamp 1586364061
transform 1 0 2484 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__097__A
timestamp 1586364061
transform 1 0 2852 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_13
timestamp 1586364061
transform 1 0 2300 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_17
timestamp 1586364061
transform 1 0 2668 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_3  FILLER_10_21
timestamp 1586364061
transform 1 0 3036 0 -1 8160
box -38 -48 314 592
use scs8hd_buf_1  _088_
timestamp 1586364061
transform 1 0 4048 0 -1 8160
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_110
timestamp 1586364061
transform 1 0 3956 0 -1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__084__A
timestamp 1586364061
transform 1 0 4508 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__098__A
timestamp 1586364061
transform 1 0 3680 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_26
timestamp 1586364061
transform 1 0 3496 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_1  FILLER_10_30
timestamp 1586364061
transform 1 0 3864 0 -1 8160
box -38 -48 130 592
use scs8hd_fill_2  FILLER_10_35
timestamp 1586364061
transform 1 0 4324 0 -1 8160
box -38 -48 222 592
use scs8hd_buf_1  _092_
timestamp 1586364061
transform 1 0 5060 0 -1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__075__B
timestamp 1586364061
transform 1 0 5520 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__091__A
timestamp 1586364061
transform 1 0 4876 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_39
timestamp 1586364061
transform 1 0 4692 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_46
timestamp 1586364061
transform 1 0 5336 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_10_50
timestamp 1586364061
transform 1 0 5704 0 -1 8160
box -38 -48 406 592
use scs8hd_buf_1  _094_
timestamp 1586364061
transform 1 0 6072 0 -1 8160
box -38 -48 314 592
use scs8hd_decap_12  FILLER_10_57
timestamp 1586364061
transform 1 0 6348 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_69
timestamp 1586364061
transform 1 0 7452 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_10_81
timestamp 1586364061
transform 1 0 8556 0 -1 8160
box -38 -48 774 592
use scs8hd_decap_3  FILLER_10_89
timestamp 1586364061
transform 1 0 9292 0 -1 8160
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_111
timestamp 1586364061
transform 1 0 9568 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_12  FILLER_10_93
timestamp 1586364061
transform 1 0 9660 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_105
timestamp 1586364061
transform 1 0 10764 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_117
timestamp 1586364061
transform 1 0 11868 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_129
timestamp 1586364061
transform 1 0 12972 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_141
timestamp 1586364061
transform 1 0 14076 0 -1 8160
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_112
timestamp 1586364061
transform 1 0 15180 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_12  FILLER_10_154
timestamp 1586364061
transform 1 0 15272 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_166
timestamp 1586364061
transform 1 0 16376 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_178
timestamp 1586364061
transform 1 0 17480 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_190
timestamp 1586364061
transform 1 0 18584 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_202
timestamp 1586364061
transform 1 0 19688 0 -1 8160
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_113
timestamp 1586364061
transform 1 0 20792 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_12  FILLER_10_215
timestamp 1586364061
transform 1 0 20884 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_10_227
timestamp 1586364061
transform 1 0 21988 0 -1 8160
box -38 -48 590 592
use scs8hd_decap_3  PHY_21
timestamp 1586364061
transform -1 0 22816 0 -1 8160
box -38 -48 314 592
use scs8hd_nor2_4  _097_
timestamp 1586364061
transform 1 0 1472 0 1 8160
box -38 -48 866 592
use scs8hd_decap_3  PHY_22
timestamp 1586364061
transform 1 0 1104 0 1 8160
box -38 -48 314 592
use scs8hd_fill_1  FILLER_11_3
timestamp 1586364061
transform 1 0 1380 0 1 8160
box -38 -48 130 592
use scs8hd_nor2_4  _095_
timestamp 1586364061
transform 1 0 3312 0 1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__097__B
timestamp 1586364061
transform 1 0 2484 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__096__B
timestamp 1586364061
transform 1 0 2852 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_13
timestamp 1586364061
transform 1 0 2300 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_17
timestamp 1586364061
transform 1 0 2668 0 1 8160
box -38 -48 222 592
use scs8hd_decap_3  FILLER_11_21
timestamp 1586364061
transform 1 0 3036 0 1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__075__A
timestamp 1586364061
transform 1 0 4324 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_33
timestamp 1586364061
transform 1 0 4140 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_37
timestamp 1586364061
transform 1 0 4508 0 1 8160
box -38 -48 222 592
use scs8hd_inv_8  _070_
timestamp 1586364061
transform 1 0 4876 0 1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__070__A
timestamp 1586364061
transform 1 0 4692 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_50
timestamp 1586364061
transform 1 0 5704 0 1 8160
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_114
timestamp 1586364061
transform 1 0 6716 0 1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__075__C
timestamp 1586364061
transform 1 0 5888 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__095__A
timestamp 1586364061
transform 1 0 6256 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_54
timestamp 1586364061
transform 1 0 6072 0 1 8160
box -38 -48 222 592
use scs8hd_decap_3  FILLER_11_58
timestamp 1586364061
transform 1 0 6440 0 1 8160
box -38 -48 314 592
use scs8hd_decap_12  FILLER_11_62
timestamp 1586364061
transform 1 0 6808 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_74
timestamp 1586364061
transform 1 0 7912 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_86
timestamp 1586364061
transform 1 0 9016 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_98
timestamp 1586364061
transform 1 0 10120 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_110
timestamp 1586364061
transform 1 0 11224 0 1 8160
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_115
timestamp 1586364061
transform 1 0 12328 0 1 8160
box -38 -48 130 592
use scs8hd_decap_12  FILLER_11_123
timestamp 1586364061
transform 1 0 12420 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_135
timestamp 1586364061
transform 1 0 13524 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_147
timestamp 1586364061
transform 1 0 14628 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_159
timestamp 1586364061
transform 1 0 15732 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_171
timestamp 1586364061
transform 1 0 16836 0 1 8160
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_116
timestamp 1586364061
transform 1 0 17940 0 1 8160
box -38 -48 130 592
use scs8hd_decap_12  FILLER_11_184
timestamp 1586364061
transform 1 0 18032 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_196
timestamp 1586364061
transform 1 0 19136 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_208
timestamp 1586364061
transform 1 0 20240 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_220
timestamp 1586364061
transform 1 0 21344 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_3  PHY_23
timestamp 1586364061
transform -1 0 22816 0 1 8160
box -38 -48 314 592
use scs8hd_fill_1  FILLER_11_232
timestamp 1586364061
transform 1 0 22448 0 1 8160
box -38 -48 130 592
use scs8hd_nor2_4  _096_
timestamp 1586364061
transform 1 0 1564 0 -1 9248
box -38 -48 866 592
use scs8hd_decap_3  PHY_24
timestamp 1586364061
transform 1 0 1104 0 -1 9248
box -38 -48 314 592
use scs8hd_fill_2  FILLER_12_3
timestamp 1586364061
transform 1 0 1380 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__087__B
timestamp 1586364061
transform 1 0 2576 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__085__A
timestamp 1586364061
transform 1 0 2944 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__085__B
timestamp 1586364061
transform 1 0 3312 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_14
timestamp 1586364061
transform 1 0 2392 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_18
timestamp 1586364061
transform 1 0 2760 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_22
timestamp 1586364061
transform 1 0 3128 0 -1 9248
box -38 -48 222 592
use scs8hd_buf_1  _084_
timestamp 1586364061
transform 1 0 4048 0 -1 9248
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_117
timestamp 1586364061
transform 1 0 3956 0 -1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__072__A
timestamp 1586364061
transform 1 0 4508 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__087__A
timestamp 1586364061
transform 1 0 3680 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_26
timestamp 1586364061
transform 1 0 3496 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_1  FILLER_12_30
timestamp 1586364061
transform 1 0 3864 0 -1 9248
box -38 -48 130 592
use scs8hd_fill_2  FILLER_12_35
timestamp 1586364061
transform 1 0 4324 0 -1 9248
box -38 -48 222 592
use scs8hd_or3_4  _075_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 5152 0 -1 9248
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__083__C
timestamp 1586364061
transform 1 0 4968 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_3  FILLER_12_39
timestamp 1586364061
transform 1 0 4692 0 -1 9248
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__071__C
timestamp 1586364061
transform 1 0 6624 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_6  FILLER_12_53
timestamp 1586364061
transform 1 0 5980 0 -1 9248
box -38 -48 590 592
use scs8hd_fill_1  FILLER_12_59
timestamp 1586364061
transform 1 0 6532 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_12  FILLER_12_62
timestamp 1586364061
transform 1 0 6808 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_74
timestamp 1586364061
transform 1 0 7912 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_12_86
timestamp 1586364061
transform 1 0 9016 0 -1 9248
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_118
timestamp 1586364061
transform 1 0 9568 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_12  FILLER_12_93
timestamp 1586364061
transform 1 0 9660 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_105
timestamp 1586364061
transform 1 0 10764 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_117
timestamp 1586364061
transform 1 0 11868 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_129
timestamp 1586364061
transform 1 0 12972 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_141
timestamp 1586364061
transform 1 0 14076 0 -1 9248
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_119
timestamp 1586364061
transform 1 0 15180 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_12  FILLER_12_154
timestamp 1586364061
transform 1 0 15272 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_166
timestamp 1586364061
transform 1 0 16376 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_178
timestamp 1586364061
transform 1 0 17480 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_190
timestamp 1586364061
transform 1 0 18584 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_202
timestamp 1586364061
transform 1 0 19688 0 -1 9248
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_120
timestamp 1586364061
transform 1 0 20792 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_12  FILLER_12_215
timestamp 1586364061
transform 1 0 20884 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_12_227
timestamp 1586364061
transform 1 0 21988 0 -1 9248
box -38 -48 590 592
use scs8hd_decap_3  PHY_25
timestamp 1586364061
transform -1 0 22816 0 -1 9248
box -38 -48 314 592
use scs8hd_buf_1  _076_
timestamp 1586364061
transform 1 0 1380 0 -1 10336
box -38 -48 314 592
use scs8hd_nor2_4  _087_
timestamp 1586364061
transform 1 0 1656 0 1 9248
box -38 -48 866 592
use scs8hd_decap_3  PHY_26
timestamp 1586364061
transform 1 0 1104 0 1 9248
box -38 -48 314 592
use scs8hd_decap_3  PHY_28
timestamp 1586364061
transform 1 0 1104 0 -1 10336
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__080__A
timestamp 1586364061
transform 1 0 1840 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__077__B
timestamp 1586364061
transform 1 0 2208 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_3  FILLER_13_3
timestamp 1586364061
transform 1 0 1380 0 1 9248
box -38 -48 314 592
use scs8hd_fill_2  FILLER_14_6
timestamp 1586364061
transform 1 0 1656 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_10
timestamp 1586364061
transform 1 0 2024 0 -1 10336
box -38 -48 222 592
use scs8hd_nor2_4  _085_
timestamp 1586364061
transform 1 0 2392 0 -1 10336
box -38 -48 866 592
use scs8hd_nor2_4  _091_
timestamp 1586364061
transform 1 0 3220 0 1 9248
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__076__A
timestamp 1586364061
transform 1 0 2668 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__091__B
timestamp 1586364061
transform 1 0 3036 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__089__B
timestamp 1586364061
transform 1 0 3404 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_15
timestamp 1586364061
transform 1 0 2484 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_19
timestamp 1586364061
transform 1 0 2852 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_23
timestamp 1586364061
transform 1 0 3220 0 -1 10336
box -38 -48 222 592
use scs8hd_buf_1  _072_
timestamp 1586364061
transform 1 0 4048 0 -1 10336
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_124
timestamp 1586364061
transform 1 0 3956 0 -1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__078__C
timestamp 1586364061
transform 1 0 4508 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__141__A
timestamp 1586364061
transform 1 0 3772 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__089__A
timestamp 1586364061
transform 1 0 4508 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_13_32
timestamp 1586364061
transform 1 0 4048 0 1 9248
box -38 -48 406 592
use scs8hd_fill_1  FILLER_13_36
timestamp 1586364061
transform 1 0 4416 0 1 9248
box -38 -48 130 592
use scs8hd_fill_2  FILLER_14_27
timestamp 1586364061
transform 1 0 3588 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_35
timestamp 1586364061
transform 1 0 4324 0 -1 10336
box -38 -48 222 592
use scs8hd_or3_4  _078_
timestamp 1586364061
transform 1 0 5060 0 -1 10336
box -38 -48 866 592
use scs8hd_or3_4  _083_
timestamp 1586364061
transform 1 0 5060 0 1 9248
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__078__B
timestamp 1586364061
transform 1 0 4876 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__083__B
timestamp 1586364061
transform 1 0 4876 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_39
timestamp 1586364061
transform 1 0 4692 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_39
timestamp 1586364061
transform 1 0 4692 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_56
timestamp 1586364061
transform 1 0 6256 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_52
timestamp 1586364061
transform 1 0 5888 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_56
timestamp 1586364061
transform 1 0 6256 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_52
timestamp 1586364061
transform 1 0 5888 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__083__A
timestamp 1586364061
transform 1 0 6072 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__067__C
timestamp 1586364061
transform 1 0 6072 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_62
timestamp 1586364061
transform 1 0 6808 0 1 9248
box -38 -48 222 592
use scs8hd_fill_1  FILLER_13_60
timestamp 1586364061
transform 1 0 6624 0 1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__078__A
timestamp 1586364061
transform 1 0 6440 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__067__D
timestamp 1586364061
transform 1 0 6440 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__071__B
timestamp 1586364061
transform 1 0 6992 0 1 9248
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_121
timestamp 1586364061
transform 1 0 6716 0 1 9248
box -38 -48 130 592
use scs8hd_or3_4  _071_
timestamp 1586364061
transform 1 0 6624 0 -1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__071__A
timestamp 1586364061
transform 1 0 7360 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_66
timestamp 1586364061
transform 1 0 7176 0 1 9248
box -38 -48 222 592
use scs8hd_decap_12  FILLER_13_70
timestamp 1586364061
transform 1 0 7544 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_69
timestamp 1586364061
transform 1 0 7452 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_82
timestamp 1586364061
transform 1 0 8648 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_14_81
timestamp 1586364061
transform 1 0 8556 0 -1 10336
box -38 -48 774 592
use scs8hd_decap_3  FILLER_14_89
timestamp 1586364061
transform 1 0 9292 0 -1 10336
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_125
timestamp 1586364061
transform 1 0 9568 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_12  FILLER_13_94
timestamp 1586364061
transform 1 0 9752 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_93
timestamp 1586364061
transform 1 0 9660 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_106
timestamp 1586364061
transform 1 0 10856 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_105
timestamp 1586364061
transform 1 0 10764 0 -1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_122
timestamp 1586364061
transform 1 0 12328 0 1 9248
box -38 -48 130 592
use scs8hd_decap_4  FILLER_13_118
timestamp 1586364061
transform 1 0 11960 0 1 9248
box -38 -48 406 592
use scs8hd_decap_12  FILLER_13_123
timestamp 1586364061
transform 1 0 12420 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_117
timestamp 1586364061
transform 1 0 11868 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_135
timestamp 1586364061
transform 1 0 13524 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_129
timestamp 1586364061
transform 1 0 12972 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_141
timestamp 1586364061
transform 1 0 14076 0 -1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_126
timestamp 1586364061
transform 1 0 15180 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_12  FILLER_13_147
timestamp 1586364061
transform 1 0 14628 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_154
timestamp 1586364061
transform 1 0 15272 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_159
timestamp 1586364061
transform 1 0 15732 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_166
timestamp 1586364061
transform 1 0 16376 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_171
timestamp 1586364061
transform 1 0 16836 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_178
timestamp 1586364061
transform 1 0 17480 0 -1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_123
timestamp 1586364061
transform 1 0 17940 0 1 9248
box -38 -48 130 592
use scs8hd_decap_12  FILLER_13_184
timestamp 1586364061
transform 1 0 18032 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_190
timestamp 1586364061
transform 1 0 18584 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_196
timestamp 1586364061
transform 1 0 19136 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_202
timestamp 1586364061
transform 1 0 19688 0 -1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_127
timestamp 1586364061
transform 1 0 20792 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_12  FILLER_13_208
timestamp 1586364061
transform 1 0 20240 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_215
timestamp 1586364061
transform 1 0 20884 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_220
timestamp 1586364061
transform 1 0 21344 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_14_227
timestamp 1586364061
transform 1 0 21988 0 -1 10336
box -38 -48 590 592
use scs8hd_decap_3  PHY_27
timestamp 1586364061
transform -1 0 22816 0 1 9248
box -38 -48 314 592
use scs8hd_decap_3  PHY_29
timestamp 1586364061
transform -1 0 22816 0 -1 10336
box -38 -48 314 592
use scs8hd_fill_1  FILLER_13_232
timestamp 1586364061
transform 1 0 22448 0 1 9248
box -38 -48 130 592
use scs8hd_nor2_4  _077_
timestamp 1586364061
transform 1 0 1380 0 1 10336
box -38 -48 866 592
use scs8hd_decap_3  PHY_30
timestamp 1586364061
transform 1 0 1104 0 1 10336
box -38 -48 314 592
use scs8hd_fill_2  FILLER_15_12
timestamp 1586364061
transform 1 0 2208 0 1 10336
box -38 -48 222 592
use scs8hd_nor2_4  _089_
timestamp 1586364061
transform 1 0 2944 0 1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__077__A
timestamp 1586364061
transform 1 0 2392 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__086__A
timestamp 1586364061
transform 1 0 2760 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_16
timestamp 1586364061
transform 1 0 2576 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__079__A
timestamp 1586364061
transform 1 0 4416 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__080__B
timestamp 1586364061
transform 1 0 3956 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_29
timestamp 1586364061
transform 1 0 3772 0 1 10336
box -38 -48 222 592
use scs8hd_decap_3  FILLER_15_33
timestamp 1586364061
transform 1 0 4140 0 1 10336
box -38 -48 314 592
use scs8hd_fill_2  FILLER_15_38
timestamp 1586364061
transform 1 0 4600 0 1 10336
box -38 -48 222 592
use scs8hd_inv_8  _074_
timestamp 1586364061
transform 1 0 4968 0 1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__074__A
timestamp 1586364061
transform 1 0 4784 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_51
timestamp 1586364061
transform 1 0 5796 0 1 10336
box -38 -48 222 592
use scs8hd_buf_1  _082_
timestamp 1586364061
transform 1 0 6808 0 1 10336
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_128
timestamp 1586364061
transform 1 0 6716 0 1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__067__A
timestamp 1586364061
transform 1 0 5980 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__067__B
timestamp 1586364061
transform 1 0 6348 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_55
timestamp 1586364061
transform 1 0 6164 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_59
timestamp 1586364061
transform 1 0 6532 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__093__C
timestamp 1586364061
transform 1 0 7268 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__133__A
timestamp 1586364061
transform 1 0 7636 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__082__A
timestamp 1586364061
transform 1 0 8004 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_65
timestamp 1586364061
transform 1 0 7084 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_69
timestamp 1586364061
transform 1 0 7452 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_73
timestamp 1586364061
transform 1 0 7820 0 1 10336
box -38 -48 222 592
use scs8hd_decap_12  FILLER_15_77
timestamp 1586364061
transform 1 0 8188 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_89
timestamp 1586364061
transform 1 0 9292 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_101
timestamp 1586364061
transform 1 0 10396 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_15_113
timestamp 1586364061
transform 1 0 11500 0 1 10336
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_129
timestamp 1586364061
transform 1 0 12328 0 1 10336
box -38 -48 130 592
use scs8hd_fill_1  FILLER_15_121
timestamp 1586364061
transform 1 0 12236 0 1 10336
box -38 -48 130 592
use scs8hd_decap_12  FILLER_15_123
timestamp 1586364061
transform 1 0 12420 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_135
timestamp 1586364061
transform 1 0 13524 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_147
timestamp 1586364061
transform 1 0 14628 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_159
timestamp 1586364061
transform 1 0 15732 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_171
timestamp 1586364061
transform 1 0 16836 0 1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_130
timestamp 1586364061
transform 1 0 17940 0 1 10336
box -38 -48 130 592
use scs8hd_decap_12  FILLER_15_184
timestamp 1586364061
transform 1 0 18032 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_196
timestamp 1586364061
transform 1 0 19136 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_208
timestamp 1586364061
transform 1 0 20240 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_220
timestamp 1586364061
transform 1 0 21344 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_3  PHY_31
timestamp 1586364061
transform -1 0 22816 0 1 10336
box -38 -48 314 592
use scs8hd_fill_1  FILLER_15_232
timestamp 1586364061
transform 1 0 22448 0 1 10336
box -38 -48 130 592
use scs8hd_nor2_4  _080_
timestamp 1586364061
transform 1 0 1380 0 -1 11424
box -38 -48 866 592
use scs8hd_decap_3  PHY_32
timestamp 1586364061
transform 1 0 1104 0 -1 11424
box -38 -48 314 592
use scs8hd_fill_2  FILLER_16_12
timestamp 1586364061
transform 1 0 2208 0 -1 11424
box -38 -48 222 592
use scs8hd_buf_1  _086_
timestamp 1586364061
transform 1 0 2944 0 -1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__073__B
timestamp 1586364061
transform 1 0 2392 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__183__A
timestamp 1586364061
transform 1 0 2760 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__090__A
timestamp 1586364061
transform 1 0 3404 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_16
timestamp 1586364061
transform 1 0 2576 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_23
timestamp 1586364061
transform 1 0 3220 0 -1 11424
box -38 -48 222 592
use scs8hd_buf_1  _079_
timestamp 1586364061
transform 1 0 4600 0 -1 11424
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_131
timestamp 1586364061
transform 1 0 3956 0 -1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__175__A
timestamp 1586364061
transform 1 0 4232 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__184__B
timestamp 1586364061
transform 1 0 3772 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_27
timestamp 1586364061
transform 1 0 3588 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_32
timestamp 1586364061
transform 1 0 4048 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_36
timestamp 1586364061
transform 1 0 4416 0 -1 11424
box -38 -48 222 592
use scs8hd_or4_4  _067_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 5704 0 -1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__106__A
timestamp 1586364061
transform 1 0 5520 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__081__D
timestamp 1586364061
transform 1 0 5152 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_3  FILLER_16_41
timestamp 1586364061
transform 1 0 4876 0 -1 11424
box -38 -48 314 592
use scs8hd_fill_2  FILLER_16_46
timestamp 1586364061
transform 1 0 5336 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__093__A
timestamp 1586364061
transform 1 0 6808 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_3  FILLER_16_59
timestamp 1586364061
transform 1 0 6532 0 -1 11424
box -38 -48 314 592
use scs8hd_decap_3  FILLER_16_64
timestamp 1586364061
transform 1 0 6992 0 -1 11424
box -38 -48 314 592
use scs8hd_buf_1  _133_
timestamp 1586364061
transform 1 0 7268 0 -1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__099__A
timestamp 1586364061
transform 1 0 7728 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__099__B
timestamp 1586364061
transform 1 0 8096 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_70
timestamp 1586364061
transform 1 0 7544 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_74
timestamp 1586364061
transform 1 0 7912 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_12  FILLER_16_78
timestamp 1586364061
transform 1 0 8280 0 -1 11424
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_132
timestamp 1586364061
transform 1 0 9568 0 -1 11424
box -38 -48 130 592
use scs8hd_fill_2  FILLER_16_90
timestamp 1586364061
transform 1 0 9384 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_12  FILLER_16_93
timestamp 1586364061
transform 1 0 9660 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_105
timestamp 1586364061
transform 1 0 10764 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_117
timestamp 1586364061
transform 1 0 11868 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_129
timestamp 1586364061
transform 1 0 12972 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_141
timestamp 1586364061
transform 1 0 14076 0 -1 11424
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_133
timestamp 1586364061
transform 1 0 15180 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_12  FILLER_16_154
timestamp 1586364061
transform 1 0 15272 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_166
timestamp 1586364061
transform 1 0 16376 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_178
timestamp 1586364061
transform 1 0 17480 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_190
timestamp 1586364061
transform 1 0 18584 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_202
timestamp 1586364061
transform 1 0 19688 0 -1 11424
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_134
timestamp 1586364061
transform 1 0 20792 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_12  FILLER_16_215
timestamp 1586364061
transform 1 0 20884 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_16_227
timestamp 1586364061
transform 1 0 21988 0 -1 11424
box -38 -48 590 592
use scs8hd_decap_3  PHY_33
timestamp 1586364061
transform -1 0 22816 0 -1 11424
box -38 -48 314 592
use scs8hd_nor2_4  _073_
timestamp 1586364061
transform 1 0 1380 0 1 11424
box -38 -48 866 592
use scs8hd_decap_3  PHY_34
timestamp 1586364061
transform 1 0 1104 0 1 11424
box -38 -48 314 592
use scs8hd_fill_2  FILLER_17_12
timestamp 1586364061
transform 1 0 2208 0 1 11424
box -38 -48 222 592
use scs8hd_nor2_4  _184_
timestamp 1586364061
transform 1 0 3036 0 1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__183__B
timestamp 1586364061
transform 1 0 2392 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__184__A
timestamp 1586364061
transform 1 0 2852 0 1 11424
box -38 -48 222 592
use scs8hd_decap_3  FILLER_17_16
timestamp 1586364061
transform 1 0 2576 0 1 11424
box -38 -48 314 592
use scs8hd_buf_1  _068_
timestamp 1586364061
transform 1 0 4600 0 1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__175__B
timestamp 1586364061
transform 1 0 4048 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__068__A
timestamp 1586364061
transform 1 0 4416 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_30
timestamp 1586364061
transform 1 0 3864 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_34
timestamp 1586364061
transform 1 0 4232 0 1 11424
box -38 -48 222 592
use scs8hd_buf_1  _106_
timestamp 1586364061
transform 1 0 5612 0 1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__081__A
timestamp 1586364061
transform 1 0 5428 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__108__D
timestamp 1586364061
transform 1 0 5060 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_41
timestamp 1586364061
transform 1 0 4876 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_45
timestamp 1586364061
transform 1 0 5244 0 1 11424
box -38 -48 222 592
use scs8hd_or4_4  _093_
timestamp 1586364061
transform 1 0 6808 0 1 11424
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_135
timestamp 1586364061
transform 1 0 6716 0 1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__081__C
timestamp 1586364061
transform 1 0 6072 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__093__D
timestamp 1586364061
transform 1 0 6532 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_52
timestamp 1586364061
transform 1 0 5888 0 1 11424
box -38 -48 222 592
use scs8hd_decap_3  FILLER_17_56
timestamp 1586364061
transform 1 0 6256 0 1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__099__C
timestamp 1586364061
transform 1 0 7820 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__099__D
timestamp 1586364061
transform 1 0 8188 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_71
timestamp 1586364061
transform 1 0 7636 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_75
timestamp 1586364061
transform 1 0 8004 0 1 11424
box -38 -48 222 592
use scs8hd_buf_1  _135_
timestamp 1586364061
transform 1 0 8372 0 1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__135__A
timestamp 1586364061
transform 1 0 8832 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_82
timestamp 1586364061
transform 1 0 8648 0 1 11424
box -38 -48 222 592
use scs8hd_decap_12  FILLER_17_86
timestamp 1586364061
transform 1 0 9016 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_98
timestamp 1586364061
transform 1 0 10120 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_110
timestamp 1586364061
transform 1 0 11224 0 1 11424
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_136
timestamp 1586364061
transform 1 0 12328 0 1 11424
box -38 -48 130 592
use scs8hd_decap_12  FILLER_17_123
timestamp 1586364061
transform 1 0 12420 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_135
timestamp 1586364061
transform 1 0 13524 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_147
timestamp 1586364061
transform 1 0 14628 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_159
timestamp 1586364061
transform 1 0 15732 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_171
timestamp 1586364061
transform 1 0 16836 0 1 11424
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_137
timestamp 1586364061
transform 1 0 17940 0 1 11424
box -38 -48 130 592
use scs8hd_decap_12  FILLER_17_184
timestamp 1586364061
transform 1 0 18032 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_196
timestamp 1586364061
transform 1 0 19136 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_208
timestamp 1586364061
transform 1 0 20240 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_220
timestamp 1586364061
transform 1 0 21344 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_3  PHY_35
timestamp 1586364061
transform -1 0 22816 0 1 11424
box -38 -48 314 592
use scs8hd_fill_1  FILLER_17_232
timestamp 1586364061
transform 1 0 22448 0 1 11424
box -38 -48 130 592
use scs8hd_buf_1  _090_
timestamp 1586364061
transform 1 0 1380 0 -1 12512
box -38 -48 314 592
use scs8hd_decap_3  PHY_36
timestamp 1586364061
transform 1 0 1104 0 -1 12512
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__073__A
timestamp 1586364061
transform 1 0 1840 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__131__A
timestamp 1586364061
transform 1 0 2208 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_6
timestamp 1586364061
transform 1 0 1656 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_10
timestamp 1586364061
transform 1 0 2024 0 -1 12512
box -38 -48 222 592
use scs8hd_nor2_4  _183_
timestamp 1586364061
transform 1 0 2392 0 -1 12512
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__171__A
timestamp 1586364061
transform 1 0 3404 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_23
timestamp 1586364061
transform 1 0 3220 0 -1 12512
box -38 -48 222 592
use scs8hd_nor2_4  _175_
timestamp 1586364061
transform 1 0 4048 0 -1 12512
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_138
timestamp 1586364061
transform 1 0 3956 0 -1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__180__A
timestamp 1586364061
transform 1 0 3772 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_27
timestamp 1586364061
transform 1 0 3588 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__108__B
timestamp 1586364061
transform 1 0 5060 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__115__A
timestamp 1586364061
transform 1 0 5428 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_41
timestamp 1586364061
transform 1 0 4876 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_45
timestamp 1586364061
transform 1 0 5244 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_3  FILLER_18_49
timestamp 1586364061
transform 1 0 5612 0 -1 12512
box -38 -48 314 592
use scs8hd_or4_4  _081_
timestamp 1586364061
transform 1 0 6072 0 -1 12512
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__081__B
timestamp 1586364061
transform 1 0 5888 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_63
timestamp 1586364061
transform 1 0 6900 0 -1 12512
box -38 -48 222 592
use scs8hd_or4_4  _099_
timestamp 1586364061
transform 1 0 7636 0 -1 12512
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__066__A
timestamp 1586364061
transform 1 0 7084 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__093__B
timestamp 1586364061
transform 1 0 7452 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_67
timestamp 1586364061
transform 1 0 7268 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_12  FILLER_18_80
timestamp 1586364061
transform 1 0 8464 0 -1 12512
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_139
timestamp 1586364061
transform 1 0 9568 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_12  FILLER_18_93
timestamp 1586364061
transform 1 0 9660 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_105
timestamp 1586364061
transform 1 0 10764 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_117
timestamp 1586364061
transform 1 0 11868 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_129
timestamp 1586364061
transform 1 0 12972 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_141
timestamp 1586364061
transform 1 0 14076 0 -1 12512
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_140
timestamp 1586364061
transform 1 0 15180 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_12  FILLER_18_154
timestamp 1586364061
transform 1 0 15272 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_166
timestamp 1586364061
transform 1 0 16376 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_178
timestamp 1586364061
transform 1 0 17480 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_190
timestamp 1586364061
transform 1 0 18584 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_202
timestamp 1586364061
transform 1 0 19688 0 -1 12512
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_141
timestamp 1586364061
transform 1 0 20792 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_12  FILLER_18_215
timestamp 1586364061
transform 1 0 20884 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_18_227
timestamp 1586364061
transform 1 0 21988 0 -1 12512
box -38 -48 590 592
use scs8hd_decap_3  PHY_37
timestamp 1586364061
transform -1 0 22816 0 -1 12512
box -38 -48 314 592
use scs8hd_fill_1  FILLER_19_3
timestamp 1586364061
transform 1 0 1380 0 1 12512
box -38 -48 130 592
use scs8hd_decap_3  PHY_40
timestamp 1586364061
transform 1 0 1104 0 -1 13600
box -38 -48 314 592
use scs8hd_decap_3  PHY_38
timestamp 1586364061
transform 1 0 1104 0 1 12512
box -38 -48 314 592
use scs8hd_buf_1  _141_
timestamp 1586364061
transform 1 0 1380 0 -1 13600
box -38 -48 314 592
use scs8hd_fill_2  FILLER_20_6
timestamp 1586364061
transform 1 0 1656 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_7
timestamp 1586364061
transform 1 0 1748 0 1 12512
box -38 -48 222 592
use scs8hd_buf_1  _131_
timestamp 1586364061
transform 1 0 1472 0 1 12512
box -38 -48 314 592
use scs8hd_fill_2  FILLER_20_10
timestamp 1586364061
transform 1 0 2024 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_11
timestamp 1586364061
transform 1 0 2116 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__181__B
timestamp 1586364061
transform 1 0 1932 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__177__B
timestamp 1586364061
transform 1 0 1840 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__182__A
timestamp 1586364061
transform 1 0 2208 0 -1 13600
box -38 -48 222 592
use scs8hd_nor2_4  _181_
timestamp 1586364061
transform 1 0 2392 0 -1 13600
box -38 -48 866 592
use scs8hd_nor2_4  _182_
timestamp 1586364061
transform 1 0 2484 0 1 12512
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__182__B
timestamp 1586364061
transform 1 0 2300 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__177__A
timestamp 1586364061
transform 1 0 3404 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_24
timestamp 1586364061
transform 1 0 3312 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_23
timestamp 1586364061
transform 1 0 3220 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_27
timestamp 1586364061
transform 1 0 3588 0 -1 13600
box -38 -48 222 592
use scs8hd_decap_3  FILLER_19_28
timestamp 1586364061
transform 1 0 3680 0 1 12512
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__181__A
timestamp 1586364061
transform 1 0 3496 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__179__A
timestamp 1586364061
transform 1 0 3772 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_32
timestamp 1586364061
transform 1 0 4048 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_33
timestamp 1586364061
transform 1 0 4140 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__115__C
timestamp 1586364061
transform 1 0 3956 0 1 12512
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_145
timestamp 1586364061
transform 1 0 3956 0 -1 13600
box -38 -48 130 592
use scs8hd_fill_2  FILLER_20_36
timestamp 1586364061
transform 1 0 4416 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_37
timestamp 1586364061
transform 1 0 4508 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__128__B
timestamp 1586364061
transform 1 0 4232 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__115__B
timestamp 1586364061
transform 1 0 4324 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__128__A
timestamp 1586364061
transform 1 0 4600 0 -1 13600
box -38 -48 222 592
use scs8hd_or4_4  _108_
timestamp 1586364061
transform 1 0 4876 0 1 12512
box -38 -48 866 592
use scs8hd_or4_4  _115_
timestamp 1586364061
transform 1 0 4784 0 -1 13600
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__108__A
timestamp 1586364061
transform 1 0 4692 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__122__C
timestamp 1586364061
transform 1 0 5796 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_50
timestamp 1586364061
transform 1 0 5704 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_49
timestamp 1586364061
transform 1 0 5612 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_53
timestamp 1586364061
transform 1 0 5980 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_54
timestamp 1586364061
transform 1 0 6072 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__122__B
timestamp 1586364061
transform 1 0 6164 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__108__C
timestamp 1586364061
transform 1 0 5888 0 1 12512
box -38 -48 222 592
use scs8hd_decap_3  FILLER_19_58
timestamp 1586364061
transform 1 0 6440 0 1 12512
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__115__D
timestamp 1586364061
transform 1 0 6256 0 1 12512
box -38 -48 222 592
use scs8hd_buf_1  _105_
timestamp 1586364061
transform 1 0 6348 0 -1 13600
box -38 -48 314 592
use scs8hd_fill_2  FILLER_20_60
timestamp 1586364061
transform 1 0 6624 0 -1 13600
box -38 -48 222 592
use scs8hd_decap_3  FILLER_19_62
timestamp 1586364061
transform 1 0 6808 0 1 12512
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__176__B
timestamp 1586364061
transform 1 0 6808 0 -1 13600
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_142
timestamp 1586364061
transform 1 0 6716 0 1 12512
box -38 -48 130 592
use scs8hd_fill_2  FILLER_20_64
timestamp 1586364061
transform 1 0 6992 0 -1 13600
box -38 -48 222 592
use scs8hd_inv_8  _065_
timestamp 1586364061
transform 1 0 7360 0 -1 13600
box -38 -48 866 592
use scs8hd_inv_8  _066_
timestamp 1586364061
transform 1 0 7084 0 1 12512
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__065__A
timestamp 1586364061
transform 1 0 8096 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__105__A
timestamp 1586364061
transform 1 0 7176 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_74
timestamp 1586364061
transform 1 0 7912 0 1 12512
box -38 -48 222 592
use scs8hd_decap_12  FILLER_20_77
timestamp 1586364061
transform 1 0 8188 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_78
timestamp 1586364061
transform 1 0 8280 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_20_89
timestamp 1586364061
transform 1 0 9292 0 -1 13600
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_146
timestamp 1586364061
transform 1 0 9568 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_12  FILLER_19_90
timestamp 1586364061
transform 1 0 9384 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_102
timestamp 1586364061
transform 1 0 10488 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_93
timestamp 1586364061
transform 1 0 9660 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_19_114
timestamp 1586364061
transform 1 0 11592 0 1 12512
box -38 -48 774 592
use scs8hd_decap_12  FILLER_20_105
timestamp 1586364061
transform 1 0 10764 0 -1 13600
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_143
timestamp 1586364061
transform 1 0 12328 0 1 12512
box -38 -48 130 592
use scs8hd_decap_12  FILLER_19_123
timestamp 1586364061
transform 1 0 12420 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_117
timestamp 1586364061
transform 1 0 11868 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_135
timestamp 1586364061
transform 1 0 13524 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_129
timestamp 1586364061
transform 1 0 12972 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_141
timestamp 1586364061
transform 1 0 14076 0 -1 13600
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_147
timestamp 1586364061
transform 1 0 15180 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_12  FILLER_19_147
timestamp 1586364061
transform 1 0 14628 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_154
timestamp 1586364061
transform 1 0 15272 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_159
timestamp 1586364061
transform 1 0 15732 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_166
timestamp 1586364061
transform 1 0 16376 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_171
timestamp 1586364061
transform 1 0 16836 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_178
timestamp 1586364061
transform 1 0 17480 0 -1 13600
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_144
timestamp 1586364061
transform 1 0 17940 0 1 12512
box -38 -48 130 592
use scs8hd_decap_12  FILLER_19_184
timestamp 1586364061
transform 1 0 18032 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_190
timestamp 1586364061
transform 1 0 18584 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_196
timestamp 1586364061
transform 1 0 19136 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_202
timestamp 1586364061
transform 1 0 19688 0 -1 13600
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_148
timestamp 1586364061
transform 1 0 20792 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_12  FILLER_19_208
timestamp 1586364061
transform 1 0 20240 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_215
timestamp 1586364061
transform 1 0 20884 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_220
timestamp 1586364061
transform 1 0 21344 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_20_227
timestamp 1586364061
transform 1 0 21988 0 -1 13600
box -38 -48 590 592
use scs8hd_decap_3  PHY_39
timestamp 1586364061
transform -1 0 22816 0 1 12512
box -38 -48 314 592
use scs8hd_decap_3  PHY_41
timestamp 1586364061
transform -1 0 22816 0 -1 13600
box -38 -48 314 592
use scs8hd_fill_1  FILLER_19_232
timestamp 1586364061
transform 1 0 22448 0 1 12512
box -38 -48 130 592
use scs8hd_nor2_4  _177_
timestamp 1586364061
transform 1 0 1380 0 1 13600
box -38 -48 866 592
use scs8hd_decap_3  PHY_42
timestamp 1586364061
transform 1 0 1104 0 1 13600
box -38 -48 314 592
use scs8hd_fill_2  FILLER_21_12
timestamp 1586364061
transform 1 0 2208 0 1 13600
box -38 -48 222 592
use scs8hd_nor2_4  _180_
timestamp 1586364061
transform 1 0 2944 0 1 13600
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__171__B
timestamp 1586364061
transform 1 0 2392 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__180__B
timestamp 1586364061
transform 1 0 2760 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_16
timestamp 1586364061
transform 1 0 2576 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__122__D
timestamp 1586364061
transform 1 0 4508 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__122__A
timestamp 1586364061
transform 1 0 4140 0 1 13600
box -38 -48 222 592
use scs8hd_decap_4  FILLER_21_29
timestamp 1586364061
transform 1 0 3772 0 1 13600
box -38 -48 406 592
use scs8hd_fill_2  FILLER_21_35
timestamp 1586364061
transform 1 0 4324 0 1 13600
box -38 -48 222 592
use scs8hd_or4_4  _122_
timestamp 1586364061
transform 1 0 5060 0 1 13600
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__128__D
timestamp 1586364061
transform 1 0 4876 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_39
timestamp 1586364061
transform 1 0 4692 0 1 13600
box -38 -48 222 592
use scs8hd_nor2_4  _176_
timestamp 1586364061
transform 1 0 6808 0 1 13600
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_149
timestamp 1586364061
transform 1 0 6716 0 1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__064__A
timestamp 1586364061
transform 1 0 6532 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__128__C
timestamp 1586364061
transform 1 0 6072 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_52
timestamp 1586364061
transform 1 0 5888 0 1 13600
box -38 -48 222 592
use scs8hd_decap_3  FILLER_21_56
timestamp 1586364061
transform 1 0 6256 0 1 13600
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__176__A
timestamp 1586364061
transform 1 0 7820 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_71
timestamp 1586364061
transform 1 0 7636 0 1 13600
box -38 -48 222 592
use scs8hd_decap_12  FILLER_21_75
timestamp 1586364061
transform 1 0 8004 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_21_87
timestamp 1586364061
transform 1 0 9108 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_21_99
timestamp 1586364061
transform 1 0 10212 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_21_111
timestamp 1586364061
transform 1 0 11316 0 1 13600
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_150
timestamp 1586364061
transform 1 0 12328 0 1 13600
box -38 -48 130 592
use scs8hd_decap_3  FILLER_21_119
timestamp 1586364061
transform 1 0 12052 0 1 13600
box -38 -48 314 592
use scs8hd_decap_12  FILLER_21_123
timestamp 1586364061
transform 1 0 12420 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_21_135
timestamp 1586364061
transform 1 0 13524 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_21_147
timestamp 1586364061
transform 1 0 14628 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_21_159
timestamp 1586364061
transform 1 0 15732 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_21_171
timestamp 1586364061
transform 1 0 16836 0 1 13600
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_151
timestamp 1586364061
transform 1 0 17940 0 1 13600
box -38 -48 130 592
use scs8hd_decap_12  FILLER_21_184
timestamp 1586364061
transform 1 0 18032 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_21_196
timestamp 1586364061
transform 1 0 19136 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_21_208
timestamp 1586364061
transform 1 0 20240 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_21_220
timestamp 1586364061
transform 1 0 21344 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_3  PHY_43
timestamp 1586364061
transform -1 0 22816 0 1 13600
box -38 -48 314 592
use scs8hd_fill_1  FILLER_21_232
timestamp 1586364061
transform 1 0 22448 0 1 13600
box -38 -48 130 592
use scs8hd_nor2_4  _171_
timestamp 1586364061
transform 1 0 2208 0 -1 14688
box -38 -48 866 592
use scs8hd_decap_3  PHY_44
timestamp 1586364061
transform 1 0 1104 0 -1 14688
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__169__B
timestamp 1586364061
transform 1 0 1748 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_22_3
timestamp 1586364061
transform 1 0 1380 0 -1 14688
box -38 -48 406 592
use scs8hd_decap_3  FILLER_22_9
timestamp 1586364061
transform 1 0 1932 0 -1 14688
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__174__B
timestamp 1586364061
transform 1 0 3220 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_21
timestamp 1586364061
transform 1 0 3036 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_22_25
timestamp 1586364061
transform 1 0 3404 0 -1 14688
box -38 -48 406 592
use scs8hd_buf_1  _179_
timestamp 1586364061
transform 1 0 4048 0 -1 14688
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_152
timestamp 1586364061
transform 1 0 3956 0 -1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__173__A
timestamp 1586364061
transform 1 0 3772 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_22_35
timestamp 1586364061
transform 1 0 4324 0 -1 14688
box -38 -48 406 592
use scs8hd_or4_4  _128_
timestamp 1586364061
transform 1 0 5060 0 -1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__160__B
timestamp 1586364061
transform 1 0 4692 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_41
timestamp 1586364061
transform 1 0 4876 0 -1 14688
box -38 -48 222 592
use scs8hd_buf_1  _064_
timestamp 1586364061
transform 1 0 6624 0 -1 14688
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__178__B
timestamp 1586364061
transform 1 0 6072 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_52
timestamp 1586364061
transform 1 0 5888 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_22_56
timestamp 1586364061
transform 1 0 6256 0 -1 14688
box -38 -48 406 592
use scs8hd_fill_2  FILLER_22_63
timestamp 1586364061
transform 1 0 6900 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__172__A
timestamp 1586364061
transform 1 0 7084 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__172__D
timestamp 1586364061
transform 1 0 7452 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_67
timestamp 1586364061
transform 1 0 7268 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_12  FILLER_22_71
timestamp 1586364061
transform 1 0 7636 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_22_83
timestamp 1586364061
transform 1 0 8740 0 -1 14688
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_153
timestamp 1586364061
transform 1 0 9568 0 -1 14688
box -38 -48 130 592
use scs8hd_fill_1  FILLER_22_91
timestamp 1586364061
transform 1 0 9476 0 -1 14688
box -38 -48 130 592
use scs8hd_decap_12  FILLER_22_93
timestamp 1586364061
transform 1 0 9660 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_105
timestamp 1586364061
transform 1 0 10764 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_117
timestamp 1586364061
transform 1 0 11868 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_129
timestamp 1586364061
transform 1 0 12972 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_141
timestamp 1586364061
transform 1 0 14076 0 -1 14688
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_154
timestamp 1586364061
transform 1 0 15180 0 -1 14688
box -38 -48 130 592
use scs8hd_decap_12  FILLER_22_154
timestamp 1586364061
transform 1 0 15272 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_166
timestamp 1586364061
transform 1 0 16376 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_178
timestamp 1586364061
transform 1 0 17480 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_190
timestamp 1586364061
transform 1 0 18584 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_202
timestamp 1586364061
transform 1 0 19688 0 -1 14688
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_155
timestamp 1586364061
transform 1 0 20792 0 -1 14688
box -38 -48 130 592
use scs8hd_decap_12  FILLER_22_215
timestamp 1586364061
transform 1 0 20884 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_22_227
timestamp 1586364061
transform 1 0 21988 0 -1 14688
box -38 -48 590 592
use scs8hd_decap_3  PHY_45
timestamp 1586364061
transform -1 0 22816 0 -1 14688
box -38 -48 314 592
use scs8hd_decap_3  PHY_46
timestamp 1586364061
transform 1 0 1104 0 1 14688
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__169__A
timestamp 1586364061
transform 1 0 1748 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__170__A
timestamp 1586364061
transform 1 0 2116 0 1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_23_3
timestamp 1586364061
transform 1 0 1380 0 1 14688
box -38 -48 406 592
use scs8hd_fill_2  FILLER_23_9
timestamp 1586364061
transform 1 0 1932 0 1 14688
box -38 -48 222 592
use scs8hd_nor2_4  _170_
timestamp 1586364061
transform 1 0 2300 0 1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__170__B
timestamp 1586364061
transform 1 0 3312 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_22
timestamp 1586364061
transform 1 0 3128 0 1 14688
box -38 -48 222 592
use scs8hd_buf_1  _173_
timestamp 1586364061
transform 1 0 3864 0 1 14688
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__160__A
timestamp 1586364061
transform 1 0 4600 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__160__D
timestamp 1586364061
transform 1 0 3680 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_26
timestamp 1586364061
transform 1 0 3496 0 1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_23_33
timestamp 1586364061
transform 1 0 4140 0 1 14688
box -38 -48 406 592
use scs8hd_fill_1  FILLER_23_37
timestamp 1586364061
transform 1 0 4508 0 1 14688
box -38 -48 130 592
use scs8hd_or4_4  _178_
timestamp 1586364061
transform 1 0 5152 0 1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__178__C
timestamp 1586364061
transform 1 0 4968 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_40
timestamp 1586364061
transform 1 0 4784 0 1 14688
box -38 -48 222 592
use scs8hd_or4_4  _172_
timestamp 1586364061
transform 1 0 6808 0 1 14688
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_156
timestamp 1586364061
transform 1 0 6716 0 1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__172__C
timestamp 1586364061
transform 1 0 6532 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__137__A
timestamp 1586364061
transform 1 0 6164 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_53
timestamp 1586364061
transform 1 0 5980 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_57
timestamp 1586364061
transform 1 0 6348 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__172__B
timestamp 1586364061
transform 1 0 7820 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_71
timestamp 1586364061
transform 1 0 7636 0 1 14688
box -38 -48 222 592
use scs8hd_decap_12  FILLER_23_75
timestamp 1586364061
transform 1 0 8004 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_87
timestamp 1586364061
transform 1 0 9108 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_99
timestamp 1586364061
transform 1 0 10212 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_23_111
timestamp 1586364061
transform 1 0 11316 0 1 14688
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_157
timestamp 1586364061
transform 1 0 12328 0 1 14688
box -38 -48 130 592
use scs8hd_decap_3  FILLER_23_119
timestamp 1586364061
transform 1 0 12052 0 1 14688
box -38 -48 314 592
use scs8hd_decap_12  FILLER_23_123
timestamp 1586364061
transform 1 0 12420 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_135
timestamp 1586364061
transform 1 0 13524 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_147
timestamp 1586364061
transform 1 0 14628 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_159
timestamp 1586364061
transform 1 0 15732 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_171
timestamp 1586364061
transform 1 0 16836 0 1 14688
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_158
timestamp 1586364061
transform 1 0 17940 0 1 14688
box -38 -48 130 592
use scs8hd_decap_12  FILLER_23_184
timestamp 1586364061
transform 1 0 18032 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_196
timestamp 1586364061
transform 1 0 19136 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_208
timestamp 1586364061
transform 1 0 20240 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_220
timestamp 1586364061
transform 1 0 21344 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_3  PHY_47
timestamp 1586364061
transform -1 0 22816 0 1 14688
box -38 -48 314 592
use scs8hd_fill_1  FILLER_23_232
timestamp 1586364061
transform 1 0 22448 0 1 14688
box -38 -48 130 592
use scs8hd_nor2_4  _169_
timestamp 1586364061
transform 1 0 1748 0 -1 15776
box -38 -48 866 592
use scs8hd_decap_3  PHY_48
timestamp 1586364061
transform 1 0 1104 0 -1 15776
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__168__A
timestamp 1586364061
transform 1 0 1564 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_3
timestamp 1586364061
transform 1 0 1380 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__164__B
timestamp 1586364061
transform 1 0 2760 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__168__B
timestamp 1586364061
transform 1 0 3128 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_16
timestamp 1586364061
transform 1 0 2576 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_20
timestamp 1586364061
transform 1 0 2944 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_24_24
timestamp 1586364061
transform 1 0 3312 0 -1 15776
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_159
timestamp 1586364061
transform 1 0 3956 0 -1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__160__C
timestamp 1586364061
transform 1 0 4508 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__161__A
timestamp 1586364061
transform 1 0 3772 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_1  FILLER_24_28
timestamp 1586364061
transform 1 0 3680 0 -1 15776
box -38 -48 130 592
use scs8hd_decap_4  FILLER_24_32
timestamp 1586364061
transform 1 0 4048 0 -1 15776
box -38 -48 406 592
use scs8hd_fill_1  FILLER_24_36
timestamp 1586364061
transform 1 0 4416 0 -1 15776
box -38 -48 130 592
use scs8hd_or4_4  _160_
timestamp 1586364061
transform 1 0 4692 0 -1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__178__A
timestamp 1586364061
transform 1 0 5704 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_48
timestamp 1586364061
transform 1 0 5520 0 -1 15776
box -38 -48 222 592
use scs8hd_inv_8  _137_
timestamp 1586364061
transform 1 0 6624 0 -1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__178__D
timestamp 1586364061
transform 1 0 6072 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__139__C
timestamp 1586364061
transform 1 0 6440 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_52
timestamp 1586364061
transform 1 0 5888 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_56
timestamp 1586364061
transform 1 0 6256 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_12  FILLER_24_69
timestamp 1586364061
transform 1 0 7452 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_24_81
timestamp 1586364061
transform 1 0 8556 0 -1 15776
box -38 -48 774 592
use scs8hd_decap_3  FILLER_24_89
timestamp 1586364061
transform 1 0 9292 0 -1 15776
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_160
timestamp 1586364061
transform 1 0 9568 0 -1 15776
box -38 -48 130 592
use scs8hd_decap_12  FILLER_24_93
timestamp 1586364061
transform 1 0 9660 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_105
timestamp 1586364061
transform 1 0 10764 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_117
timestamp 1586364061
transform 1 0 11868 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_129
timestamp 1586364061
transform 1 0 12972 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_141
timestamp 1586364061
transform 1 0 14076 0 -1 15776
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_161
timestamp 1586364061
transform 1 0 15180 0 -1 15776
box -38 -48 130 592
use scs8hd_decap_12  FILLER_24_154
timestamp 1586364061
transform 1 0 15272 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_166
timestamp 1586364061
transform 1 0 16376 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_178
timestamp 1586364061
transform 1 0 17480 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_190
timestamp 1586364061
transform 1 0 18584 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_202
timestamp 1586364061
transform 1 0 19688 0 -1 15776
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_162
timestamp 1586364061
transform 1 0 20792 0 -1 15776
box -38 -48 130 592
use scs8hd_decap_12  FILLER_24_215
timestamp 1586364061
transform 1 0 20884 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_24_227
timestamp 1586364061
transform 1 0 21988 0 -1 15776
box -38 -48 590 592
use scs8hd_decap_3  PHY_49
timestamp 1586364061
transform -1 0 22816 0 -1 15776
box -38 -48 314 592
use scs8hd_nor2_4  _168_
timestamp 1586364061
transform 1 0 1564 0 1 15776
box -38 -48 866 592
use scs8hd_decap_3  PHY_50
timestamp 1586364061
transform 1 0 1104 0 1 15776
box -38 -48 314 592
use scs8hd_fill_2  FILLER_25_3
timestamp 1586364061
transform 1 0 1380 0 1 15776
box -38 -48 222 592
use scs8hd_nor2_4  _174_
timestamp 1586364061
transform 1 0 3128 0 1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__164__A
timestamp 1586364061
transform 1 0 2576 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__174__A
timestamp 1586364061
transform 1 0 2944 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_14
timestamp 1586364061
transform 1 0 2392 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_18
timestamp 1586364061
transform 1 0 2760 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__166__B
timestamp 1586364061
transform 1 0 4508 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__166__A
timestamp 1586364061
transform 1 0 4140 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_31
timestamp 1586364061
transform 1 0 3956 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_35
timestamp 1586364061
transform 1 0 4324 0 1 15776
box -38 -48 222 592
use scs8hd_or4_4  _166_
timestamp 1586364061
transform 1 0 4692 0 1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__139__A
timestamp 1586364061
transform 1 0 5704 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_48
timestamp 1586364061
transform 1 0 5520 0 1 15776
box -38 -48 222 592
use scs8hd_buf_1  _107_
timestamp 1586364061
transform 1 0 6808 0 1 15776
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_163
timestamp 1586364061
transform 1 0 6716 0 1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__139__B
timestamp 1586364061
transform 1 0 6072 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__166__D
timestamp 1586364061
transform 1 0 6440 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_52
timestamp 1586364061
transform 1 0 5888 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_56
timestamp 1586364061
transform 1 0 6256 0 1 15776
box -38 -48 222 592
use scs8hd_fill_1  FILLER_25_60
timestamp 1586364061
transform 1 0 6624 0 1 15776
box -38 -48 130 592
use scs8hd_buf_1  _138_
timestamp 1586364061
transform 1 0 7820 0 1 15776
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__114__A
timestamp 1586364061
transform 1 0 7268 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__107__A
timestamp 1586364061
transform 1 0 7636 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_65
timestamp 1586364061
transform 1 0 7084 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_69
timestamp 1586364061
transform 1 0 7452 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_76
timestamp 1586364061
transform 1 0 8096 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__138__A
timestamp 1586364061
transform 1 0 8280 0 1 15776
box -38 -48 222 592
use scs8hd_decap_12  FILLER_25_80
timestamp 1586364061
transform 1 0 8464 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_92
timestamp 1586364061
transform 1 0 9568 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_104
timestamp 1586364061
transform 1 0 10672 0 1 15776
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_164
timestamp 1586364061
transform 1 0 12328 0 1 15776
box -38 -48 130 592
use scs8hd_decap_6  FILLER_25_116
timestamp 1586364061
transform 1 0 11776 0 1 15776
box -38 -48 590 592
use scs8hd_decap_12  FILLER_25_123
timestamp 1586364061
transform 1 0 12420 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_135
timestamp 1586364061
transform 1 0 13524 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_147
timestamp 1586364061
transform 1 0 14628 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_159
timestamp 1586364061
transform 1 0 15732 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_171
timestamp 1586364061
transform 1 0 16836 0 1 15776
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_165
timestamp 1586364061
transform 1 0 17940 0 1 15776
box -38 -48 130 592
use scs8hd_decap_12  FILLER_25_184
timestamp 1586364061
transform 1 0 18032 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_196
timestamp 1586364061
transform 1 0 19136 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_208
timestamp 1586364061
transform 1 0 20240 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_220
timestamp 1586364061
transform 1 0 21344 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_3  PHY_51
timestamp 1586364061
transform -1 0 22816 0 1 15776
box -38 -48 314 592
use scs8hd_fill_1  FILLER_25_232
timestamp 1586364061
transform 1 0 22448 0 1 15776
box -38 -48 130 592
use scs8hd_nor2_4  _163_
timestamp 1586364061
transform 1 0 1380 0 1 16864
box -38 -48 866 592
use scs8hd_nor2_4  _164_
timestamp 1586364061
transform 1 0 2024 0 -1 16864
box -38 -48 866 592
use scs8hd_decap_3  PHY_52
timestamp 1586364061
transform 1 0 1104 0 -1 16864
box -38 -48 314 592
use scs8hd_decap_3  PHY_54
timestamp 1586364061
transform 1 0 1104 0 1 16864
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__163__A
timestamp 1586364061
transform 1 0 1564 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_3
timestamp 1586364061
transform 1 0 1380 0 -1 16864
box -38 -48 222 592
use scs8hd_decap_3  FILLER_26_7
timestamp 1586364061
transform 1 0 1748 0 -1 16864
box -38 -48 314 592
use scs8hd_fill_2  FILLER_27_12
timestamp 1586364061
transform 1 0 2208 0 1 16864
box -38 -48 222 592
use scs8hd_nor2_4  _165_
timestamp 1586364061
transform 1 0 3036 0 1 16864
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__165__A
timestamp 1586364061
transform 1 0 2852 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__162__A
timestamp 1586364061
transform 1 0 2392 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__165__B
timestamp 1586364061
transform 1 0 3036 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__162__B
timestamp 1586364061
transform 1 0 3404 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_19
timestamp 1586364061
transform 1 0 2852 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_23
timestamp 1586364061
transform 1 0 3220 0 -1 16864
box -38 -48 222 592
use scs8hd_decap_3  FILLER_27_16
timestamp 1586364061
transform 1 0 2576 0 1 16864
box -38 -48 314 592
use scs8hd_buf_1  _161_
timestamp 1586364061
transform 1 0 4048 0 -1 16864
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_166
timestamp 1586364061
transform 1 0 3956 0 -1 16864
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__154__A
timestamp 1586364061
transform 1 0 4600 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__142__A
timestamp 1586364061
transform 1 0 4232 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__167__A
timestamp 1586364061
transform 1 0 3772 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_27
timestamp 1586364061
transform 1 0 3588 0 -1 16864
box -38 -48 222 592
use scs8hd_decap_4  FILLER_26_35
timestamp 1586364061
transform 1 0 4324 0 -1 16864
box -38 -48 406 592
use scs8hd_decap_4  FILLER_27_30
timestamp 1586364061
transform 1 0 3864 0 1 16864
box -38 -48 406 592
use scs8hd_fill_2  FILLER_27_36
timestamp 1586364061
transform 1 0 4416 0 1 16864
box -38 -48 222 592
use scs8hd_or4_4  _139_
timestamp 1586364061
transform 1 0 5152 0 -1 16864
box -38 -48 866 592
use scs8hd_or4_4  _142_
timestamp 1586364061
transform 1 0 5152 0 1 16864
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__142__B
timestamp 1586364061
transform 1 0 4968 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__166__C
timestamp 1586364061
transform 1 0 4692 0 -1 16864
box -38 -48 222 592
use scs8hd_decap_3  FILLER_26_41
timestamp 1586364061
transform 1 0 4876 0 -1 16864
box -38 -48 314 592
use scs8hd_fill_2  FILLER_27_40
timestamp 1586364061
transform 1 0 4784 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_57
timestamp 1586364061
transform 1 0 6348 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_53
timestamp 1586364061
transform 1 0 5980 0 1 16864
box -38 -48 222 592
use scs8hd_decap_4  FILLER_26_57
timestamp 1586364061
transform 1 0 6348 0 -1 16864
box -38 -48 406 592
use scs8hd_fill_2  FILLER_26_53
timestamp 1586364061
transform 1 0 5980 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__139__D
timestamp 1586364061
transform 1 0 6164 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__154__B
timestamp 1586364061
transform 1 0 6164 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__062__A
timestamp 1586364061
transform 1 0 6532 0 1 16864
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_170
timestamp 1586364061
transform 1 0 6716 0 1 16864
box -38 -48 130 592
use scs8hd_buf_1  _121_
timestamp 1586364061
transform 1 0 6808 0 1 16864
box -38 -48 314 592
use scs8hd_buf_1  _114_
timestamp 1586364061
transform 1 0 6716 0 -1 16864
box -38 -48 314 592
use scs8hd_decap_12  FILLER_26_64
timestamp 1586364061
transform 1 0 6992 0 -1 16864
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA__121__A
timestamp 1586364061
transform 1 0 7268 0 1 16864
box -38 -48 222 592
use scs8hd_decap_12  FILLER_26_76
timestamp 1586364061
transform 1 0 8096 0 -1 16864
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_27_65
timestamp 1586364061
transform 1 0 7084 0 1 16864
box -38 -48 222 592
use scs8hd_decap_12  FILLER_27_69
timestamp 1586364061
transform 1 0 7452 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_26_88
timestamp 1586364061
transform 1 0 9200 0 -1 16864
box -38 -48 406 592
use scs8hd_decap_12  FILLER_27_81
timestamp 1586364061
transform 1 0 8556 0 1 16864
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_167
timestamp 1586364061
transform 1 0 9568 0 -1 16864
box -38 -48 130 592
use scs8hd_decap_12  FILLER_26_93
timestamp 1586364061
transform 1 0 9660 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_93
timestamp 1586364061
transform 1 0 9660 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_26_105
timestamp 1586364061
transform 1 0 10764 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_105
timestamp 1586364061
transform 1 0 10764 0 1 16864
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_171
timestamp 1586364061
transform 1 0 12328 0 1 16864
box -38 -48 130 592
use scs8hd_decap_12  FILLER_26_117
timestamp 1586364061
transform 1 0 11868 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_27_117
timestamp 1586364061
transform 1 0 11868 0 1 16864
box -38 -48 406 592
use scs8hd_fill_1  FILLER_27_121
timestamp 1586364061
transform 1 0 12236 0 1 16864
box -38 -48 130 592
use scs8hd_decap_12  FILLER_27_123
timestamp 1586364061
transform 1 0 12420 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_26_129
timestamp 1586364061
transform 1 0 12972 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_26_141
timestamp 1586364061
transform 1 0 14076 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_135
timestamp 1586364061
transform 1 0 13524 0 1 16864
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_168
timestamp 1586364061
transform 1 0 15180 0 -1 16864
box -38 -48 130 592
use scs8hd_decap_12  FILLER_26_154
timestamp 1586364061
transform 1 0 15272 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_147
timestamp 1586364061
transform 1 0 14628 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_26_166
timestamp 1586364061
transform 1 0 16376 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_159
timestamp 1586364061
transform 1 0 15732 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_26_178
timestamp 1586364061
transform 1 0 17480 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_171
timestamp 1586364061
transform 1 0 16836 0 1 16864
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_172
timestamp 1586364061
transform 1 0 17940 0 1 16864
box -38 -48 130 592
use scs8hd_decap_12  FILLER_26_190
timestamp 1586364061
transform 1 0 18584 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_184
timestamp 1586364061
transform 1 0 18032 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_26_202
timestamp 1586364061
transform 1 0 19688 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_196
timestamp 1586364061
transform 1 0 19136 0 1 16864
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_169
timestamp 1586364061
transform 1 0 20792 0 -1 16864
box -38 -48 130 592
use scs8hd_decap_12  FILLER_26_215
timestamp 1586364061
transform 1 0 20884 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_208
timestamp 1586364061
transform 1 0 20240 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_26_227
timestamp 1586364061
transform 1 0 21988 0 -1 16864
box -38 -48 590 592
use scs8hd_decap_12  FILLER_27_220
timestamp 1586364061
transform 1 0 21344 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_3  PHY_53
timestamp 1586364061
transform -1 0 22816 0 -1 16864
box -38 -48 314 592
use scs8hd_decap_3  PHY_55
timestamp 1586364061
transform -1 0 22816 0 1 16864
box -38 -48 314 592
use scs8hd_fill_1  FILLER_27_232
timestamp 1586364061
transform 1 0 22448 0 1 16864
box -38 -48 130 592
use scs8hd_nor2_4  _162_
timestamp 1586364061
transform 1 0 1380 0 -1 17952
box -38 -48 866 592
use scs8hd_decap_3  PHY_56
timestamp 1586364061
transform 1 0 1104 0 -1 17952
box -38 -48 314 592
use scs8hd_fill_2  FILLER_28_12
timestamp 1586364061
transform 1 0 2208 0 -1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__159__B
timestamp 1586364061
transform 1 0 3312 0 -1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__157__B
timestamp 1586364061
transform 1 0 2392 0 -1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__163__B
timestamp 1586364061
transform 1 0 2760 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_16
timestamp 1586364061
transform 1 0 2576 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_4  FILLER_28_20
timestamp 1586364061
transform 1 0 2944 0 -1 17952
box -38 -48 406 592
use scs8hd_buf_1  _167_
timestamp 1586364061
transform 1 0 4048 0 -1 17952
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_173
timestamp 1586364061
transform 1 0 3956 0 -1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__142__D
timestamp 1586364061
transform 1 0 4508 0 -1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__158__B
timestamp 1586364061
transform 1 0 3772 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_3  FILLER_28_26
timestamp 1586364061
transform 1 0 3496 0 -1 17952
box -38 -48 314 592
use scs8hd_fill_2  FILLER_28_35
timestamp 1586364061
transform 1 0 4324 0 -1 17952
box -38 -48 222 592
use scs8hd_or4_4  _154_
timestamp 1586364061
transform 1 0 5060 0 -1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__154__D
timestamp 1586364061
transform 1 0 4876 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_39
timestamp 1586364061
transform 1 0 4692 0 -1 17952
box -38 -48 222 592
use scs8hd_inv_8  _062_
timestamp 1586364061
transform 1 0 6624 0 -1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__154__C
timestamp 1586364061
transform 1 0 6072 0 -1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__142__C
timestamp 1586364061
transform 1 0 6440 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_52
timestamp 1586364061
transform 1 0 5888 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_56
timestamp 1586364061
transform 1 0 6256 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_12  FILLER_28_69
timestamp 1586364061
transform 1 0 7452 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_28_81
timestamp 1586364061
transform 1 0 8556 0 -1 17952
box -38 -48 774 592
use scs8hd_decap_3  FILLER_28_89
timestamp 1586364061
transform 1 0 9292 0 -1 17952
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_174
timestamp 1586364061
transform 1 0 9568 0 -1 17952
box -38 -48 130 592
use scs8hd_decap_12  FILLER_28_93
timestamp 1586364061
transform 1 0 9660 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_105
timestamp 1586364061
transform 1 0 10764 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_117
timestamp 1586364061
transform 1 0 11868 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_129
timestamp 1586364061
transform 1 0 12972 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_141
timestamp 1586364061
transform 1 0 14076 0 -1 17952
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_175
timestamp 1586364061
transform 1 0 15180 0 -1 17952
box -38 -48 130 592
use scs8hd_decap_12  FILLER_28_154
timestamp 1586364061
transform 1 0 15272 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_166
timestamp 1586364061
transform 1 0 16376 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_178
timestamp 1586364061
transform 1 0 17480 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_190
timestamp 1586364061
transform 1 0 18584 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_202
timestamp 1586364061
transform 1 0 19688 0 -1 17952
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_176
timestamp 1586364061
transform 1 0 20792 0 -1 17952
box -38 -48 130 592
use scs8hd_decap_12  FILLER_28_215
timestamp 1586364061
transform 1 0 20884 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_28_227
timestamp 1586364061
transform 1 0 21988 0 -1 17952
box -38 -48 590 592
use scs8hd_decap_3  PHY_57
timestamp 1586364061
transform -1 0 22816 0 -1 17952
box -38 -48 314 592
use scs8hd_nor2_4  _157_
timestamp 1586364061
transform 1 0 1748 0 1 17952
box -38 -48 866 592
use scs8hd_decap_3  PHY_58
timestamp 1586364061
transform 1 0 1104 0 1 17952
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__157__A
timestamp 1586364061
transform 1 0 1564 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_3
timestamp 1586364061
transform 1 0 1380 0 1 17952
box -38 -48 222 592
use scs8hd_nor2_4  _159_
timestamp 1586364061
transform 1 0 3312 0 1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__159__A
timestamp 1586364061
transform 1 0 3128 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__156__A
timestamp 1586364061
transform 1 0 2760 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_16
timestamp 1586364061
transform 1 0 2576 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_20
timestamp 1586364061
transform 1 0 2944 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__158__A
timestamp 1586364061
transform 1 0 4324 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_33
timestamp 1586364061
transform 1 0 4140 0 1 17952
box -38 -48 222 592
use scs8hd_decap_4  FILLER_29_37
timestamp 1586364061
transform 1 0 4508 0 1 17952
box -38 -48 406 592
use scs8hd_or4_4  _148_
timestamp 1586364061
transform 1 0 5152 0 1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__148__A
timestamp 1586364061
transform 1 0 4968 0 1 17952
box -38 -48 222 592
use scs8hd_fill_1  FILLER_29_41
timestamp 1586364061
transform 1 0 4876 0 1 17952
box -38 -48 130 592
use scs8hd_buf_1  _063_
timestamp 1586364061
transform 1 0 6808 0 1 17952
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_177
timestamp 1586364061
transform 1 0 6716 0 1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__148__D
timestamp 1586364061
transform 1 0 6164 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__155__A
timestamp 1586364061
transform 1 0 6532 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_53
timestamp 1586364061
transform 1 0 5980 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_57
timestamp 1586364061
transform 1 0 6348 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__063__A
timestamp 1586364061
transform 1 0 7268 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_65
timestamp 1586364061
transform 1 0 7084 0 1 17952
box -38 -48 222 592
use scs8hd_decap_12  FILLER_29_69
timestamp 1586364061
transform 1 0 7452 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_81
timestamp 1586364061
transform 1 0 8556 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_93
timestamp 1586364061
transform 1 0 9660 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_105
timestamp 1586364061
transform 1 0 10764 0 1 17952
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_178
timestamp 1586364061
transform 1 0 12328 0 1 17952
box -38 -48 130 592
use scs8hd_decap_4  FILLER_29_117
timestamp 1586364061
transform 1 0 11868 0 1 17952
box -38 -48 406 592
use scs8hd_fill_1  FILLER_29_121
timestamp 1586364061
transform 1 0 12236 0 1 17952
box -38 -48 130 592
use scs8hd_decap_12  FILLER_29_123
timestamp 1586364061
transform 1 0 12420 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_135
timestamp 1586364061
transform 1 0 13524 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_147
timestamp 1586364061
transform 1 0 14628 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_159
timestamp 1586364061
transform 1 0 15732 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_171
timestamp 1586364061
transform 1 0 16836 0 1 17952
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_179
timestamp 1586364061
transform 1 0 17940 0 1 17952
box -38 -48 130 592
use scs8hd_decap_12  FILLER_29_184
timestamp 1586364061
transform 1 0 18032 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_196
timestamp 1586364061
transform 1 0 19136 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_208
timestamp 1586364061
transform 1 0 20240 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_220
timestamp 1586364061
transform 1 0 21344 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_3  PHY_59
timestamp 1586364061
transform -1 0 22816 0 1 17952
box -38 -48 314 592
use scs8hd_fill_1  FILLER_29_232
timestamp 1586364061
transform 1 0 22448 0 1 17952
box -38 -48 130 592
use scs8hd_nor2_4  _156_
timestamp 1586364061
transform 1 0 1656 0 -1 19040
box -38 -48 866 592
use scs8hd_decap_3  PHY_60
timestamp 1586364061
transform 1 0 1104 0 -1 19040
box -38 -48 314 592
use scs8hd_decap_3  FILLER_30_3
timestamp 1586364061
transform 1 0 1380 0 -1 19040
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__145__B
timestamp 1586364061
transform 1 0 3128 0 -1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__156__B
timestamp 1586364061
transform 1 0 2668 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_15
timestamp 1586364061
transform 1 0 2484 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_3  FILLER_30_19
timestamp 1586364061
transform 1 0 2852 0 -1 19040
box -38 -48 314 592
use scs8hd_decap_4  FILLER_30_24
timestamp 1586364061
transform 1 0 3312 0 -1 19040
box -38 -48 406 592
use scs8hd_nor2_4  _158_
timestamp 1586364061
transform 1 0 4048 0 -1 19040
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_180
timestamp 1586364061
transform 1 0 3956 0 -1 19040
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__153__B
timestamp 1586364061
transform 1 0 3772 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_1  FILLER_30_28
timestamp 1586364061
transform 1 0 3680 0 -1 19040
box -38 -48 130 592
use scs8hd_buf_1  _155_
timestamp 1586364061
transform 1 0 5612 0 -1 19040
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__148__B
timestamp 1586364061
transform 1 0 5152 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_3  FILLER_30_41
timestamp 1586364061
transform 1 0 4876 0 -1 19040
box -38 -48 314 592
use scs8hd_decap_3  FILLER_30_46
timestamp 1586364061
transform 1 0 5336 0 -1 19040
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__148__C
timestamp 1586364061
transform 1 0 6072 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_52
timestamp 1586364061
transform 1 0 5888 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_12  FILLER_30_56
timestamp 1586364061
transform 1 0 6256 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_68
timestamp 1586364061
transform 1 0 7360 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_80
timestamp 1586364061
transform 1 0 8464 0 -1 19040
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_181
timestamp 1586364061
transform 1 0 9568 0 -1 19040
box -38 -48 130 592
use scs8hd_decap_12  FILLER_30_93
timestamp 1586364061
transform 1 0 9660 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_105
timestamp 1586364061
transform 1 0 10764 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_117
timestamp 1586364061
transform 1 0 11868 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_129
timestamp 1586364061
transform 1 0 12972 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_141
timestamp 1586364061
transform 1 0 14076 0 -1 19040
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_182
timestamp 1586364061
transform 1 0 15180 0 -1 19040
box -38 -48 130 592
use scs8hd_decap_12  FILLER_30_154
timestamp 1586364061
transform 1 0 15272 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_166
timestamp 1586364061
transform 1 0 16376 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_178
timestamp 1586364061
transform 1 0 17480 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_190
timestamp 1586364061
transform 1 0 18584 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_202
timestamp 1586364061
transform 1 0 19688 0 -1 19040
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_183
timestamp 1586364061
transform 1 0 20792 0 -1 19040
box -38 -48 130 592
use scs8hd_decap_12  FILLER_30_215
timestamp 1586364061
transform 1 0 20884 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_30_227
timestamp 1586364061
transform 1 0 21988 0 -1 19040
box -38 -48 590 592
use scs8hd_decap_3  PHY_61
timestamp 1586364061
transform -1 0 22816 0 -1 19040
box -38 -48 314 592
use scs8hd_decap_3  PHY_62
timestamp 1586364061
transform 1 0 1104 0 1 19040
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__152__A
timestamp 1586364061
transform 1 0 1564 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__152__B
timestamp 1586364061
transform 1 0 1932 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_3
timestamp 1586364061
transform 1 0 1380 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_7
timestamp 1586364061
transform 1 0 1748 0 1 19040
box -38 -48 222 592
use scs8hd_decap_8  FILLER_31_11
timestamp 1586364061
transform 1 0 2116 0 1 19040
box -38 -48 774 592
use scs8hd_nor2_4  _145_
timestamp 1586364061
transform 1 0 3128 0 1 19040
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__145__A
timestamp 1586364061
transform 1 0 2944 0 1 19040
box -38 -48 222 592
use scs8hd_fill_1  FILLER_31_19
timestamp 1586364061
transform 1 0 2852 0 1 19040
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__153__A
timestamp 1586364061
transform 1 0 4508 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__140__A
timestamp 1586364061
transform 1 0 4140 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_31
timestamp 1586364061
transform 1 0 3956 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_35
timestamp 1586364061
transform 1 0 4324 0 1 19040
box -38 -48 222 592
use scs8hd_nor2_4  _140_
timestamp 1586364061
transform 1 0 4876 0 1 19040
box -38 -48 866 592
use scs8hd_fill_2  FILLER_31_39
timestamp 1586364061
transform 1 0 4692 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_50
timestamp 1586364061
transform 1 0 5704 0 1 19040
box -38 -48 222 592
use scs8hd_buf_1  _143_
timestamp 1586364061
transform 1 0 6808 0 1 19040
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_184
timestamp 1586364061
transform 1 0 6716 0 1 19040
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__140__B
timestamp 1586364061
transform 1 0 5888 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__149__A
timestamp 1586364061
transform 1 0 6256 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_54
timestamp 1586364061
transform 1 0 6072 0 1 19040
box -38 -48 222 592
use scs8hd_decap_3  FILLER_31_58
timestamp 1586364061
transform 1 0 6440 0 1 19040
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__143__A
timestamp 1586364061
transform 1 0 7268 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_65
timestamp 1586364061
transform 1 0 7084 0 1 19040
box -38 -48 222 592
use scs8hd_decap_12  FILLER_31_69
timestamp 1586364061
transform 1 0 7452 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_81
timestamp 1586364061
transform 1 0 8556 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_93
timestamp 1586364061
transform 1 0 9660 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_105
timestamp 1586364061
transform 1 0 10764 0 1 19040
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_185
timestamp 1586364061
transform 1 0 12328 0 1 19040
box -38 -48 130 592
use scs8hd_decap_4  FILLER_31_117
timestamp 1586364061
transform 1 0 11868 0 1 19040
box -38 -48 406 592
use scs8hd_fill_1  FILLER_31_121
timestamp 1586364061
transform 1 0 12236 0 1 19040
box -38 -48 130 592
use scs8hd_decap_12  FILLER_31_123
timestamp 1586364061
transform 1 0 12420 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_135
timestamp 1586364061
transform 1 0 13524 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_147
timestamp 1586364061
transform 1 0 14628 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_159
timestamp 1586364061
transform 1 0 15732 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_171
timestamp 1586364061
transform 1 0 16836 0 1 19040
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_186
timestamp 1586364061
transform 1 0 17940 0 1 19040
box -38 -48 130 592
use scs8hd_decap_12  FILLER_31_184
timestamp 1586364061
transform 1 0 18032 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_196
timestamp 1586364061
transform 1 0 19136 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_208
timestamp 1586364061
transform 1 0 20240 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_220
timestamp 1586364061
transform 1 0 21344 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_3  PHY_63
timestamp 1586364061
transform -1 0 22816 0 1 19040
box -38 -48 314 592
use scs8hd_fill_1  FILLER_31_232
timestamp 1586364061
transform 1 0 22448 0 1 19040
box -38 -48 130 592
use scs8hd_nor2_4  _152_
timestamp 1586364061
transform 1 0 1472 0 -1 20128
box -38 -48 866 592
use scs8hd_decap_3  PHY_64
timestamp 1586364061
transform 1 0 1104 0 -1 20128
box -38 -48 314 592
use scs8hd_fill_1  FILLER_32_3
timestamp 1586364061
transform 1 0 1380 0 -1 20128
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__144__A
timestamp 1586364061
transform 1 0 3036 0 -1 20128
box -38 -48 222 592
use scs8hd_decap_8  FILLER_32_13
timestamp 1586364061
transform 1 0 2300 0 -1 20128
box -38 -48 774 592
use scs8hd_decap_8  FILLER_32_23
timestamp 1586364061
transform 1 0 3220 0 -1 20128
box -38 -48 774 592
use scs8hd_nor2_4  _153_
timestamp 1586364061
transform 1 0 4508 0 -1 20128
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_187
timestamp 1586364061
transform 1 0 3956 0 -1 20128
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__146__B
timestamp 1586364061
transform 1 0 4232 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_32
timestamp 1586364061
transform 1 0 4048 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_1  FILLER_32_36
timestamp 1586364061
transform 1 0 4416 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_8  FILLER_32_46
timestamp 1586364061
transform 1 0 5336 0 -1 20128
box -38 -48 774 592
use scs8hd_buf_1  _149_
timestamp 1586364061
transform 1 0 6072 0 -1 20128
box -38 -48 314 592
use scs8hd_decap_12  FILLER_32_57
timestamp 1586364061
transform 1 0 6348 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_69
timestamp 1586364061
transform 1 0 7452 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_32_81
timestamp 1586364061
transform 1 0 8556 0 -1 20128
box -38 -48 774 592
use scs8hd_decap_3  FILLER_32_89
timestamp 1586364061
transform 1 0 9292 0 -1 20128
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_188
timestamp 1586364061
transform 1 0 9568 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_12  FILLER_32_93
timestamp 1586364061
transform 1 0 9660 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_105
timestamp 1586364061
transform 1 0 10764 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_117
timestamp 1586364061
transform 1 0 11868 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_129
timestamp 1586364061
transform 1 0 12972 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_141
timestamp 1586364061
transform 1 0 14076 0 -1 20128
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_189
timestamp 1586364061
transform 1 0 15180 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_12  FILLER_32_154
timestamp 1586364061
transform 1 0 15272 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_166
timestamp 1586364061
transform 1 0 16376 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_178
timestamp 1586364061
transform 1 0 17480 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_190
timestamp 1586364061
transform 1 0 18584 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_202
timestamp 1586364061
transform 1 0 19688 0 -1 20128
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_190
timestamp 1586364061
transform 1 0 20792 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_12  FILLER_32_215
timestamp 1586364061
transform 1 0 20884 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_32_227
timestamp 1586364061
transform 1 0 21988 0 -1 20128
box -38 -48 590 592
use scs8hd_decap_3  PHY_65
timestamp 1586364061
transform -1 0 22816 0 -1 20128
box -38 -48 314 592
use scs8hd_nor2_4  _150_
timestamp 1586364061
transform 1 0 1380 0 -1 21216
box -38 -48 866 592
use scs8hd_nor2_4  _151_
timestamp 1586364061
transform 1 0 1380 0 1 20128
box -38 -48 866 592
use scs8hd_decap_3  PHY_66
timestamp 1586364061
transform 1 0 1104 0 1 20128
box -38 -48 314 592
use scs8hd_decap_3  PHY_68
timestamp 1586364061
transform 1 0 1104 0 -1 21216
box -38 -48 314 592
use scs8hd_fill_2  FILLER_33_12
timestamp 1586364061
transform 1 0 2208 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_34_12
timestamp 1586364061
transform 1 0 2208 0 -1 21216
box -38 -48 222 592
use scs8hd_decap_4  FILLER_34_16
timestamp 1586364061
transform 1 0 2576 0 -1 21216
box -38 -48 406 592
use scs8hd_fill_2  FILLER_33_16
timestamp 1586364061
transform 1 0 2576 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__150__B
timestamp 1586364061
transform 1 0 2392 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__150__A
timestamp 1586364061
transform 1 0 2760 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__151__A
timestamp 1586364061
transform 1 0 2392 0 1 20128
box -38 -48 222 592
use scs8hd_fill_1  FILLER_34_20
timestamp 1586364061
transform 1 0 2944 0 -1 21216
box -38 -48 130 592
use scs8hd_fill_1  FILLER_33_20
timestamp 1586364061
transform 1 0 2944 0 1 20128
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__144__B
timestamp 1586364061
transform 1 0 3036 0 -1 21216
box -38 -48 222 592
use scs8hd_decap_8  FILLER_34_23
timestamp 1586364061
transform 1 0 3220 0 -1 21216
box -38 -48 774 592
use scs8hd_nor2_4  _144_
timestamp 1586364061
transform 1 0 3036 0 1 20128
box -38 -48 866 592
use scs8hd_nor2_4  _146_
timestamp 1586364061
transform 1 0 4048 0 -1 21216
box -38 -48 866 592
use scs8hd_nor2_4  _147_
timestamp 1586364061
transform 1 0 4600 0 1 20128
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_194
timestamp 1586364061
transform 1 0 3956 0 -1 21216
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__146__A
timestamp 1586364061
transform 1 0 4048 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__147__A
timestamp 1586364061
transform 1 0 4416 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_30
timestamp 1586364061
transform 1 0 3864 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_34
timestamp 1586364061
transform 1 0 4232 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__147__B
timestamp 1586364061
transform 1 0 5060 0 -1 21216
box -38 -48 222 592
use scs8hd_decap_12  FILLER_33_47
timestamp 1586364061
transform 1 0 5428 0 1 20128
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_34_41
timestamp 1586364061
transform 1 0 4876 0 -1 21216
box -38 -48 222 592
use scs8hd_decap_12  FILLER_34_45
timestamp 1586364061
transform 1 0 5244 0 -1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_191
timestamp 1586364061
transform 1 0 6716 0 1 20128
box -38 -48 130 592
use scs8hd_fill_2  FILLER_33_59
timestamp 1586364061
transform 1 0 6532 0 1 20128
box -38 -48 222 592
use scs8hd_decap_12  FILLER_33_62
timestamp 1586364061
transform 1 0 6808 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_57
timestamp 1586364061
transform 1 0 6348 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_74
timestamp 1586364061
transform 1 0 7912 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_69
timestamp 1586364061
transform 1 0 7452 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_86
timestamp 1586364061
transform 1 0 9016 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_34_81
timestamp 1586364061
transform 1 0 8556 0 -1 21216
box -38 -48 774 592
use scs8hd_decap_3  FILLER_34_89
timestamp 1586364061
transform 1 0 9292 0 -1 21216
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_195
timestamp 1586364061
transform 1 0 9568 0 -1 21216
box -38 -48 130 592
use scs8hd_decap_12  FILLER_33_98
timestamp 1586364061
transform 1 0 10120 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_93
timestamp 1586364061
transform 1 0 9660 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_110
timestamp 1586364061
transform 1 0 11224 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_105
timestamp 1586364061
transform 1 0 10764 0 -1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_192
timestamp 1586364061
transform 1 0 12328 0 1 20128
box -38 -48 130 592
use scs8hd_decap_12  FILLER_33_123
timestamp 1586364061
transform 1 0 12420 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_117
timestamp 1586364061
transform 1 0 11868 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_135
timestamp 1586364061
transform 1 0 13524 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_129
timestamp 1586364061
transform 1 0 12972 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_141
timestamp 1586364061
transform 1 0 14076 0 -1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_196
timestamp 1586364061
transform 1 0 15180 0 -1 21216
box -38 -48 130 592
use scs8hd_decap_12  FILLER_33_147
timestamp 1586364061
transform 1 0 14628 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_154
timestamp 1586364061
transform 1 0 15272 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_159
timestamp 1586364061
transform 1 0 15732 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_166
timestamp 1586364061
transform 1 0 16376 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_171
timestamp 1586364061
transform 1 0 16836 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_178
timestamp 1586364061
transform 1 0 17480 0 -1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_193
timestamp 1586364061
transform 1 0 17940 0 1 20128
box -38 -48 130 592
use scs8hd_decap_12  FILLER_33_184
timestamp 1586364061
transform 1 0 18032 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_190
timestamp 1586364061
transform 1 0 18584 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_196
timestamp 1586364061
transform 1 0 19136 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_202
timestamp 1586364061
transform 1 0 19688 0 -1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_197
timestamp 1586364061
transform 1 0 20792 0 -1 21216
box -38 -48 130 592
use scs8hd_decap_12  FILLER_33_208
timestamp 1586364061
transform 1 0 20240 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_215
timestamp 1586364061
transform 1 0 20884 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_220
timestamp 1586364061
transform 1 0 21344 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_34_227
timestamp 1586364061
transform 1 0 21988 0 -1 21216
box -38 -48 590 592
use scs8hd_decap_3  PHY_67
timestamp 1586364061
transform -1 0 22816 0 1 20128
box -38 -48 314 592
use scs8hd_decap_3  PHY_69
timestamp 1586364061
transform -1 0 22816 0 -1 21216
box -38 -48 314 592
use scs8hd_fill_1  FILLER_33_232
timestamp 1586364061
transform 1 0 22448 0 1 20128
box -38 -48 130 592
use scs8hd_decap_3  PHY_70
timestamp 1586364061
transform 1 0 1104 0 1 21216
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__151__B
timestamp 1586364061
transform 1 0 1564 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_3
timestamp 1586364061
transform 1 0 1380 0 1 21216
box -38 -48 222 592
use scs8hd_decap_12  FILLER_35_7
timestamp 1586364061
transform 1 0 1748 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_19
timestamp 1586364061
transform 1 0 2852 0 1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_198
timestamp 1586364061
transform 1 0 3956 0 1 21216
box -38 -48 130 592
use scs8hd_decap_12  FILLER_35_32
timestamp 1586364061
transform 1 0 4048 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_44
timestamp 1586364061
transform 1 0 5152 0 1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_199
timestamp 1586364061
transform 1 0 6808 0 1 21216
box -38 -48 130 592
use scs8hd_decap_6  FILLER_35_56
timestamp 1586364061
transform 1 0 6256 0 1 21216
box -38 -48 590 592
use scs8hd_decap_12  FILLER_35_63
timestamp 1586364061
transform 1 0 6900 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_75
timestamp 1586364061
transform 1 0 8004 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_35_87
timestamp 1586364061
transform 1 0 9108 0 1 21216
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_200
timestamp 1586364061
transform 1 0 9660 0 1 21216
box -38 -48 130 592
use scs8hd_decap_12  FILLER_35_94
timestamp 1586364061
transform 1 0 9752 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_106
timestamp 1586364061
transform 1 0 10856 0 1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_201
timestamp 1586364061
transform 1 0 12512 0 1 21216
box -38 -48 130 592
use scs8hd_decap_6  FILLER_35_118
timestamp 1586364061
transform 1 0 11960 0 1 21216
box -38 -48 590 592
use scs8hd_decap_12  FILLER_35_125
timestamp 1586364061
transform 1 0 12604 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_137
timestamp 1586364061
transform 1 0 13708 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_35_149
timestamp 1586364061
transform 1 0 14812 0 1 21216
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_202
timestamp 1586364061
transform 1 0 15364 0 1 21216
box -38 -48 130 592
use scs8hd_decap_12  FILLER_35_156
timestamp 1586364061
transform 1 0 15456 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_168
timestamp 1586364061
transform 1 0 16560 0 1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_203
timestamp 1586364061
transform 1 0 18216 0 1 21216
box -38 -48 130 592
use scs8hd_decap_6  FILLER_35_180
timestamp 1586364061
transform 1 0 17664 0 1 21216
box -38 -48 590 592
use scs8hd_decap_12  FILLER_35_187
timestamp 1586364061
transform 1 0 18308 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_199
timestamp 1586364061
transform 1 0 19412 0 1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_204
timestamp 1586364061
transform 1 0 21068 0 1 21216
box -38 -48 130 592
use scs8hd_decap_6  FILLER_35_211
timestamp 1586364061
transform 1 0 20516 0 1 21216
box -38 -48 590 592
use scs8hd_decap_12  FILLER_35_218
timestamp 1586364061
transform 1 0 21160 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_35_230
timestamp 1586364061
transform 1 0 22264 0 1 21216
box -38 -48 314 592
use scs8hd_decap_3  PHY_71
timestamp 1586364061
transform -1 0 22816 0 1 21216
box -38 -48 314 592
<< labels >>
rlabel metal2 s 1950 23520 2006 24000 6 address[0]
port 0 nsew default input
rlabel metal2 s 5906 23520 5962 24000 6 address[1]
port 1 nsew default input
rlabel metal2 s 9954 23520 10010 24000 6 address[2]
port 2 nsew default input
rlabel metal2 s 13910 23520 13966 24000 6 address[3]
port 3 nsew default input
rlabel metal2 s 17958 23520 18014 24000 6 address[4]
port 4 nsew default input
rlabel metal2 s 21914 23520 21970 24000 6 address[5]
port 5 nsew default input
rlabel metal3 s 0 144 480 264 6 data_out[0]
port 6 nsew default tristate
rlabel metal3 s 0 3952 480 4072 6 data_out[10]
port 7 nsew default tristate
rlabel metal3 s 0 4360 480 4480 6 data_out[11]
port 8 nsew default tristate
rlabel metal3 s 0 4768 480 4888 6 data_out[12]
port 9 nsew default tristate
rlabel metal3 s 0 5176 480 5296 6 data_out[13]
port 10 nsew default tristate
rlabel metal3 s 0 5584 480 5704 6 data_out[14]
port 11 nsew default tristate
rlabel metal3 s 0 5992 480 6112 6 data_out[15]
port 12 nsew default tristate
rlabel metal3 s 0 6400 480 6520 6 data_out[16]
port 13 nsew default tristate
rlabel metal3 s 0 6808 480 6928 6 data_out[17]
port 14 nsew default tristate
rlabel metal3 s 0 7080 480 7200 6 data_out[18]
port 15 nsew default tristate
rlabel metal3 s 0 7488 480 7608 6 data_out[19]
port 16 nsew default tristate
rlabel metal3 s 0 416 480 536 6 data_out[1]
port 17 nsew default tristate
rlabel metal3 s 0 7896 480 8016 6 data_out[20]
port 18 nsew default tristate
rlabel metal3 s 0 8304 480 8424 6 data_out[21]
port 19 nsew default tristate
rlabel metal3 s 0 8712 480 8832 6 data_out[22]
port 20 nsew default tristate
rlabel metal3 s 0 9120 480 9240 6 data_out[23]
port 21 nsew default tristate
rlabel metal3 s 0 9528 480 9648 6 data_out[24]
port 22 nsew default tristate
rlabel metal3 s 0 9936 480 10056 6 data_out[25]
port 23 nsew default tristate
rlabel metal3 s 0 10344 480 10464 6 data_out[26]
port 24 nsew default tristate
rlabel metal3 s 0 10616 480 10736 6 data_out[27]
port 25 nsew default tristate
rlabel metal3 s 0 11024 480 11144 6 data_out[28]
port 26 nsew default tristate
rlabel metal3 s 0 11432 480 11552 6 data_out[29]
port 27 nsew default tristate
rlabel metal3 s 0 824 480 944 6 data_out[2]
port 28 nsew default tristate
rlabel metal3 s 0 11840 480 11960 6 data_out[30]
port 29 nsew default tristate
rlabel metal3 s 0 12248 480 12368 6 data_out[31]
port 30 nsew default tristate
rlabel metal3 s 0 12656 480 12776 6 data_out[32]
port 31 nsew default tristate
rlabel metal3 s 0 13064 480 13184 6 data_out[33]
port 32 nsew default tristate
rlabel metal3 s 0 13472 480 13592 6 data_out[34]
port 33 nsew default tristate
rlabel metal3 s 0 13744 480 13864 6 data_out[35]
port 34 nsew default tristate
rlabel metal3 s 0 14152 480 14272 6 data_out[36]
port 35 nsew default tristate
rlabel metal3 s 0 14560 480 14680 6 data_out[37]
port 36 nsew default tristate
rlabel metal3 s 0 14968 480 15088 6 data_out[38]
port 37 nsew default tristate
rlabel metal3 s 0 15376 480 15496 6 data_out[39]
port 38 nsew default tristate
rlabel metal3 s 0 1232 480 1352 6 data_out[3]
port 39 nsew default tristate
rlabel metal3 s 0 15784 480 15904 6 data_out[40]
port 40 nsew default tristate
rlabel metal3 s 0 16192 480 16312 6 data_out[41]
port 41 nsew default tristate
rlabel metal3 s 0 16600 480 16720 6 data_out[42]
port 42 nsew default tristate
rlabel metal3 s 0 17008 480 17128 6 data_out[43]
port 43 nsew default tristate
rlabel metal3 s 0 17280 480 17400 6 data_out[44]
port 44 nsew default tristate
rlabel metal3 s 0 17688 480 17808 6 data_out[45]
port 45 nsew default tristate
rlabel metal3 s 0 18096 480 18216 6 data_out[46]
port 46 nsew default tristate
rlabel metal3 s 0 18504 480 18624 6 data_out[47]
port 47 nsew default tristate
rlabel metal3 s 0 18912 480 19032 6 data_out[48]
port 48 nsew default tristate
rlabel metal3 s 0 19320 480 19440 6 data_out[49]
port 49 nsew default tristate
rlabel metal3 s 0 1640 480 1760 6 data_out[4]
port 50 nsew default tristate
rlabel metal3 s 0 19728 480 19848 6 data_out[50]
port 51 nsew default tristate
rlabel metal3 s 0 20136 480 20256 6 data_out[51]
port 52 nsew default tristate
rlabel metal3 s 0 20544 480 20664 6 data_out[52]
port 53 nsew default tristate
rlabel metal3 s 0 20816 480 20936 6 data_out[53]
port 54 nsew default tristate
rlabel metal3 s 0 21224 480 21344 6 data_out[54]
port 55 nsew default tristate
rlabel metal3 s 0 21632 480 21752 6 data_out[55]
port 56 nsew default tristate
rlabel metal3 s 0 22040 480 22160 6 data_out[56]
port 57 nsew default tristate
rlabel metal3 s 0 22448 480 22568 6 data_out[57]
port 58 nsew default tristate
rlabel metal3 s 0 22856 480 22976 6 data_out[58]
port 59 nsew default tristate
rlabel metal3 s 0 23264 480 23384 6 data_out[59]
port 60 nsew default tristate
rlabel metal3 s 0 2048 480 2168 6 data_out[5]
port 61 nsew default tristate
rlabel metal3 s 0 23672 480 23792 6 data_out[60]
port 62 nsew default tristate
rlabel metal3 s 0 2456 480 2576 6 data_out[6]
port 63 nsew default tristate
rlabel metal3 s 0 2864 480 2984 6 data_out[7]
port 64 nsew default tristate
rlabel metal3 s 0 3272 480 3392 6 data_out[8]
port 65 nsew default tristate
rlabel metal3 s 0 3544 480 3664 6 data_out[9]
port 66 nsew default tristate
rlabel metal2 s 11978 0 12034 480 6 enable
port 67 nsew default input
rlabel metal4 s 4944 2128 5264 21808 6 vpwr
port 68 nsew default input
rlabel metal4 s 8944 2128 9264 21808 6 vgnd
port 69 nsew default input
<< end >>
