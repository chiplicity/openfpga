* NGSPICE file created from sb_0__2_.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_12 abstract view
.subckt sky130_fd_sc_hd__decap_12 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A X VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxbp_1 abstract view
.subckt sky130_fd_sc_hd__dfxbp_1 D Q Q_N CLK VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S X VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_1 abstract view
.subckt sky130_fd_sc_hd__buf_1 A X VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
.subckt sky130_fd_sc_hd__conb_1 HI LO VGND VNB VPB VPWR
.ends

.subckt sb_0__2_ bottom_left_grid_pin_1_ ccff_head ccff_tail chanx_right_in[0] chanx_right_in[10]
+ chanx_right_in[11] chanx_right_in[12] chanx_right_in[13] chanx_right_in[14] chanx_right_in[15]
+ chanx_right_in[16] chanx_right_in[17] chanx_right_in[18] chanx_right_in[19] chanx_right_in[1]
+ chanx_right_in[2] chanx_right_in[3] chanx_right_in[4] chanx_right_in[5] chanx_right_in[6]
+ chanx_right_in[7] chanx_right_in[8] chanx_right_in[9] chanx_right_out[0] chanx_right_out[10]
+ chanx_right_out[11] chanx_right_out[12] chanx_right_out[13] chanx_right_out[14]
+ chanx_right_out[15] chanx_right_out[16] chanx_right_out[17] chanx_right_out[18]
+ chanx_right_out[19] chanx_right_out[1] chanx_right_out[2] chanx_right_out[3] chanx_right_out[4]
+ chanx_right_out[5] chanx_right_out[6] chanx_right_out[7] chanx_right_out[8] chanx_right_out[9]
+ chany_bottom_in[0] chany_bottom_in[10] chany_bottom_in[11] chany_bottom_in[12] chany_bottom_in[13]
+ chany_bottom_in[14] chany_bottom_in[15] chany_bottom_in[16] chany_bottom_in[17]
+ chany_bottom_in[18] chany_bottom_in[19] chany_bottom_in[1] chany_bottom_in[2] chany_bottom_in[3]
+ chany_bottom_in[4] chany_bottom_in[5] chany_bottom_in[6] chany_bottom_in[7] chany_bottom_in[8]
+ chany_bottom_in[9] chany_bottom_out[0] chany_bottom_out[10] chany_bottom_out[11]
+ chany_bottom_out[12] chany_bottom_out[13] chany_bottom_out[14] chany_bottom_out[15]
+ chany_bottom_out[16] chany_bottom_out[17] chany_bottom_out[18] chany_bottom_out[19]
+ chany_bottom_out[1] chany_bottom_out[2] chany_bottom_out[3] chany_bottom_out[4]
+ chany_bottom_out[5] chany_bottom_out[6] chany_bottom_out[7] chany_bottom_out[8]
+ chany_bottom_out[9] prog_clk right_top_grid_pin_1_ VPWR VGND
XFILLER_13_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mem_bottom_track_1.sky130_fd_sc_hd__dfxbp_1_1__D mux_bottom_track_1.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_right_track_4.mux_l1_in_0__A1 right_top_grid_pin_1_ VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_15_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_49_ chany_bottom_in[3] chanx_right_out[15] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_20_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_48_ chany_bottom_in[2] chanx_right_out[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_20_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mem_bottom_track_9.sky130_fd_sc_hd__dfxbp_1_1__CLK prog_clk VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mem_right_track_0.sky130_fd_sc_hd__dfxbp_1_1__CLK prog_clk VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_47_ chany_bottom_in[1] chanx_right_out[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_20_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmem_bottom_track_5.sky130_fd_sc_hd__dfxbp_1_1_ mux_bottom_track_5.mux_l1_in_0_/S
+ mux_bottom_track_5.mux_l2_in_0_/S mem_bottom_track_5.sky130_fd_sc_hd__dfxbp_1_1_/Q_N
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_18_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mem_right_track_24.sky130_fd_sc_hd__dfxbp_1_1__CLK prog_clk VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_46_ chany_bottom_in[0] chanx_right_out[18] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
Xmem_bottom_track_5.sky130_fd_sc_hd__dfxbp_1_0_ mux_bottom_track_1.mux_l2_in_0_/S
+ mux_bottom_track_5.mux_l1_in_0_/S mem_bottom_track_5.sky130_fd_sc_hd__dfxbp_1_0_/Q_N
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_18_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_29_ chanx_right_in[3] chany_bottom_out[15] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_4_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__20__A _20_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_mux_bottom_track_5.sky130_fd_sc_hd__buf_4_0__A mux_bottom_track_5.mux_l2_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_45_ chany_bottom_in[19] chanx_right_out[19] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_20_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__23__A chany_bottom_in[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28_ chanx_right_in[2] chany_bottom_out[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_37_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__18__A chany_bottom_in[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_right_track_8.mux_l2_in_0_ _15_/HI mux_right_track_8.mux_l1_in_0_/X mux_right_track_8.mux_l2_in_0_/S
+ mux_right_track_8.mux_l2_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_24_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__31__A chanx_right_in[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_bottom_track_9.mux_l2_in_0__S mux_bottom_track_9.mux_l2_in_0_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__26__A chanx_right_in[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mem_bottom_track_5.sky130_fd_sc_hd__dfxbp_1_0__D mux_bottom_track_1.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_44_ _44_/A chany_bottom_out[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_20_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_mem_right_track_4.sky130_fd_sc_hd__dfxbp_1_1__CLK prog_clk VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_27_ chanx_right_in[1] chany_bottom_out[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_20_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__34__A chanx_right_in[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__29__A chanx_right_in[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_0 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mux_bottom_track_25.mux_l1_in_0__A0 bottom_left_grid_pin_1_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_right_track_8.mux_l1_in_0_ chany_bottom_in[14] right_top_grid_pin_1_ mux_right_track_8.mux_l1_in_0_/S
+ mux_right_track_8.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_12_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__42__A _42_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_bottom_track_9.mux_l2_in_0__A0 _11_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mem_bottom_track_1.sky130_fd_sc_hd__dfxbp_1_0__CLK prog_clk VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_right_track_8.sky130_fd_sc_hd__buf_4_0_ mux_right_track_8.mux_l2_in_0_/X _20_/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_1
XANTENNA__37__A chanx_right_in[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_43_ chanx_right_in[17] chany_bottom_out[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_1_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_26_ chanx_right_in[0] chany_bottom_out[18] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_37_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mux_right_track_0.sky130_fd_sc_hd__buf_4_0__A mux_right_track_0.mux_l2_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__50__A chany_bottom_in[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09_ _09_/HI _09_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XFILLER_40_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__45__A chany_bottom_in[19] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mux_bottom_track_25.mux_l1_in_0__A1 chanx_right_in[6] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_12_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_right_track_24.mux_l2_in_0__A0 _13_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_bottom_track_9.mux_l2_in_0__A1 mux_bottom_track_9.mux_l1_in_0_/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_bottom_track_5.mux_l2_in_0__S mux_bottom_track_5.mux_l2_in_0_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__53__A chany_bottom_in[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_bottom_track_25.mux_l2_in_0_ _09_/HI mux_bottom_track_25.mux_l1_in_0_/X ccff_tail
+ mux_bottom_track_25.mux_l2_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
X_42_ _42_/A chany_bottom_out[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_18_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__48__A chany_bottom_in[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25_ chanx_right_in[19] chany_bottom_out[19] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_37_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmux_bottom_track_9.mux_l2_in_0_ _11_/HI mux_bottom_track_9.mux_l1_in_0_/X mux_bottom_track_9.mux_l2_in_0_/S
+ mux_bottom_track_9.mux_l2_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_34_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08_ _08_/HI _08_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XFILLER_33_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_mux_right_track_0.mux_l1_in_0__A0 chany_bottom_in[18] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_39_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_mux_right_track_24.mux_l2_in_0__A1 mux_right_track_24.mux_l1_in_0_/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_41_ chanx_right_in[15] chany_bottom_out[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_1_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mem_right_track_8.sky130_fd_sc_hd__dfxbp_1_1__CLK prog_clk VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
X_24_ _24_/A chanx_right_out[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_37_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_bottom_track_25.mux_l1_in_0_ bottom_left_grid_pin_1_ chanx_right_in[6] mux_bottom_track_25.mux_l1_in_0_/S
+ mux_bottom_track_25.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_3_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_mux_right_track_0.mux_l1_in_0__A1 right_top_grid_pin_1_ VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XPHY_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_bottom_track_9.mux_l1_in_0_ bottom_left_grid_pin_1_ chanx_right_in[14] mux_bottom_track_9.mux_l1_in_0_/S
+ mux_bottom_track_9.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_42_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_bottom_track_9.sky130_fd_sc_hd__buf_4_0_ mux_bottom_track_9.mux_l2_in_0_/X _40_/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_1
XFILLER_35_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_right_track_24.mux_l1_in_0__S mux_right_track_24.mux_l1_in_0_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_40_ _40_/A chany_bottom_out[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_1_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mem_bottom_track_5.sky130_fd_sc_hd__dfxbp_1_0__CLK prog_clk VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmem_right_track_0.sky130_fd_sc_hd__dfxbp_1_1_ mux_right_track_0.mux_l1_in_0_/S mux_right_track_0.mux_l2_in_0_/S
+ mem_right_track_0.sky130_fd_sc_hd__dfxbp_1_1_/Q_N prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_40_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_bottom_track_1.mux_l2_in_0__S mux_bottom_track_1.mux_l2_in_0_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23_ chany_bottom_in[17] chanx_right_out[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_37_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mem_right_track_4.sky130_fd_sc_hd__dfxbp_1_1__D mux_right_track_4.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_bottom_track_25.mux_l2_in_0__S ccff_tail VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_right_track_0.sky130_fd_sc_hd__dfxbp_1_0_ ccff_head mux_right_track_0.mux_l1_in_0_/S
+ mem_right_track_0.sky130_fd_sc_hd__dfxbp_1_0_/Q_N prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
X_22_ _22_/A chanx_right_out[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_3_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_right_track_8.mux_l2_in_0__S mux_right_track_8.mux_l2_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mem_bottom_track_25.sky130_fd_sc_hd__dfxbp_1_1__D mux_bottom_track_25.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_right_track_4.mux_l2_in_0_ _14_/HI mux_right_track_4.mux_l1_in_0_/X mux_right_track_4.mux_l2_in_0_/S
+ mux_right_track_4.mux_l2_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
X_21_ chany_bottom_in[15] chanx_right_out[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_10_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmem_right_track_24.sky130_fd_sc_hd__dfxbp_1_1_ mux_right_track_24.mux_l1_in_0_/S
+ mux_right_track_24.mux_l2_in_0_/S mem_right_track_24.sky130_fd_sc_hd__dfxbp_1_1_/Q_N
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XPHY_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20_ _20_/A chanx_right_out[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XANTENNA_mem_bottom_track_9.sky130_fd_sc_hd__dfxbp_1_0__CLK prog_clk VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_right_track_4.mux_l1_in_0_ chany_bottom_in[16] right_top_grid_pin_1_ mux_right_track_4.mux_l1_in_0_/S
+ mux_right_track_4.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XPHY_116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmux_right_track_4.sky130_fd_sc_hd__buf_4_0_ mux_right_track_4.mux_l2_in_0_/X _22_/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_1
XFILLER_24_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmem_right_track_24.sky130_fd_sc_hd__dfxbp_1_0_ mux_right_track_8.mux_l2_in_0_/S mux_right_track_24.mux_l1_in_0_/S
+ mem_right_track_24.sky130_fd_sc_hd__dfxbp_1_0_/Q_N prog_clk VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__dfxbp_1
XPHY_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_right_track_4.mux_l2_in_0__S mux_right_track_4.mux_l2_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_right_track_24.sky130_fd_sc_hd__buf_4_0__A mux_right_track_24.mux_l2_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mem_right_track_0.sky130_fd_sc_hd__dfxbp_1_0__CLK prog_clk VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmem_bottom_track_1.sky130_fd_sc_hd__dfxbp_1_1_ mux_bottom_track_1.mux_l1_in_0_/S
+ mux_bottom_track_1.mux_l2_in_0_/S mem_bottom_track_1.sky130_fd_sc_hd__dfxbp_1_1_/Q_N
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_24_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_bottom_track_9.mux_l1_in_0__S mux_bottom_track_9.mux_l1_in_0_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_right_track_24.sky130_fd_sc_hd__dfxbp_1_0__CLK prog_clk VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_bottom_track_5.mux_l2_in_0_ _10_/HI mux_bottom_track_5.mux_l1_in_0_/X mux_bottom_track_5.mux_l2_in_0_/S
+ mux_bottom_track_5.mux_l2_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_9_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmem_bottom_track_1.sky130_fd_sc_hd__dfxbp_1_0_ mux_right_track_24.mux_l2_in_0_/S
+ mux_bottom_track_1.mux_l1_in_0_/S mem_bottom_track_1.sky130_fd_sc_hd__dfxbp_1_0_/Q_N
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_40_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mem_right_track_8.sky130_fd_sc_hd__dfxbp_1_0__D mux_right_track_4.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_bottom_track_5.mux_l2_in_0__A0 _10_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_bottom_track_1.sky130_fd_sc_hd__buf_4_0__A mux_bottom_track_1.mux_l2_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_right_track_0.mux_l2_in_0__S mux_right_track_0.mux_l2_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_bottom_track_5.sky130_fd_sc_hd__buf_4_0_ mux_bottom_track_5.mux_l2_in_0_/X _42_/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_1
XFILLER_39_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_bottom_track_5.mux_l1_in_0_ bottom_left_grid_pin_1_ chanx_right_in[16] mux_bottom_track_5.mux_l1_in_0_/S
+ mux_bottom_track_5.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_42_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_bottom_track_5.mux_l2_in_0__A1 mux_bottom_track_5.mux_l1_in_0_/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_right_track_8.mux_l2_in_0__A0 _15_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21__A chany_bottom_in[15] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mem_right_track_0.sky130_fd_sc_hd__dfxbp_1_0__D ccff_head VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__16__A chany_bottom_in[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mem_right_track_24.sky130_fd_sc_hd__dfxbp_1_0__D mux_right_track_8.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_mem_right_track_4.sky130_fd_sc_hd__dfxbp_1_0__CLK prog_clk VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_bottom_track_5.mux_l1_in_0__S mux_bottom_track_5.mux_l1_in_0_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24__A _24_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19__A chany_bottom_in[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_right_track_8.mux_l2_in_0__A1 mux_right_track_8.mux_l1_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_bottom_track_9.mux_l1_in_0__A0 bottom_left_grid_pin_1_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__32__A _32_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__27__A chanx_right_in[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_bottom_track_5.sky130_fd_sc_hd__dfxbp_1_1__D mux_bottom_track_5.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__40__A _40_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_90 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_mux_right_track_24.mux_l1_in_0__A0 chany_bottom_in[6] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_21_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__35__A chanx_right_in[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_bottom_track_9.mux_l1_in_0__A1 chanx_right_in[14] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_16_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_right_track_0.mux_l2_in_0_ _12_/HI mux_right_track_0.mux_l1_in_0_/X mux_right_track_0.mux_l2_in_0_/S
+ mux_right_track_0.mux_l2_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_16_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__43__A chanx_right_in[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__38__A chanx_right_in[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_bottom_track_1.mux_l1_in_0__S mux_bottom_track_1.mux_l1_in_0_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_91 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_mux_right_track_24.mux_l1_in_0__A1 right_top_grid_pin_1_ VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_24_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__51__A chany_bottom_in[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_bottom_track_25.mux_l1_in_0__S mux_bottom_track_25.mux_l1_in_0_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__46__A chany_bottom_in[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_bottom_track_25.sky130_fd_sc_hd__dfxbp_1_1__CLK prog_clk VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XPHY_261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmux_right_track_0.sky130_fd_sc_hd__buf_4_0_ mux_right_track_0.mux_l2_in_0_/X _24_/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_1
XFILLER_13_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmux_right_track_0.mux_l1_in_0_ chany_bottom_in[18] right_top_grid_pin_1_ mux_right_track_0.mux_l1_in_0_/S
+ mux_right_track_0.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_24_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_right_track_24.mux_l2_in_0_ _13_/HI mux_right_track_24.mux_l1_in_0_/X mux_right_track_24.mux_l2_in_0_/S
+ mux_right_track_24.mux_l2_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA__54__A chany_bottom_in[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mem_right_track_8.sky130_fd_sc_hd__dfxbp_1_0__CLK prog_clk VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__49__A chany_bottom_in[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_92 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_39_ chanx_right_in[13] chany_bottom_out[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_37_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mux_right_track_8.mux_l1_in_0__S mux_right_track_8.mux_l1_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_right_track_8.sky130_fd_sc_hd__buf_4_0__A mux_right_track_8.mux_l2_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_93 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_55_ chany_bottom_in[9] chanx_right_out[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
Xmux_right_track_24.mux_l1_in_0_ chany_bottom_in[6] right_top_grid_pin_1_ mux_right_track_24.mux_l1_in_0_/S
+ mux_right_track_24.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_24_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_42_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_38_ chanx_right_in[12] chany_bottom_out[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_37_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_bottom_track_1.mux_l2_in_0_ _08_/HI mux_bottom_track_1.mux_l1_in_0_/X mux_bottom_track_1.mux_l2_in_0_/S
+ mux_bottom_track_1.mux_l2_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_7_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_94 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_54_ chany_bottom_in[8] chanx_right_out[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_17_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_37_ chanx_right_in[11] chany_bottom_out[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_20_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_bottom_track_1.sky130_fd_sc_hd__buf_4_0_ mux_bottom_track_1.mux_l2_in_0_/X _44_/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_1
XFILLER_11_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_right_track_4.mux_l1_in_0__S mux_right_track_4.mux_l1_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_bottom_track_1.mux_l1_in_0_ bottom_left_grid_pin_1_ chanx_right_in[18] mux_bottom_track_1.mux_l1_in_0_/S
+ mux_bottom_track_1.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_0_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mem_bottom_track_9.sky130_fd_sc_hd__dfxbp_1_0__D mux_bottom_track_5.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_95 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_53_ chany_bottom_in[7] chanx_right_out[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_2_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_36_ chanx_right_in[10] chany_bottom_out[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_28_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_19_ chany_bottom_in[13] chanx_right_out[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_17_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_bottom_track_1.mux_l2_in_0__A0 _08_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_right_track_8.sky130_fd_sc_hd__dfxbp_1_1_ mux_right_track_8.mux_l1_in_0_/S mux_right_track_8.mux_l2_in_0_/S
+ mem_right_track_8.sky130_fd_sc_hd__dfxbp_1_1_/Q_N prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_0_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_96 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_52_ _52_/A chanx_right_out[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_2_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mem_bottom_track_1.sky130_fd_sc_hd__dfxbp_1_0__D mux_right_track_24.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_35_ chanx_right_in[9] chany_bottom_out[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_37_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18_ chany_bottom_in[12] chanx_right_out[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_31_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_right_track_8.sky130_fd_sc_hd__dfxbp_1_0_ mux_right_track_4.mux_l2_in_0_/S mux_right_track_8.mux_l1_in_0_/S
+ mem_right_track_8.sky130_fd_sc_hd__dfxbp_1_0_/Q_N prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_0_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_bottom_track_1.mux_l2_in_0__A1 mux_bottom_track_1.mux_l1_in_0_/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_track_0.mux_l1_in_0__S mux_right_track_0.mux_l1_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_4.mux_l2_in_0__A0 _14_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmem_bottom_track_25.sky130_fd_sc_hd__dfxbp_1_1_ mux_bottom_track_25.mux_l1_in_0_/S
+ ccff_tail mem_bottom_track_25.sky130_fd_sc_hd__dfxbp_1_1_/Q_N prog_clk VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_27_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_97 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_86 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_51_ chany_bottom_in[5] chanx_right_out[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_2_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_34_ chanx_right_in[8] chany_bottom_out[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_37_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_17_ chany_bottom_in[11] chanx_right_out[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_33_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_right_track_4.mux_l2_in_0__A1 mux_right_track_4.mux_l1_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_bottom_track_5.mux_l1_in_0__A0 bottom_left_grid_pin_1_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmem_bottom_track_25.sky130_fd_sc_hd__dfxbp_1_0_ mux_bottom_track_9.mux_l2_in_0_/S
+ mux_bottom_track_25.mux_l1_in_0_/S mem_bottom_track_25.sky130_fd_sc_hd__dfxbp_1_0_/Q_N
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_4_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_98 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_87 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_50_ chany_bottom_in[4] chanx_right_out[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_17_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_33_ chanx_right_in[7] chany_bottom_out[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_9_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_16_ chany_bottom_in[10] chanx_right_out[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_26_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_bottom_track_5.mux_l1_in_0__A1 chanx_right_in[16] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_29_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_right_track_8.mux_l1_in_0__A0 chany_bottom_in[14] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_26_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_99 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_88 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_32_ _32_/A chany_bottom_out[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_20_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_right_track_8.sky130_fd_sc_hd__dfxbp_1_1__D mux_right_track_8.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15_ _15_/HI _15_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XFILLER_25_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmem_bottom_track_9.sky130_fd_sc_hd__dfxbp_1_1_ mux_bottom_track_9.mux_l1_in_0_/S
+ mux_bottom_track_9.mux_l2_in_0_/S mem_bottom_track_9.sky130_fd_sc_hd__dfxbp_1_1_/Q_N
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_28_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_bottom_track_25.sky130_fd_sc_hd__buf_4_0_ mux_bottom_track_25.mux_l2_in_0_/X
+ _32_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_1
XFILLER_38_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_right_track_8.mux_l1_in_0__A1 right_top_grid_pin_1_ VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_6_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_89 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_31_ chanx_right_in[5] chany_bottom_out[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_20_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14_ _14_/HI _14_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XFILLER_33_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__22__A _22_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mem_right_track_0.sky130_fd_sc_hd__dfxbp_1_1__D mux_right_track_0.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_right_track_24.sky130_fd_sc_hd__buf_4_0_ mux_right_track_24.mux_l2_in_0_/X _52_/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_1
XFILLER_15_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmem_bottom_track_9.sky130_fd_sc_hd__dfxbp_1_0_ mux_bottom_track_5.mux_l2_in_0_/S
+ mux_bottom_track_9.mux_l1_in_0_/S mem_bottom_track_9.sky130_fd_sc_hd__dfxbp_1_0_/Q_N
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_21_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__17__A chany_bottom_in[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mem_right_track_24.sky130_fd_sc_hd__dfxbp_1_1__D mux_right_track_24.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_bottom_track_9.sky130_fd_sc_hd__buf_4_0__A mux_bottom_track_9.mux_l2_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__30__A chanx_right_in[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__25__A chanx_right_in[19] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_30_ chanx_right_in[4] chany_bottom_out[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_13_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13_ _13_/HI _13_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XFILLER_33_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__33__A chanx_right_in[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__28__A chanx_right_in[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__41__A chanx_right_in[15] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__36__A chanx_right_in[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12_ _12_/HI _12_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XFILLER_17_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_mem_bottom_track_25.sky130_fd_sc_hd__dfxbp_1_0__CLK prog_clk VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__44__A _44_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__39__A chanx_right_in[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__52__A _52_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11_ _11_/HI _11_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XANTENNA_mem_bottom_track_1.sky130_fd_sc_hd__dfxbp_1_1__CLK prog_clk VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_bottom_track_25.mux_l2_in_0__A0 _09_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__47__A chany_bottom_in[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_right_track_4.sky130_fd_sc_hd__buf_4_0__A mux_right_track_4.mux_l2_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__55__A chany_bottom_in[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_10_ _10_/HI _10_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XFILLER_18_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_bottom_track_25.mux_l2_in_0__A1 mux_bottom_track_25.mux_l1_in_0_/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_right_track_0.mux_l2_in_0__A0 _12_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mem_right_track_4.sky130_fd_sc_hd__dfxbp_1_0__D mux_right_track_0.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_right_track_0.mux_l2_in_0__A1 mux_right_track_0.mux_l1_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_bottom_track_1.mux_l1_in_0__A0 bottom_left_grid_pin_1_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_mem_bottom_track_5.sky130_fd_sc_hd__dfxbp_1_1__CLK prog_clk VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmem_right_track_4.sky130_fd_sc_hd__dfxbp_1_1_ mux_right_track_4.mux_l1_in_0_/S mux_right_track_4.mux_l2_in_0_/S
+ mem_right_track_4.sky130_fd_sc_hd__dfxbp_1_1_/Q_N prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_7_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_bottom_track_9.sky130_fd_sc_hd__dfxbp_1_1__D mux_bottom_track_9.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_bottom_track_1.mux_l1_in_0__A1 chanx_right_in[18] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_38_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_mem_bottom_track_25.sky130_fd_sc_hd__dfxbp_1_0__D mux_bottom_track_9.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_right_track_4.mux_l1_in_0__A0 chany_bottom_in[16] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_23_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmem_right_track_4.sky130_fd_sc_hd__dfxbp_1_0_ mux_right_track_0.mux_l2_in_0_/S mux_right_track_4.mux_l1_in_0_/S
+ mem_right_track_4.sky130_fd_sc_hd__dfxbp_1_0_/Q_N prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_11_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_bottom_track_25.sky130_fd_sc_hd__buf_4_0__A mux_bottom_track_25.mux_l2_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_mux_right_track_24.mux_l2_in_0__S mux_right_track_24.mux_l2_in_0_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
.ends

