magic
tech sky130A
magscale 1 2
timestamp 1608157820
<< obsli1 >>
rect 1104 2159 21620 20145
<< obsm1 >>
rect 198 1300 22618 20176
<< metal2 >>
rect 202 0 258 800
rect 570 0 626 800
rect 1030 0 1086 800
rect 1490 0 1546 800
rect 1950 0 2006 800
rect 2318 0 2374 800
rect 2778 0 2834 800
rect 3238 0 3294 800
rect 3698 0 3754 800
rect 4066 0 4122 800
rect 4526 0 4582 800
rect 4986 0 5042 800
rect 5446 0 5502 800
rect 5906 0 5962 800
rect 6274 0 6330 800
rect 6734 0 6790 800
rect 7194 0 7250 800
rect 7654 0 7710 800
rect 8022 0 8078 800
rect 8482 0 8538 800
rect 8942 0 8998 800
rect 9402 0 9458 800
rect 9770 0 9826 800
rect 10230 0 10286 800
rect 10690 0 10746 800
rect 11150 0 11206 800
rect 11610 0 11666 800
rect 11978 0 12034 800
rect 12438 0 12494 800
rect 12898 0 12954 800
rect 13358 0 13414 800
rect 13726 0 13782 800
rect 14186 0 14242 800
rect 14646 0 14702 800
rect 15106 0 15162 800
rect 15474 0 15530 800
rect 15934 0 15990 800
rect 16394 0 16450 800
rect 16854 0 16910 800
rect 17314 0 17370 800
rect 17682 0 17738 800
rect 18142 0 18198 800
rect 18602 0 18658 800
rect 19062 0 19118 800
rect 19430 0 19486 800
rect 19890 0 19946 800
rect 20350 0 20406 800
rect 20810 0 20866 800
rect 21178 0 21234 800
rect 21638 0 21694 800
rect 22098 0 22154 800
rect 22558 0 22614 800
<< obsm2 >>
rect 204 856 22612 22545
rect 314 167 514 856
rect 682 167 974 856
rect 1142 167 1434 856
rect 1602 167 1894 856
rect 2062 167 2262 856
rect 2430 167 2722 856
rect 2890 167 3182 856
rect 3350 167 3642 856
rect 3810 167 4010 856
rect 4178 167 4470 856
rect 4638 167 4930 856
rect 5098 167 5390 856
rect 5558 167 5850 856
rect 6018 167 6218 856
rect 6386 167 6678 856
rect 6846 167 7138 856
rect 7306 167 7598 856
rect 7766 167 7966 856
rect 8134 167 8426 856
rect 8594 167 8886 856
rect 9054 167 9346 856
rect 9514 167 9714 856
rect 9882 167 10174 856
rect 10342 167 10634 856
rect 10802 167 11094 856
rect 11262 167 11554 856
rect 11722 167 11922 856
rect 12090 167 12382 856
rect 12550 167 12842 856
rect 13010 167 13302 856
rect 13470 167 13670 856
rect 13838 167 14130 856
rect 14298 167 14590 856
rect 14758 167 15050 856
rect 15218 167 15418 856
rect 15586 167 15878 856
rect 16046 167 16338 856
rect 16506 167 16798 856
rect 16966 167 17258 856
rect 17426 167 17626 856
rect 17794 167 18086 856
rect 18254 167 18546 856
rect 18714 167 19006 856
rect 19174 167 19374 856
rect 19542 167 19834 856
rect 20002 167 20294 856
rect 20462 167 20754 856
rect 20922 167 21122 856
rect 21290 167 21582 856
rect 21750 167 22042 856
rect 22210 167 22502 856
<< metal3 >>
rect 0 22448 800 22568
rect 0 22040 800 22160
rect 0 21496 800 21616
rect 0 21088 800 21208
rect 0 20544 800 20664
rect 0 20136 800 20256
rect 0 19728 800 19848
rect 0 19184 800 19304
rect 0 18776 800 18896
rect 0 18232 800 18352
rect 0 17824 800 17944
rect 0 17280 800 17400
rect 22000 17144 22800 17264
rect 0 16872 800 16992
rect 0 16464 800 16584
rect 0 15920 800 16040
rect 0 15512 800 15632
rect 0 14968 800 15088
rect 0 14560 800 14680
rect 0 14016 800 14136
rect 0 13608 800 13728
rect 0 13200 800 13320
rect 0 12656 800 12776
rect 0 12248 800 12368
rect 0 11704 800 11824
rect 0 11296 800 11416
rect 0 10752 800 10872
rect 0 10344 800 10464
rect 0 9936 800 10056
rect 0 9392 800 9512
rect 0 8984 800 9104
rect 0 8440 800 8560
rect 0 8032 800 8152
rect 0 7488 800 7608
rect 0 7080 800 7200
rect 0 6672 800 6792
rect 0 6128 800 6248
rect 0 5720 800 5840
rect 22000 5720 22800 5840
rect 0 5176 800 5296
rect 0 4768 800 4888
rect 0 4224 800 4344
rect 0 3816 800 3936
rect 0 3408 800 3528
rect 0 2864 800 2984
rect 0 2456 800 2576
rect 0 1912 800 2032
rect 0 1504 800 1624
rect 0 960 800 1080
rect 0 552 800 672
rect 0 144 800 264
<< obsm3 >>
rect 880 22368 22000 22541
rect 800 22240 22000 22368
rect 880 21960 22000 22240
rect 800 21696 22000 21960
rect 880 21416 22000 21696
rect 800 21288 22000 21416
rect 880 21008 22000 21288
rect 800 20744 22000 21008
rect 880 20464 22000 20744
rect 800 20336 22000 20464
rect 880 20056 22000 20336
rect 800 19928 22000 20056
rect 880 19648 22000 19928
rect 800 19384 22000 19648
rect 880 19104 22000 19384
rect 800 18976 22000 19104
rect 880 18696 22000 18976
rect 800 18432 22000 18696
rect 880 18152 22000 18432
rect 800 18024 22000 18152
rect 880 17744 22000 18024
rect 800 17480 22000 17744
rect 880 17344 22000 17480
rect 880 17200 21920 17344
rect 800 17072 21920 17200
rect 880 17064 21920 17072
rect 880 16792 22000 17064
rect 800 16664 22000 16792
rect 880 16384 22000 16664
rect 800 16120 22000 16384
rect 880 15840 22000 16120
rect 800 15712 22000 15840
rect 880 15432 22000 15712
rect 800 15168 22000 15432
rect 880 14888 22000 15168
rect 800 14760 22000 14888
rect 880 14480 22000 14760
rect 800 14216 22000 14480
rect 880 13936 22000 14216
rect 800 13808 22000 13936
rect 880 13528 22000 13808
rect 800 13400 22000 13528
rect 880 13120 22000 13400
rect 800 12856 22000 13120
rect 880 12576 22000 12856
rect 800 12448 22000 12576
rect 880 12168 22000 12448
rect 800 11904 22000 12168
rect 880 11624 22000 11904
rect 800 11496 22000 11624
rect 880 11216 22000 11496
rect 800 10952 22000 11216
rect 880 10672 22000 10952
rect 800 10544 22000 10672
rect 880 10264 22000 10544
rect 800 10136 22000 10264
rect 880 9856 22000 10136
rect 800 9592 22000 9856
rect 880 9312 22000 9592
rect 800 9184 22000 9312
rect 880 8904 22000 9184
rect 800 8640 22000 8904
rect 880 8360 22000 8640
rect 800 8232 22000 8360
rect 880 7952 22000 8232
rect 800 7688 22000 7952
rect 880 7408 22000 7688
rect 800 7280 22000 7408
rect 880 7000 22000 7280
rect 800 6872 22000 7000
rect 880 6592 22000 6872
rect 800 6328 22000 6592
rect 880 6048 22000 6328
rect 800 5920 22000 6048
rect 880 5640 21920 5920
rect 800 5376 22000 5640
rect 880 5096 22000 5376
rect 800 4968 22000 5096
rect 880 4688 22000 4968
rect 800 4424 22000 4688
rect 880 4144 22000 4424
rect 800 4016 22000 4144
rect 880 3736 22000 4016
rect 800 3608 22000 3736
rect 880 3328 22000 3608
rect 800 3064 22000 3328
rect 880 2784 22000 3064
rect 800 2656 22000 2784
rect 880 2376 22000 2656
rect 800 2112 22000 2376
rect 880 1832 22000 2112
rect 800 1704 22000 1832
rect 880 1424 22000 1704
rect 800 1160 22000 1424
rect 880 880 22000 1160
rect 800 752 22000 880
rect 880 472 22000 752
rect 800 344 22000 472
rect 880 171 22000 344
<< metal4 >>
rect 4376 2128 4696 20176
rect 7808 2128 8128 20176
<< obsm4 >>
rect 11240 2128 18424 20176
<< labels >>
rlabel metal2 s 21638 0 21694 800 6 SC_IN_BOT
port 1 nsew default input
rlabel metal2 s 22098 0 22154 800 6 SC_OUT_BOT
port 2 nsew default output
rlabel metal2 s 202 0 258 800 6 bottom_left_grid_pin_42_
port 3 nsew default input
rlabel metal2 s 570 0 626 800 6 bottom_left_grid_pin_43_
port 4 nsew default input
rlabel metal2 s 1030 0 1086 800 6 bottom_left_grid_pin_44_
port 5 nsew default input
rlabel metal2 s 1490 0 1546 800 6 bottom_left_grid_pin_45_
port 6 nsew default input
rlabel metal2 s 1950 0 2006 800 6 bottom_left_grid_pin_46_
port 7 nsew default input
rlabel metal2 s 2318 0 2374 800 6 bottom_left_grid_pin_47_
port 8 nsew default input
rlabel metal2 s 2778 0 2834 800 6 bottom_left_grid_pin_48_
port 9 nsew default input
rlabel metal2 s 3238 0 3294 800 6 bottom_left_grid_pin_49_
port 10 nsew default input
rlabel metal2 s 21178 0 21234 800 6 bottom_right_grid_pin_1_
port 11 nsew default input
rlabel metal3 s 22000 5720 22800 5840 6 ccff_head
port 12 nsew default input
rlabel metal3 s 22000 17144 22800 17264 6 ccff_tail
port 13 nsew default output
rlabel metal3 s 0 3816 800 3936 6 chanx_left_in[0]
port 14 nsew default input
rlabel metal3 s 0 8440 800 8560 6 chanx_left_in[10]
port 15 nsew default input
rlabel metal3 s 0 8984 800 9104 6 chanx_left_in[11]
port 16 nsew default input
rlabel metal3 s 0 9392 800 9512 6 chanx_left_in[12]
port 17 nsew default input
rlabel metal3 s 0 9936 800 10056 6 chanx_left_in[13]
port 18 nsew default input
rlabel metal3 s 0 10344 800 10464 6 chanx_left_in[14]
port 19 nsew default input
rlabel metal3 s 0 10752 800 10872 6 chanx_left_in[15]
port 20 nsew default input
rlabel metal3 s 0 11296 800 11416 6 chanx_left_in[16]
port 21 nsew default input
rlabel metal3 s 0 11704 800 11824 6 chanx_left_in[17]
port 22 nsew default input
rlabel metal3 s 0 12248 800 12368 6 chanx_left_in[18]
port 23 nsew default input
rlabel metal3 s 0 12656 800 12776 6 chanx_left_in[19]
port 24 nsew default input
rlabel metal3 s 0 4224 800 4344 6 chanx_left_in[1]
port 25 nsew default input
rlabel metal3 s 0 4768 800 4888 6 chanx_left_in[2]
port 26 nsew default input
rlabel metal3 s 0 5176 800 5296 6 chanx_left_in[3]
port 27 nsew default input
rlabel metal3 s 0 5720 800 5840 6 chanx_left_in[4]
port 28 nsew default input
rlabel metal3 s 0 6128 800 6248 6 chanx_left_in[5]
port 29 nsew default input
rlabel metal3 s 0 6672 800 6792 6 chanx_left_in[6]
port 30 nsew default input
rlabel metal3 s 0 7080 800 7200 6 chanx_left_in[7]
port 31 nsew default input
rlabel metal3 s 0 7488 800 7608 6 chanx_left_in[8]
port 32 nsew default input
rlabel metal3 s 0 8032 800 8152 6 chanx_left_in[9]
port 33 nsew default input
rlabel metal3 s 0 13200 800 13320 6 chanx_left_out[0]
port 34 nsew default output
rlabel metal3 s 0 17824 800 17944 6 chanx_left_out[10]
port 35 nsew default output
rlabel metal3 s 0 18232 800 18352 6 chanx_left_out[11]
port 36 nsew default output
rlabel metal3 s 0 18776 800 18896 6 chanx_left_out[12]
port 37 nsew default output
rlabel metal3 s 0 19184 800 19304 6 chanx_left_out[13]
port 38 nsew default output
rlabel metal3 s 0 19728 800 19848 6 chanx_left_out[14]
port 39 nsew default output
rlabel metal3 s 0 20136 800 20256 6 chanx_left_out[15]
port 40 nsew default output
rlabel metal3 s 0 20544 800 20664 6 chanx_left_out[16]
port 41 nsew default output
rlabel metal3 s 0 21088 800 21208 6 chanx_left_out[17]
port 42 nsew default output
rlabel metal3 s 0 21496 800 21616 6 chanx_left_out[18]
port 43 nsew default output
rlabel metal3 s 0 22040 800 22160 6 chanx_left_out[19]
port 44 nsew default output
rlabel metal3 s 0 13608 800 13728 6 chanx_left_out[1]
port 45 nsew default output
rlabel metal3 s 0 14016 800 14136 6 chanx_left_out[2]
port 46 nsew default output
rlabel metal3 s 0 14560 800 14680 6 chanx_left_out[3]
port 47 nsew default output
rlabel metal3 s 0 14968 800 15088 6 chanx_left_out[4]
port 48 nsew default output
rlabel metal3 s 0 15512 800 15632 6 chanx_left_out[5]
port 49 nsew default output
rlabel metal3 s 0 15920 800 16040 6 chanx_left_out[6]
port 50 nsew default output
rlabel metal3 s 0 16464 800 16584 6 chanx_left_out[7]
port 51 nsew default output
rlabel metal3 s 0 16872 800 16992 6 chanx_left_out[8]
port 52 nsew default output
rlabel metal3 s 0 17280 800 17400 6 chanx_left_out[9]
port 53 nsew default output
rlabel metal2 s 3698 0 3754 800 6 chany_bottom_in[0]
port 54 nsew default input
rlabel metal2 s 8022 0 8078 800 6 chany_bottom_in[10]
port 55 nsew default input
rlabel metal2 s 8482 0 8538 800 6 chany_bottom_in[11]
port 56 nsew default input
rlabel metal2 s 8942 0 8998 800 6 chany_bottom_in[12]
port 57 nsew default input
rlabel metal2 s 9402 0 9458 800 6 chany_bottom_in[13]
port 58 nsew default input
rlabel metal2 s 9770 0 9826 800 6 chany_bottom_in[14]
port 59 nsew default input
rlabel metal2 s 10230 0 10286 800 6 chany_bottom_in[15]
port 60 nsew default input
rlabel metal2 s 10690 0 10746 800 6 chany_bottom_in[16]
port 61 nsew default input
rlabel metal2 s 11150 0 11206 800 6 chany_bottom_in[17]
port 62 nsew default input
rlabel metal2 s 11610 0 11666 800 6 chany_bottom_in[18]
port 63 nsew default input
rlabel metal2 s 11978 0 12034 800 6 chany_bottom_in[19]
port 64 nsew default input
rlabel metal2 s 4066 0 4122 800 6 chany_bottom_in[1]
port 65 nsew default input
rlabel metal2 s 4526 0 4582 800 6 chany_bottom_in[2]
port 66 nsew default input
rlabel metal2 s 4986 0 5042 800 6 chany_bottom_in[3]
port 67 nsew default input
rlabel metal2 s 5446 0 5502 800 6 chany_bottom_in[4]
port 68 nsew default input
rlabel metal2 s 5906 0 5962 800 6 chany_bottom_in[5]
port 69 nsew default input
rlabel metal2 s 6274 0 6330 800 6 chany_bottom_in[6]
port 70 nsew default input
rlabel metal2 s 6734 0 6790 800 6 chany_bottom_in[7]
port 71 nsew default input
rlabel metal2 s 7194 0 7250 800 6 chany_bottom_in[8]
port 72 nsew default input
rlabel metal2 s 7654 0 7710 800 6 chany_bottom_in[9]
port 73 nsew default input
rlabel metal2 s 12438 0 12494 800 6 chany_bottom_out[0]
port 74 nsew default output
rlabel metal2 s 16854 0 16910 800 6 chany_bottom_out[10]
port 75 nsew default output
rlabel metal2 s 17314 0 17370 800 6 chany_bottom_out[11]
port 76 nsew default output
rlabel metal2 s 17682 0 17738 800 6 chany_bottom_out[12]
port 77 nsew default output
rlabel metal2 s 18142 0 18198 800 6 chany_bottom_out[13]
port 78 nsew default output
rlabel metal2 s 18602 0 18658 800 6 chany_bottom_out[14]
port 79 nsew default output
rlabel metal2 s 19062 0 19118 800 6 chany_bottom_out[15]
port 80 nsew default output
rlabel metal2 s 19430 0 19486 800 6 chany_bottom_out[16]
port 81 nsew default output
rlabel metal2 s 19890 0 19946 800 6 chany_bottom_out[17]
port 82 nsew default output
rlabel metal2 s 20350 0 20406 800 6 chany_bottom_out[18]
port 83 nsew default output
rlabel metal2 s 20810 0 20866 800 6 chany_bottom_out[19]
port 84 nsew default output
rlabel metal2 s 12898 0 12954 800 6 chany_bottom_out[1]
port 85 nsew default output
rlabel metal2 s 13358 0 13414 800 6 chany_bottom_out[2]
port 86 nsew default output
rlabel metal2 s 13726 0 13782 800 6 chany_bottom_out[3]
port 87 nsew default output
rlabel metal2 s 14186 0 14242 800 6 chany_bottom_out[4]
port 88 nsew default output
rlabel metal2 s 14646 0 14702 800 6 chany_bottom_out[5]
port 89 nsew default output
rlabel metal2 s 15106 0 15162 800 6 chany_bottom_out[6]
port 90 nsew default output
rlabel metal2 s 15474 0 15530 800 6 chany_bottom_out[7]
port 91 nsew default output
rlabel metal2 s 15934 0 15990 800 6 chany_bottom_out[8]
port 92 nsew default output
rlabel metal2 s 16394 0 16450 800 6 chany_bottom_out[9]
port 93 nsew default output
rlabel metal3 s 0 144 800 264 6 left_bottom_grid_pin_34_
port 94 nsew default input
rlabel metal3 s 0 552 800 672 6 left_bottom_grid_pin_35_
port 95 nsew default input
rlabel metal3 s 0 960 800 1080 6 left_bottom_grid_pin_36_
port 96 nsew default input
rlabel metal3 s 0 1504 800 1624 6 left_bottom_grid_pin_37_
port 97 nsew default input
rlabel metal3 s 0 1912 800 2032 6 left_bottom_grid_pin_38_
port 98 nsew default input
rlabel metal3 s 0 2456 800 2576 6 left_bottom_grid_pin_39_
port 99 nsew default input
rlabel metal3 s 0 2864 800 2984 6 left_bottom_grid_pin_40_
port 100 nsew default input
rlabel metal3 s 0 3408 800 3528 6 left_bottom_grid_pin_41_
port 101 nsew default input
rlabel metal3 s 0 22448 800 22568 6 left_top_grid_pin_1_
port 102 nsew default input
rlabel metal2 s 22558 0 22614 800 6 prog_clk_0_S_in
port 103 nsew default input
rlabel metal4 s 4376 2128 4696 20176 6 VPWR
port 104 nsew power input
rlabel metal4 s 7808 2128 8128 20176 6 VGND
port 105 nsew ground input
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 22800 22568
string LEFview TRUE
<< end >>
