* NGSPICE file created from sb_1__0_.ext - technology: EFS8A

* Black-box entry subcircuit for scs8hd_fill_2 abstract view
.subckt scs8hd_fill_2 vpwr vgnd
.ends

* Black-box entry subcircuit for scs8hd_decap_4 abstract view
.subckt scs8hd_decap_4 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_diode_2 abstract view
.subckt scs8hd_diode_2 DIODE vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_decap_12 abstract view
.subckt scs8hd_decap_12 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_inv_1 abstract view
.subckt scs8hd_inv_1 A Y vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_ebufn_2 abstract view
.subckt scs8hd_ebufn_2 A TEB Z vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_buf_2 abstract view
.subckt scs8hd_buf_2 A X vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_nor2_4 abstract view
.subckt scs8hd_nor2_4 A B Y vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_decap_3 abstract view
.subckt scs8hd_decap_3 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_decap_6 abstract view
.subckt scs8hd_decap_6 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_lpflow_inputisolatch_1 abstract view
.subckt scs8hd_lpflow_inputisolatch_1 D Q SLEEPB vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_fill_1 abstract view
.subckt scs8hd_fill_1 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_tapvpwrvgnd_1 abstract view
.subckt scs8hd_tapvpwrvgnd_1 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_decap_8 abstract view
.subckt scs8hd_decap_8 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_buf_1 abstract view
.subckt scs8hd_buf_1 A X vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_conb_1 abstract view
.subckt scs8hd_conb_1 HI LO vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_or3_4 abstract view
.subckt scs8hd_or3_4 A B C X vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_or2_4 abstract view
.subckt scs8hd_or2_4 A B X vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_inv_8 abstract view
.subckt scs8hd_inv_8 A Y vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_nor4_4 abstract view
.subckt scs8hd_nor4_4 A B C D Y vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_nor3_4 abstract view
.subckt scs8hd_nor3_4 A B C Y vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_or4_4 abstract view
.subckt scs8hd_or4_4 A B C D X vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_nand3_4 abstract view
.subckt scs8hd_nand3_4 A B C Y vgnd vpwr
.ends

.subckt sb_1__0_ address[0] address[1] address[2] address[3] address[4] address[5]
+ address[6] chanx_left_in[0] chanx_left_in[1] chanx_left_in[2] chanx_left_in[3] chanx_left_in[4]
+ chanx_left_in[5] chanx_left_in[6] chanx_left_in[7] chanx_left_in[8] chanx_left_out[0]
+ chanx_left_out[1] chanx_left_out[2] chanx_left_out[3] chanx_left_out[4] chanx_left_out[5]
+ chanx_left_out[6] chanx_left_out[7] chanx_left_out[8] chanx_right_in[0] chanx_right_in[1]
+ chanx_right_in[2] chanx_right_in[3] chanx_right_in[4] chanx_right_in[5] chanx_right_in[6]
+ chanx_right_in[7] chanx_right_in[8] chanx_right_out[0] chanx_right_out[1] chanx_right_out[2]
+ chanx_right_out[3] chanx_right_out[4] chanx_right_out[5] chanx_right_out[6] chanx_right_out[7]
+ chanx_right_out[8] chany_top_in[0] chany_top_in[1] chany_top_in[2] chany_top_in[3]
+ chany_top_in[4] chany_top_in[5] chany_top_in[6] chany_top_in[7] chany_top_in[8]
+ chany_top_out[0] chany_top_out[1] chany_top_out[2] chany_top_out[3] chany_top_out[4]
+ chany_top_out[5] chany_top_out[6] chany_top_out[7] chany_top_out[8] data_in enable
+ left_bottom_grid_pin_11_ left_bottom_grid_pin_13_ left_bottom_grid_pin_15_ left_bottom_grid_pin_1_
+ left_bottom_grid_pin_3_ left_bottom_grid_pin_5_ left_bottom_grid_pin_7_ left_bottom_grid_pin_9_
+ left_top_grid_pin_10_ right_bottom_grid_pin_11_ right_bottom_grid_pin_13_ right_bottom_grid_pin_15_
+ right_bottom_grid_pin_1_ right_bottom_grid_pin_3_ right_bottom_grid_pin_5_ right_bottom_grid_pin_7_
+ right_bottom_grid_pin_9_ right_top_grid_pin_10_ top_left_grid_pin_13_ top_right_grid_pin_11_
+ vpwr vgnd
XFILLER_39_222 vpwr vgnd scs8hd_fill_2
XFILLER_36_19 vpwr vgnd scs8hd_fill_2
XFILLER_22_111 vgnd vpwr scs8hd_decap_4
XANTENNA_mem_top_track_2.LATCH_1_.latch_SLEEPB _159_/Y vgnd vpwr scs8hd_diode_2
XFILLER_7_7 vgnd vpwr scs8hd_decap_12
XFILLER_9_159 vgnd vpwr scs8hd_decap_12
XANTENNA__113__B _110_/X vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_track_0.LATCH_3_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_36_236 vgnd vpwr scs8hd_decap_12
Xmux_top_track_8.INVTX1_0_.scs8hd_inv_1 chanx_right_in[6] mux_top_track_8.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_27_258 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_9.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_left_track_9.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_6_129 vgnd vpwr scs8hd_decap_12
XFILLER_12_32 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_top_track_16.LATCH_0_.latch_SLEEPB _172_/Y vgnd vpwr scs8hd_diode_2
XFILLER_37_73 vpwr vgnd scs8hd_fill_2
XFILLER_37_62 vpwr vgnd scs8hd_fill_2
XANTENNA__108__B _106_/B vgnd vpwr scs8hd_diode_2
XANTENNA__124__A _124_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_16.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB mem_right_track_16.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_5_184 vgnd vpwr scs8hd_decap_12
XFILLER_24_206 vpwr vgnd scs8hd_fill_2
XFILLER_24_228 vgnd vpwr scs8hd_decap_4
Xmux_left_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_left_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ mem_left_track_1.LATCH_3_.latch/Q mux_left_track_1.tap_buf4_0_.scs8hd_inv_1/A vgnd
+ vpwr scs8hd_ebufn_2
X_200_ chanx_left_in[0] chanx_right_out[1] vgnd vpwr scs8hd_buf_2
XANTENNA_mem_right_track_16.LATCH_4_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA__209__A _209_/A vgnd vpwr scs8hd_diode_2
XFILLER_15_217 vgnd vpwr scs8hd_decap_12
XFILLER_23_20 vgnd vpwr scs8hd_decap_4
XFILLER_23_261 vgnd vpwr scs8hd_decap_12
X_131_ _113_/A _132_/B _131_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_2_154 vgnd vpwr scs8hd_decap_12
XANTENNA__119__A address[4] vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_track_16.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_18_53 vpwr vgnd scs8hd_fill_2
XFILLER_34_96 vpwr vgnd scs8hd_fill_2
XFILLER_34_52 vpwr vgnd scs8hd_fill_2
XFILLER_11_220 vgnd vpwr scs8hd_decap_12
XFILLER_11_253 vpwr vgnd scs8hd_fill_2
X_114_ _124_/A _110_/X _114_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_7_257 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_top_track_0.LATCH_2_.latch_SLEEPB _155_/Y vgnd vpwr scs8hd_diode_2
Xmux_right_track_16.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_right_track_16.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2/Z
+ mem_right_track_16.LATCH_4_.latch/Q mux_right_track_16.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA__121__B _125_/B vgnd vpwr scs8hd_diode_2
Xmux_left_track_9.INVTX1_3_.scs8hd_inv_1 chanx_right_in[1] mux_left_track_9.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_22_7 vgnd vpwr scs8hd_decap_3
Xmux_top_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_top_track_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ mem_top_track_0.LATCH_4_.latch/Q mux_top_track_0.tap_buf4_0_.scs8hd_inv_1/A vgnd
+ vpwr scs8hd_ebufn_2
Xmux_right_track_8.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2 mux_right_track_8.INVTX1_5_.scs8hd_inv_1/Y
+ mem_right_track_8.LATCH_2_.latch/Q mux_right_track_8.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_right_track_16.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_right_track_16.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_4_227 vgnd vpwr scs8hd_decap_12
XFILLER_20_43 vpwr vgnd scs8hd_fill_2
XANTENNA__116__B _110_/X vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_16.INVTX1_7_.scs8hd_inv_1_A chanx_left_in[6] vgnd vpwr scs8hd_diode_2
XFILLER_6_56 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_top_track_14.LATCH_1_.latch_SLEEPB _163_/Y vgnd vpwr scs8hd_diode_2
XANTENNA__132__A _124_/A vgnd vpwr scs8hd_diode_2
XFILLER_26_109 vgnd vpwr scs8hd_decap_6
Xmem_right_track_8.LATCH_1_.latch data_in mem_right_track_8.LATCH_1_.latch/Q _106_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_34_142 vgnd vpwr scs8hd_decap_4
XFILLER_1_208 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A _179_/HI vgnd vpwr
+ scs8hd_diode_2
XFILLER_40_101 vgnd vpwr scs8hd_fill_1
XFILLER_25_142 vgnd vpwr scs8hd_decap_4
XFILLER_25_175 vpwr vgnd scs8hd_fill_2
XFILLER_31_53 vpwr vgnd scs8hd_fill_2
XFILLER_15_87 vpwr vgnd scs8hd_fill_2
XFILLER_0_263 vgnd vpwr scs8hd_decap_12
XFILLER_31_156 vgnd vpwr scs8hd_fill_1
XFILLER_31_112 vpwr vgnd scs8hd_fill_2
XPHY_170 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mem_left_track_9.LATCH_4_.latch_SLEEPB _130_/Y vgnd vpwr scs8hd_diode_2
XANTENNA__127__A address[4] vgnd vpwr scs8hd_diode_2
XPHY_181 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_192 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_39_245 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_left_track_1.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A mux_left_track_1.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_26_97 vgnd vpwr scs8hd_fill_1
XFILLER_26_86 vgnd vpwr scs8hd_decap_6
XFILLER_13_123 vpwr vgnd scs8hd_fill_2
XFILLER_13_145 vgnd vpwr scs8hd_decap_8
XFILLER_13_156 vgnd vpwr scs8hd_decap_4
XFILLER_42_63 vgnd vpwr scs8hd_decap_12
XFILLER_36_248 vgnd vpwr scs8hd_decap_12
Xmux_left_track_9.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_left_track_9.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2/Z
+ mem_left_track_9.LATCH_5_.latch/Q mux_left_track_9.tap_buf4_0_.scs8hd_inv_1/A vgnd
+ vpwr scs8hd_ebufn_2
Xmux_top_track_0.INVTX1_3_.scs8hd_inv_1 chanx_left_in[0] mux_top_track_0.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_27_226 vgnd vpwr scs8hd_decap_12
XFILLER_42_218 vgnd vpwr scs8hd_decap_12
Xmux_left_track_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 mux_left_track_1.INVTX1_4_.scs8hd_inv_1/Y
+ mem_left_track_1.LATCH_1_.latch/Q mux_left_track_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_right_track_0.INVTX1_4_.scs8hd_inv_1_A right_bottom_grid_pin_5_ vgnd
+ vpwr scs8hd_diode_2
XFILLER_12_66 vgnd vpwr scs8hd_decap_4
XFILLER_37_41 vgnd vpwr scs8hd_decap_3
Xmux_left_track_17.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2 mux_left_track_17.INVTX1_7_.scs8hd_inv_1/Y
+ mem_left_track_17.LATCH_1_.latch/Q mux_left_track_17.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_left_track_17.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_left_track_17.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__124__B _125_/B vgnd vpwr scs8hd_diode_2
XFILLER_5_196 vgnd vpwr scs8hd_decap_12
XANTENNA__140__A _124_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_0.INVTX1_0_.scs8hd_inv_1_A top_left_grid_pin_13_ vgnd vpwr
+ scs8hd_diode_2
Xmux_right_track_8.INVTX1_4_.scs8hd_inv_1 right_bottom_grid_pin_7_ mux_right_track_8.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_right_track_8.INVTX1_6_.scs8hd_inv_1_A chanx_left_in[1] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_9.INVTX1_0_.scs8hd_inv_1_A chany_top_in[2] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_right_track_0.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_15_229 vgnd vpwr scs8hd_decap_12
X_130_ _112_/A _132_/B _130_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA_mux_right_track_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_right_track_0.LATCH_5_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_23_273 vgnd vpwr scs8hd_decap_4
XANTENNA_mem_right_track_0.LATCH_4_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_23_98 vpwr vgnd scs8hd_fill_2
Xmux_right_track_16.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2 mux_right_track_16.INVTX1_5_.scs8hd_inv_1/Y
+ mem_right_track_16.LATCH_2_.latch/Q mux_right_track_16.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_right_track_16.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB mem_right_track_16.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_2_166 vgnd vpwr scs8hd_decap_12
XANTENNA__119__B address[3] vgnd vpwr scs8hd_diode_2
XANTENNA__135__A _095_/A vgnd vpwr scs8hd_diode_2
XFILLER_9_45 vgnd vpwr scs8hd_decap_12
XFILLER_9_34 vgnd vpwr scs8hd_decap_8
XFILLER_14_251 vgnd vpwr scs8hd_decap_12
XFILLER_20_276 vgnd vpwr scs8hd_fill_1
XFILLER_34_64 vgnd vpwr scs8hd_decap_4
X_113_ _113_/A _110_/X _113_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_11_232 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_left_track_1.LATCH_0_.latch_SLEEPB _126_/Y vgnd vpwr scs8hd_diode_2
XFILLER_7_269 vgnd vpwr scs8hd_decap_8
XFILLER_38_129 vgnd vpwr scs8hd_decap_6
Xmux_left_track_1.INVTX1_6_.scs8hd_inv_1 left_bottom_grid_pin_5_ mux_left_track_1.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_left_track_9.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A mux_left_track_9.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_37_184 vpwr vgnd scs8hd_fill_2
XFILLER_37_173 vpwr vgnd scs8hd_fill_2
XFILLER_4_239 vgnd vpwr scs8hd_decap_12
XFILLER_20_88 vgnd vpwr scs8hd_decap_4
XFILLER_20_99 vpwr vgnd scs8hd_fill_2
XFILLER_29_53 vpwr vgnd scs8hd_fill_2
XFILLER_28_184 vgnd vpwr scs8hd_fill_1
XFILLER_6_68 vgnd vpwr scs8hd_decap_12
XANTENNA__132__B _132_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_track_16.LATCH_0_.latch_SLEEPB _116_/Y vgnd vpwr scs8hd_diode_2
XFILLER_19_184 vgnd vpwr scs8hd_decap_3
XFILLER_34_165 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_1.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_TEB mem_left_track_1.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_top_track_0.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_top_track_16.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_25_132 vgnd vpwr scs8hd_decap_4
XFILLER_40_179 vgnd vpwr scs8hd_decap_8
XFILLER_40_168 vgnd vpwr scs8hd_decap_8
XFILLER_40_157 vgnd vpwr scs8hd_decap_3
XFILLER_31_21 vpwr vgnd scs8hd_fill_2
XFILLER_15_77 vpwr vgnd scs8hd_fill_2
XFILLER_15_99 vgnd vpwr scs8hd_decap_4
XFILLER_31_87 vpwr vgnd scs8hd_fill_2
XFILLER_0_242 vgnd vpwr scs8hd_decap_6
XFILLER_0_275 vpwr vgnd scs8hd_fill_2
Xmux_right_track_16.INVTX1_0_.scs8hd_inv_1 chany_top_in[1] mux_right_track_16.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
Xmux_left_track_17.INVTX1_1_.scs8hd_inv_1 chany_top_in[4] mux_left_track_17.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_31_179 vpwr vgnd scs8hd_fill_2
XPHY_160 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_16_154 vpwr vgnd scs8hd_fill_2
XFILLER_16_187 vpwr vgnd scs8hd_fill_2
XPHY_171 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_182 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_193 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__127__B _109_/B vgnd vpwr scs8hd_diode_2
XANTENNA__143__A _143_/A vgnd vpwr scs8hd_diode_2
XFILLER_30_190 vpwr vgnd scs8hd_fill_2
Xmux_top_track_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_top_track_2.INVTX1_1_.scs8hd_inv_1/Y
+ _144_/Y mux_top_track_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XFILLER_26_10 vpwr vgnd scs8hd_fill_2
XFILLER_26_32 vgnd vpwr scs8hd_decap_4
XANTENNA_mem_left_track_1.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_13_102 vgnd vpwr scs8hd_decap_12
XFILLER_13_168 vpwr vgnd scs8hd_fill_2
XFILLER_26_65 vgnd vpwr scs8hd_decap_4
XFILLER_42_75 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_16.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A mux_right_track_16.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_36_205 vgnd vpwr scs8hd_decap_3
XANTENNA__138__A _112_/A vgnd vpwr scs8hd_diode_2
XFILLER_12_190 vgnd vpwr scs8hd_decap_12
XFILLER_27_238 vgnd vpwr scs8hd_decap_6
XFILLER_10_105 vgnd vpwr scs8hd_decap_12
XFILLER_12_23 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_left_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_left_track_9.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_37_86 vgnd vpwr scs8hd_decap_12
XFILLER_37_53 vgnd vpwr scs8hd_decap_8
XFILLER_37_31 vgnd vpwr scs8hd_decap_8
XFILLER_37_20 vgnd vpwr scs8hd_decap_4
XFILLER_26_271 vgnd vpwr scs8hd_decap_4
XFILLER_18_205 vgnd vpwr scs8hd_fill_1
XANTENNA__140__B _136_/X vgnd vpwr scs8hd_diode_2
XFILLER_32_274 vgnd vpwr scs8hd_fill_1
Xmux_right_track_0.INVTX1_7_.scs8hd_inv_1 chanx_left_in[4] mux_right_track_0.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_15_208 vgnd vpwr scs8hd_decap_6
XFILLER_23_77 vpwr vgnd scs8hd_fill_2
XFILLER_3_3 vgnd vpwr scs8hd_decap_12
XFILLER_2_178 vgnd vpwr scs8hd_decap_12
XFILLER_0_15 vgnd vpwr scs8hd_decap_12
XFILLER_14_263 vgnd vpwr scs8hd_decap_12
XANTENNA__119__C address[5] vgnd vpwr scs8hd_diode_2
X_189_ chanx_right_in[2] chanx_left_out[3] vgnd vpwr scs8hd_buf_2
XFILLER_9_57 vgnd vpwr scs8hd_decap_4
XANTENNA__135__B address[3] vgnd vpwr scs8hd_diode_2
XFILLER_36_3 vgnd vpwr scs8hd_decap_3
XANTENNA__151__A _150_/X vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _144_/Y vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_right_track_16.INVTX1_2_.scs8hd_inv_1_A chany_top_in[7] vgnd vpwr scs8hd_diode_2
XFILLER_34_32 vgnd vpwr scs8hd_decap_8
XFILLER_34_21 vpwr vgnd scs8hd_fill_2
XFILLER_18_88 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_top_track_16.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A _181_/HI vgnd vpwr
+ scs8hd_diode_2
X_112_ _112_/A _110_/X _112_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA__146__A _146_/A vgnd vpwr scs8hd_diode_2
XFILLER_37_152 vpwr vgnd scs8hd_fill_2
XFILLER_20_23 vpwr vgnd scs8hd_fill_2
XFILLER_29_65 vpwr vgnd scs8hd_fill_2
XFILLER_29_32 vpwr vgnd scs8hd_fill_2
XFILLER_28_196 vpwr vgnd scs8hd_fill_2
XFILLER_34_100 vgnd vpwr scs8hd_decap_8
XFILLER_19_130 vpwr vgnd scs8hd_fill_2
XFILLER_19_152 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A mux_right_track_0.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_34_188 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_left_track_17.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_left_track_17.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_40_136 vgnd vpwr scs8hd_decap_4
XFILLER_25_100 vgnd vpwr scs8hd_decap_3
XFILLER_25_199 vpwr vgnd scs8hd_fill_2
XFILLER_0_221 vpwr vgnd scs8hd_fill_2
XFILLER_16_122 vgnd vpwr scs8hd_decap_4
Xmux_right_track_0.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2 _176_/HI mem_right_track_0.LATCH_2_.latch/Q
+ mux_right_track_0.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XFILLER_31_136 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_right_track_8.LATCH_5_.latch_SLEEPB _098_/Y vgnd vpwr scs8hd_diode_2
XPHY_150 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_161 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_172 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mem_left_track_9.LATCH_4_.latch_D data_in vgnd vpwr scs8hd_diode_2
XPHY_183 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_194 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__127__C address[5] vgnd vpwr scs8hd_diode_2
XFILLER_39_258 vpwr vgnd scs8hd_fill_2
XFILLER_39_214 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_top_track_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB mem_top_track_0.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_26_55 vpwr vgnd scs8hd_fill_2
XFILLER_42_87 vgnd vpwr scs8hd_decap_6
XFILLER_42_32 vgnd vpwr scs8hd_decap_12
XFILLER_13_114 vgnd vpwr scs8hd_decap_6
XFILLER_21_180 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_right_track_8.INVTX1_1_.scs8hd_inv_1_A chany_top_in[3] vgnd vpwr scs8hd_diode_2
XFILLER_3_59 vpwr vgnd scs8hd_fill_2
XFILLER_3_15 vgnd vpwr scs8hd_decap_12
XANTENNA__138__B _136_/X vgnd vpwr scs8hd_diode_2
XANTENNA__154__A _113_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_17.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_left_track_17.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_10_117 vgnd vpwr scs8hd_decap_12
XFILLER_12_13 vgnd vpwr scs8hd_fill_1
XFILLER_41_220 vgnd vpwr scs8hd_decap_12
XFILLER_37_98 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_top_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A _183_/HI vgnd vpwr
+ scs8hd_diode_2
XFILLER_18_228 vgnd vpwr scs8hd_decap_12
XFILLER_5_110 vgnd vpwr scs8hd_decap_12
XFILLER_38_7 vpwr vgnd scs8hd_fill_2
Xmem_top_track_0.LATCH_0_.latch data_in mem_top_track_0.LATCH_0_.latch/Q _157_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_left_track_17.INVTX1_5_.scs8hd_inv_1_A left_bottom_grid_pin_3_ vgnd vpwr
+ scs8hd_diode_2
XANTENNA__149__A _118_/A vgnd vpwr scs8hd_diode_2
XFILLER_4_80 vgnd vpwr scs8hd_decap_12
XFILLER_23_231 vpwr vgnd scs8hd_fill_2
XFILLER_23_12 vpwr vgnd scs8hd_fill_2
XFILLER_23_56 vpwr vgnd scs8hd_fill_2
XFILLER_23_253 vpwr vgnd scs8hd_fill_2
XFILLER_0_27 vgnd vpwr scs8hd_decap_4
Xmem_left_track_17.LATCH_3_.latch data_in mem_left_track_17.LATCH_3_.latch/Q _139_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA__119__D _118_/X vgnd vpwr scs8hd_diode_2
X_188_ _188_/A chanx_left_out[4] vgnd vpwr scs8hd_buf_2
XANTENNA__135__C address[5] vgnd vpwr scs8hd_diode_2
XFILLER_29_3 vpwr vgnd scs8hd_fill_2
XFILLER_18_12 vgnd vpwr scs8hd_decap_4
XFILLER_18_23 vpwr vgnd scs8hd_fill_2
XFILLER_18_67 vgnd vpwr scs8hd_decap_6
XFILLER_34_88 vgnd vpwr scs8hd_decap_4
X_111_ _111_/A _110_/X _111_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_11_245 vgnd vpwr scs8hd_decap_8
XANTENNA_mem_right_track_0.LATCH_1_.latch_SLEEPB _090_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_2.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB _144_/A vgnd vpwr
+ scs8hd_diode_2
XANTENNA__162__A _096_/B vgnd vpwr scs8hd_diode_2
XFILLER_6_271 vgnd vpwr scs8hd_decap_4
XFILLER_37_142 vgnd vpwr scs8hd_fill_1
XFILLER_37_197 vgnd vpwr scs8hd_decap_8
XANTENNA__072__A address[6] vgnd vpwr scs8hd_diode_2
XFILLER_29_22 vgnd vpwr scs8hd_decap_4
XFILLER_20_68 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_right_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_right_track_8.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_29_88 vpwr vgnd scs8hd_fill_2
XFILLER_6_15 vgnd vpwr scs8hd_decap_12
XFILLER_10_90 vpwr vgnd scs8hd_fill_2
XFILLER_13_6 vpwr vgnd scs8hd_fill_2
XFILLER_19_175 vpwr vgnd scs8hd_fill_2
XANTENNA__157__A _108_/A vgnd vpwr scs8hd_diode_2
Xmux_top_track_2.INVTX1_0_.scs8hd_inv_1 top_right_grid_pin_11_ mux_top_track_2.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_right_track_16.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_16.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_40_104 vgnd vpwr scs8hd_decap_8
XANTENNA__067__A address[1] vgnd vpwr scs8hd_diode_2
XFILLER_15_35 vpwr vgnd scs8hd_fill_2
XFILLER_15_57 vpwr vgnd scs8hd_fill_2
XFILLER_0_233 vpwr vgnd scs8hd_fill_2
XFILLER_31_104 vpwr vgnd scs8hd_fill_2
XPHY_140 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_151 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_162 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_173 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_184 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__127__D _118_/X vgnd vpwr scs8hd_diode_2
XPHY_195 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_39_226 vgnd vpwr scs8hd_decap_12
XFILLER_22_126 vpwr vgnd scs8hd_fill_2
Xmem_left_track_1.LATCH_1_.latch data_in mem_left_track_1.LATCH_1_.latch/Q _125_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_left_track_17.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_left_track_17.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_26_23 vpwr vgnd scs8hd_fill_2
XFILLER_42_44 vgnd vpwr scs8hd_decap_12
XFILLER_3_27 vgnd vpwr scs8hd_decap_12
XFILLER_8_141 vgnd vpwr scs8hd_decap_12
XANTENNA__154__B _157_/B vgnd vpwr scs8hd_diode_2
XANTENNA__170__A _103_/A vgnd vpwr scs8hd_diode_2
XFILLER_35_262 vgnd vpwr scs8hd_decap_12
XFILLER_27_218 vpwr vgnd scs8hd_fill_2
XFILLER_27_207 vpwr vgnd scs8hd_fill_2
Xmem_right_track_16.LATCH_2_.latch data_in mem_right_track_16.LATCH_2_.latch/Q _114_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_10_129 vgnd vpwr scs8hd_decap_12
XFILLER_12_36 vgnd vpwr scs8hd_decap_6
XANTENNA__080__A _076_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_track_16.LATCH_4_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_41_232 vgnd vpwr scs8hd_decap_12
XANTENNA__149__B address[6] vgnd vpwr scs8hd_diode_2
XFILLER_32_276 vgnd vpwr scs8hd_fill_1
XANTENNA__165__A address[4] vgnd vpwr scs8hd_diode_2
XFILLER_23_243 vgnd vpwr scs8hd_fill_1
XANTENNA_mem_top_track_8.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA__075__A _074_/X vgnd vpwr scs8hd_diode_2
XFILLER_23_35 vpwr vgnd scs8hd_fill_2
XFILLER_14_210 vgnd vpwr scs8hd_decap_4
XFILLER_14_276 vgnd vpwr scs8hd_fill_1
X_187_ chanx_right_in[4] chanx_left_out[5] vgnd vpwr scs8hd_buf_2
XANTENNA__135__D _118_/X vgnd vpwr scs8hd_diode_2
Xmux_right_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_right_track_8.INVTX1_1_.scs8hd_inv_1/Y
+ mem_right_track_8.LATCH_1_.latch/Q mux_right_track_8.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
Xmux_left_track_9.INVTX1_0_.scs8hd_inv_1 chany_top_in[2] mux_left_track_9.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_20_213 vgnd vpwr scs8hd_fill_1
XFILLER_20_224 vgnd vpwr scs8hd_decap_12
XFILLER_18_57 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_right_track_0.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_0.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
X_110_ _110_/A _110_/X vgnd vpwr scs8hd_buf_1
XFILLER_34_56 vgnd vpwr scs8hd_decap_6
XFILLER_11_257 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_17.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A mux_left_track_17.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__162__B _158_/X vgnd vpwr scs8hd_diode_2
XFILLER_37_132 vgnd vpwr scs8hd_decap_4
XFILLER_37_121 vgnd vpwr scs8hd_fill_1
XFILLER_20_47 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_top_track_16.tap_buf4_0_.scs8hd_inv_1_A mux_top_track_16.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_28_176 vgnd vpwr scs8hd_decap_8
XFILLER_28_165 vpwr vgnd scs8hd_fill_2
XFILLER_6_27 vgnd vpwr scs8hd_decap_4
XFILLER_3_220 vgnd vpwr scs8hd_decap_12
XFILLER_19_121 vgnd vpwr scs8hd_fill_1
XFILLER_19_165 vpwr vgnd scs8hd_fill_2
XFILLER_34_146 vgnd vpwr scs8hd_fill_1
XANTENNA__157__B _157_/B vgnd vpwr scs8hd_diode_2
XFILLER_19_198 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_left_track_9.LATCH_1_.latch_SLEEPB _133_/Y vgnd vpwr scs8hd_diode_2
XFILLER_25_146 vgnd vpwr scs8hd_fill_1
XFILLER_40_116 vgnd vpwr scs8hd_decap_12
XANTENNA__067__B _078_/B vgnd vpwr scs8hd_diode_2
XANTENNA__083__A _082_/X vgnd vpwr scs8hd_diode_2
XFILLER_25_179 vpwr vgnd scs8hd_fill_2
XFILLER_31_57 vpwr vgnd scs8hd_fill_2
XFILLER_31_149 vgnd vpwr scs8hd_decap_4
XFILLER_31_116 vgnd vpwr scs8hd_decap_4
XPHY_130 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_141 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_152 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_16_102 vgnd vpwr scs8hd_decap_3
XANTENNA_mem_left_track_17.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XPHY_163 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_174 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_185 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_196 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_39_238 vgnd vpwr scs8hd_decap_6
XANTENNA__168__A _099_/A vgnd vpwr scs8hd_diode_2
XFILLER_22_149 vpwr vgnd scs8hd_fill_2
Xmux_left_track_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_left_track_1.INVTX1_0_.scs8hd_inv_1/Y
+ mem_left_track_1.LATCH_0_.latch/Q mux_left_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_left_track_17.INVTX1_0_.scs8hd_inv_1_A chany_top_in[1] vgnd vpwr scs8hd_diode_2
Xmux_top_track_0.INVTX1_0_.scs8hd_inv_1 top_left_grid_pin_13_ mux_top_track_0.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_38_271 vgnd vpwr scs8hd_decap_4
XFILLER_13_127 vgnd vpwr scs8hd_decap_3
XANTENNA__078__A address[1] vgnd vpwr scs8hd_diode_2
XFILLER_42_56 vgnd vpwr scs8hd_decap_6
XFILLER_21_193 vpwr vgnd scs8hd_fill_2
Xmux_left_track_17.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 mux_left_track_17.INVTX1_3_.scs8hd_inv_1/Y
+ mem_left_track_17.LATCH_0_.latch/Q mux_left_track_17.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_3_39 vgnd vpwr scs8hd_decap_12
XANTENNA__170__B _167_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_17.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB mem_left_track_17.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_35_274 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_right_track_8.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A mux_right_track_8.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_16.INVTX1_2_.scs8hd_inv_1_A chanx_left_in[1] vgnd vpwr scs8hd_diode_2
XANTENNA__080__B _099_/A vgnd vpwr scs8hd_diode_2
Xmux_right_track_8.INVTX1_1_.scs8hd_inv_1 chany_top_in[3] mux_right_track_8.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_18_208 vgnd vpwr scs8hd_decap_4
XFILLER_26_241 vgnd vpwr scs8hd_decap_12
Xmem_right_track_0.LATCH_1_.latch data_in mem_right_track_0.LATCH_1_.latch/Q _090_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
Xmux_right_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_right_track_16.INVTX1_1_.scs8hd_inv_1/Y
+ mem_right_track_16.LATCH_1_.latch/Q mux_right_track_16.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
Xmem_top_track_8.LATCH_1_.latch data_in _145_/A _161_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_5_123 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_8.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_TEB mem_right_track_8.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xmux_top_track_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_top_track_0.INVTX1_1_.scs8hd_inv_1/Y
+ mem_top_track_0.LATCH_1_.latch/Q mux_top_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_17_241 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_right_track_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB mem_right_track_0.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__149__C address[5] vgnd vpwr scs8hd_diode_2
XANTENNA__165__B address[3] vgnd vpwr scs8hd_diode_2
XFILLER_4_93 vgnd vpwr scs8hd_decap_12
XANTENNA__091__A address[1] vgnd vpwr scs8hd_diode_2
X_186_ chanx_right_in[5] chanx_left_out[6] vgnd vpwr scs8hd_buf_2
XFILLER_20_203 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_16.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_top_track_16.LATCH_4_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_top_track_0.LATCH_5_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_20_236 vgnd vpwr scs8hd_decap_12
Xmux_left_track_1.INVTX1_3_.scs8hd_inv_1 chanx_right_in[0] mux_left_track_1.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_18_36 vpwr vgnd scs8hd_fill_2
XFILLER_34_68 vgnd vpwr scs8hd_fill_1
XFILLER_11_269 vgnd vpwr scs8hd_decap_8
XANTENNA__086__A _085_/X vgnd vpwr scs8hd_diode_2
XFILLER_1_3 vgnd vpwr scs8hd_decap_12
XANTENNA__162__C _162_/C vgnd vpwr scs8hd_diode_2
XFILLER_6_251 vgnd vpwr scs8hd_decap_4
X_169_ _084_/B _167_/B _169_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_34_3 vgnd vpwr scs8hd_decap_3
XFILLER_37_177 vgnd vpwr scs8hd_decap_4
XANTENNA_mem_right_track_8.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_20_15 vpwr vgnd scs8hd_fill_2
XFILLER_20_59 vgnd vpwr scs8hd_decap_3
XFILLER_29_57 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_top_track_16.LATCH_5_.latch_SLEEPB _167_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mem_left_track_1.LATCH_3_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_10_70 vgnd vpwr scs8hd_decap_12
XFILLER_3_232 vgnd vpwr scs8hd_decap_12
Xmux_left_track_9.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_left_track_9.INVTX1_2_.scs8hd_inv_1/Y
+ mem_left_track_9.LATCH_2_.latch/Q mux_left_track_9.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_42_180 vgnd vpwr scs8hd_decap_6
XFILLER_34_169 vgnd vpwr scs8hd_decap_4
XFILLER_34_125 vpwr vgnd scs8hd_fill_2
XANTENNA__067__C _161_/C vgnd vpwr scs8hd_diode_2
XFILLER_25_114 vgnd vpwr scs8hd_decap_3
XFILLER_25_158 vpwr vgnd scs8hd_fill_2
XFILLER_40_128 vgnd vpwr scs8hd_decap_4
XFILLER_33_180 vgnd vpwr scs8hd_fill_1
XFILLER_31_36 vpwr vgnd scs8hd_fill_2
XFILLER_31_25 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_9.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_left_track_9.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_31_69 vpwr vgnd scs8hd_fill_2
XPHY_131 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_120 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_142 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_153 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_16_158 vgnd vpwr scs8hd_fill_1
XPHY_164 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_175 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_186 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmux_right_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ mem_right_track_0.LATCH_3_.latch/Q mux_right_track_0.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XPHY_197 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_39_206 vpwr vgnd scs8hd_fill_2
XPHY_0 vgnd vpwr scs8hd_decap_3
XANTENNA__168__B _167_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_left_track_1.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__184__A _184_/A vgnd vpwr scs8hd_diode_2
Xmem_left_track_9.LATCH_2_.latch data_in mem_left_track_9.LATCH_2_.latch/Q _132_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA__078__B _078_/B vgnd vpwr scs8hd_diode_2
XANTENNA__094__A address[4] vgnd vpwr scs8hd_diode_2
XFILLER_21_161 vpwr vgnd scs8hd_fill_2
XFILLER_21_172 vpwr vgnd scs8hd_fill_2
Xmem_top_track_14.LATCH_0_.latch data_in _148_/A _164_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_8_154 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _143_/Y vgnd vpwr
+ scs8hd_diode_2
XFILLER_35_253 vpwr vgnd scs8hd_fill_2
XFILLER_12_16 vgnd vpwr scs8hd_decap_4
XFILLER_26_253 vpwr vgnd scs8hd_fill_2
XANTENNA__089__A _088_/X vgnd vpwr scs8hd_diode_2
Xmem_top_track_16.LATCH_3_.latch data_in mem_top_track_16.LATCH_3_.latch/Q _169_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
Xmux_right_track_0.INVTX1_4_.scs8hd_inv_1 right_bottom_grid_pin_5_ mux_right_track_0.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_41_245 vgnd vpwr scs8hd_decap_12
XFILLER_5_135 vgnd vpwr scs8hd_decap_12
Xmux_top_track_14.tap_buf4_0_.scs8hd_inv_1 mux_top_track_14.tap_buf4_0_.scs8hd_inv_1/A
+ _203_/A vgnd vpwr scs8hd_inv_1
XFILLER_32_223 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_1.INVTX1_4_.scs8hd_inv_1_A chanx_right_in[4] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_left_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XANTENNA__165__C _096_/A vgnd vpwr scs8hd_diode_2
XFILLER_4_190 vgnd vpwr scs8hd_decap_12
XFILLER_23_201 vpwr vgnd scs8hd_fill_2
XFILLER_23_245 vgnd vpwr scs8hd_decap_4
XFILLER_2_105 vgnd vpwr scs8hd_decap_12
XANTENNA__091__B address[2] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_0.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB mem_right_track_0.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
X_185_ chanx_right_in[6] chanx_left_out[7] vgnd vpwr scs8hd_buf_2
XANTENNA_mux_left_track_9.INVTX1_6_.scs8hd_inv_1_A left_bottom_grid_pin_7_ vgnd vpwr
+ scs8hd_diode_2
XFILLER_1_171 vgnd vpwr scs8hd_decap_12
XFILLER_20_248 vgnd vpwr scs8hd_decap_12
XANTENNA__192__A _192_/A vgnd vpwr scs8hd_diode_2
XFILLER_34_25 vpwr vgnd scs8hd_fill_2
XFILLER_7_208 vgnd vpwr scs8hd_decap_12
XFILLER_40_90 vpwr vgnd scs8hd_fill_2
X_168_ _099_/A _167_/B _168_/Y vgnd vpwr scs8hd_nor2_4
X_099_ _099_/A _112_/A vgnd vpwr scs8hd_buf_1
XFILLER_27_3 vpwr vgnd scs8hd_fill_2
XFILLER_37_156 vpwr vgnd scs8hd_fill_2
XANTENNA__187__A chanx_right_in[4] vgnd vpwr scs8hd_diode_2
XFILLER_1_62 vgnd vpwr scs8hd_decap_12
Xmux_left_track_9.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2 mux_left_track_9.INVTX1_6_.scs8hd_inv_1/Y
+ mem_left_track_9.LATCH_0_.latch/Q mux_left_track_9.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
Xmux_right_track_8.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_right_track_8.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2/Z
+ mem_right_track_8.LATCH_5_.latch/Q mux_right_track_8.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_20_27 vpwr vgnd scs8hd_fill_2
XFILLER_29_69 vpwr vgnd scs8hd_fill_2
XFILLER_28_145 vpwr vgnd scs8hd_fill_2
XFILLER_28_112 vpwr vgnd scs8hd_fill_2
XANTENNA__097__A _096_/X vgnd vpwr scs8hd_diode_2
XFILLER_10_93 vgnd vpwr scs8hd_decap_12
XFILLER_10_82 vgnd vpwr scs8hd_decap_8
Xmux_right_track_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 mux_right_track_0.INVTX1_4_.scs8hd_inv_1/Y
+ mem_right_track_0.LATCH_1_.latch/Q mux_right_track_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_19_134 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_right_track_8.LATCH_2_.latch_SLEEPB _104_/Y vgnd vpwr scs8hd_diode_2
XFILLER_15_16 vpwr vgnd scs8hd_fill_2
XFILLER_0_225 vgnd vpwr scs8hd_decap_8
XPHY_132 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_121 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_110 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_143 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_154 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_165 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_176 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_187 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_198 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_39_218 vpwr vgnd scs8hd_fill_2
XFILLER_11_6 vpwr vgnd scs8hd_fill_2
XPHY_1 vgnd vpwr scs8hd_decap_3
XFILLER_22_107 vpwr vgnd scs8hd_fill_2
XANTENNA__078__C _162_/C vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_14.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_top_track_14.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_26_59 vgnd vpwr scs8hd_decap_4
XANTENNA_mem_left_track_1.LATCH_5_.latch_SLEEPB _121_/Y vgnd vpwr scs8hd_diode_2
XFILLER_8_166 vgnd vpwr scs8hd_decap_12
XFILLER_35_243 vgnd vpwr scs8hd_fill_1
XANTENNA__195__A chanx_left_in[5] vgnd vpwr scs8hd_diode_2
Xmux_left_track_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_left_track_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ mem_left_track_1.LATCH_4_.latch/Q mux_left_track_1.tap_buf4_0_.scs8hd_inv_1/A vgnd
+ vpwr scs8hd_ebufn_2
XFILLER_37_69 vpwr vgnd scs8hd_fill_2
Xmem_right_track_8.LATCH_2_.latch data_in mem_right_track_8.LATCH_2_.latch/Q _104_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_26_276 vgnd vpwr scs8hd_fill_1
XFILLER_41_257 vgnd vpwr scs8hd_decap_12
XFILLER_5_147 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_right_track_16.LATCH_5_.latch_SLEEPB _111_/Y vgnd vpwr scs8hd_diode_2
XFILLER_32_235 vgnd vpwr scs8hd_decap_12
XFILLER_32_213 vgnd vpwr scs8hd_fill_1
XFILLER_23_16 vpwr vgnd scs8hd_fill_2
XFILLER_23_235 vgnd vpwr scs8hd_decap_8
XFILLER_23_257 vpwr vgnd scs8hd_fill_2
XFILLER_2_117 vgnd vpwr scs8hd_decap_12
XANTENNA__091__C _162_/C vgnd vpwr scs8hd_diode_2
Xmux_right_track_16.INVTX1_5_.scs8hd_inv_1 right_bottom_grid_pin_15_ mux_right_track_16.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
Xmux_left_track_17.INVTX1_6_.scs8hd_inv_1 left_bottom_grid_pin_9_ mux_left_track_17.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
Xmux_right_track_16.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_right_track_16.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2/Z
+ mem_right_track_16.LATCH_5_.latch/Q mux_right_track_16.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
X_184_ _184_/A chanx_left_out[8] vgnd vpwr scs8hd_buf_2
XFILLER_13_71 vpwr vgnd scs8hd_fill_2
XFILLER_13_82 vpwr vgnd scs8hd_fill_2
XFILLER_13_93 vgnd vpwr scs8hd_decap_6
XANTENNA_mem_right_track_16.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
Xmux_top_track_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2 _179_/HI mem_top_track_0.LATCH_5_.latch/Q
+ mux_top_track_0.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XFILLER_18_27 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_top_track_14.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_41_6 vpwr vgnd scs8hd_fill_2
X_098_ _111_/A _106_/B _098_/Y vgnd vpwr scs8hd_nor2_4
X_167_ _167_/A _167_/B _167_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_37_113 vpwr vgnd scs8hd_fill_2
XFILLER_1_74 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_17.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_left_track_17.LATCH_4_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_20_39 vpwr vgnd scs8hd_fill_2
XFILLER_28_135 vgnd vpwr scs8hd_fill_1
XANTENNA_mem_top_track_8.LATCH_0_.latch_SLEEPB _162_/Y vgnd vpwr scs8hd_diode_2
XFILLER_3_245 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_left_track_17.LATCH_3_.latch_SLEEPB _139_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A mux_left_track_1.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_19_113 vpwr vgnd scs8hd_fill_2
XFILLER_34_149 vpwr vgnd scs8hd_fill_2
XFILLER_34_138 vpwr vgnd scs8hd_fill_2
XFILLER_19_92 vpwr vgnd scs8hd_fill_2
XFILLER_19_179 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_17.tap_buf4_0_.scs8hd_inv_1_A mux_left_track_17.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XANTENNA__198__A chanx_left_in[2] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_16.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_TEB mem_right_track_16.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_15_39 vgnd vpwr scs8hd_decap_3
XFILLER_25_138 vpwr vgnd scs8hd_fill_2
XFILLER_0_215 vpwr vgnd scs8hd_fill_2
XFILLER_0_259 vpwr vgnd scs8hd_fill_2
XPHY_100 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_31_108 vpwr vgnd scs8hd_fill_2
XPHY_133 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_122 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_111 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_144 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_155 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_166 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_177 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_188 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_199 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_21_82 vpwr vgnd scs8hd_fill_2
XPHY_2 vgnd vpwr scs8hd_decap_3
XFILLER_15_193 vpwr vgnd scs8hd_fill_2
XFILLER_30_174 vgnd vpwr scs8hd_decap_3
XFILLER_7_62 vgnd vpwr scs8hd_decap_12
Xmux_left_track_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2 mux_left_track_1.INVTX1_5_.scs8hd_inv_1/Y
+ mem_left_track_1.LATCH_2_.latch/Q mux_left_track_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_right_track_0.INVTX1_5_.scs8hd_inv_1_A right_bottom_grid_pin_11_ vgnd
+ vpwr scs8hd_diode_2
XFILLER_26_27 vpwr vgnd scs8hd_fill_2
XFILLER_42_15 vgnd vpwr scs8hd_decap_12
Xmux_left_track_17.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2 _174_/HI mem_left_track_17.LATCH_2_.latch/Q
+ mux_left_track_17.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XFILLER_8_178 vgnd vpwr scs8hd_decap_12
XFILLER_12_152 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_top_track_0.INVTX1_1_.scs8hd_inv_1_A chanx_right_in[1] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_8.INVTX1_7_.scs8hd_inv_1_A chanx_left_in[5] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_9.INVTX1_1_.scs8hd_inv_1_A chany_top_in[5] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_16.tap_buf4_0_.scs8hd_inv_1_A mux_right_track_16.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_41_269 vgnd vpwr scs8hd_decap_8
XFILLER_5_159 vgnd vpwr scs8hd_decap_12
XFILLER_32_258 vgnd vpwr scs8hd_decap_12
XFILLER_32_247 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_top_track_16.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_top_track_16.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xmux_left_track_1.tap_buf4_0_.scs8hd_inv_1 mux_left_track_1.tap_buf4_0_.scs8hd_inv_1/A
+ _192_/A vgnd vpwr scs8hd_inv_1
XFILLER_23_214 vpwr vgnd scs8hd_fill_2
XFILLER_23_39 vpwr vgnd scs8hd_fill_2
XFILLER_2_129 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_left_track_9.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_9_19 vgnd vpwr scs8hd_decap_12
Xmux_top_track_2.tap_buf4_0_.scs8hd_inv_1 mux_top_track_2.tap_buf4_0_.scs8hd_inv_1/A
+ _209_/A vgnd vpwr scs8hd_inv_1
X_183_ _183_/HI _183_/LO vgnd vpwr scs8hd_conb_1
XFILLER_1_184 vgnd vpwr scs8hd_decap_12
XFILLER_38_80 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_right_track_0.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_8.tap_buf4_0_.scs8hd_inv_1_A mux_top_track_8.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
Xmux_top_track_16.INVTX1_1_.scs8hd_inv_1 chanx_right_in[3] mux_top_track_16.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_left_track_9.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A _175_/HI vgnd vpwr
+ scs8hd_diode_2
X_097_ _096_/X _106_/B vgnd vpwr scs8hd_buf_1
XFILLER_6_276 vgnd vpwr scs8hd_fill_1
X_166_ _165_/X _167_/B vgnd vpwr scs8hd_buf_1
XANTENNA_mem_left_track_17.LATCH_4_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_37_169 vpwr vgnd scs8hd_fill_2
XFILLER_1_86 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_left_track_9.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_29_49 vpwr vgnd scs8hd_fill_2
XFILLER_28_169 vgnd vpwr scs8hd_decap_4
XFILLER_28_125 vpwr vgnd scs8hd_fill_2
XFILLER_3_257 vgnd vpwr scs8hd_decap_12
XFILLER_19_71 vpwr vgnd scs8hd_fill_2
XFILLER_19_147 vgnd vpwr scs8hd_decap_3
XFILLER_35_92 vgnd vpwr scs8hd_fill_1
XFILLER_19_169 vgnd vpwr scs8hd_decap_4
X_149_ _118_/A address[6] address[5] _158_/A vgnd vpwr scs8hd_or3_4
XFILLER_33_172 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_16.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_right_track_16.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_0_238 vpwr vgnd scs8hd_fill_2
XFILLER_0_249 vgnd vpwr scs8hd_decap_6
XPHY_134 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_123 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_112 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_101 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_16_128 vpwr vgnd scs8hd_fill_2
XPHY_145 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_156 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_167 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_178 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_189 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_183 vgnd vpwr scs8hd_fill_1
XPHY_3 vgnd vpwr scs8hd_decap_3
XFILLER_30_186 vpwr vgnd scs8hd_fill_2
XFILLER_7_74 vgnd vpwr scs8hd_decap_12
XFILLER_42_27 vgnd vpwr scs8hd_decap_4
XFILLER_21_197 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_top_track_0.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_29_231 vgnd vpwr scs8hd_decap_12
XFILLER_16_50 vgnd vpwr scs8hd_fill_1
XFILLER_16_83 vpwr vgnd scs8hd_fill_2
XFILLER_32_71 vpwr vgnd scs8hd_fill_2
XFILLER_35_245 vgnd vpwr scs8hd_decap_8
XFILLER_35_223 vpwr vgnd scs8hd_fill_2
XFILLER_35_212 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_right_track_16.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_16.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_37_27 vpwr vgnd scs8hd_fill_2
XFILLER_37_16 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_8.tap_buf4_0_.scs8hd_inv_1_A mux_right_track_8.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_27_93 vpwr vgnd scs8hd_fill_2
XFILLER_17_201 vpwr vgnd scs8hd_fill_2
XFILLER_17_245 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_right_track_8.LATCH_4_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_16.INVTX1_3_.scs8hd_inv_1_A right_bottom_grid_pin_3_ vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mux_top_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_top_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
X_182_ _182_/HI _182_/LO vgnd vpwr scs8hd_conb_1
Xmux_left_track_1.INVTX1_0_.scs8hd_inv_1 chany_top_in[0] mux_left_track_1.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_14_215 vgnd vpwr scs8hd_decap_12
XFILLER_1_196 vgnd vpwr scs8hd_decap_12
XANTENNA__100__A _112_/A vgnd vpwr scs8hd_diode_2
XFILLER_9_263 vgnd vpwr scs8hd_decap_12
XFILLER_20_207 vgnd vpwr scs8hd_decap_6
XFILLER_18_18 vpwr vgnd scs8hd_fill_2
XFILLER_34_17 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_right_track_0.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_10_251 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_top_track_16.LATCH_2_.latch_SLEEPB _170_/Y vgnd vpwr scs8hd_diode_2
X_165_ address[4] address[3] _096_/A _165_/X vgnd vpwr scs8hd_or3_4
XFILLER_40_93 vgnd vpwr scs8hd_decap_8
X_096_ _096_/A _096_/B _096_/X vgnd vpwr scs8hd_or2_4
XFILLER_1_98 vgnd vpwr scs8hd_decap_12
Xmem_top_track_0.LATCH_1_.latch data_in mem_top_track_0.LATCH_1_.latch/Q _156_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_20_19 vpwr vgnd scs8hd_fill_2
XFILLER_29_28 vpwr vgnd scs8hd_fill_2
XFILLER_3_269 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_right_track_0.INVTX1_0_.scs8hd_inv_1_A chany_top_in[2] vgnd vpwr scs8hd_diode_2
XFILLER_19_126 vpwr vgnd scs8hd_fill_2
XFILLER_42_140 vgnd vpwr scs8hd_decap_12
XFILLER_35_71 vgnd vpwr scs8hd_decap_4
XFILLER_27_170 vgnd vpwr scs8hd_decap_3
Xmux_top_track_14.INVTX1_1_.scs8hd_inv_1 chanx_left_in[8] mux_top_track_14.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_left_track_9.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB mem_left_track_9.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_left_track_1.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
X_148_ _148_/A _148_/Y vgnd vpwr scs8hd_inv_8
X_079_ _078_/X _099_/A vgnd vpwr scs8hd_buf_1
XFILLER_25_3 vgnd vpwr scs8hd_decap_3
XFILLER_33_195 vpwr vgnd scs8hd_fill_2
Xmem_left_track_17.LATCH_4_.latch data_in mem_left_track_17.LATCH_4_.latch/Q _138_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_right_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XPHY_135 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_124 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_113 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_102 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_146 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_157 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_16_107 vgnd vpwr scs8hd_decap_4
XFILLER_24_151 vpwr vgnd scs8hd_fill_2
XFILLER_24_195 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_8.INVTX1_2_.scs8hd_inv_1_A chany_top_in[6] vgnd vpwr scs8hd_diode_2
XPHY_168 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_179 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_21_62 vgnd vpwr scs8hd_decap_4
XFILLER_21_95 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_top_track_0.LATCH_4_.latch_SLEEPB _153_/Y vgnd vpwr scs8hd_diode_2
XFILLER_30_154 vgnd vpwr scs8hd_decap_3
XFILLER_30_143 vpwr vgnd scs8hd_fill_2
XFILLER_30_110 vgnd vpwr scs8hd_fill_1
Xmux_left_track_9.INVTX1_5_.scs8hd_inv_1 left_bottom_grid_pin_1_ mux_left_track_9.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XPHY_4 vgnd vpwr scs8hd_decap_3
XFILLER_15_151 vpwr vgnd scs8hd_fill_2
XFILLER_7_86 vgnd vpwr scs8hd_decap_12
XFILLER_7_31 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_left_track_9.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_38_276 vgnd vpwr scs8hd_fill_1
XFILLER_21_132 vpwr vgnd scs8hd_fill_2
XFILLER_21_143 vpwr vgnd scs8hd_fill_2
XFILLER_21_165 vpwr vgnd scs8hd_fill_2
XFILLER_21_176 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_top_track_2.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB _144_/Y vgnd vpwr
+ scs8hd_diode_2
XFILLER_29_243 vgnd vpwr scs8hd_fill_1
XFILLER_12_154 vgnd vpwr scs8hd_decap_12
XFILLER_16_62 vpwr vgnd scs8hd_fill_2
XFILLER_32_50 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_17.INVTX1_6_.scs8hd_inv_1_A left_bottom_grid_pin_9_ vgnd vpwr
+ scs8hd_diode_2
XANTENNA__103__A _103_/A vgnd vpwr scs8hd_diode_2
Xmux_right_track_0.INVTX1_1_.scs8hd_inv_1 chany_top_in[5] mux_right_track_0.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_26_202 vgnd vpwr scs8hd_decap_12
XFILLER_32_205 vpwr vgnd scs8hd_fill_2
XFILLER_17_257 vgnd vpwr scs8hd_decap_12
XFILLER_27_72 vpwr vgnd scs8hd_fill_2
XFILLER_4_32 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_9.tap_buf4_0_.scs8hd_inv_1_A mux_left_track_9.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_23_249 vgnd vpwr scs8hd_fill_1
XFILLER_14_227 vgnd vpwr scs8hd_decap_12
X_181_ _181_/HI _181_/LO vgnd vpwr scs8hd_conb_1
XFILLER_13_30 vpwr vgnd scs8hd_fill_2
XFILLER_22_271 vgnd vpwr scs8hd_decap_4
XFILLER_38_93 vgnd vpwr scs8hd_decap_8
Xmem_left_track_1.LATCH_2_.latch data_in mem_left_track_1.LATCH_2_.latch/Q _124_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA__100__B _106_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_17.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_left_track_17.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_9_275 vpwr vgnd scs8hd_fill_2
XFILLER_9_253 vpwr vgnd scs8hd_fill_2
XFILLER_9_220 vgnd vpwr scs8hd_decap_12
XFILLER_34_29 vpwr vgnd scs8hd_fill_2
XFILLER_11_208 vgnd vpwr scs8hd_decap_12
XANTENNA__201__A _201_/A vgnd vpwr scs8hd_diode_2
Xmem_right_track_16.LATCH_3_.latch data_in mem_right_track_16.LATCH_3_.latch/Q _113_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
Xmux_right_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_0.INVTX1_0_.scs8hd_inv_1/Y
+ mem_right_track_0.LATCH_0_.latch/Q mux_right_track_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_right_track_16.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_16.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
X_095_ _095_/A address[3] _096_/B vgnd vpwr scs8hd_or2_4
XFILLER_10_263 vgnd vpwr scs8hd_decap_12
XFILLER_24_84 vgnd vpwr scs8hd_decap_8
X_164_ _095_/A _109_/B _158_/X _162_/C _164_/Y vgnd vpwr scs8hd_nor4_4
XFILLER_27_7 vgnd vpwr scs8hd_decap_3
XANTENNA__111__A _111_/A vgnd vpwr scs8hd_diode_2
XFILLER_37_138 vpwr vgnd scs8hd_fill_2
XFILLER_1_33 vpwr vgnd scs8hd_fill_2
XFILLER_29_18 vpwr vgnd scs8hd_fill_2
Xmux_right_track_8.INVTX1_6_.scs8hd_inv_1 chanx_left_in[1] mux_right_track_8.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_28_149 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_16.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_top_track_16.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_34_119 vgnd vpwr scs8hd_decap_4
XFILLER_42_152 vgnd vpwr scs8hd_decap_3
XANTENNA__106__A _125_/A vgnd vpwr scs8hd_diode_2
X_147_ _147_/A _147_/Y vgnd vpwr scs8hd_inv_8
XANTENNA_mux_top_track_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A mux_top_track_0.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
X_078_ address[1] _078_/B _162_/C _078_/X vgnd vpwr scs8hd_or3_4
XFILLER_25_119 vgnd vpwr scs8hd_decap_3
XANTENNA_mem_top_track_0.LATCH_2_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_0_207 vgnd vpwr scs8hd_decap_8
XPHY_136 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_125 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_114 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_103 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_147 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_158 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_169 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_130 vgnd vpwr scs8hd_decap_6
XFILLER_24_163 vgnd vpwr scs8hd_decap_3
Xmux_top_track_16.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_top_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ mem_top_track_16.LATCH_3_.latch/Q mux_top_track_16.tap_buf4_0_.scs8hd_inv_1/A vgnd
+ vpwr scs8hd_ebufn_2
XANTENNA_mem_left_track_1.LATCH_2_.latch_SLEEPB _124_/Y vgnd vpwr scs8hd_diode_2
XPHY_5 vgnd vpwr scs8hd_decap_3
XFILLER_15_130 vpwr vgnd scs8hd_fill_2
XFILLER_30_166 vgnd vpwr scs8hd_decap_8
XFILLER_30_122 vpwr vgnd scs8hd_fill_2
XFILLER_7_43 vgnd vpwr scs8hd_decap_12
XFILLER_7_98 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_16.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_top_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_16_41 vgnd vpwr scs8hd_decap_3
Xmux_left_track_17.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_left_track_17.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ mem_left_track_17.LATCH_3_.latch/Q mux_left_track_17.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_12_166 vgnd vpwr scs8hd_decap_12
XFILLER_32_84 vgnd vpwr scs8hd_decap_6
XANTENNA_mem_right_track_16.LATCH_3_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_35_258 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_right_track_16.LATCH_2_.latch_SLEEPB _114_/Y vgnd vpwr scs8hd_diode_2
XANTENNA__204__A chanx_left_in[4] vgnd vpwr scs8hd_diode_2
XFILLER_17_214 vpwr vgnd scs8hd_fill_2
XFILLER_17_225 vpwr vgnd scs8hd_fill_2
XFILLER_17_269 vgnd vpwr scs8hd_decap_8
XFILLER_27_62 vgnd vpwr scs8hd_fill_1
XANTENNA_mem_top_track_16.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_0.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__114__A _124_/A vgnd vpwr scs8hd_diode_2
Xmux_left_track_17.INVTX1_3_.scs8hd_inv_1 chanx_right_in[2] mux_left_track_17.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
Xmux_right_track_16.INVTX1_2_.scs8hd_inv_1 chany_top_in[7] mux_right_track_16.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_4_44 vgnd vpwr scs8hd_decap_12
Xmux_right_track_8.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_right_track_8.INVTX1_2_.scs8hd_inv_1/Y
+ mem_right_track_8.LATCH_2_.latch/Q mux_right_track_8.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_left_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_left_track_17.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_14_239 vgnd vpwr scs8hd_decap_12
XFILLER_13_20 vgnd vpwr scs8hd_decap_3
XFILLER_13_53 vpwr vgnd scs8hd_fill_2
X_180_ _180_/HI _180_/LO vgnd vpwr scs8hd_conb_1
XFILLER_13_75 vgnd vpwr scs8hd_decap_4
XFILLER_13_86 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_top_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_top_track_8.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_1_110 vgnd vpwr scs8hd_decap_12
XFILLER_38_61 vgnd vpwr scs8hd_fill_1
XFILLER_9_232 vgnd vpwr scs8hd_decap_12
XANTENNA__109__A _095_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_17.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A mux_left_track_17.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_17.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB mem_left_track_17.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_24_41 vpwr vgnd scs8hd_fill_2
XFILLER_6_202 vgnd vpwr scs8hd_decap_12
X_094_ address[4] _095_/A vgnd vpwr scs8hd_inv_8
X_163_ _095_/A _109_/B _158_/X _161_/C _163_/Y vgnd vpwr scs8hd_nor4_4
XANTENNA__111__B _110_/X vgnd vpwr scs8hd_diode_2
XFILLER_37_117 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_left_track_17.LATCH_0_.latch_SLEEPB _142_/Y vgnd vpwr scs8hd_diode_2
Xmem_right_track_0.LATCH_2_.latch data_in mem_right_track_0.LATCH_2_.latch/Q _087_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_36_183 vgnd vpwr scs8hd_fill_1
XFILLER_19_52 vpwr vgnd scs8hd_fill_2
XFILLER_19_96 vpwr vgnd scs8hd_fill_2
XFILLER_19_117 vgnd vpwr scs8hd_decap_4
XFILLER_35_95 vgnd vpwr scs8hd_fill_1
X_146_ _146_/A _146_/Y vgnd vpwr scs8hd_inv_8
XANTENNA__106__B _106_/B vgnd vpwr scs8hd_diode_2
X_077_ address[0] _162_/C vgnd vpwr scs8hd_buf_1
XANTENNA__122__A _112_/A vgnd vpwr scs8hd_diode_2
XFILLER_32_6 vgnd vpwr scs8hd_decap_4
XFILLER_33_153 vgnd vpwr scs8hd_fill_1
XFILLER_18_161 vgnd vpwr scs8hd_decap_4
Xmux_left_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_left_track_1.INVTX1_1_.scs8hd_inv_1/Y
+ mem_left_track_1.LATCH_1_.latch/Q mux_left_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_left_track_17.INVTX1_1_.scs8hd_inv_1_A chany_top_in[4] vgnd vpwr scs8hd_diode_2
XPHY_137 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_126 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_115 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_104 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_148 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_159 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__207__A chanx_right_in[5] vgnd vpwr scs8hd_diode_2
XFILLER_24_175 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_right_track_8.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xmux_left_track_17.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 mux_left_track_17.INVTX1_4_.scs8hd_inv_1/Y
+ mem_left_track_17.LATCH_1_.latch/Q mux_left_track_17.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_21_42 vpwr vgnd scs8hd_fill_2
XFILLER_21_53 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_16.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_top_track_16.LATCH_5_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XPHY_6 vgnd vpwr scs8hd_decap_3
XFILLER_15_164 vpwr vgnd scs8hd_fill_2
XFILLER_15_175 vpwr vgnd scs8hd_fill_2
XFILLER_7_55 vgnd vpwr scs8hd_decap_6
XFILLER_15_197 vpwr vgnd scs8hd_fill_2
XANTENNA__117__A enable vgnd vpwr scs8hd_diode_2
XFILLER_30_3 vgnd vpwr scs8hd_decap_3
X_129_ _111_/A _132_/B _129_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA_mux_top_track_16.INVTX1_3_.scs8hd_inv_1_A chanx_left_in[7] vgnd vpwr scs8hd_diode_2
XFILLER_29_245 vgnd vpwr scs8hd_decap_12
Xmux_right_track_16.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_right_track_16.INVTX1_2_.scs8hd_inv_1/Y
+ mem_right_track_16.LATCH_2_.latch/Q mux_right_track_16.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_8_105 vgnd vpwr scs8hd_decap_12
XFILLER_12_134 vgnd vpwr scs8hd_decap_12
XFILLER_12_178 vgnd vpwr scs8hd_decap_12
Xmux_top_track_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_top_track_0.INVTX1_2_.scs8hd_inv_1/Y
+ mem_top_track_0.LATCH_2_.latch/Q mux_top_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_right_track_8.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A _178_/HI vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mem_right_track_0.LATCH_3_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_7_171 vgnd vpwr scs8hd_decap_12
XFILLER_34_270 vgnd vpwr scs8hd_decap_4
XFILLER_26_259 vgnd vpwr scs8hd_decap_12
Xmux_right_track_8.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_8.INVTX1_6_.scs8hd_inv_1/Y
+ mem_right_track_8.LATCH_0_.latch/Q mux_right_track_8.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_32_218 vgnd vpwr scs8hd_decap_3
XANTENNA__114__B _110_/X vgnd vpwr scs8hd_diode_2
XFILLER_4_141 vgnd vpwr scs8hd_decap_12
XFILLER_4_56 vgnd vpwr scs8hd_decap_12
XANTENNA__130__A _112_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_9.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_left_track_9.LATCH_4_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_23_218 vpwr vgnd scs8hd_fill_2
XFILLER_31_262 vpwr vgnd scs8hd_fill_2
XFILLER_22_240 vgnd vpwr scs8hd_decap_12
XFILLER_13_10 vgnd vpwr scs8hd_decap_4
Xmem_left_track_9.LATCH_3_.latch data_in mem_left_track_9.LATCH_3_.latch/Q _131_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_38_84 vgnd vpwr scs8hd_decap_8
XANTENNA__109__B _109_/B vgnd vpwr scs8hd_diode_2
XFILLER_13_262 vgnd vpwr scs8hd_decap_12
Xmem_top_track_14.LATCH_1_.latch data_in _147_/A _163_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA__125__A _125_/A vgnd vpwr scs8hd_diode_2
XFILLER_39_192 vgnd vpwr scs8hd_decap_8
X_162_ _096_/B _158_/X _162_/C _162_/Y vgnd vpwr scs8hd_nor3_4
XFILLER_24_53 vgnd vpwr scs8hd_fill_1
XFILLER_10_276 vgnd vpwr scs8hd_fill_1
X_093_ _076_/B _172_/A _093_/Y vgnd vpwr scs8hd_nor2_4
Xmem_top_track_16.LATCH_4_.latch data_in mem_top_track_16.LATCH_4_.latch/Q _168_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_left_track_17.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB mem_left_track_17.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_28_129 vgnd vpwr scs8hd_decap_6
XFILLER_36_195 vgnd vpwr scs8hd_decap_8
XFILLER_27_184 vgnd vpwr scs8hd_decap_3
XFILLER_19_75 vgnd vpwr scs8hd_decap_4
XFILLER_42_187 vgnd vpwr scs8hd_decap_12
X_145_ _145_/A _145_/Y vgnd vpwr scs8hd_inv_8
Xmux_right_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_right_track_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ mem_right_track_0.LATCH_4_.latch/Q mux_right_track_0.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
X_076_ _111_/A _076_/B _076_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA__122__B _125_/B vgnd vpwr scs8hd_diode_2
XFILLER_33_176 vgnd vpwr scs8hd_decap_4
XFILLER_33_132 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_14.INVTX1_0_.scs8hd_inv_1_A chanx_left_in[2] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_0.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_TEB mem_right_track_0.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XPHY_116 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_105 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_138 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_127 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_149 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_30_102 vpwr vgnd scs8hd_fill_2
XPHY_7 vgnd vpwr scs8hd_decap_3
XFILLER_15_143 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_right_track_0.LATCH_3_.latch_SLEEPB _084_/Y vgnd vpwr scs8hd_diode_2
X_128_ _127_/X _132_/B vgnd vpwr scs8hd_buf_1
XANTENNA__133__A _125_/A vgnd vpwr scs8hd_diode_2
Xmux_right_track_16.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_16.INVTX1_6_.scs8hd_inv_1/Y
+ mem_right_track_16.LATCH_0_.latch/Q mux_right_track_16.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_38_235 vgnd vpwr scs8hd_decap_12
XFILLER_38_224 vgnd vpwr scs8hd_decap_8
XFILLER_38_213 vgnd vpwr scs8hd_fill_1
XFILLER_29_257 vgnd vpwr scs8hd_decap_12
XFILLER_29_202 vpwr vgnd scs8hd_fill_2
XFILLER_16_87 vgnd vpwr scs8hd_decap_3
XFILLER_8_117 vgnd vpwr scs8hd_decap_12
XFILLER_12_146 vgnd vpwr scs8hd_decap_6
XANTENNA_mux_left_track_1.INVTX1_5_.scs8hd_inv_1_A left_top_grid_pin_10_ vgnd vpwr
+ scs8hd_diode_2
XFILLER_35_227 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_2.tap_buf4_0_.scs8hd_inv_1_A mux_top_track_2.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XANTENNA__128__A _127_/X vgnd vpwr scs8hd_diode_2
Xmux_top_track_2.INVTX1_2_.scs8hd_inv_1 chanx_right_in[8] mux_top_track_2.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_41_208 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_right_track_8.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_27_42 vpwr vgnd scs8hd_fill_2
XFILLER_27_53 vpwr vgnd scs8hd_fill_2
XFILLER_40_274 vgnd vpwr scs8hd_fill_1
XFILLER_40_230 vgnd vpwr scs8hd_decap_12
XFILLER_27_97 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_9.INVTX1_7_.scs8hd_inv_1_A left_bottom_grid_pin_13_ vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mem_top_track_2.LATCH_0_.latch_SLEEPB _160_/Y vgnd vpwr scs8hd_diode_2
XFILLER_4_68 vgnd vpwr scs8hd_decap_12
XANTENNA__130__B _132_/B vgnd vpwr scs8hd_diode_2
XFILLER_16_271 vgnd vpwr scs8hd_decap_4
XFILLER_31_274 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_top_track_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_top_track_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_22_252 vgnd vpwr scs8hd_decap_3
XFILLER_13_99 vgnd vpwr scs8hd_fill_1
XFILLER_38_30 vgnd vpwr scs8hd_fill_1
XFILLER_1_123 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_left_track_1.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__125__B _125_/B vgnd vpwr scs8hd_diode_2
XANTENNA__109__C _096_/A vgnd vpwr scs8hd_diode_2
XFILLER_9_245 vgnd vpwr scs8hd_decap_8
XFILLER_13_274 vgnd vpwr scs8hd_decap_3
XANTENNA__141__A _125_/A vgnd vpwr scs8hd_diode_2
Xmux_left_track_9.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2 mux_left_track_9.INVTX1_7_.scs8hd_inv_1/Y
+ mem_left_track_9.LATCH_1_.latch/Q mux_left_track_9.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
X_161_ _096_/B _158_/X _161_/C _161_/Y vgnd vpwr scs8hd_nor3_4
XFILLER_6_215 vgnd vpwr scs8hd_decap_12
XFILLER_24_65 vpwr vgnd scs8hd_fill_2
XFILLER_6_259 vgnd vpwr scs8hd_decap_12
X_092_ _091_/X _172_/A vgnd vpwr scs8hd_buf_1
Xmux_right_track_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2 mux_right_track_0.INVTX1_5_.scs8hd_inv_1/Y
+ mem_right_track_0.LATCH_2_.latch/Q mux_right_track_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
Xmem_right_track_8.LATCH_3_.latch data_in mem_right_track_8.LATCH_3_.latch/Q _102_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA__136__A _136_/A vgnd vpwr scs8hd_diode_2
XFILLER_36_141 vpwr vgnd scs8hd_fill_2
XFILLER_28_108 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_left_track_9.LATCH_3_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_35_53 vpwr vgnd scs8hd_fill_2
XFILLER_27_196 vpwr vgnd scs8hd_fill_2
XFILLER_27_163 vpwr vgnd scs8hd_fill_2
XFILLER_42_199 vgnd vpwr scs8hd_decap_12
X_144_ _144_/A _144_/Y vgnd vpwr scs8hd_inv_8
X_075_ _074_/X _076_/B vgnd vpwr scs8hd_buf_1
XFILLER_2_251 vgnd vpwr scs8hd_decap_12
XFILLER_18_174 vgnd vpwr scs8hd_decap_12
XFILLER_33_199 vgnd vpwr scs8hd_decap_3
XANTENNA_mem_top_track_0.LATCH_1_.latch_SLEEPB _156_/Y vgnd vpwr scs8hd_diode_2
XPHY_128 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_117 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_106 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_139 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_left_track_9.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_left_track_9.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
Xmux_left_track_9.INVTX1_2_.scs8hd_inv_1 chany_top_in[8] mux_left_track_9.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_24_122 vpwr vgnd scs8hd_fill_2
XFILLER_24_199 vgnd vpwr scs8hd_decap_4
XFILLER_21_66 vgnd vpwr scs8hd_fill_1
XFILLER_21_99 vpwr vgnd scs8hd_fill_2
XFILLER_30_147 vgnd vpwr scs8hd_decap_4
XPHY_8 vgnd vpwr scs8hd_decap_3
XANTENNA__133__B _132_/B vgnd vpwr scs8hd_diode_2
X_127_ address[4] _109_/B address[5] _118_/X _127_/X vgnd vpwr scs8hd_or4_4
XFILLER_38_247 vgnd vpwr scs8hd_decap_12
XFILLER_21_114 vpwr vgnd scs8hd_fill_2
XFILLER_21_136 vpwr vgnd scs8hd_fill_2
XFILLER_21_147 vgnd vpwr scs8hd_decap_3
Xmux_left_track_1.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_left_track_1.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2/Z
+ mem_left_track_1.LATCH_5_.latch/Q mux_left_track_1.tap_buf4_0_.scs8hd_inv_1/A vgnd
+ vpwr scs8hd_ebufn_2
XFILLER_29_269 vgnd vpwr scs8hd_decap_8
XANTENNA_mem_top_track_14.LATCH_0_.latch_SLEEPB _164_/Y vgnd vpwr scs8hd_diode_2
XFILLER_16_66 vpwr vgnd scs8hd_fill_2
XFILLER_32_54 vgnd vpwr scs8hd_decap_4
XFILLER_32_32 vgnd vpwr scs8hd_decap_4
XFILLER_8_129 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_17.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_left_track_17.LATCH_5_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_35_239 vgnd vpwr scs8hd_decap_4
XFILLER_35_217 vgnd vpwr scs8hd_decap_3
XANTENNA__144__A _144_/A vgnd vpwr scs8hd_diode_2
XFILLER_7_184 vgnd vpwr scs8hd_decap_12
Xmux_top_track_14.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_top_track_14.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ _147_/A mux_top_track_14.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XANTENNA_mem_left_track_9.LATCH_3_.latch_SLEEPB _131_/Y vgnd vpwr scs8hd_diode_2
XFILLER_32_209 vgnd vpwr scs8hd_decap_4
XFILLER_27_21 vpwr vgnd scs8hd_fill_2
XFILLER_27_76 vpwr vgnd scs8hd_fill_2
XFILLER_40_242 vgnd vpwr scs8hd_decap_12
XFILLER_4_154 vgnd vpwr scs8hd_decap_12
XFILLER_31_253 vpwr vgnd scs8hd_fill_2
XANTENNA__139__A _113_/A vgnd vpwr scs8hd_diode_2
XFILLER_13_45 vpwr vgnd scs8hd_fill_2
Xmux_top_track_0.INVTX1_2_.scs8hd_inv_1 chanx_right_in[7] mux_top_track_0.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_38_53 vgnd vpwr scs8hd_decap_8
XFILLER_38_42 vpwr vgnd scs8hd_fill_2
XFILLER_1_135 vgnd vpwr scs8hd_decap_12
XFILLER_13_220 vgnd vpwr scs8hd_decap_12
XFILLER_13_253 vpwr vgnd scs8hd_fill_2
XANTENNA__141__B _136_/X vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_left_track_1.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_track_0.LATCH_5_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_39_150 vgnd vpwr scs8hd_decap_4
Xmux_right_track_8.INVTX1_3_.scs8hd_inv_1 right_bottom_grid_pin_1_ mux_right_track_8.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_40_32 vgnd vpwr scs8hd_decap_12
X_160_ _074_/A _158_/X _162_/C _160_/Y vgnd vpwr scs8hd_nor3_4
XFILLER_6_227 vgnd vpwr scs8hd_decap_12
X_091_ address[1] address[2] _162_/C _091_/X vgnd vpwr scs8hd_or3_4
XANTENNA_mem_top_track_2.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_1_15 vgnd vpwr scs8hd_decap_12
XFILLER_1_37 vgnd vpwr scs8hd_decap_12
XANTENNA__152__A _167_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_1.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A mux_left_track_1.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_36_175 vgnd vpwr scs8hd_decap_8
XFILLER_36_164 vpwr vgnd scs8hd_fill_2
XFILLER_36_120 vgnd vpwr scs8hd_decap_3
XFILLER_10_46 vgnd vpwr scs8hd_decap_12
XFILLER_10_35 vgnd vpwr scs8hd_decap_8
XFILLER_3_208 vgnd vpwr scs8hd_decap_12
XFILLER_27_142 vgnd vpwr scs8hd_decap_4
XFILLER_19_11 vpwr vgnd scs8hd_fill_2
XFILLER_19_109 vpwr vgnd scs8hd_fill_2
XFILLER_42_156 vgnd vpwr scs8hd_decap_12
XFILLER_42_112 vgnd vpwr scs8hd_fill_1
XFILLER_27_175 vpwr vgnd scs8hd_fill_2
X_143_ _143_/A _143_/Y vgnd vpwr scs8hd_inv_8
X_074_ _074_/A _096_/A _074_/X vgnd vpwr scs8hd_or2_4
XFILLER_2_263 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_2.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A mux_top_track_2.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_33_112 vpwr vgnd scs8hd_fill_2
XFILLER_33_101 vpwr vgnd scs8hd_fill_2
XFILLER_18_120 vgnd vpwr scs8hd_decap_6
XFILLER_18_197 vpwr vgnd scs8hd_fill_2
XFILLER_33_156 vgnd vpwr scs8hd_decap_3
XANTENNA__147__A _147_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_1.INVTX1_0_.scs8hd_inv_1_A chany_top_in[0] vgnd vpwr scs8hd_diode_2
XFILLER_2_80 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_0.INVTX1_6_.scs8hd_inv_1_A chanx_left_in[0] vgnd vpwr scs8hd_diode_2
Xmux_left_track_1.INVTX1_5_.scs8hd_inv_1 left_top_grid_pin_10_ mux_left_track_1.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XPHY_129 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_118 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_107 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_145 vgnd vpwr scs8hd_decap_4
XFILLER_21_12 vpwr vgnd scs8hd_fill_2
XFILLER_21_78 vpwr vgnd scs8hd_fill_2
XPHY_9 vgnd vpwr scs8hd_decap_3
XFILLER_30_126 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_top_track_16.LATCH_3_.latch_D data_in vgnd vpwr scs8hd_diode_2
X_126_ _108_/A _125_/B _126_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_38_259 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_0.INVTX1_2_.scs8hd_inv_1_A chanx_right_in[7] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_9.INVTX1_2_.scs8hd_inv_1_A chany_top_in[8] vgnd vpwr scs8hd_diode_2
XFILLER_16_12 vpwr vgnd scs8hd_fill_2
XFILLER_16_23 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_9.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_left_track_9.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__160__A _074_/A vgnd vpwr scs8hd_diode_2
X_109_ _095_/A _109_/B _096_/A _110_/A vgnd vpwr scs8hd_or3_4
XFILLER_7_196 vgnd vpwr scs8hd_decap_12
XFILLER_26_229 vgnd vpwr scs8hd_decap_12
XFILLER_26_218 vgnd vpwr scs8hd_decap_8
Xmux_left_track_17.INVTX1_0_.scs8hd_inv_1 chany_top_in[1] mux_left_track_17.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_top_track_14.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_top_track_14.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__070__A address[3] vgnd vpwr scs8hd_diode_2
XFILLER_17_218 vpwr vgnd scs8hd_fill_2
XFILLER_17_229 vgnd vpwr scs8hd_decap_12
XFILLER_40_276 vgnd vpwr scs8hd_fill_1
XFILLER_40_254 vgnd vpwr scs8hd_decap_12
XFILLER_4_166 vgnd vpwr scs8hd_decap_12
XFILLER_4_15 vgnd vpwr scs8hd_decap_12
XFILLER_31_243 vgnd vpwr scs8hd_fill_1
XANTENNA__155__A _124_/A vgnd vpwr scs8hd_diode_2
XANTENNA__139__B _136_/X vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_9.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A mux_left_track_9.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_13_57 vpwr vgnd scs8hd_fill_2
XANTENNA__065__A address[2] vgnd vpwr scs8hd_diode_2
XFILLER_22_276 vgnd vpwr scs8hd_fill_1
XFILLER_1_147 vgnd vpwr scs8hd_decap_12
XFILLER_38_76 vpwr vgnd scs8hd_fill_2
XFILLER_38_65 vgnd vpwr scs8hd_decap_8
XFILLER_38_32 vgnd vpwr scs8hd_decap_6
XFILLER_13_232 vgnd vpwr scs8hd_decap_12
XFILLER_0_180 vgnd vpwr scs8hd_decap_6
XFILLER_0_191 vpwr vgnd scs8hd_fill_2
XFILLER_39_173 vgnd vpwr scs8hd_decap_3
XFILLER_24_23 vpwr vgnd scs8hd_fill_2
XFILLER_24_45 vpwr vgnd scs8hd_fill_2
XFILLER_40_66 vgnd vpwr scs8hd_decap_12
XFILLER_40_55 vgnd vpwr scs8hd_decap_8
XFILLER_40_44 vgnd vpwr scs8hd_decap_8
XFILLER_10_202 vgnd vpwr scs8hd_decap_12
XFILLER_6_239 vgnd vpwr scs8hd_decap_12
X_090_ _076_/B _090_/B _090_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_6_3 vgnd vpwr scs8hd_decap_12
Xmux_top_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_top_track_16.INVTX1_0_.scs8hd_inv_1/Y
+ mem_top_track_16.LATCH_0_.latch/Q mux_top_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
Xmux_right_track_0.INVTX1_6_.scs8hd_inv_1 chanx_left_in[0] mux_right_track_0.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_1_27 vgnd vpwr scs8hd_decap_3
XFILLER_1_49 vgnd vpwr scs8hd_decap_12
XANTENNA__152__B _157_/B vgnd vpwr scs8hd_diode_2
XFILLER_36_154 vgnd vpwr scs8hd_fill_1
XANTENNA_mem_left_track_17.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_10_58 vgnd vpwr scs8hd_decap_12
XFILLER_35_22 vpwr vgnd scs8hd_fill_2
Xmux_left_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_left_track_17.INVTX1_0_.scs8hd_inv_1/Y
+ mem_left_track_17.LATCH_0_.latch/Q mux_left_track_17.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_27_132 vgnd vpwr scs8hd_decap_4
XFILLER_19_34 vgnd vpwr scs8hd_decap_3
XFILLER_19_56 vgnd vpwr scs8hd_decap_3
XFILLER_42_168 vgnd vpwr scs8hd_decap_12
XFILLER_35_88 vgnd vpwr scs8hd_decap_4
XFILLER_35_77 vpwr vgnd scs8hd_fill_2
X_142_ _108_/A _136_/X _142_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA_mux_right_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_right_track_16.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
X_073_ enable _118_/B address[5] _096_/A vgnd vpwr scs8hd_nand3_4
XFILLER_33_168 vpwr vgnd scs8hd_fill_2
XFILLER_18_132 vgnd vpwr scs8hd_decap_4
XANTENNA__163__A _095_/A vgnd vpwr scs8hd_diode_2
XFILLER_24_102 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_top_track_2.INVTX1_0_.scs8hd_inv_1_A top_right_grid_pin_11_ vgnd vpwr
+ scs8hd_diode_2
XPHY_119 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_108 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_168 vgnd vpwr scs8hd_decap_3
XFILLER_24_179 vgnd vpwr scs8hd_decap_4
XFILLER_21_46 vpwr vgnd scs8hd_fill_2
XFILLER_21_57 vpwr vgnd scs8hd_fill_2
XANTENNA__073__A enable vgnd vpwr scs8hd_diode_2
XFILLER_15_168 vpwr vgnd scs8hd_fill_2
X_125_ _125_/A _125_/B _125_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_15_179 vpwr vgnd scs8hd_fill_2
XANTENNA__158__A _158_/A vgnd vpwr scs8hd_diode_2
XANTENNA__068__A _067_/X vgnd vpwr scs8hd_diode_2
XFILLER_16_46 vpwr vgnd scs8hd_fill_2
XFILLER_32_67 vpwr vgnd scs8hd_fill_2
XFILLER_32_23 vpwr vgnd scs8hd_fill_2
XFILLER_32_12 vpwr vgnd scs8hd_fill_2
XFILLER_12_105 vgnd vpwr scs8hd_decap_12
XFILLER_16_79 vpwr vgnd scs8hd_fill_2
Xmem_top_track_0.LATCH_2_.latch data_in mem_top_track_0.LATCH_2_.latch/Q _155_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_20_182 vgnd vpwr scs8hd_decap_4
X_108_ _108_/A _106_/B _108_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_11_171 vgnd vpwr scs8hd_decap_12
XANTENNA__160__B _158_/X vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_16.INVTX1_4_.scs8hd_inv_1_A right_bottom_grid_pin_9_ vgnd
+ vpwr scs8hd_diode_2
XFILLER_34_274 vgnd vpwr scs8hd_fill_1
Xmux_top_track_8.tap_buf4_0_.scs8hd_inv_1 mux_top_track_8.tap_buf4_0_.scs8hd_inv_1/A
+ _206_/A vgnd vpwr scs8hd_inv_1
XANTENNA_mem_right_track_8.LATCH_4_.latch_SLEEPB _100_/Y vgnd vpwr scs8hd_diode_2
XFILLER_8_80 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_9.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB mem_left_track_9.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_left_track_1.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xmem_left_track_17.LATCH_5_.latch data_in mem_left_track_17.LATCH_5_.latch/Q _137_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_27_89 vpwr vgnd scs8hd_fill_2
XFILLER_25_252 vgnd vpwr scs8hd_decap_3
XFILLER_40_266 vgnd vpwr scs8hd_decap_8
XFILLER_4_178 vgnd vpwr scs8hd_decap_12
XFILLER_4_27 vgnd vpwr scs8hd_decap_4
XFILLER_16_230 vgnd vpwr scs8hd_decap_12
XPHY_280 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_31_266 vgnd vpwr scs8hd_decap_8
XANTENNA__155__B _157_/B vgnd vpwr scs8hd_diode_2
XANTENNA__171__A _090_/B vgnd vpwr scs8hd_diode_2
XFILLER_22_200 vgnd vpwr scs8hd_decap_4
XFILLER_22_211 vgnd vpwr scs8hd_decap_3
XFILLER_22_222 vpwr vgnd scs8hd_fill_2
XFILLER_38_11 vgnd vpwr scs8hd_decap_4
XANTENNA_mem_right_track_8.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_8_7 vgnd vpwr scs8hd_decap_12
XFILLER_1_159 vgnd vpwr scs8hd_decap_12
XANTENNA__081__A address[1] vgnd vpwr scs8hd_diode_2
XFILLER_9_259 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_left_track_1.LATCH_2_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA__166__A _165_/X vgnd vpwr scs8hd_diode_2
XANTENNA__076__A _111_/A vgnd vpwr scs8hd_diode_2
XFILLER_40_78 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_0.INVTX1_1_.scs8hd_inv_1_A chany_top_in[5] vgnd vpwr scs8hd_diode_2
XFILLER_36_100 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_right_track_8.INVTX1_3_.scs8hd_inv_1_A right_bottom_grid_pin_1_ vgnd
+ vpwr scs8hd_diode_2
X_210_ _210_/A chany_top_out[0] vgnd vpwr scs8hd_buf_2
X_141_ _125_/A _136_/X _141_/Y vgnd vpwr scs8hd_nor2_4
X_072_ address[6] _118_/B vgnd vpwr scs8hd_inv_8
Xmux_right_track_16.INVTX1_7_.scs8hd_inv_1 chanx_left_in[6] mux_right_track_16.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
Xmux_top_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_top_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ _145_/A mux_top_track_8.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XFILLER_2_276 vgnd vpwr scs8hd_fill_1
XFILLER_33_136 vpwr vgnd scs8hd_fill_2
XANTENNA__163__B _109_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_right_track_8.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xmem_left_track_1.LATCH_3_.latch data_in mem_left_track_1.LATCH_3_.latch/Q _123_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mem_right_track_0.LATCH_0_.latch_SLEEPB _093_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_17.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_left_track_17.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_2_93 vgnd vpwr scs8hd_decap_12
XPHY_109 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__073__B _118_/B vgnd vpwr scs8hd_diode_2
XFILLER_21_25 vpwr vgnd scs8hd_fill_2
XFILLER_30_106 vgnd vpwr scs8hd_decap_4
XFILLER_15_114 vpwr vgnd scs8hd_fill_2
XFILLER_15_147 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_17.INVTX1_7_.scs8hd_inv_1_A left_bottom_grid_pin_15_ vgnd
+ vpwr scs8hd_diode_2
X_124_ _124_/A _125_/B _124_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_30_139 vpwr vgnd scs8hd_fill_2
XFILLER_16_6 vgnd vpwr scs8hd_decap_4
Xmem_right_track_16.LATCH_4_.latch data_in mem_right_track_16.LATCH_4_.latch/Q _112_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_29_206 vpwr vgnd scs8hd_fill_2
XFILLER_12_117 vgnd vpwr scs8hd_decap_12
XANTENNA__084__A _076_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_9.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A mux_left_track_9.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_left_track_17.LATCH_5_.latch_SLEEPB _137_/Y vgnd vpwr scs8hd_diode_2
XFILLER_7_110 vgnd vpwr scs8hd_decap_12
X_107_ _172_/A _108_/A vgnd vpwr scs8hd_buf_1
XANTENNA__160__C _162_/C vgnd vpwr scs8hd_diode_2
XANTENNA__169__A _084_/B vgnd vpwr scs8hd_diode_2
XANTENNA__079__A _078_/X vgnd vpwr scs8hd_diode_2
XFILLER_27_57 vpwr vgnd scs8hd_fill_2
XFILLER_16_242 vgnd vpwr scs8hd_decap_12
XPHY_281 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_270 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_top_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _146_/A vgnd vpwr
+ scs8hd_diode_2
XFILLER_31_245 vgnd vpwr scs8hd_decap_8
XFILLER_31_223 vpwr vgnd scs8hd_fill_2
XFILLER_31_212 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_left_track_9.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB mem_left_track_9.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__171__B _167_/B vgnd vpwr scs8hd_diode_2
Xmux_left_track_9.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 mux_left_track_9.INVTX1_3_.scs8hd_inv_1/Y
+ mem_left_track_9.LATCH_0_.latch/Q mux_left_track_9.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_left_track_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB mem_left_track_1.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_16.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_13_26 vpwr vgnd scs8hd_fill_2
Xmux_right_track_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_right_track_0.INVTX1_1_.scs8hd_inv_1/Y
+ mem_right_track_0.LATCH_1_.latch/Q mux_right_track_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_right_track_8.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_right_track_8.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_13_245 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_top_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_top_track_0.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_16.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A mux_right_track_16.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_10_215 vgnd vpwr scs8hd_decap_12
XANTENNA__076__B _076_/B vgnd vpwr scs8hd_diode_2
XFILLER_24_69 vgnd vpwr scs8hd_decap_4
XANTENNA__092__A _091_/X vgnd vpwr scs8hd_diode_2
XFILLER_36_145 vpwr vgnd scs8hd_fill_2
XFILLER_27_101 vpwr vgnd scs8hd_fill_2
XFILLER_35_57 vpwr vgnd scs8hd_fill_2
XFILLER_35_35 vpwr vgnd scs8hd_fill_2
XANTENNA__087__A _076_/B vgnd vpwr scs8hd_diode_2
X_140_ _124_/A _136_/X _140_/Y vgnd vpwr scs8hd_nor2_4
X_071_ address[4] _109_/B _074_/A vgnd vpwr scs8hd_or2_4
Xmux_top_track_16.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_top_track_16.INVTX1_3_.scs8hd_inv_1/Y
+ mem_top_track_16.LATCH_4_.latch/Q mux_top_track_16.tap_buf4_0_.scs8hd_inv_1/A vgnd
+ vpwr scs8hd_ebufn_2
XFILLER_18_145 vgnd vpwr scs8hd_decap_8
XPHY_90 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_25_90 vgnd vpwr scs8hd_decap_4
XANTENNA__163__C _158_/X vgnd vpwr scs8hd_diode_2
XFILLER_24_126 vpwr vgnd scs8hd_fill_2
XFILLER_32_192 vpwr vgnd scs8hd_fill_2
XANTENNA__073__C address[5] vgnd vpwr scs8hd_diode_2
Xmux_left_track_17.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_left_track_17.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2/Z
+ mem_left_track_17.LATCH_4_.latch/Q mux_left_track_17.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
Xmux_top_track_16.INVTX1_3_.scs8hd_inv_1 chanx_left_in[7] mux_top_track_16.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_15_126 vpwr vgnd scs8hd_fill_2
X_123_ _113_/A _125_/B _123_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_38_207 vgnd vpwr scs8hd_decap_6
XFILLER_14_181 vgnd vpwr scs8hd_decap_3
XFILLER_21_118 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_17.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB mem_left_track_17.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__190__A chanx_right_in[1] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_0.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_12_129 vgnd vpwr scs8hd_decap_3
Xmem_right_track_0.LATCH_3_.latch data_in mem_right_track_0.LATCH_3_.latch/Q _084_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_32_36 vgnd vpwr scs8hd_fill_1
XANTENNA__084__B _084_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mem_left_track_9.LATCH_0_.latch_SLEEPB _134_/Y vgnd vpwr scs8hd_diode_2
X_106_ _125_/A _106_/B _106_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_11_184 vgnd vpwr scs8hd_decap_12
XFILLER_22_91 vgnd vpwr scs8hd_fill_1
XANTENNA__169__B _167_/B vgnd vpwr scs8hd_diode_2
XFILLER_34_276 vgnd vpwr scs8hd_fill_1
XANTENNA__185__A chanx_right_in[6] vgnd vpwr scs8hd_diode_2
XFILLER_19_262 vgnd vpwr scs8hd_decap_12
XFILLER_8_93 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_14.tap_buf4_0_.scs8hd_inv_1_A mux_top_track_14.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_25_221 vgnd vpwr scs8hd_decap_4
XFILLER_25_232 vpwr vgnd scs8hd_fill_2
XFILLER_27_25 vpwr vgnd scs8hd_fill_2
XFILLER_40_202 vgnd vpwr scs8hd_decap_12
XANTENNA__095__A _095_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_0.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A mux_right_track_0.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_track_14.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_17.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A mux_left_track_17.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_16_254 vgnd vpwr scs8hd_fill_1
XFILLER_16_276 vgnd vpwr scs8hd_fill_1
XPHY_282 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_271 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_260 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_13_16 vpwr vgnd scs8hd_fill_2
XFILLER_13_49 vpwr vgnd scs8hd_fill_2
XFILLER_38_46 vgnd vpwr scs8hd_decap_4
Xmux_right_track_8.INVTX1_0_.scs8hd_inv_1 chany_top_in[0] mux_right_track_8.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_39_132 vpwr vgnd scs8hd_fill_2
XFILLER_10_227 vgnd vpwr scs8hd_decap_12
XFILLER_5_253 vpwr vgnd scs8hd_fill_2
XFILLER_5_220 vgnd vpwr scs8hd_decap_12
XFILLER_36_168 vgnd vpwr scs8hd_decap_4
Xmux_left_track_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_left_track_1.INVTX1_2_.scs8hd_inv_1/Y
+ mem_left_track_1.LATCH_2_.latch/Q mux_left_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA__193__A _193_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_17.INVTX1_2_.scs8hd_inv_1_A chany_top_in[7] vgnd vpwr scs8hd_diode_2
XFILLER_19_15 vpwr vgnd scs8hd_fill_2
XFILLER_42_116 vgnd vpwr scs8hd_decap_8
XFILLER_27_179 vpwr vgnd scs8hd_fill_2
XANTENNA__087__B _103_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_9.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_left_track_9.LATCH_5_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xmux_left_track_17.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2 mux_left_track_17.INVTX1_5_.scs8hd_inv_1/Y
+ mem_left_track_17.LATCH_2_.latch/Q mux_left_track_17.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
X_070_ address[3] _109_/B vgnd vpwr scs8hd_inv_8
XFILLER_4_3 vgnd vpwr scs8hd_decap_12
Xmux_left_track_1.INVTX1_2_.scs8hd_inv_1 chany_top_in[6] mux_left_track_1.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_33_116 vgnd vpwr scs8hd_decap_4
XFILLER_33_105 vpwr vgnd scs8hd_fill_2
XFILLER_18_157 vpwr vgnd scs8hd_fill_2
XPHY_80 vgnd vpwr scs8hd_decap_3
XFILLER_33_149 vgnd vpwr scs8hd_decap_4
XPHY_91 vgnd vpwr scs8hd_tapvpwrvgnd_1
X_199_ chanx_left_in[1] chanx_right_out[2] vgnd vpwr scs8hd_buf_2
Xmem_left_track_9.LATCH_4_.latch data_in mem_left_track_9.LATCH_4_.latch/Q _130_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
Xmux_top_track_14.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_top_track_14.INVTX1_0_.scs8hd_inv_1/Y
+ _148_/A mux_top_track_14.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A vgnd vpwr scs8hd_ebufn_2
XANTENNA__163__D _161_/C vgnd vpwr scs8hd_diode_2
XFILLER_37_3 vpwr vgnd scs8hd_fill_2
XANTENNA__188__A _188_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_8.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A mux_right_track_8.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__098__A _111_/A vgnd vpwr scs8hd_diode_2
X_122_ _112_/A _125_/B _122_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA_mem_top_track_16.LATCH_4_.latch_SLEEPB _168_/Y vgnd vpwr scs8hd_diode_2
Xmem_top_track_16.LATCH_5_.latch data_in mem_top_track_16.LATCH_5_.latch/Q _167_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_29_219 vgnd vpwr scs8hd_decap_12
XFILLER_16_27 vpwr vgnd scs8hd_fill_2
XFILLER_20_141 vgnd vpwr scs8hd_decap_6
Xmux_right_track_8.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2 mux_right_track_8.INVTX1_7_.scs8hd_inv_1/Y
+ mem_right_track_8.LATCH_1_.latch/Q mux_right_track_8.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_28_274 vgnd vpwr scs8hd_fill_1
XFILLER_28_230 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_17.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB mem_left_track_17.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_7_123 vgnd vpwr scs8hd_decap_12
XFILLER_11_196 vgnd vpwr scs8hd_decap_12
X_105_ _090_/B _125_/A vgnd vpwr scs8hd_buf_1
XFILLER_22_70 vpwr vgnd scs8hd_fill_2
XFILLER_22_81 vpwr vgnd scs8hd_fill_2
XFILLER_19_274 vgnd vpwr scs8hd_decap_3
XFILLER_34_222 vgnd vpwr scs8hd_decap_12
XANTENNA__095__B address[3] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_top_track_16.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XPHY_261 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_250 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_31_258 vpwr vgnd scs8hd_fill_2
XPHY_283 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_272 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmux_left_track_9.INVTX1_7_.scs8hd_inv_1 left_bottom_grid_pin_13_ mux_left_track_9.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA__196__A chanx_left_in[4] vgnd vpwr scs8hd_diode_2
XANTENNA_mem_left_track_17.LATCH_3_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_16.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_right_track_16.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_13_258 vpwr vgnd scs8hd_fill_2
XFILLER_28_80 vpwr vgnd scs8hd_fill_2
XFILLER_0_195 vgnd vpwr scs8hd_decap_12
Xmux_right_track_0.INVTX1_3_.scs8hd_inv_1 right_top_grid_pin_10_ mux_right_track_0.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_8_251 vgnd vpwr scs8hd_decap_12
XFILLER_5_62 vgnd vpwr scs8hd_decap_12
XFILLER_5_51 vgnd vpwr scs8hd_decap_8
XFILLER_39_111 vpwr vgnd scs8hd_fill_2
XFILLER_39_188 vpwr vgnd scs8hd_fill_2
XFILLER_24_27 vpwr vgnd scs8hd_fill_2
XFILLER_24_49 vpwr vgnd scs8hd_fill_2
XFILLER_10_239 vgnd vpwr scs8hd_decap_12
Xmux_left_track_1.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2 mux_left_track_1.INVTX1_6_.scs8hd_inv_1/Y
+ mem_left_track_1.LATCH_0_.latch/Q mux_left_track_1.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
Xmux_right_track_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_right_track_0.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2/Z
+ mem_right_track_0.LATCH_5_.latch/Q mux_right_track_0.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_right_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_right_track_8.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_5_232 vgnd vpwr scs8hd_decap_12
XFILLER_14_93 vgnd vpwr scs8hd_decap_6
XFILLER_39_7 vpwr vgnd scs8hd_fill_2
XFILLER_36_125 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_top_track_14.INVTX1_1_.scs8hd_inv_1_A chanx_left_in[8] vgnd vpwr scs8hd_diode_2
XFILLER_27_114 vpwr vgnd scs8hd_fill_2
XFILLER_42_128 vgnd vpwr scs8hd_decap_12
XFILLER_42_106 vgnd vpwr scs8hd_decap_6
XFILLER_2_202 vgnd vpwr scs8hd_decap_12
XFILLER_18_103 vpwr vgnd scs8hd_fill_2
XPHY_81 vgnd vpwr scs8hd_decap_3
XPHY_70 vgnd vpwr scs8hd_decap_3
XPHY_92 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmux_right_track_16.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2 mux_right_track_16.INVTX1_7_.scs8hd_inv_1/Y
+ mem_right_track_16.LATCH_1_.latch/Q mux_right_track_16.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
X_198_ chanx_left_in[2] chanx_right_out[3] vgnd vpwr scs8hd_buf_2
XANTENNA_mux_left_track_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_left_track_1.LATCH_4_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__098__B _106_/B vgnd vpwr scs8hd_diode_2
X_121_ _111_/A _125_/B _121_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_7_19 vgnd vpwr scs8hd_decap_12
XFILLER_11_72 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_1.INVTX1_6_.scs8hd_inv_1_A left_bottom_grid_pin_5_ vgnd vpwr
+ scs8hd_diode_2
XFILLER_14_161 vgnd vpwr scs8hd_decap_6
XANTENNA_mux_left_track_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_left_track_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XANTENNA__199__A chanx_left_in[1] vgnd vpwr scs8hd_diode_2
XFILLER_37_242 vpwr vgnd scs8hd_fill_2
XFILLER_37_231 vgnd vpwr scs8hd_fill_1
Xmem_right_track_8.LATCH_4_.latch data_in mem_right_track_8.LATCH_4_.latch/Q _100_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_32_27 vpwr vgnd scs8hd_fill_2
XFILLER_20_186 vgnd vpwr scs8hd_fill_1
XANTENNA_mem_right_track_8.LATCH_3_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_track_8.LATCH_1_.latch_SLEEPB _106_/Y vgnd vpwr scs8hd_diode_2
XFILLER_28_242 vgnd vpwr scs8hd_decap_12
X_104_ _124_/A _106_/B _104_/Y vgnd vpwr scs8hd_nor2_4
Xmem_top_track_2.LATCH_0_.latch data_in _144_/A _160_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
Xmem_left_track_17.LATCH_0_.latch data_in mem_left_track_17.LATCH_0_.latch/Q _142_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_7_135 vgnd vpwr scs8hd_decap_12
XFILLER_11_120 vpwr vgnd scs8hd_fill_2
XFILLER_22_93 vgnd vpwr scs8hd_decap_4
XFILLER_34_234 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_left_track_1.LATCH_5_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_14_6 vpwr vgnd scs8hd_fill_2
XFILLER_19_242 vpwr vgnd scs8hd_fill_2
XFILLER_19_253 vpwr vgnd scs8hd_fill_2
XFILLER_21_7 vgnd vpwr scs8hd_decap_3
XFILLER_6_190 vgnd vpwr scs8hd_decap_12
XFILLER_27_38 vpwr vgnd scs8hd_fill_2
XFILLER_4_105 vgnd vpwr scs8hd_decap_12
XFILLER_16_212 vpwr vgnd scs8hd_fill_2
XPHY_284 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_273 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_262 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_251 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_240 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_17_71 vgnd vpwr scs8hd_decap_4
XANTENNA_mem_left_track_1.LATCH_4_.latch_SLEEPB _122_/Y vgnd vpwr scs8hd_diode_2
XFILLER_3_171 vgnd vpwr scs8hd_decap_12
Xmux_left_track_9.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2 _175_/HI mem_left_track_9.LATCH_2_.latch/Q
+ mux_left_track_9.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XFILLER_22_204 vgnd vpwr scs8hd_fill_1
XFILLER_22_259 vgnd vpwr scs8hd_decap_12
XFILLER_9_208 vgnd vpwr scs8hd_decap_12
Xmux_top_track_2.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 mux_top_track_2.INVTX1_2_.scs8hd_inv_1/Y
+ _144_/A mux_top_track_2.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XFILLER_8_263 vgnd vpwr scs8hd_decap_12
XFILLER_5_74 vgnd vpwr scs8hd_decap_12
XFILLER_39_178 vgnd vpwr scs8hd_decap_3
XFILLER_39_156 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_right_track_16.LATCH_4_.latch_SLEEPB _112_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_8.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_8.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_30_71 vpwr vgnd scs8hd_fill_2
XFILLER_36_137 vpwr vgnd scs8hd_fill_2
Xmux_right_track_16.INVTX1_4_.scs8hd_inv_1 right_bottom_grid_pin_9_ mux_right_track_16.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
Xmux_left_track_17.INVTX1_5_.scs8hd_inv_1 left_bottom_grid_pin_3_ mux_left_track_17.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_10_19 vgnd vpwr scs8hd_decap_12
XFILLER_19_28 vgnd vpwr scs8hd_decap_4
XFILLER_27_159 vpwr vgnd scs8hd_fill_2
XFILLER_19_39 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_14.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A _180_/HI vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_right_track_8.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB mem_right_track_8.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_right_track_0.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XPHY_82 vgnd vpwr scs8hd_decap_3
XPHY_71 vgnd vpwr scs8hd_decap_3
XPHY_60 vgnd vpwr scs8hd_decap_3
XFILLER_41_184 vgnd vpwr scs8hd_decap_12
XFILLER_41_151 vpwr vgnd scs8hd_fill_2
XPHY_93 vgnd vpwr scs8hd_tapvpwrvgnd_1
X_197_ _197_/A chanx_right_out[4] vgnd vpwr scs8hd_buf_2
XFILLER_24_107 vpwr vgnd scs8hd_fill_2
Xmux_top_track_16.tap_buf4_0_.scs8hd_inv_1 mux_top_track_16.tap_buf4_0_.scs8hd_inv_1/A
+ _202_/A vgnd vpwr scs8hd_inv_1
XFILLER_21_29 vpwr vgnd scs8hd_fill_2
XFILLER_15_118 vpwr vgnd scs8hd_fill_2
XFILLER_23_140 vpwr vgnd scs8hd_fill_2
X_120_ _119_/X _125_/B vgnd vpwr scs8hd_buf_1
XFILLER_23_151 vpwr vgnd scs8hd_fill_2
XFILLER_23_184 vpwr vgnd scs8hd_fill_2
XFILLER_11_40 vpwr vgnd scs8hd_fill_2
XFILLER_11_51 vpwr vgnd scs8hd_fill_2
XFILLER_11_62 vgnd vpwr scs8hd_decap_8
XFILLER_11_84 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _145_/A vgnd vpwr
+ scs8hd_diode_2
XFILLER_36_70 vgnd vpwr scs8hd_decap_3
Xmux_top_track_14.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 _180_/HI _147_/Y mux_top_track_14.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_42_3 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_left_track_17.LATCH_2_.latch_SLEEPB _140_/Y vgnd vpwr scs8hd_diode_2
XFILLER_37_221 vpwr vgnd scs8hd_fill_2
XFILLER_20_154 vpwr vgnd scs8hd_fill_2
XFILLER_20_165 vgnd vpwr scs8hd_decap_8
XFILLER_28_254 vgnd vpwr scs8hd_decap_12
XFILLER_28_276 vgnd vpwr scs8hd_fill_1
XFILLER_7_147 vgnd vpwr scs8hd_decap_12
X_103_ _103_/A _124_/A vgnd vpwr scs8hd_buf_1
XFILLER_34_246 vgnd vpwr scs8hd_decap_12
XFILLER_34_202 vpwr vgnd scs8hd_fill_2
XFILLER_19_221 vpwr vgnd scs8hd_fill_2
XFILLER_25_257 vgnd vpwr scs8hd_decap_12
XFILLER_4_117 vgnd vpwr scs8hd_decap_12
XPHY_285 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_274 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_263 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_252 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_241 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_33_60 vgnd vpwr scs8hd_fill_1
XFILLER_31_227 vgnd vpwr scs8hd_decap_12
XPHY_230 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_17_94 vpwr vgnd scs8hd_fill_2
XFILLER_38_38 vgnd vpwr scs8hd_fill_1
Xmux_top_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_top_track_8.INVTX1_0_.scs8hd_inv_1/Y
+ _146_/A mux_top_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_left_track_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A mux_left_track_1.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_0_120 vgnd vpwr scs8hd_decap_4
XFILLER_28_93 vpwr vgnd scs8hd_fill_2
XFILLER_12_271 vgnd vpwr scs8hd_decap_4
XFILLER_5_86 vgnd vpwr scs8hd_decap_12
XFILLER_40_17 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_top_track_2.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_track_0.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_14_84 vgnd vpwr scs8hd_decap_8
Xmux_right_track_8.tap_buf4_0_.scs8hd_inv_1 mux_right_track_8.tap_buf4_0_.scs8hd_inv_1/A
+ _197_/A vgnd vpwr scs8hd_inv_1
XFILLER_5_245 vgnd vpwr scs8hd_decap_8
XFILLER_36_149 vpwr vgnd scs8hd_fill_2
XANTENNA__101__A _084_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_0.INVTX1_7_.scs8hd_inv_1_A chanx_left_in[4] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_1.INVTX1_1_.scs8hd_inv_1_A chany_top_in[3] vgnd vpwr scs8hd_diode_2
XFILLER_35_39 vgnd vpwr scs8hd_decap_3
XFILLER_27_138 vpwr vgnd scs8hd_fill_2
XFILLER_2_215 vgnd vpwr scs8hd_decap_12
XPHY_83 vgnd vpwr scs8hd_decap_3
XPHY_72 vgnd vpwr scs8hd_decap_3
XPHY_61 vgnd vpwr scs8hd_decap_3
XPHY_94 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_50 vgnd vpwr scs8hd_decap_3
XFILLER_41_196 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_0.INVTX1_3_.scs8hd_inv_1_A chanx_left_in[0] vgnd vpwr scs8hd_diode_2
X_196_ chanx_left_in[4] chanx_right_out[5] vgnd vpwr scs8hd_buf_2
XFILLER_2_32 vgnd vpwr scs8hd_decap_12
Xmux_top_track_16.INVTX1_0_.scs8hd_inv_1 chanx_right_in[0] mux_top_track_16.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_left_track_9.INVTX1_3_.scs8hd_inv_1_A chanx_right_in[1] vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_track_16.LATCH_2_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_2_3 vgnd vpwr scs8hd_decap_12
XFILLER_11_96 vgnd vpwr scs8hd_decap_12
X_179_ _179_/HI _179_/LO vgnd vpwr scs8hd_conb_1
XFILLER_35_3 vgnd vpwr scs8hd_decap_4
XFILLER_20_122 vpwr vgnd scs8hd_fill_2
XFILLER_28_266 vgnd vpwr scs8hd_decap_8
XFILLER_28_200 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_left_track_9.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_left_track_9.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
X_102_ _113_/A _106_/B _102_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_7_159 vgnd vpwr scs8hd_decap_12
XFILLER_22_62 vpwr vgnd scs8hd_fill_2
XFILLER_34_258 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_right_track_16.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_25_203 vgnd vpwr scs8hd_decap_3
XFILLER_25_236 vgnd vpwr scs8hd_decap_8
XFILLER_25_269 vgnd vpwr scs8hd_decap_8
XFILLER_4_129 vgnd vpwr scs8hd_decap_12
XFILLER_31_217 vgnd vpwr scs8hd_decap_3
XFILLER_17_40 vpwr vgnd scs8hd_fill_2
XPHY_275 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_264 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_253 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_242 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_31_239 vgnd vpwr scs8hd_decap_4
XPHY_231 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_220 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__104__A _124_/A vgnd vpwr scs8hd_diode_2
XFILLER_3_184 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_right_track_0.LATCH_5_.latch_SLEEPB _076_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_9.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_left_track_9.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
Xmux_top_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_top_track_16.INVTX1_1_.scs8hd_inv_1/Y
+ mem_top_track_16.LATCH_1_.latch/Q mux_top_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_28_61 vpwr vgnd scs8hd_fill_2
XFILLER_8_276 vgnd vpwr scs8hd_fill_1
Xmem_top_track_0.LATCH_3_.latch data_in mem_top_track_0.LATCH_3_.latch/Q _154_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_5_98 vgnd vpwr scs8hd_decap_12
XFILLER_39_169 vpwr vgnd scs8hd_fill_2
XFILLER_39_136 vgnd vpwr scs8hd_decap_3
XFILLER_24_19 vpwr vgnd scs8hd_fill_2
XFILLER_40_29 vpwr vgnd scs8hd_fill_2
Xmux_left_track_17.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_left_track_17.INVTX1_1_.scs8hd_inv_1/Y
+ mem_left_track_17.LATCH_1_.latch/Q mux_left_track_17.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_38_191 vpwr vgnd scs8hd_fill_2
XFILLER_38_180 vgnd vpwr scs8hd_decap_8
XFILLER_14_52 vpwr vgnd scs8hd_fill_2
XFILLER_30_84 vpwr vgnd scs8hd_fill_2
XFILLER_5_257 vgnd vpwr scs8hd_decap_12
XFILLER_39_82 vpwr vgnd scs8hd_fill_2
XFILLER_39_71 vpwr vgnd scs8hd_fill_2
XFILLER_36_106 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_left_track_9.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB mem_left_track_9.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_left_track_1.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_35_18 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_2.INVTX1_1_.scs8hd_inv_1_A chanx_right_in[2] vgnd vpwr scs8hd_diode_2
XANTENNA__202__A _202_/A vgnd vpwr scs8hd_diode_2
XFILLER_2_227 vgnd vpwr scs8hd_decap_12
Xmux_top_track_8.INVTX1_1_.scs8hd_inv_1 chanx_left_in[6] mux_top_track_8.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_18_128 vpwr vgnd scs8hd_fill_2
XPHY_84 vgnd vpwr scs8hd_decap_3
XPHY_73 vgnd vpwr scs8hd_decap_3
XPHY_62 vgnd vpwr scs8hd_decap_3
XFILLER_26_172 vgnd vpwr scs8hd_decap_4
XFILLER_26_150 vgnd vpwr scs8hd_decap_3
XPHY_95 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_40 vgnd vpwr scs8hd_decap_3
XFILLER_25_73 vpwr vgnd scs8hd_fill_2
XPHY_51 vgnd vpwr scs8hd_decap_3
X_195_ chanx_left_in[5] chanx_right_out[6] vgnd vpwr scs8hd_buf_2
XANTENNA__112__A _112_/A vgnd vpwr scs8hd_diode_2
XFILLER_2_44 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_16.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_right_track_16.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_track_16.LATCH_1_.latch_SLEEPB _171_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_track_0.LATCH_2_.latch_D data_in vgnd vpwr scs8hd_diode_2
Xmux_right_track_8.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_8.INVTX1_3_.scs8hd_inv_1/Y
+ mem_right_track_8.LATCH_0_.latch/Q mux_right_track_8.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
Xmem_top_track_16.LATCH_0_.latch data_in mem_top_track_16.LATCH_0_.latch/Q _172_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_23_164 vpwr vgnd scs8hd_fill_2
XFILLER_23_175 vpwr vgnd scs8hd_fill_2
XFILLER_23_197 vpwr vgnd scs8hd_fill_2
XANTENNA__107__A _172_/A vgnd vpwr scs8hd_diode_2
XFILLER_14_186 vgnd vpwr scs8hd_decap_12
X_178_ _178_/HI _178_/LO vgnd vpwr scs8hd_conb_1
XFILLER_37_245 vgnd vpwr scs8hd_decap_12
XFILLER_37_234 vgnd vpwr scs8hd_decap_8
XFILLER_28_3 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_right_track_16.INVTX1_5_.scs8hd_inv_1_A right_bottom_grid_pin_15_ vgnd
+ vpwr scs8hd_diode_2
Xmux_top_track_14.INVTX1_0_.scs8hd_inv_1 chanx_left_in[2] mux_top_track_14.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_20_189 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_top_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_top_track_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_28_212 vpwr vgnd scs8hd_fill_2
XFILLER_11_123 vgnd vpwr scs8hd_decap_12
X_101_ _084_/B _113_/A vgnd vpwr scs8hd_buf_1
XFILLER_22_41 vpwr vgnd scs8hd_fill_2
XFILLER_22_85 vgnd vpwr scs8hd_decap_6
XFILLER_19_234 vgnd vpwr scs8hd_decap_8
XFILLER_19_245 vgnd vpwr scs8hd_decap_8
XFILLER_8_32 vgnd vpwr scs8hd_decap_12
XFILLER_25_248 vpwr vgnd scs8hd_fill_2
XFILLER_40_218 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_top_track_0.LATCH_3_.latch_SLEEPB _154_/Y vgnd vpwr scs8hd_diode_2
Xmux_left_track_9.INVTX1_4_.scs8hd_inv_1 chanx_right_in[5] mux_left_track_9.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
Xmem_left_track_1.LATCH_4_.latch data_in mem_left_track_1.LATCH_4_.latch/Q _122_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA__210__A _210_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_right_track_8.LATCH_4_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XPHY_243 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_232 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_221 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_210 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_16_204 vgnd vpwr scs8hd_decap_8
XFILLER_16_259 vgnd vpwr scs8hd_decap_12
XPHY_276 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_265 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_254 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_33_84 vpwr vgnd scs8hd_fill_2
XANTENNA__104__B _106_/B vgnd vpwr scs8hd_diode_2
XFILLER_3_196 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_16.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB mem_right_track_16.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__120__A _119_/X vgnd vpwr scs8hd_diode_2
Xmux_left_track_9.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_left_track_9.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ mem_left_track_9.LATCH_3_.latch/Q mux_left_track_9.tap_buf4_0_.scs8hd_inv_1/A vgnd
+ vpwr scs8hd_ebufn_2
XFILLER_22_207 vpwr vgnd scs8hd_fill_2
XFILLER_22_218 vpwr vgnd scs8hd_fill_2
XFILLER_22_229 vgnd vpwr scs8hd_decap_8
XFILLER_38_18 vgnd vpwr scs8hd_decap_12
Xmem_right_track_16.LATCH_5_.latch data_in mem_right_track_16.LATCH_5_.latch/Q _111_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
Xmux_right_track_0.INVTX1_0_.scs8hd_inv_1 chany_top_in[2] mux_right_track_0.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_right_track_0.INVTX1_2_.scs8hd_inv_1_A chany_top_in[8] vgnd vpwr scs8hd_diode_2
XANTENNA__205__A chanx_left_in[5] vgnd vpwr scs8hd_diode_2
XFILLER_28_84 vgnd vpwr scs8hd_decap_8
XFILLER_12_251 vgnd vpwr scs8hd_decap_4
XANTENNA__115__A _125_/A vgnd vpwr scs8hd_diode_2
XFILLER_39_115 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_right_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_right_track_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_8.INVTX1_4_.scs8hd_inv_1_A right_bottom_grid_pin_7_ vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mem_left_track_9.LATCH_5_.latch_SLEEPB _129_/Y vgnd vpwr scs8hd_diode_2
Xmux_top_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 _183_/HI _145_/Y mux_top_track_8.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_30_63 vpwr vgnd scs8hd_fill_2
XFILLER_30_52 vpwr vgnd scs8hd_fill_2
XFILLER_5_269 vgnd vpwr scs8hd_decap_8
Xmux_right_track_16.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_16.INVTX1_3_.scs8hd_inv_1/Y
+ mem_right_track_16.LATCH_0_.latch/Q mux_right_track_16.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
Xmux_top_track_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 mux_top_track_0.INVTX1_3_.scs8hd_inv_1/Y
+ mem_top_track_0.LATCH_0_.latch/Q mux_top_track_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_top_track_8.INVTX1_0_.scs8hd_inv_1_A chanx_right_in[6] vgnd vpwr scs8hd_diode_2
XFILLER_27_118 vpwr vgnd scs8hd_fill_2
XFILLER_35_195 vgnd vpwr scs8hd_decap_6
XFILLER_35_162 vpwr vgnd scs8hd_fill_2
XFILLER_35_140 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_top_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _146_/Y vgnd vpwr
+ scs8hd_diode_2
XFILLER_2_239 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_9.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB mem_left_track_9.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB mem_left_track_1.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xmux_top_track_0.INVTX1_4_.scs8hd_inv_1 chanx_left_in[3] mux_top_track_0.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XPHY_30 vgnd vpwr scs8hd_decap_3
XFILLER_18_107 vgnd vpwr scs8hd_decap_4
XPHY_85 vgnd vpwr scs8hd_decap_3
XFILLER_41_132 vpwr vgnd scs8hd_fill_2
XFILLER_41_110 vgnd vpwr scs8hd_fill_1
XPHY_74 vgnd vpwr scs8hd_decap_3
XPHY_63 vgnd vpwr scs8hd_decap_3
XPHY_96 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_41 vgnd vpwr scs8hd_decap_3
XFILLER_25_96 vpwr vgnd scs8hd_fill_2
XPHY_52 vgnd vpwr scs8hd_decap_3
XFILLER_41_62 vgnd vpwr scs8hd_decap_12
X_194_ chanx_left_in[6] chanx_right_out[7] vgnd vpwr scs8hd_buf_2
XANTENNA__112__B _110_/X vgnd vpwr scs8hd_diode_2
XFILLER_2_56 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_9.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A mux_left_track_9.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_32_165 vpwr vgnd scs8hd_fill_2
XFILLER_32_110 vgnd vpwr scs8hd_decap_4
XFILLER_17_184 vpwr vgnd scs8hd_fill_2
XFILLER_11_10 vpwr vgnd scs8hd_fill_2
Xmux_right_track_8.INVTX1_5_.scs8hd_inv_1 right_bottom_grid_pin_13_ mux_right_track_8.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_36_84 vgnd vpwr scs8hd_decap_8
XFILLER_36_62 vgnd vpwr scs8hd_decap_8
X_177_ _177_/HI _177_/LO vgnd vpwr scs8hd_conb_1
XFILLER_14_198 vgnd vpwr scs8hd_decap_12
XANTENNA__123__A _113_/A vgnd vpwr scs8hd_diode_2
XFILLER_37_257 vgnd vpwr scs8hd_decap_12
X_100_ _112_/A _106_/B _100_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_11_135 vgnd vpwr scs8hd_decap_12
XANTENNA__208__A chanx_right_in[4] vgnd vpwr scs8hd_diode_2
XFILLER_22_97 vgnd vpwr scs8hd_fill_1
XFILLER_19_202 vpwr vgnd scs8hd_fill_2
XANTENNA__118__A _118_/A vgnd vpwr scs8hd_diode_2
XFILLER_10_190 vgnd vpwr scs8hd_decap_12
XFILLER_8_44 vgnd vpwr scs8hd_decap_12
Xmux_left_track_9.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 mux_left_track_9.INVTX1_4_.scs8hd_inv_1/Y
+ mem_left_track_9.LATCH_1_.latch/Q mux_left_track_9.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mem_left_track_1.LATCH_1_.latch_SLEEPB _125_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_14.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _148_/A vgnd vpwr
+ scs8hd_diode_2
Xmux_left_track_1.INVTX1_7_.scs8hd_inv_1 left_bottom_grid_pin_11_ mux_left_track_1.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
Xmux_right_track_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_right_track_0.INVTX1_2_.scs8hd_inv_1/Y
+ mem_right_track_0.LATCH_2_.latch/Q mux_right_track_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XPHY_277 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_266 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_255 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_244 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_33_52 vpwr vgnd scs8hd_fill_2
XPHY_233 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_222 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_17_53 vpwr vgnd scs8hd_fill_2
XPHY_200 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_271 vgnd vpwr scs8hd_decap_4
XPHY_211 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_right_track_16.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A mux_right_track_16.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_12_7 vgnd vpwr scs8hd_decap_6
XFILLER_30_274 vgnd vpwr scs8hd_fill_1
XFILLER_30_230 vgnd vpwr scs8hd_decap_12
XFILLER_13_208 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_right_track_0.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_track_16.LATCH_1_.latch_SLEEPB _115_/Y vgnd vpwr scs8hd_diode_2
XFILLER_0_112 vgnd vpwr scs8hd_fill_1
XFILLER_0_145 vpwr vgnd scs8hd_fill_2
XFILLER_0_156 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_left_track_9.LATCH_2_.latch_D data_in vgnd vpwr scs8hd_diode_2
Xmem_right_track_0.LATCH_4_.latch data_in mem_right_track_0.LATCH_4_.latch/Q _080_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA__115__B _110_/X vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A mux_top_track_0.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__131__A _113_/A vgnd vpwr scs8hd_diode_2
Xmux_right_track_16.INVTX1_1_.scs8hd_inv_1 chany_top_in[4] mux_right_track_16.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
Xmux_left_track_17.INVTX1_2_.scs8hd_inv_1 chany_top_in[7] mux_left_track_17.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_14_10 vpwr vgnd scs8hd_fill_2
XFILLER_14_32 vpwr vgnd scs8hd_fill_2
Xmux_top_track_16.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2 _181_/HI mem_top_track_16.LATCH_5_.latch/Q
+ mux_top_track_16.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XFILLER_39_62 vpwr vgnd scs8hd_fill_2
XANTENNA__126__A _108_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_16.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_top_track_16.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_16.INVTX1_0_.scs8hd_inv_1_A chany_top_in[1] vgnd vpwr scs8hd_diode_2
XPHY_64 vgnd vpwr scs8hd_decap_3
XPHY_53 vgnd vpwr scs8hd_decap_3
XFILLER_26_185 vpwr vgnd scs8hd_fill_2
Xmux_left_track_17.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_left_track_17.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2/Z
+ mem_left_track_17.LATCH_5_.latch/Q mux_left_track_17.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XPHY_20 vgnd vpwr scs8hd_decap_3
XPHY_31 vgnd vpwr scs8hd_decap_3
XPHY_42 vgnd vpwr scs8hd_decap_3
XFILLER_25_20 vpwr vgnd scs8hd_fill_2
XFILLER_25_53 vpwr vgnd scs8hd_fill_2
XFILLER_41_155 vgnd vpwr scs8hd_decap_12
XFILLER_41_74 vgnd vpwr scs8hd_decap_12
X_193_ _193_/A chanx_right_out[8] vgnd vpwr scs8hd_buf_2
XPHY_75 vgnd vpwr scs8hd_decap_3
XPHY_86 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_97 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_2_68 vgnd vpwr scs8hd_decap_12
XFILLER_32_188 vpwr vgnd scs8hd_fill_2
XFILLER_32_177 vpwr vgnd scs8hd_fill_2
XFILLER_17_141 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_1.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB mem_left_track_1.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_top_track_0.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_11_55 vgnd vpwr scs8hd_decap_6
XFILLER_36_96 vpwr vgnd scs8hd_fill_2
XFILLER_14_177 vpwr vgnd scs8hd_fill_2
X_176_ _176_/HI _176_/LO vgnd vpwr scs8hd_conb_1
XANTENNA__123__B _125_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A mux_right_track_0.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_37_269 vgnd vpwr scs8hd_decap_8
XFILLER_37_225 vgnd vpwr scs8hd_decap_6
XFILLER_20_103 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_17.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_left_track_17.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_11_147 vgnd vpwr scs8hd_decap_12
XFILLER_0_3 vgnd vpwr scs8hd_decap_12
XFILLER_34_206 vgnd vpwr scs8hd_decap_8
XFILLER_19_258 vpwr vgnd scs8hd_fill_2
XFILLER_42_261 vgnd vpwr scs8hd_decap_12
XANTENNA__118__B _118_/B vgnd vpwr scs8hd_diode_2
XFILLER_8_56 vgnd vpwr scs8hd_decap_12
X_159_ _074_/A _158_/X _161_/C _159_/Y vgnd vpwr scs8hd_nor3_4
XANTENNA__134__A _108_/A vgnd vpwr scs8hd_diode_2
Xmux_right_track_0.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_0.INVTX1_6_.scs8hd_inv_1/Y
+ mem_right_track_0.LATCH_0_.latch/Q mux_right_track_0.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_25_217 vpwr vgnd scs8hd_fill_2
XFILLER_25_228 vpwr vgnd scs8hd_fill_2
Xmem_left_track_9.LATCH_5_.latch data_in mem_left_track_9.LATCH_5_.latch/Q _129_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_left_track_17.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A _174_/HI vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mem_top_track_0.LATCH_4_.latch_D data_in vgnd vpwr scs8hd_diode_2
XPHY_278 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_267 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_256 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_245 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_33_31 vpwr vgnd scs8hd_fill_2
XPHY_234 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_223 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_212 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_17_98 vgnd vpwr scs8hd_decap_4
XPHY_201 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_3_110 vgnd vpwr scs8hd_decap_12
XANTENNA__129__A _111_/A vgnd vpwr scs8hd_diode_2
XFILLER_30_242 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_top_track_2.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_21_231 vgnd vpwr scs8hd_decap_6
XFILLER_21_253 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_top_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_0_168 vgnd vpwr scs8hd_decap_12
XFILLER_28_97 vpwr vgnd scs8hd_fill_2
XFILLER_8_202 vgnd vpwr scs8hd_decap_12
XANTENNA__131__B _132_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_17.INVTX1_3_.scs8hd_inv_1_A chanx_right_in[2] vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_track_16.LATCH_5_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_17.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_TEB mem_left_track_17.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_14_99 vgnd vpwr scs8hd_fill_1
XFILLER_30_32 vgnd vpwr scs8hd_decap_3
XFILLER_30_21 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_8.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_right_track_8.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xmux_top_track_14.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_top_track_14.INVTX1_1_.scs8hd_inv_1/Y
+ _148_/Y mux_top_track_14.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A vgnd vpwr scs8hd_ebufn_2
XANTENNA__126__B _125_/B vgnd vpwr scs8hd_diode_2
XANTENNA__142__A _108_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_track_16.LATCH_2_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_35_175 vpwr vgnd scs8hd_fill_2
XFILLER_41_123 vpwr vgnd scs8hd_fill_2
XPHY_76 vgnd vpwr scs8hd_decap_3
XPHY_65 vgnd vpwr scs8hd_decap_3
XFILLER_26_164 vpwr vgnd scs8hd_fill_2
XPHY_21 vgnd vpwr scs8hd_decap_3
XPHY_10 vgnd vpwr scs8hd_decap_3
XPHY_98 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_87 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_32 vgnd vpwr scs8hd_decap_3
XPHY_43 vgnd vpwr scs8hd_decap_3
XFILLER_25_32 vpwr vgnd scs8hd_fill_2
XPHY_54 vgnd vpwr scs8hd_decap_3
XFILLER_41_167 vgnd vpwr scs8hd_decap_12
XFILLER_41_86 vgnd vpwr scs8hd_decap_12
X_192_ _192_/A chanx_left_out[0] vgnd vpwr scs8hd_buf_2
XFILLER_17_164 vpwr vgnd scs8hd_fill_2
XFILLER_32_145 vpwr vgnd scs8hd_fill_2
XFILLER_17_175 vpwr vgnd scs8hd_fill_2
XFILLER_17_197 vpwr vgnd scs8hd_fill_2
XANTENNA__137__A _111_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_16.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_right_track_16.LATCH_4_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_23_123 vpwr vgnd scs8hd_fill_2
Xmux_right_track_8.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2 _178_/HI mem_right_track_8.LATCH_2_.latch/Q
+ mux_right_track_8.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_right_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_8.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_14_134 vpwr vgnd scs8hd_fill_2
XFILLER_14_145 vgnd vpwr scs8hd_decap_8
XFILLER_14_167 vgnd vpwr scs8hd_fill_1
X_175_ _175_/HI _175_/LO vgnd vpwr scs8hd_conb_1
XFILLER_9_171 vgnd vpwr scs8hd_decap_12
XFILLER_20_137 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_8.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_right_track_8.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_11_159 vgnd vpwr scs8hd_decap_12
XFILLER_22_66 vpwr vgnd scs8hd_fill_2
XFILLER_34_218 vpwr vgnd scs8hd_fill_2
XFILLER_42_273 vgnd vpwr scs8hd_decap_4
XFILLER_8_68 vgnd vpwr scs8hd_decap_12
X_158_ _158_/A _158_/X vgnd vpwr scs8hd_buf_1
XFILLER_6_141 vgnd vpwr scs8hd_decap_12
X_089_ _088_/X _090_/B vgnd vpwr scs8hd_buf_1
XANTENNA__134__B _132_/B vgnd vpwr scs8hd_diode_2
XANTENNA__150__A address[4] vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_track_0.LATCH_2_.latch_SLEEPB _087_/Y vgnd vpwr scs8hd_diode_2
XFILLER_16_218 vgnd vpwr scs8hd_decap_12
XFILLER_17_77 vgnd vpwr scs8hd_decap_4
XPHY_279 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_268 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_257 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_246 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_33_65 vpwr vgnd scs8hd_fill_2
XPHY_235 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_224 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_213 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_202 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_left_track_1.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_left_track_1.LATCH_5_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__129__B _132_/B vgnd vpwr scs8hd_diode_2
XANTENNA__145__A _145_/A vgnd vpwr scs8hd_diode_2
XFILLER_30_276 vgnd vpwr scs8hd_fill_1
XFILLER_30_254 vgnd vpwr scs8hd_decap_12
XFILLER_21_210 vgnd vpwr scs8hd_decap_4
XFILLER_21_243 vgnd vpwr scs8hd_fill_1
Xmux_left_track_1.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2 mux_left_track_1.INVTX1_7_.scs8hd_inv_1/Y
+ mem_left_track_1.LATCH_1_.latch/Q mux_left_track_1.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
Xmem_right_track_8.LATCH_5_.latch data_in mem_right_track_8.LATCH_5_.latch/Q _098_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_28_65 vpwr vgnd scs8hd_fill_2
XFILLER_28_32 vgnd vpwr scs8hd_decap_3
XFILLER_28_21 vgnd vpwr scs8hd_decap_4
XFILLER_0_125 vgnd vpwr scs8hd_decap_12
Xmux_top_track_2.INVTX1_1_.scs8hd_inv_1 chanx_right_in[2] mux_top_track_2.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
Xmux_top_track_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_top_track_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ _143_/A mux_top_track_2.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XFILLER_12_276 vgnd vpwr scs8hd_fill_1
Xmem_top_track_2.LATCH_1_.latch data_in _143_/A _159_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
Xmem_left_track_17.LATCH_1_.latch data_in mem_left_track_17.LATCH_1_.latch/Q _141_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mem_right_track_0.LATCH_5_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_38_195 vgnd vpwr scs8hd_decap_12
XFILLER_14_23 vpwr vgnd scs8hd_fill_2
XFILLER_14_56 vgnd vpwr scs8hd_decap_4
XFILLER_30_88 vgnd vpwr scs8hd_decap_4
XFILLER_39_86 vgnd vpwr scs8hd_decap_12
XFILLER_39_75 vgnd vpwr scs8hd_decap_4
XFILLER_39_53 vpwr vgnd scs8hd_fill_2
XFILLER_29_184 vgnd vpwr scs8hd_decap_4
XFILLER_29_162 vpwr vgnd scs8hd_fill_2
XFILLER_29_140 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_top_track_0.tap_buf4_0_.scs8hd_inv_1_A mux_top_track_0.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
Xmux_right_track_16.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2 _177_/HI mem_right_track_16.LATCH_2_.latch/Q
+ mux_right_track_16.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XANTENNA__142__B _136_/X vgnd vpwr scs8hd_diode_2
XFILLER_35_132 vpwr vgnd scs8hd_fill_2
XFILLER_41_179 vgnd vpwr scs8hd_decap_4
XPHY_77 vgnd vpwr scs8hd_decap_3
XPHY_66 vgnd vpwr scs8hd_decap_3
XPHY_55 vgnd vpwr scs8hd_decap_3
XFILLER_26_154 vgnd vpwr scs8hd_fill_1
XFILLER_26_132 vgnd vpwr scs8hd_decap_4
XPHY_11 vgnd vpwr scs8hd_decap_3
XPHY_99 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_88 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_22 vgnd vpwr scs8hd_decap_3
XPHY_33 vgnd vpwr scs8hd_decap_3
XPHY_44 vgnd vpwr scs8hd_decap_3
XFILLER_25_77 vpwr vgnd scs8hd_fill_2
XFILLER_41_98 vgnd vpwr scs8hd_decap_12
XFILLER_41_10 vgnd vpwr scs8hd_decap_12
X_191_ chanx_right_in[0] chanx_left_out[1] vgnd vpwr scs8hd_buf_2
XANTENNA_mux_left_track_1.INVTX1_7_.scs8hd_inv_1_A left_bottom_grid_pin_11_ vgnd vpwr
+ scs8hd_diode_2
XFILLER_1_220 vgnd vpwr scs8hd_decap_12
XFILLER_2_15 vgnd vpwr scs8hd_decap_12
XFILLER_32_102 vgnd vpwr scs8hd_decap_6
XFILLER_40_190 vgnd vpwr scs8hd_decap_12
XFILLER_32_135 vgnd vpwr scs8hd_fill_1
XANTENNA__137__B _136_/X vgnd vpwr scs8hd_diode_2
XANTENNA__153__A _112_/A vgnd vpwr scs8hd_diode_2
XFILLER_23_102 vgnd vpwr scs8hd_decap_3
XFILLER_23_168 vpwr vgnd scs8hd_fill_2
XFILLER_23_179 vpwr vgnd scs8hd_fill_2
XFILLER_36_32 vgnd vpwr scs8hd_decap_4
XFILLER_14_157 vpwr vgnd scs8hd_fill_2
X_174_ _174_/HI _174_/LO vgnd vpwr scs8hd_conb_1
XFILLER_37_205 vgnd vpwr scs8hd_fill_1
XANTENNA__148__A _148_/A vgnd vpwr scs8hd_diode_2
XFILLER_20_149 vpwr vgnd scs8hd_fill_2
XFILLER_36_260 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_top_track_2.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_22_23 vgnd vpwr scs8hd_decap_3
XFILLER_22_45 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_top_track_0.LATCH_0_.latch_SLEEPB _157_/Y vgnd vpwr scs8hd_diode_2
XFILLER_42_230 vgnd vpwr scs8hd_decap_12
X_157_ _108_/A _157_/B _157_/Y vgnd vpwr scs8hd_nor2_4
Xmux_left_track_9.INVTX1_1_.scs8hd_inv_1 chany_top_in[5] mux_left_track_9.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_40_6 vgnd vpwr scs8hd_decap_8
X_088_ address[1] address[2] _161_/C _088_/X vgnd vpwr scs8hd_or3_4
XANTENNA__150__B address[3] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_8.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB mem_right_track_8.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_33_230 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_right_track_0.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_left_track_1.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XPHY_225 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_214 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_17_23 vpwr vgnd scs8hd_fill_2
XPHY_203 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_269 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_258 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_247 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_33_88 vpwr vgnd scs8hd_fill_2
Xmem_right_track_16.LATCH_0_.latch data_in mem_right_track_16.LATCH_0_.latch/Q _116_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_33_11 vpwr vgnd scs8hd_fill_2
XPHY_236 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmux_top_track_2.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 _182_/HI _144_/Y mux_top_track_2.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_3_123 vgnd vpwr scs8hd_decap_12
XFILLER_15_241 vgnd vpwr scs8hd_decap_3
XFILLER_15_263 vgnd vpwr scs8hd_decap_12
XFILLER_30_266 vgnd vpwr scs8hd_decap_8
XANTENNA__161__A _096_/B vgnd vpwr scs8hd_diode_2
X_209_ _209_/A chany_top_out[1] vgnd vpwr scs8hd_buf_2
XANTENNA_mux_right_track_0.tap_buf4_0_.scs8hd_inv_1_A mux_right_track_0.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_8.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_8.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_0_70 vgnd vpwr scs8hd_decap_4
XFILLER_0_81 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _145_/Y vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_top_track_16.INVTX1_0_.scs8hd_inv_1_A chanx_right_in[0] vgnd vpwr scs8hd_diode_2
XANTENNA__071__A address[4] vgnd vpwr scs8hd_diode_2
XFILLER_28_44 vpwr vgnd scs8hd_fill_2
XFILLER_0_137 vgnd vpwr scs8hd_decap_4
XFILLER_8_215 vgnd vpwr scs8hd_decap_12
XFILLER_5_15 vgnd vpwr scs8hd_decap_12
XFILLER_39_119 vgnd vpwr scs8hd_fill_1
XFILLER_5_59 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_left_track_9.LATCH_2_.latch_SLEEPB _132_/Y vgnd vpwr scs8hd_diode_2
XFILLER_10_7 vgnd vpwr scs8hd_decap_12
XANTENNA__156__A _125_/A vgnd vpwr scs8hd_diode_2
XFILLER_38_163 vpwr vgnd scs8hd_fill_2
XANTENNA__066__A address[0] vgnd vpwr scs8hd_diode_2
XFILLER_30_67 vpwr vgnd scs8hd_fill_2
XFILLER_39_98 vpwr vgnd scs8hd_fill_2
XFILLER_4_251 vgnd vpwr scs8hd_decap_12
Xmux_top_track_0.INVTX1_1_.scs8hd_inv_1 chanx_right_in[1] mux_top_track_0.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_35_144 vgnd vpwr scs8hd_fill_1
XFILLER_35_111 vpwr vgnd scs8hd_fill_2
XFILLER_6_80 vgnd vpwr scs8hd_decap_12
XPHY_12 vgnd vpwr scs8hd_decap_3
XFILLER_41_136 vgnd vpwr scs8hd_decap_12
XFILLER_41_114 vpwr vgnd scs8hd_fill_2
XFILLER_41_22 vgnd vpwr scs8hd_decap_12
XPHY_78 vgnd vpwr scs8hd_decap_3
XPHY_67 vgnd vpwr scs8hd_decap_3
XPHY_56 vgnd vpwr scs8hd_decap_3
XPHY_89 vgnd vpwr scs8hd_tapvpwrvgnd_1
X_190_ chanx_right_in[1] chanx_left_out[2] vgnd vpwr scs8hd_buf_2
XPHY_23 vgnd vpwr scs8hd_decap_3
XPHY_34 vgnd vpwr scs8hd_decap_3
XPHY_45 vgnd vpwr scs8hd_decap_3
XFILLER_2_27 vgnd vpwr scs8hd_decap_4
XFILLER_1_232 vgnd vpwr scs8hd_decap_12
XFILLER_32_125 vpwr vgnd scs8hd_fill_2
XFILLER_32_169 vgnd vpwr scs8hd_decap_8
XANTENNA__153__B _157_/B vgnd vpwr scs8hd_diode_2
Xmux_right_track_8.INVTX1_2_.scs8hd_inv_1 chany_top_in[6] mux_right_track_8.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_top_track_14.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _147_/A vgnd vpwr
+ scs8hd_diode_2
XFILLER_23_114 vpwr vgnd scs8hd_fill_2
XFILLER_23_136 vpwr vgnd scs8hd_fill_2
XFILLER_23_147 vpwr vgnd scs8hd_fill_2
XFILLER_11_14 vgnd vpwr scs8hd_decap_6
XFILLER_11_25 vpwr vgnd scs8hd_fill_2
XFILLER_11_36 vpwr vgnd scs8hd_fill_2
XFILLER_11_47 vpwr vgnd scs8hd_fill_2
XFILLER_14_103 vpwr vgnd scs8hd_fill_2
X_173_ _173_/HI _173_/LO vgnd vpwr scs8hd_conb_1
XFILLER_37_217 vpwr vgnd scs8hd_fill_2
Xmux_left_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_left_track_9.INVTX1_0_.scs8hd_inv_1/Y
+ mem_left_track_9.LATCH_0_.latch/Q mux_left_track_9.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_9_184 vgnd vpwr scs8hd_decap_12
XANTENNA__164__A _095_/A vgnd vpwr scs8hd_diode_2
XFILLER_36_272 vgnd vpwr scs8hd_decap_3
XANTENNA__074__A _074_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mem_left_track_9.LATCH_5_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_19_217 vpwr vgnd scs8hd_fill_2
XFILLER_42_242 vgnd vpwr scs8hd_decap_6
Xmux_left_track_1.INVTX1_4_.scs8hd_inv_1 chanx_right_in[4] mux_left_track_1.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_6_154 vgnd vpwr scs8hd_decap_12
X_156_ _125_/A _157_/B _156_/Y vgnd vpwr scs8hd_nor2_4
X_087_ _076_/B _103_/A _087_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA__150__C _158_/A vgnd vpwr scs8hd_diode_2
XANTENNA__159__A _074_/A vgnd vpwr scs8hd_diode_2
XFILLER_18_272 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_left_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_left_track_1.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_33_242 vpwr vgnd scs8hd_fill_2
XANTENNA__069__A _167_/A vgnd vpwr scs8hd_diode_2
XPHY_259 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_248 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_237 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_226 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_215 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_17_57 vpwr vgnd scs8hd_fill_2
XPHY_204 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_33_56 vgnd vpwr scs8hd_decap_4
Xmux_top_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_top_track_8.INVTX1_1_.scs8hd_inv_1/Y
+ _146_/Y mux_top_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A vgnd vpwr scs8hd_ebufn_2
XFILLER_3_135 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_8.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB mem_right_track_8.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_15_275 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB mem_right_track_0.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__161__B _158_/X vgnd vpwr scs8hd_diode_2
X_208_ chanx_right_in[4] chany_top_out[2] vgnd vpwr scs8hd_buf_2
X_139_ _113_/A _136_/X _139_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_31_3 vpwr vgnd scs8hd_fill_2
XFILLER_2_190 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_1.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A _173_/HI vgnd vpwr
+ scs8hd_diode_2
XFILLER_21_245 vgnd vpwr scs8hd_decap_8
XFILLER_0_116 vpwr vgnd scs8hd_fill_2
XFILLER_0_149 vgnd vpwr scs8hd_decap_6
XANTENNA__071__B _109_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_1.tap_buf4_0_.scs8hd_inv_1_A mux_left_track_1.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_8_227 vgnd vpwr scs8hd_decap_12
XFILLER_5_27 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_2.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A _182_/HI vgnd vpwr
+ scs8hd_diode_2
XANTENNA__172__A _172_/A vgnd vpwr scs8hd_diode_2
XANTENNA__156__B _157_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_1.INVTX1_2_.scs8hd_inv_1_A chany_top_in[6] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_top_track_0.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_14_36 vgnd vpwr scs8hd_decap_3
XFILLER_14_69 vgnd vpwr scs8hd_decap_12
XFILLER_5_208 vgnd vpwr scs8hd_decap_12
XANTENNA__082__A _082_/A vgnd vpwr scs8hd_diode_2
XFILLER_39_66 vpwr vgnd scs8hd_fill_2
XFILLER_39_33 vgnd vpwr scs8hd_decap_12
XFILLER_39_22 vgnd vpwr scs8hd_decap_4
XFILLER_39_11 vpwr vgnd scs8hd_fill_2
XFILLER_29_120 vpwr vgnd scs8hd_fill_2
XFILLER_29_175 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_0.INVTX1_4_.scs8hd_inv_1_A chanx_left_in[3] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_16.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_right_track_16.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_4_263 vgnd vpwr scs8hd_decap_12
XANTENNA__167__A _167_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_9.INVTX1_4_.scs8hd_inv_1_A chanx_right_in[5] vgnd vpwr scs8hd_diode_2
XFILLER_26_189 vpwr vgnd scs8hd_fill_2
XFILLER_26_145 vgnd vpwr scs8hd_decap_3
XPHY_13 vgnd vpwr scs8hd_decap_3
XPHY_24 vgnd vpwr scs8hd_decap_3
XANTENNA__077__A address[0] vgnd vpwr scs8hd_diode_2
XPHY_35 vgnd vpwr scs8hd_decap_3
XPHY_46 vgnd vpwr scs8hd_decap_3
XFILLER_25_24 vpwr vgnd scs8hd_fill_2
XFILLER_41_34 vgnd vpwr scs8hd_decap_12
XPHY_79 vgnd vpwr scs8hd_decap_3
XPHY_68 vgnd vpwr scs8hd_decap_3
XPHY_57 vgnd vpwr scs8hd_decap_3
XFILLER_25_57 vpwr vgnd scs8hd_fill_2
XFILLER_9_3 vpwr vgnd scs8hd_fill_2
XFILLER_17_123 vgnd vpwr scs8hd_decap_3
XFILLER_17_145 vpwr vgnd scs8hd_fill_2
Xmux_right_track_0.INVTX1_5_.scs8hd_inv_1 right_bottom_grid_pin_11_ mux_right_track_0.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_31_170 vgnd vpwr scs8hd_decap_3
Xmem_top_track_0.LATCH_4_.latch data_in mem_top_track_0.LATCH_4_.latch/Q _153_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
Xmux_right_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_8.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ mem_right_track_8.LATCH_3_.latch/Q mux_right_track_8.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_top_track_14.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_top_track_14.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_36_45 vpwr vgnd scs8hd_fill_2
XFILLER_36_23 vgnd vpwr scs8hd_decap_3
X_172_ _172_/A _167_/B _172_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_20_118 vpwr vgnd scs8hd_fill_2
XANTENNA__164__B _109_/B vgnd vpwr scs8hd_diode_2
XFILLER_9_196 vgnd vpwr scs8hd_decap_12
XFILLER_28_218 vgnd vpwr scs8hd_decap_12
XANTENNA__074__B _096_/A vgnd vpwr scs8hd_diode_2
XFILLER_22_58 vpwr vgnd scs8hd_fill_2
Xmem_left_track_9.LATCH_0_.latch data_in mem_left_track_9.LATCH_0_.latch/Q _134_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA__090__A _076_/B vgnd vpwr scs8hd_diode_2
XFILLER_27_262 vgnd vpwr scs8hd_decap_12
XFILLER_6_166 vgnd vpwr scs8hd_decap_12
XFILLER_12_91 vgnd vpwr scs8hd_fill_1
X_155_ _124_/A _157_/B _155_/Y vgnd vpwr scs8hd_nor2_4
X_086_ _085_/X _103_/A vgnd vpwr scs8hd_buf_1
XFILLER_33_7 vpwr vgnd scs8hd_fill_2
XFILLER_26_6 vpwr vgnd scs8hd_fill_2
XANTENNA__159__B _158_/X vgnd vpwr scs8hd_diode_2
XFILLER_18_240 vgnd vpwr scs8hd_decap_12
XFILLER_17_36 vpwr vgnd scs8hd_fill_2
XPHY_249 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_238 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_33_35 vpwr vgnd scs8hd_fill_2
XPHY_227 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_216 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmux_top_track_16.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_top_track_16.INVTX1_2_.scs8hd_inv_1/Y
+ mem_top_track_16.LATCH_2_.latch/Q mux_top_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA__085__A _082_/A vgnd vpwr scs8hd_diode_2
XFILLER_24_210 vgnd vpwr scs8hd_decap_4
XFILLER_24_276 vgnd vpwr scs8hd_fill_1
XPHY_205 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_3_147 vgnd vpwr scs8hd_decap_12
Xmem_top_track_16.LATCH_1_.latch data_in mem_top_track_16.LATCH_1_.latch/Q _171_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_30_213 vgnd vpwr scs8hd_fill_1
X_207_ chanx_right_in[5] chany_top_out[3] vgnd vpwr scs8hd_buf_2
XANTENNA__161__C _161_/C vgnd vpwr scs8hd_diode_2
X_069_ _167_/A _111_/A vgnd vpwr scs8hd_buf_1
X_138_ _112_/A _136_/X _138_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_24_3 vgnd vpwr scs8hd_decap_3
XFILLER_0_94 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_top_track_16.LATCH_5_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_21_257 vgnd vpwr scs8hd_decap_12
Xmux_left_track_17.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_left_track_17.INVTX1_2_.scs8hd_inv_1/Y
+ mem_left_track_17.LATCH_2_.latch/Q mux_left_track_17.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_0_106 vgnd vpwr scs8hd_decap_6
XFILLER_8_239 vgnd vpwr scs8hd_decap_12
XFILLER_12_202 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_right_track_8.LATCH_3_.latch_SLEEPB _102_/Y vgnd vpwr scs8hd_diode_2
XFILLER_5_39 vgnd vpwr scs8hd_decap_12
XANTENNA__172__B _167_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_track_8.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_38_121 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_2.INVTX1_2_.scs8hd_inv_1_A chanx_right_in[8] vgnd vpwr scs8hd_diode_2
XFILLER_30_25 vpwr vgnd scs8hd_fill_2
XANTENNA__082__B address[2] vgnd vpwr scs8hd_diode_2
XFILLER_39_45 vgnd vpwr scs8hd_decap_4
XFILLER_29_132 vpwr vgnd scs8hd_fill_2
Xmem_left_track_1.LATCH_5_.latch data_in mem_left_track_1.LATCH_5_.latch/Q _121_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
Xmux_right_track_16.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_16.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ mem_right_track_16.LATCH_3_.latch/Q mux_right_track_16.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_35_179 vpwr vgnd scs8hd_fill_2
XANTENNA__167__B _167_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_8.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_right_track_8.LATCH_5_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_6_93 vgnd vpwr scs8hd_decap_12
Xmux_top_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_top_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ mem_top_track_0.LATCH_3_.latch/Q mux_top_track_0.tap_buf4_0_.scs8hd_inv_1/A vgnd
+ vpwr scs8hd_ebufn_2
Xmux_top_track_0.tap_buf4_0_.scs8hd_inv_1 mux_top_track_0.tap_buf4_0_.scs8hd_inv_1/A
+ _210_/A vgnd vpwr scs8hd_inv_1
XFILLER_41_127 vgnd vpwr scs8hd_fill_1
Xmux_right_track_8.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 mux_right_track_8.INVTX1_4_.scs8hd_inv_1/Y
+ mem_right_track_8.LATCH_1_.latch/Q mux_right_track_8.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XPHY_69 vgnd vpwr scs8hd_decap_3
XPHY_58 vgnd vpwr scs8hd_decap_3
XFILLER_26_168 vpwr vgnd scs8hd_fill_2
XPHY_14 vgnd vpwr scs8hd_decap_3
XPHY_25 vgnd vpwr scs8hd_decap_3
XPHY_36 vgnd vpwr scs8hd_decap_3
XPHY_47 vgnd vpwr scs8hd_decap_3
XFILLER_41_46 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_16.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB mem_right_track_16.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__093__A _076_/B vgnd vpwr scs8hd_diode_2
XFILLER_1_245 vgnd vpwr scs8hd_decap_12
XFILLER_17_102 vgnd vpwr scs8hd_fill_1
XFILLER_32_149 vpwr vgnd scs8hd_fill_2
XFILLER_15_91 vpwr vgnd scs8hd_fill_2
XFILLER_17_168 vpwr vgnd scs8hd_fill_2
XFILLER_17_179 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_16.INVTX1_6_.scs8hd_inv_1_A chanx_left_in[2] vgnd vpwr scs8hd_diode_2
XANTENNA__088__A address[1] vgnd vpwr scs8hd_diode_2
XFILLER_14_138 vpwr vgnd scs8hd_fill_2
X_171_ _090_/B _167_/B _171_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_13_160 vgnd vpwr scs8hd_fill_1
XFILLER_13_182 vgnd vpwr scs8hd_fill_1
XANTENNA__164__C _158_/X vgnd vpwr scs8hd_diode_2
Xmux_right_track_16.INVTX1_6_.scs8hd_inv_1 chanx_left_in[2] mux_right_track_16.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
Xmux_left_track_17.INVTX1_7_.scs8hd_inv_1 left_bottom_grid_pin_15_ mux_left_track_17.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_28_208 vpwr vgnd scs8hd_fill_2
XFILLER_11_108 vgnd vpwr scs8hd_decap_12
XANTENNA__090__B _090_/B vgnd vpwr scs8hd_diode_2
XFILLER_42_211 vgnd vpwr scs8hd_decap_6
XANTENNA_mem_left_track_17.LATCH_2_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_27_274 vgnd vpwr scs8hd_decap_3
XFILLER_10_141 vgnd vpwr scs8hd_decap_12
XFILLER_6_178 vgnd vpwr scs8hd_decap_12
X_154_ _113_/A _157_/B _154_/Y vgnd vpwr scs8hd_nor2_4
X_085_ _082_/A address[2] _162_/C _085_/X vgnd vpwr scs8hd_or3_4
XANTENNA__159__C _161_/C vgnd vpwr scs8hd_diode_2
XFILLER_18_252 vgnd vpwr scs8hd_decap_12
Xmux_left_track_9.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_left_track_9.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2/Z
+ mem_left_track_9.LATCH_4_.latch/Q mux_left_track_9.tap_buf4_0_.scs8hd_inv_1/A vgnd
+ vpwr scs8hd_ebufn_2
XANTENNA_mux_left_track_9.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_TEB mem_left_track_9.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB mem_left_track_1.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__191__A chanx_right_in[0] vgnd vpwr scs8hd_diode_2
XPHY_239 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_33_69 vpwr vgnd scs8hd_fill_2
XPHY_228 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_217 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__085__B address[2] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_0.INVTX1_3_.scs8hd_inv_1_A right_top_grid_pin_10_ vgnd vpwr
+ scs8hd_diode_2
Xmux_left_track_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 mux_left_track_1.INVTX1_3_.scs8hd_inv_1/Y
+ mem_left_track_1.LATCH_0_.latch/Q mux_left_track_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XPHY_206 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_3_159 vgnd vpwr scs8hd_decap_12
Xmem_right_track_8.LATCH_0_.latch data_in mem_right_track_8.LATCH_0_.latch/Q _108_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_30_203 vpwr vgnd scs8hd_fill_2
X_206_ _206_/A chany_top_out[4] vgnd vpwr scs8hd_buf_2
Xmux_left_track_17.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2 mux_left_track_17.INVTX1_6_.scs8hd_inv_1/Y
+ mem_left_track_17.LATCH_0_.latch/Q mux_left_track_17.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
X_137_ _111_/A _136_/X _137_/Y vgnd vpwr scs8hd_nor2_4
X_068_ _067_/X _167_/A vgnd vpwr scs8hd_buf_1
XFILLER_17_3 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_top_track_8.LATCH_1_.latch_SLEEPB _161_/Y vgnd vpwr scs8hd_diode_2
XANTENNA__186__A chanx_right_in[5] vgnd vpwr scs8hd_diode_2
XFILLER_21_214 vgnd vpwr scs8hd_fill_1
XFILLER_21_269 vgnd vpwr scs8hd_decap_8
XANTENNA_mem_left_track_17.LATCH_4_.latch_SLEEPB _138_/Y vgnd vpwr scs8hd_diode_2
Xmux_left_track_17.tap_buf4_0_.scs8hd_inv_1 mux_left_track_17.tap_buf4_0_.scs8hd_inv_1/A
+ _184_/A vgnd vpwr scs8hd_inv_1
XANTENNA_mux_right_track_8.INVTX1_5_.scs8hd_inv_1_A right_bottom_grid_pin_13_ vgnd
+ vpwr scs8hd_diode_2
XANTENNA__096__A _096_/A vgnd vpwr scs8hd_diode_2
Xmux_right_track_16.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 mux_right_track_16.INVTX1_4_.scs8hd_inv_1/Y
+ mem_right_track_16.LATCH_1_.latch/Q mux_right_track_16.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
Xmux_top_track_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 mux_top_track_0.INVTX1_4_.scs8hd_inv_1/Y
+ mem_top_track_0.LATCH_1_.latch/Q mux_top_track_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_top_track_8.INVTX1_1_.scs8hd_inv_1_A chanx_left_in[6] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_17.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_left_track_17.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_14_27 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_left_track_9.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_30_48 vpwr vgnd scs8hd_fill_2
XANTENNA__082__C _161_/C vgnd vpwr scs8hd_diode_2
XFILLER_39_57 vpwr vgnd scs8hd_fill_2
XFILLER_29_188 vgnd vpwr scs8hd_fill_1
XFILLER_29_144 vgnd vpwr scs8hd_fill_1
XFILLER_4_276 vgnd vpwr scs8hd_fill_1
XFILLER_35_158 vpwr vgnd scs8hd_fill_2
XFILLER_35_136 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_14.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _148_/Y vgnd vpwr
+ scs8hd_diode_2
Xmux_left_track_9.tap_buf4_0_.scs8hd_inv_1 mux_left_track_9.tap_buf4_0_.scs8hd_inv_1/A
+ _188_/A vgnd vpwr scs8hd_inv_1
XPHY_59 vgnd vpwr scs8hd_decap_3
XPHY_15 vgnd vpwr scs8hd_decap_3
XPHY_26 vgnd vpwr scs8hd_decap_3
XPHY_37 vgnd vpwr scs8hd_decap_3
XPHY_48 vgnd vpwr scs8hd_decap_3
XFILLER_41_58 vgnd vpwr scs8hd_decap_3
XANTENNA__093__B _172_/A vgnd vpwr scs8hd_diode_2
XFILLER_1_257 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_9.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A mux_left_track_9.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_17_114 vpwr vgnd scs8hd_fill_2
XFILLER_15_81 vgnd vpwr scs8hd_decap_3
XANTENNA_mem_right_track_8.LATCH_2_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_31_91 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_right_track_0.LATCH_4_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__194__A chanx_left_in[6] vgnd vpwr scs8hd_diode_2
XFILLER_16_191 vpwr vgnd scs8hd_fill_2
Xmem_right_track_0.LATCH_5_.latch data_in mem_right_track_0.LATCH_5_.latch/Q _076_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_right_track_16.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB mem_right_track_16.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_left_track_1.LATCH_4_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA__088__B address[2] vgnd vpwr scs8hd_diode_2
X_170_ _103_/A _167_/B _170_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_22_183 vpwr vgnd scs8hd_fill_2
Xmux_left_track_9.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2 mux_left_track_9.INVTX1_5_.scs8hd_inv_1/Y
+ mem_left_track_9.LATCH_2_.latch/Q mux_left_track_9.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_9_110 vgnd vpwr scs8hd_decap_12
XFILLER_13_172 vpwr vgnd scs8hd_fill_2
XANTENNA__164__D _162_/C vgnd vpwr scs8hd_diode_2
XANTENNA__189__A chanx_right_in[2] vgnd vpwr scs8hd_diode_2
XFILLER_3_62 vgnd vpwr scs8hd_decap_12
XFILLER_3_51 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_right_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_right_track_16.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__099__A _099_/A vgnd vpwr scs8hd_diode_2
XFILLER_27_253 vpwr vgnd scs8hd_fill_2
Xmux_top_track_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_top_track_2.INVTX1_0_.scs8hd_inv_1/Y
+ _144_/A mux_top_track_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
X_153_ _112_/A _157_/B _153_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_12_93 vgnd vpwr scs8hd_decap_12
X_084_ _076_/B _084_/B _084_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_19_7 vpwr vgnd scs8hd_fill_2
XFILLER_33_245 vgnd vpwr scs8hd_decap_12
Xmux_top_track_16.INVTX1_2_.scs8hd_inv_1 chanx_left_in[1] mux_top_track_16.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_18_264 vgnd vpwr scs8hd_decap_8
XPHY_207 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_right_track_16.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A _177_/HI vgnd vpwr
+ scs8hd_diode_2
XFILLER_33_15 vgnd vpwr scs8hd_decap_3
XPHY_229 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_218 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_top_track_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_top_track_0.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__085__C _162_/C vgnd vpwr scs8hd_diode_2
XFILLER_15_245 vgnd vpwr scs8hd_decap_8
X_136_ _136_/A _136_/X vgnd vpwr scs8hd_buf_1
X_205_ chanx_left_in[5] chany_top_out[5] vgnd vpwr scs8hd_buf_2
XANTENNA_mux_left_track_1.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB mem_left_track_1.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_top_track_16.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_top_track_0.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_23_81 vpwr vgnd scs8hd_fill_2
X_067_ address[1] _078_/B _161_/C _067_/X vgnd vpwr scs8hd_or3_4
XFILLER_28_48 vpwr vgnd scs8hd_fill_2
XANTENNA__096__B _096_/B vgnd vpwr scs8hd_diode_2
XFILLER_12_215 vgnd vpwr scs8hd_decap_12
XFILLER_12_259 vgnd vpwr scs8hd_decap_12
XFILLER_34_80 vpwr vgnd scs8hd_fill_2
X_119_ address[4] address[3] address[5] _118_/X _119_/X vgnd vpwr scs8hd_or4_4
XFILLER_38_145 vgnd vpwr scs8hd_decap_8
XFILLER_38_167 vgnd vpwr scs8hd_decap_4
XANTENNA__197__A _197_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_16.INVTX1_1_.scs8hd_inv_1_A chany_top_in[4] vgnd vpwr scs8hd_diode_2
XFILLER_29_112 vpwr vgnd scs8hd_fill_2
XFILLER_29_101 vpwr vgnd scs8hd_fill_2
XFILLER_20_71 vpwr vgnd scs8hd_fill_2
XFILLER_20_93 vgnd vpwr scs8hd_decap_3
XFILLER_35_115 vgnd vpwr scs8hd_decap_4
XFILLER_41_118 vpwr vgnd scs8hd_fill_2
XPHY_16 vgnd vpwr scs8hd_decap_3
XPHY_27 vgnd vpwr scs8hd_decap_3
XPHY_38 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_right_track_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_right_track_0.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XPHY_49 vgnd vpwr scs8hd_decap_3
XFILLER_1_269 vgnd vpwr scs8hd_decap_8
XFILLER_32_129 vgnd vpwr scs8hd_decap_6
XFILLER_17_137 vpwr vgnd scs8hd_fill_2
XFILLER_40_162 vgnd vpwr scs8hd_decap_3
XFILLER_40_151 vpwr vgnd scs8hd_fill_2
XFILLER_40_140 vgnd vpwr scs8hd_fill_1
XFILLER_16_170 vgnd vpwr scs8hd_decap_8
XFILLER_23_118 vpwr vgnd scs8hd_fill_2
XFILLER_31_195 vpwr vgnd scs8hd_fill_2
XFILLER_11_29 vgnd vpwr scs8hd_decap_4
XFILLER_39_262 vgnd vpwr scs8hd_decap_12
XFILLER_36_15 vpwr vgnd scs8hd_fill_2
XFILLER_14_107 vgnd vpwr scs8hd_decap_12
XANTENNA__088__C _161_/C vgnd vpwr scs8hd_diode_2
XFILLER_22_173 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_right_track_0.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A _176_/HI vgnd vpwr
+ scs8hd_diode_2
XFILLER_7_3 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _144_/A vgnd vpwr
+ scs8hd_diode_2
Xmux_right_track_0.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2 mux_right_track_0.INVTX1_7_.scs8hd_inv_1/Y
+ mem_right_track_0.LATCH_1_.latch/Q mux_right_track_0.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_left_track_17.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A mux_left_track_17.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_13_184 vgnd vpwr scs8hd_decap_12
XFILLER_3_74 vgnd vpwr scs8hd_decap_12
Xmux_left_track_1.INVTX1_1_.scs8hd_inv_1 chany_top_in[3] mux_left_track_1.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_36_276 vgnd vpwr scs8hd_fill_1
XFILLER_36_210 vgnd vpwr scs8hd_decap_4
XFILLER_22_28 vgnd vpwr scs8hd_decap_3
XFILLER_10_154 vgnd vpwr scs8hd_decap_12
XFILLER_8_19 vgnd vpwr scs8hd_decap_12
X_083_ _082_/X _084_/B vgnd vpwr scs8hd_buf_1
X_152_ _167_/A _157_/B _152_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA_mux_right_track_8.INVTX1_0_.scs8hd_inv_1_A chany_top_in[0] vgnd vpwr scs8hd_diode_2
XFILLER_18_276 vgnd vpwr scs8hd_fill_1
XFILLER_33_257 vgnd vpwr scs8hd_decap_12
XFILLER_33_213 vgnd vpwr scs8hd_decap_6
XPHY_219 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_208 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mem_top_track_16.LATCH_3_.latch_SLEEPB _169_/Y vgnd vpwr scs8hd_diode_2
XFILLER_24_224 vpwr vgnd scs8hd_fill_2
XFILLER_24_235 vgnd vpwr scs8hd_decap_12
XFILLER_33_27 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_16.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_right_track_16.LATCH_5_.latch/Q
+ vgnd vpwr scs8hd_diode_2
X_204_ chanx_left_in[4] chany_top_out[6] vgnd vpwr scs8hd_buf_2
XANTENNA_mem_top_track_0.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
X_066_ address[0] _161_/C vgnd vpwr scs8hd_inv_8
XFILLER_23_60 vgnd vpwr scs8hd_fill_1
X_135_ _095_/A address[3] address[5] _118_/X _136_/A vgnd vpwr scs8hd_or4_4
XFILLER_31_7 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_left_track_17.INVTX1_4_.scs8hd_inv_1_A chanx_right_in[6] vgnd vpwr scs8hd_diode_2
XFILLER_9_62 vgnd vpwr scs8hd_decap_12
XFILLER_21_227 vpwr vgnd scs8hd_fill_2
XFILLER_28_27 vpwr vgnd scs8hd_fill_2
XFILLER_12_227 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB mem_top_track_0.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_20_260 vgnd vpwr scs8hd_decap_12
XFILLER_18_93 vgnd vpwr scs8hd_fill_1
XFILLER_7_220 vgnd vpwr scs8hd_decap_12
X_118_ _118_/A _118_/B _118_/X vgnd vpwr scs8hd_or2_4
XFILLER_38_135 vgnd vpwr scs8hd_fill_1
XFILLER_22_3 vpwr vgnd scs8hd_fill_2
XFILLER_30_17 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_right_track_16.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_29_179 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_top_track_0.LATCH_5_.latch_SLEEPB _152_/Y vgnd vpwr scs8hd_diode_2
Xmux_left_track_9.INVTX1_6_.scs8hd_inv_1 left_bottom_grid_pin_7_ mux_left_track_9.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_35_105 vgnd vpwr scs8hd_decap_4
XPHY_17 vgnd vpwr scs8hd_decap_3
XPHY_28 vgnd vpwr scs8hd_decap_3
XPHY_39 vgnd vpwr scs8hd_decap_3
XFILLER_25_28 vpwr vgnd scs8hd_fill_2
XFILLER_9_7 vgnd vpwr scs8hd_decap_12
Xmux_right_track_0.INVTX1_2_.scs8hd_inv_1 chany_top_in[8] mux_right_track_0.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_17_149 vpwr vgnd scs8hd_fill_2
XFILLER_39_274 vgnd vpwr scs8hd_decap_3
XFILLER_36_49 vgnd vpwr scs8hd_decap_4
XFILLER_14_119 vgnd vpwr scs8hd_decap_6
Xmem_left_track_17.LATCH_2_.latch data_in mem_left_track_17.LATCH_2_.latch/Q _140_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_top_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_top_track_16.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_22_130 vgnd vpwr scs8hd_decap_4
XFILLER_26_93 vgnd vpwr scs8hd_decap_4
XFILLER_26_82 vpwr vgnd scs8hd_fill_2
XFILLER_9_123 vgnd vpwr scs8hd_decap_12
XFILLER_13_141 vpwr vgnd scs8hd_fill_2
XFILLER_26_71 vpwr vgnd scs8hd_fill_2
XFILLER_13_196 vgnd vpwr scs8hd_decap_12
XFILLER_3_86 vgnd vpwr scs8hd_decap_12
XFILLER_27_222 vpwr vgnd scs8hd_fill_2
XFILLER_27_211 vgnd vpwr scs8hd_decap_4
XFILLER_27_200 vgnd vpwr scs8hd_decap_4
XFILLER_10_166 vgnd vpwr scs8hd_decap_12
X_151_ _150_/X _157_/B vgnd vpwr scs8hd_buf_1
XFILLER_12_51 vgnd vpwr scs8hd_decap_8
XFILLER_12_62 vpwr vgnd scs8hd_fill_2
XFILLER_12_73 vgnd vpwr scs8hd_decap_12
X_082_ _082_/A address[2] _161_/C _082_/X vgnd vpwr scs8hd_or3_4
XFILLER_33_269 vgnd vpwr scs8hd_decap_8
XFILLER_33_39 vpwr vgnd scs8hd_fill_2
XPHY_209 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_247 vgnd vpwr scs8hd_decap_8
Xmux_left_track_1.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2 _173_/HI mem_left_track_1.LATCH_2_.latch/Q
+ mux_left_track_1.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XFILLER_15_214 vgnd vpwr scs8hd_fill_1
Xmux_top_track_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_top_track_2.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ _143_/Y mux_top_track_2.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
X_203_ _203_/A chany_top_out[7] vgnd vpwr scs8hd_buf_2
Xmux_right_track_8.INVTX1_7_.scs8hd_inv_1 chanx_left_in[5] mux_right_track_8.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
X_065_ address[2] _078_/B vgnd vpwr scs8hd_inv_8
X_134_ _108_/A _132_/B _134_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_23_94 vpwr vgnd scs8hd_fill_2
XFILLER_0_32 vgnd vpwr scs8hd_decap_12
XFILLER_21_217 vgnd vpwr scs8hd_fill_1
XANTENNA_mem_right_track_8.LATCH_0_.latch_SLEEPB _108_/Y vgnd vpwr scs8hd_diode_2
XFILLER_9_74 vgnd vpwr scs8hd_decap_12
XFILLER_21_239 vgnd vpwr scs8hd_decap_4
XFILLER_28_17 vpwr vgnd scs8hd_fill_2
XFILLER_12_239 vgnd vpwr scs8hd_decap_12
XFILLER_20_272 vgnd vpwr scs8hd_decap_3
XFILLER_18_61 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_left_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_left_track_17.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_7_232 vgnd vpwr scs8hd_decap_12
X_117_ enable _118_/A vgnd vpwr scs8hd_inv_8
XFILLER_38_125 vpwr vgnd scs8hd_fill_2
Xmem_left_track_1.LATCH_0_.latch data_in mem_left_track_1.LATCH_0_.latch/Q _126_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_15_3 vpwr vgnd scs8hd_fill_2
XFILLER_30_29 vpwr vgnd scs8hd_fill_2
Xmux_right_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_8.INVTX1_0_.scs8hd_inv_1/Y
+ mem_right_track_8.LATCH_0_.latch/Q mux_right_track_8.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_29_136 vpwr vgnd scs8hd_fill_2
XFILLER_29_158 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_left_track_1.LATCH_3_.latch_SLEEPB _123_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_8.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB mem_right_track_8.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_top_track_8.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_track_0.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_4_202 vgnd vpwr scs8hd_decap_12
XFILLER_20_84 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_right_track_0.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xmem_right_track_16.LATCH_1_.latch data_in mem_right_track_16.LATCH_1_.latch/Q _115_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_left_track_1.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_left_track_1.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_26_128 vpwr vgnd scs8hd_fill_2
XPHY_18 vgnd vpwr scs8hd_decap_3
XPHY_29 vgnd vpwr scs8hd_decap_3
XFILLER_34_183 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_left_track_17.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A mux_left_track_17.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_left_track_17.LATCH_5_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_15_73 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_right_track_16.LATCH_3_.latch_SLEEPB _113_/Y vgnd vpwr scs8hd_diode_2
XFILLER_15_95 vpwr vgnd scs8hd_fill_2
XANTENNA__102__A _113_/A vgnd vpwr scs8hd_diode_2
XFILLER_31_175 vpwr vgnd scs8hd_fill_2
XFILLER_31_153 vgnd vpwr scs8hd_fill_1
XFILLER_39_253 vpwr vgnd scs8hd_fill_2
XFILLER_36_28 vgnd vpwr scs8hd_decap_3
Xmux_left_track_17.INVTX1_4_.scs8hd_inv_1 chanx_right_in[6] mux_left_track_17.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
Xmux_right_track_16.INVTX1_3_.scs8hd_inv_1 right_bottom_grid_pin_3_ mux_right_track_16.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_9_135 vgnd vpwr scs8hd_decap_12
XFILLER_13_153 vgnd vpwr scs8hd_fill_1
XFILLER_13_164 vpwr vgnd scs8hd_fill_2
XFILLER_3_98 vgnd vpwr scs8hd_decap_12
XFILLER_8_190 vgnd vpwr scs8hd_decap_12
XFILLER_22_19 vpwr vgnd scs8hd_fill_2
XFILLER_27_245 vgnd vpwr scs8hd_decap_8
X_150_ address[4] address[3] _158_/A _150_/X vgnd vpwr scs8hd_or3_4
XANTENNA_mux_right_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_8.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_10_178 vgnd vpwr scs8hd_decap_12
XFILLER_6_105 vgnd vpwr scs8hd_decap_12
XFILLER_12_85 vgnd vpwr scs8hd_decap_6
X_081_ address[1] _082_/A vgnd vpwr scs8hd_inv_8
XFILLER_18_201 vgnd vpwr scs8hd_decap_4
XFILLER_5_171 vgnd vpwr scs8hd_decap_12
XFILLER_17_19 vpwr vgnd scs8hd_fill_2
XFILLER_32_270 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_top_track_16.INVTX1_1_.scs8hd_inv_1_A chanx_right_in[3] vgnd vpwr scs8hd_diode_2
XFILLER_24_259 vgnd vpwr scs8hd_decap_12
XANTENNA__200__A chanx_left_in[0] vgnd vpwr scs8hd_diode_2
XFILLER_15_204 vpwr vgnd scs8hd_fill_2
XFILLER_15_259 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_left_track_17.LATCH_1_.latch_SLEEPB _141_/Y vgnd vpwr scs8hd_diode_2
X_202_ _202_/A chany_top_out[8] vgnd vpwr scs8hd_buf_2
XFILLER_30_218 vgnd vpwr scs8hd_decap_12
XFILLER_30_207 vgnd vpwr scs8hd_decap_6
X_133_ _125_/A _132_/B _133_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_23_62 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_right_track_8.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A mux_right_track_8.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xmux_right_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_16.INVTX1_0_.scs8hd_inv_1/Y
+ mem_right_track_16.LATCH_0_.latch/Q mux_right_track_16.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_2_141 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_14.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _147_/Y vgnd vpwr
+ scs8hd_diode_2
XANTENNA__110__A _110_/A vgnd vpwr scs8hd_diode_2
XFILLER_0_44 vgnd vpwr scs8hd_decap_12
XFILLER_17_7 vgnd vpwr scs8hd_decap_3
XFILLER_24_8 vpwr vgnd scs8hd_fill_2
XFILLER_9_42 vgnd vpwr scs8hd_fill_1
XFILLER_9_31 vgnd vpwr scs8hd_fill_1
XFILLER_0_66 vpwr vgnd scs8hd_fill_2
XFILLER_0_77 vpwr vgnd scs8hd_fill_2
Xmux_top_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_top_track_0.INVTX1_0_.scs8hd_inv_1/Y
+ mem_top_track_0.LATCH_0_.latch/Q mux_top_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_9_86 vgnd vpwr scs8hd_decap_12
XFILLER_18_40 vpwr vgnd scs8hd_fill_2
XFILLER_18_84 vpwr vgnd scs8hd_fill_2
X_116_ _108_/A _110_/X _116_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA__105__A _090_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_track_8.LATCH_5_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_38_104 vgnd vpwr scs8hd_decap_8
XFILLER_6_32 vgnd vpwr scs8hd_decap_12
XFILLER_34_173 vgnd vpwr scs8hd_fill_1
XPHY_19 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_right_track_8.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB mem_right_track_8.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xmem_top_track_8.LATCH_0_.latch data_in _146_/A _162_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
Xmem_right_track_0.LATCH_0_.latch data_in mem_right_track_0.LATCH_0_.latch/Q _093_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_right_track_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB mem_right_track_0.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_17_118 vpwr vgnd scs8hd_fill_2
XFILLER_40_143 vgnd vpwr scs8hd_decap_8
XFILLER_25_162 vpwr vgnd scs8hd_fill_2
XFILLER_25_195 vpwr vgnd scs8hd_fill_2
XFILLER_31_73 vgnd vpwr scs8hd_decap_3
XFILLER_31_40 vpwr vgnd scs8hd_fill_2
Xmux_left_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_left_track_9.INVTX1_1_.scs8hd_inv_1/Y
+ mem_left_track_9.LATCH_1_.latch/Q mux_left_track_9.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA__102__B _106_/B vgnd vpwr scs8hd_diode_2
XFILLER_31_132 vpwr vgnd scs8hd_fill_2
XPHY_190 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_39_210 vgnd vpwr scs8hd_decap_4
XFILLER_22_143 vgnd vpwr scs8hd_decap_4
XFILLER_22_154 vpwr vgnd scs8hd_fill_2
XFILLER_22_165 vgnd vpwr scs8hd_decap_8
XFILLER_22_187 vpwr vgnd scs8hd_fill_2
XANTENNA__203__A _203_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_16.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_top_track_16.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_top_track_0.LATCH_4_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_42_94 vgnd vpwr scs8hd_decap_12
XFILLER_9_147 vgnd vpwr scs8hd_decap_12
XFILLER_13_176 vgnd vpwr scs8hd_decap_6
XANTENNA__113__A _113_/A vgnd vpwr scs8hd_diode_2
XFILLER_36_224 vgnd vpwr scs8hd_decap_12
XFILLER_42_249 vgnd vpwr scs8hd_decap_12
XFILLER_6_117 vgnd vpwr scs8hd_decap_12
X_080_ _076_/B _099_/A _080_/Y vgnd vpwr scs8hd_nor2_4
Xmux_right_track_0.tap_buf4_0_.scs8hd_inv_1 mux_right_track_0.tap_buf4_0_.scs8hd_inv_1/A
+ _201_/A vgnd vpwr scs8hd_inv_1
XFILLER_5_3 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A mux_left_track_1.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_18_224 vpwr vgnd scs8hd_fill_2
XANTENNA__108__A _108_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mem_left_track_9.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_top_track_2.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
X_201_ _201_/A chanx_right_out[0] vgnd vpwr scs8hd_buf_2
Xmem_top_track_0.LATCH_5_.latch data_in mem_top_track_0.LATCH_5_.latch/Q _152_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_23_52 vpwr vgnd scs8hd_fill_2
X_132_ _124_/A _132_/B _132_/Y vgnd vpwr scs8hd_nor2_4
Xmux_right_track_16.tap_buf4_0_.scs8hd_inv_1 mux_right_track_16.tap_buf4_0_.scs8hd_inv_1/A
+ _193_/A vgnd vpwr scs8hd_inv_1
XFILLER_0_56 vgnd vpwr scs8hd_decap_6
XFILLER_9_98 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_1.INVTX1_3_.scs8hd_inv_1_A chanx_right_in[0] vgnd vpwr scs8hd_diode_2
XFILLER_34_84 vpwr vgnd scs8hd_fill_2
XFILLER_34_40 vgnd vpwr scs8hd_fill_1
X_115_ _125_/A _110_/X _115_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_7_245 vgnd vpwr scs8hd_decap_12
XANTENNA__121__A _111_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_9.INVTX1_5_.scs8hd_inv_1_A left_bottom_grid_pin_1_ vgnd vpwr
+ scs8hd_diode_2
Xmem_left_track_9.LATCH_1_.latch data_in mem_left_track_9.LATCH_1_.latch/Q _133_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_39_29 vpwr vgnd scs8hd_fill_2
XFILLER_39_18 vpwr vgnd scs8hd_fill_2
XFILLER_29_116 vpwr vgnd scs8hd_fill_2
XFILLER_29_105 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_right_track_0.LATCH_4_.latch_SLEEPB _080_/Y vgnd vpwr scs8hd_diode_2
XANTENNA__206__A _206_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _143_/A vgnd vpwr
+ scs8hd_diode_2
XFILLER_4_215 vgnd vpwr scs8hd_decap_12
XFILLER_20_64 vgnd vpwr scs8hd_decap_4
XFILLER_35_119 vgnd vpwr scs8hd_fill_1
XFILLER_29_84 vpwr vgnd scs8hd_fill_2
XANTENNA__116__A _108_/A vgnd vpwr scs8hd_diode_2
XFILLER_6_44 vgnd vpwr scs8hd_decap_12
Xmem_top_track_16.LATCH_2_.latch data_in mem_top_track_16.LATCH_2_.latch/Q _170_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_20_3 vgnd vpwr scs8hd_decap_3
Xmux_right_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_right_track_8.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ mem_right_track_8.LATCH_4_.latch/Q mux_right_track_8.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_15_20 vpwr vgnd scs8hd_fill_2
XFILLER_15_53 vpwr vgnd scs8hd_fill_2
Xmux_right_track_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_0.INVTX1_3_.scs8hd_inv_1/Y
+ mem_right_track_0.LATCH_0_.latch/Q mux_right_track_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_16_141 vgnd vpwr scs8hd_decap_12
XFILLER_31_199 vpwr vgnd scs8hd_fill_2
XFILLER_31_166 vpwr vgnd scs8hd_fill_2
XPHY_180 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_191 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_right_track_0.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB mem_right_track_0.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_39_200 vpwr vgnd scs8hd_fill_2
.ends

