magic
tech EFS8A
magscale 1 2
timestamp 1602088566
<< locali >>
rect 11799 18921 11805 18955
rect 11799 18853 11833 18921
rect 2231 17833 2237 17867
rect 15663 17833 15669 17867
rect 17503 17833 17509 17867
rect 2231 17765 2265 17833
rect 15663 17765 15697 17833
rect 17503 17765 17537 17833
rect 9631 16609 9758 16643
rect 15427 16609 15554 16643
rect 10971 15895 11005 15963
rect 10971 15861 10977 15895
rect 15663 15657 15669 15691
rect 15663 15589 15697 15657
rect 4663 15521 4790 15555
rect 13403 15521 13530 15555
rect 19895 14807 19929 14875
rect 19895 14773 19901 14807
rect 2599 14569 2605 14603
rect 4439 14569 4445 14603
rect 2599 14501 2633 14569
rect 4439 14501 4473 14569
rect 6469 13787 6503 14025
rect 19435 13719 19469 13787
rect 19435 13685 19441 13719
rect 19435 13481 19441 13515
rect 19435 13413 19469 13481
rect 11931 13345 11966 13379
rect 5675 12733 5710 12767
rect 14651 12631 14685 12699
rect 14651 12597 14657 12631
rect 8343 12257 8378 12291
rect 6469 11543 6503 11849
rect 7199 11543 7233 11611
rect 7199 11509 7205 11543
rect 3985 10523 4019 10761
rect 1863 10217 1869 10251
rect 4439 10217 4445 10251
rect 15755 10217 15761 10251
rect 1863 10149 1897 10217
rect 4439 10149 4473 10217
rect 15755 10149 15789 10217
rect 19947 9129 20085 9163
rect 13679 8993 13714 9027
rect 18797 8279 18831 8449
rect 4439 8041 4445 8075
rect 4439 7973 4473 8041
rect 19291 7973 19336 8007
rect 8251 7905 8286 7939
rect 15243 7905 15370 7939
rect 11529 6817 11690 6851
rect 11529 6783 11563 6817
rect 12449 5083 12483 5253
rect 15847 4777 15853 4811
rect 18975 4777 18981 4811
rect 15847 4709 15881 4777
rect 18975 4709 19009 4777
rect 13415 3689 13461 3723
<< viali >>
rect 5825 20553 5859 20587
rect 8125 20553 8159 20587
rect 10885 20553 10919 20587
rect 15301 20553 15335 20587
rect 19441 20553 19475 20587
rect 1547 20417 1581 20451
rect 1460 20349 1494 20383
rect 5641 20349 5675 20383
rect 6193 20349 6227 20383
rect 7941 20349 7975 20383
rect 10701 20349 10735 20383
rect 15117 20349 15151 20383
rect 15669 20349 15703 20383
rect 19257 20349 19291 20383
rect 19809 20349 19843 20383
rect 1869 20213 1903 20247
rect 8493 20213 8527 20247
rect 11345 20213 11379 20247
rect 17325 20009 17359 20043
rect 9756 19873 9790 19907
rect 17141 19873 17175 19907
rect 9827 19669 9861 19703
rect 10241 19669 10275 19703
rect 21051 19465 21085 19499
rect 20948 19261 20982 19295
rect 21373 19261 21407 19295
rect 8861 19193 8895 19227
rect 9689 19193 9723 19227
rect 9965 19193 9999 19227
rect 10057 19193 10091 19227
rect 10609 19193 10643 19227
rect 9413 19125 9447 19159
rect 17233 19125 17267 19159
rect 10609 18921 10643 18955
rect 11805 18921 11839 18955
rect 21097 18921 21131 18955
rect 1547 18853 1581 18887
rect 10051 18853 10085 18887
rect 1460 18785 1494 18819
rect 6929 18785 6963 18819
rect 7113 18785 7147 18819
rect 15336 18785 15370 18819
rect 16589 18785 16623 18819
rect 17049 18785 17083 18819
rect 20913 18785 20947 18819
rect 7205 18717 7239 18751
rect 9689 18717 9723 18751
rect 11437 18717 11471 18751
rect 17325 18717 17359 18751
rect 19441 18717 19475 18751
rect 4905 18581 4939 18615
rect 8309 18581 8343 18615
rect 12357 18581 12391 18615
rect 12633 18581 12667 18615
rect 15439 18581 15473 18615
rect 15761 18581 15795 18615
rect 16129 18581 16163 18615
rect 18797 18581 18831 18615
rect 9689 18377 9723 18411
rect 11529 18377 11563 18411
rect 12265 18377 12299 18411
rect 20361 18377 20395 18411
rect 7021 18309 7055 18343
rect 14335 18309 14369 18343
rect 4997 18241 5031 18275
rect 5365 18241 5399 18275
rect 8585 18241 8619 18275
rect 10517 18241 10551 18275
rect 10793 18241 10827 18275
rect 12541 18241 12575 18275
rect 12817 18241 12851 18275
rect 15393 18241 15427 18275
rect 18797 18241 18831 18275
rect 20637 18241 20671 18275
rect 20913 18241 20947 18275
rect 3433 18173 3467 18207
rect 3893 18173 3927 18207
rect 9873 18173 9907 18207
rect 10333 18173 10367 18207
rect 14264 18173 14298 18207
rect 14657 18173 14691 18207
rect 3249 18105 3283 18139
rect 4077 18105 4111 18139
rect 5089 18105 5123 18139
rect 8309 18105 8343 18139
rect 8401 18105 8435 18139
rect 9321 18105 9355 18139
rect 12633 18105 12667 18139
rect 15485 18105 15519 18139
rect 16037 18105 16071 18139
rect 19118 18105 19152 18139
rect 20729 18105 20763 18139
rect 1685 18037 1719 18071
rect 1961 18037 1995 18071
rect 4445 18037 4479 18071
rect 4813 18037 4847 18071
rect 7481 18037 7515 18071
rect 8033 18037 8067 18071
rect 11805 18037 11839 18071
rect 15209 18037 15243 18071
rect 16681 18037 16715 18071
rect 17049 18037 17083 18071
rect 18613 18037 18647 18071
rect 19717 18037 19751 18071
rect 21557 18037 21591 18071
rect 2237 17833 2271 17867
rect 3433 17833 3467 17867
rect 5181 17833 5215 17867
rect 15669 17833 15703 17867
rect 16221 17833 16255 17867
rect 17509 17833 17543 17867
rect 18981 17833 19015 17867
rect 20545 17833 20579 17867
rect 21097 17833 21131 17867
rect 4582 17765 4616 17799
rect 7567 17765 7601 17799
rect 11345 17765 11379 17799
rect 12633 17765 12667 17799
rect 4261 17697 4295 17731
rect 6044 17697 6078 17731
rect 7205 17697 7239 17731
rect 10885 17697 10919 17731
rect 11069 17697 11103 17731
rect 14048 17697 14082 17731
rect 17141 17697 17175 17731
rect 18889 17697 18923 17731
rect 19349 17697 19383 17731
rect 20913 17697 20947 17731
rect 1869 17629 1903 17663
rect 12541 17629 12575 17663
rect 12817 17629 12851 17663
rect 14151 17629 14185 17663
rect 15301 17629 15335 17663
rect 1777 17493 1811 17527
rect 2789 17493 2823 17527
rect 6147 17493 6181 17527
rect 8125 17493 8159 17527
rect 9873 17493 9907 17527
rect 10517 17493 10551 17527
rect 18061 17493 18095 17527
rect 18429 17493 18463 17527
rect 19901 17493 19935 17527
rect 1961 17289 1995 17323
rect 3893 17289 3927 17323
rect 6009 17289 6043 17323
rect 9551 17289 9585 17323
rect 16681 17289 16715 17323
rect 17877 17289 17911 17323
rect 19441 17289 19475 17323
rect 20913 17289 20947 17323
rect 2881 17221 2915 17255
rect 7389 17221 7423 17255
rect 2329 17153 2363 17187
rect 3249 17153 3283 17187
rect 5089 17153 5123 17187
rect 6975 17153 7009 17187
rect 7941 17153 7975 17187
rect 8861 17153 8895 17187
rect 12541 17153 12575 17187
rect 12817 17153 12851 17187
rect 14841 17153 14875 17187
rect 15761 17153 15795 17187
rect 18153 17153 18187 17187
rect 18797 17153 18831 17187
rect 19993 17153 20027 17187
rect 6888 17085 6922 17119
rect 9480 17085 9514 17119
rect 10701 17085 10735 17119
rect 10885 17085 10919 17119
rect 11437 17085 11471 17119
rect 14105 17085 14139 17119
rect 14565 17085 14599 17119
rect 2421 17017 2455 17051
rect 4445 17017 4479 17051
rect 4537 17017 4571 17051
rect 8033 17017 8067 17051
rect 8585 17017 8619 17051
rect 10333 17017 10367 17051
rect 11161 17017 11195 17051
rect 12633 17017 12667 17051
rect 13645 17017 13679 17051
rect 15853 17017 15887 17051
rect 16405 17017 16439 17051
rect 18245 17017 18279 17051
rect 19717 17017 19751 17051
rect 19809 17017 19843 17051
rect 4169 16949 4203 16983
rect 5365 16949 5399 16983
rect 7757 16949 7791 16983
rect 9965 16949 9999 16983
rect 11805 16949 11839 16983
rect 12265 16949 12299 16983
rect 13921 16949 13955 16983
rect 15393 16949 15427 16983
rect 17141 16949 17175 16983
rect 19073 16949 19107 16983
rect 1869 16745 1903 16779
rect 2789 16745 2823 16779
rect 4997 16745 5031 16779
rect 7205 16745 7239 16779
rect 7941 16745 7975 16779
rect 10701 16745 10735 16779
rect 12357 16745 12391 16779
rect 12725 16745 12759 16779
rect 14197 16745 14231 16779
rect 15945 16745 15979 16779
rect 16313 16745 16347 16779
rect 17969 16745 18003 16779
rect 19441 16745 19475 16779
rect 19809 16745 19843 16779
rect 4398 16677 4432 16711
rect 5733 16677 5767 16711
rect 5917 16677 5951 16711
rect 6009 16677 6043 16711
rect 8217 16677 8251 16711
rect 11758 16677 11792 16711
rect 13369 16677 13403 16711
rect 18842 16677 18876 16711
rect 1777 16609 1811 16643
rect 2329 16609 2363 16643
rect 9597 16609 9631 16643
rect 13001 16609 13035 16643
rect 15393 16609 15427 16643
rect 17233 16609 17267 16643
rect 17417 16609 17451 16643
rect 20913 16609 20947 16643
rect 4077 16541 4111 16575
rect 6193 16541 6227 16575
rect 8125 16541 8159 16575
rect 8401 16541 8435 16575
rect 11437 16541 11471 16575
rect 13277 16541 13311 16575
rect 13553 16541 13587 16575
rect 17693 16541 17727 16575
rect 18521 16541 18555 16575
rect 21097 16473 21131 16507
rect 6929 16405 6963 16439
rect 9827 16405 9861 16439
rect 15623 16405 15657 16439
rect 18337 16405 18371 16439
rect 3801 16201 3835 16235
rect 4169 16201 4203 16235
rect 4813 16201 4847 16235
rect 5917 16201 5951 16235
rect 6193 16201 6227 16235
rect 6561 16201 6595 16235
rect 10517 16201 10551 16235
rect 11529 16201 11563 16235
rect 12173 16201 12207 16235
rect 12587 16201 12621 16235
rect 13645 16201 13679 16235
rect 15485 16201 15519 16235
rect 19073 16201 19107 16235
rect 19441 16201 19475 16235
rect 1593 16133 1627 16167
rect 9045 16133 9079 16167
rect 11897 16133 11931 16167
rect 13277 16133 13311 16167
rect 16405 16133 16439 16167
rect 2513 16065 2547 16099
rect 3341 16065 3375 16099
rect 7205 16065 7239 16099
rect 8493 16065 8527 16099
rect 14841 16065 14875 16099
rect 15853 16065 15887 16099
rect 18153 16065 18187 16099
rect 18429 16065 18463 16099
rect 1409 15997 1443 16031
rect 2605 15997 2639 16031
rect 3157 15997 3191 16031
rect 4537 15997 4571 16031
rect 4997 15997 5031 16031
rect 10149 15997 10183 16031
rect 10609 15997 10643 16031
rect 12516 15997 12550 16031
rect 2053 15929 2087 15963
rect 5318 15929 5352 15963
rect 6929 15929 6963 15963
rect 7021 15929 7055 15963
rect 7941 15929 7975 15963
rect 8309 15929 8343 15963
rect 8585 15929 8619 15963
rect 15209 15929 15243 15963
rect 15945 15929 15979 15963
rect 17877 15929 17911 15963
rect 18245 15929 18279 15963
rect 20913 15929 20947 15963
rect 9689 15861 9723 15895
rect 10977 15861 11011 15895
rect 13001 15861 13035 15895
rect 16957 15861 16991 15895
rect 17417 15861 17451 15895
rect 1961 15657 1995 15691
rect 4859 15657 4893 15691
rect 8769 15657 8803 15691
rect 9137 15657 9171 15691
rect 10241 15657 10275 15691
rect 15669 15657 15703 15691
rect 16221 15657 16255 15691
rect 17187 15657 17221 15691
rect 21051 15657 21085 15691
rect 1547 15589 1581 15623
rect 5273 15589 5307 15623
rect 8211 15589 8245 15623
rect 18346 15589 18380 15623
rect 18889 15589 18923 15623
rect 1460 15521 1494 15555
rect 4629 15521 4663 15555
rect 6009 15521 6043 15555
rect 6193 15521 6227 15555
rect 10241 15521 10275 15555
rect 10425 15521 10459 15555
rect 11964 15521 11998 15555
rect 13369 15521 13403 15555
rect 17116 15521 17150 15555
rect 20948 15521 20982 15555
rect 6469 15453 6503 15487
rect 7849 15453 7883 15487
rect 12541 15453 12575 15487
rect 15301 15453 15335 15487
rect 18245 15453 18279 15487
rect 2237 15385 2271 15419
rect 7205 15385 7239 15419
rect 12035 15385 12069 15419
rect 13599 15385 13633 15419
rect 2605 15317 2639 15351
rect 7573 15317 7607 15351
rect 12817 15317 12851 15351
rect 14013 15317 14047 15351
rect 16497 15317 16531 15351
rect 19533 15317 19567 15351
rect 3065 15113 3099 15147
rect 7297 15113 7331 15147
rect 9413 15113 9447 15147
rect 13553 15113 13587 15147
rect 16957 15113 16991 15147
rect 18245 15113 18279 15147
rect 20913 15113 20947 15147
rect 6193 14977 6227 15011
rect 8033 14977 8067 15011
rect 12541 14977 12575 15011
rect 2329 14909 2363 14943
rect 2605 14909 2639 14943
rect 3617 14909 3651 14943
rect 4169 14909 4203 14943
rect 5457 14909 5491 14943
rect 5641 14909 5675 14943
rect 7665 14909 7699 14943
rect 7941 14909 7975 14943
rect 9045 14909 9079 14943
rect 9505 14909 9539 14943
rect 9965 14909 9999 14943
rect 10517 14909 10551 14943
rect 11253 14909 11287 14943
rect 11380 14909 11414 14943
rect 14013 14909 14047 14943
rect 14565 14909 14599 14943
rect 16037 14909 16071 14943
rect 19533 14909 19567 14943
rect 2789 14841 2823 14875
rect 6653 14841 6687 14875
rect 10241 14841 10275 14875
rect 12633 14841 12667 14875
rect 13185 14841 13219 14875
rect 13921 14841 13955 14875
rect 14749 14841 14783 14875
rect 16358 14841 16392 14875
rect 17233 14841 17267 14875
rect 1961 14773 1995 14807
rect 3433 14773 3467 14807
rect 3893 14773 3927 14807
rect 4813 14773 4847 14807
rect 5457 14773 5491 14807
rect 8585 14773 8619 14807
rect 11483 14773 11517 14807
rect 11989 14773 12023 14807
rect 15301 14773 15335 14807
rect 15853 14773 15887 14807
rect 18705 14773 18739 14807
rect 19441 14773 19475 14807
rect 19901 14773 19935 14807
rect 20453 14773 20487 14807
rect 21281 14773 21315 14807
rect 2605 14569 2639 14603
rect 3617 14569 3651 14603
rect 4445 14569 4479 14603
rect 5365 14569 5399 14603
rect 7849 14569 7883 14603
rect 8723 14569 8757 14603
rect 15485 14569 15519 14603
rect 19579 14569 19613 14603
rect 2145 14501 2179 14535
rect 7021 14501 7055 14535
rect 10603 14501 10637 14535
rect 12173 14501 12207 14535
rect 12265 14501 12299 14535
rect 13829 14501 13863 14535
rect 15853 14501 15887 14535
rect 16405 14501 16439 14535
rect 18613 14501 18647 14535
rect 21005 14501 21039 14535
rect 21097 14501 21131 14535
rect 4077 14433 4111 14467
rect 8652 14433 8686 14467
rect 10241 14433 10275 14467
rect 17877 14433 17911 14467
rect 18337 14433 18371 14467
rect 19508 14433 19542 14467
rect 2237 14365 2271 14399
rect 6929 14365 6963 14399
rect 12449 14365 12483 14399
rect 13737 14365 13771 14399
rect 14013 14365 14047 14399
rect 15761 14365 15795 14399
rect 21281 14365 21315 14399
rect 3157 14297 3191 14331
rect 7481 14297 7515 14331
rect 11161 14297 11195 14331
rect 1593 14229 1627 14263
rect 4997 14229 5031 14263
rect 6653 14229 6687 14263
rect 10057 14229 10091 14263
rect 19073 14229 19107 14263
rect 2605 14025 2639 14059
rect 2881 14025 2915 14059
rect 3617 14025 3651 14059
rect 4721 14025 4755 14059
rect 6469 14025 6503 14059
rect 6561 14025 6595 14059
rect 9597 14025 9631 14059
rect 10333 14025 10367 14059
rect 11897 14025 11931 14059
rect 16129 14025 16163 14059
rect 16451 14025 16485 14059
rect 17877 14025 17911 14059
rect 20729 14025 20763 14059
rect 22201 14025 22235 14059
rect 2145 13957 2179 13991
rect 5089 13957 5123 13991
rect 6285 13957 6319 13991
rect 1593 13889 1627 13923
rect 3801 13889 3835 13923
rect 5800 13821 5834 13855
rect 11345 13957 11379 13991
rect 12173 13957 12207 13991
rect 13645 13957 13679 13991
rect 15853 13957 15887 13991
rect 6837 13889 6871 13923
rect 9965 13889 9999 13923
rect 12817 13889 12851 13923
rect 15485 13889 15519 13923
rect 19073 13889 19107 13923
rect 20361 13889 20395 13923
rect 21281 13889 21315 13923
rect 10425 13821 10459 13855
rect 14749 13821 14783 13855
rect 15209 13821 15243 13855
rect 16380 13821 16414 13855
rect 16865 13821 16899 13855
rect 18096 13821 18130 13855
rect 18521 13821 18555 13855
rect 1685 13753 1719 13787
rect 3893 13753 3927 13787
rect 4445 13753 4479 13787
rect 6469 13753 6503 13787
rect 7158 13753 7192 13787
rect 10787 13753 10821 13787
rect 12541 13753 12575 13787
rect 12633 13753 12667 13787
rect 20913 13753 20947 13787
rect 21005 13753 21039 13787
rect 21833 13753 21867 13787
rect 5871 13685 5905 13719
rect 7757 13685 7791 13719
rect 8033 13685 8067 13719
rect 8677 13685 8711 13719
rect 14013 13685 14047 13719
rect 14565 13685 14599 13719
rect 17509 13685 17543 13719
rect 18199 13685 18233 13719
rect 18889 13685 18923 13719
rect 19441 13685 19475 13719
rect 19993 13685 20027 13719
rect 2329 13481 2363 13515
rect 2605 13481 2639 13515
rect 3801 13481 3835 13515
rect 6055 13481 6089 13515
rect 6745 13481 6779 13515
rect 12817 13481 12851 13515
rect 14749 13481 14783 13515
rect 18521 13481 18555 13515
rect 19441 13481 19475 13515
rect 19993 13481 20027 13515
rect 1771 13413 1805 13447
rect 4537 13413 4571 13447
rect 7113 13413 7147 13447
rect 10425 13413 10459 13447
rect 10701 13413 10735 13447
rect 12035 13413 12069 13447
rect 16037 13413 16071 13447
rect 21097 13413 21131 13447
rect 5984 13345 6018 13379
rect 9689 13345 9723 13379
rect 10149 13345 10183 13379
rect 11897 13345 11931 13379
rect 13737 13345 13771 13379
rect 14197 13345 14231 13379
rect 17509 13345 17543 13379
rect 18061 13345 18095 13379
rect 1409 13277 1443 13311
rect 4445 13277 4479 13311
rect 4721 13277 4755 13311
rect 7021 13277 7055 13311
rect 7297 13277 7331 13311
rect 14289 13277 14323 13311
rect 15945 13277 15979 13311
rect 18245 13277 18279 13311
rect 19073 13277 19107 13311
rect 21005 13277 21039 13311
rect 21281 13277 21315 13311
rect 16497 13209 16531 13243
rect 6469 13141 6503 13175
rect 8677 13141 8711 13175
rect 12449 13141 12483 13175
rect 16865 13141 16899 13175
rect 20637 13141 20671 13175
rect 3617 12937 3651 12971
rect 5089 12937 5123 12971
rect 6469 12937 6503 12971
rect 11345 12937 11379 12971
rect 12587 12937 12621 12971
rect 15209 12937 15243 12971
rect 15577 12937 15611 12971
rect 15945 12937 15979 12971
rect 20913 12937 20947 12971
rect 21925 12937 21959 12971
rect 4721 12869 4755 12903
rect 7481 12869 7515 12903
rect 11897 12869 11931 12903
rect 13277 12869 13311 12903
rect 17417 12869 17451 12903
rect 17785 12869 17819 12903
rect 21465 12869 21499 12903
rect 2145 12801 2179 12835
rect 2789 12801 2823 12835
rect 4169 12801 4203 12835
rect 5457 12801 5491 12835
rect 5779 12801 5813 12835
rect 6929 12801 6963 12835
rect 8493 12801 8527 12835
rect 14289 12801 14323 12835
rect 16129 12801 16163 12835
rect 18797 12801 18831 12835
rect 1685 12733 1719 12767
rect 1961 12733 1995 12767
rect 3132 12733 3166 12767
rect 5641 12733 5675 12767
rect 8677 12733 8711 12767
rect 9045 12733 9079 12767
rect 10149 12733 10183 12767
rect 10609 12733 10643 12767
rect 10793 12733 10827 12767
rect 12484 12733 12518 12767
rect 12909 12733 12943 12767
rect 18061 12733 18095 12767
rect 18521 12733 18555 12767
rect 21281 12733 21315 12767
rect 3985 12665 4019 12699
rect 4261 12665 4295 12699
rect 7021 12665 7055 12699
rect 11069 12665 11103 12699
rect 16221 12665 16255 12699
rect 16773 12665 16807 12699
rect 19809 12665 19843 12699
rect 19901 12665 19935 12699
rect 20453 12665 20487 12699
rect 2513 12597 2547 12631
rect 3203 12597 3237 12631
rect 6193 12597 6227 12631
rect 7849 12597 7883 12631
rect 8861 12597 8895 12631
rect 9689 12597 9723 12631
rect 13737 12597 13771 12631
rect 14197 12597 14231 12631
rect 14657 12597 14691 12631
rect 17141 12597 17175 12631
rect 19073 12597 19107 12631
rect 19625 12597 19659 12631
rect 1409 12393 1443 12427
rect 2237 12393 2271 12427
rect 3893 12393 3927 12427
rect 6285 12393 6319 12427
rect 7849 12393 7883 12427
rect 8447 12393 8481 12427
rect 8861 12393 8895 12427
rect 10793 12393 10827 12427
rect 14289 12393 14323 12427
rect 15945 12393 15979 12427
rect 19073 12393 19107 12427
rect 20269 12393 20303 12427
rect 21051 12393 21085 12427
rect 21373 12393 21407 12427
rect 1869 12325 1903 12359
rect 4261 12325 4295 12359
rect 6929 12325 6963 12359
rect 9873 12325 9907 12359
rect 11574 12325 11608 12359
rect 13185 12325 13219 12359
rect 16221 12325 16255 12359
rect 17785 12325 17819 12359
rect 19441 12325 19475 12359
rect 2421 12257 2455 12291
rect 2881 12257 2915 12291
rect 5784 12257 5818 12291
rect 8309 12257 8343 12291
rect 10425 12257 10459 12291
rect 16773 12257 16807 12291
rect 20948 12257 20982 12291
rect 3157 12189 3191 12223
rect 4169 12189 4203 12223
rect 4629 12189 4663 12223
rect 5871 12189 5905 12223
rect 6837 12189 6871 12223
rect 7113 12189 7147 12223
rect 9781 12189 9815 12223
rect 11253 12189 11287 12223
rect 13093 12189 13127 12223
rect 16129 12189 16163 12223
rect 17693 12189 17727 12223
rect 17969 12189 18003 12223
rect 19349 12189 19383 12223
rect 13645 12121 13679 12155
rect 19901 12121 19935 12155
rect 5273 12053 5307 12087
rect 6561 12053 6595 12087
rect 12173 12053 12207 12087
rect 12541 12053 12575 12087
rect 18613 12053 18647 12087
rect 2973 11849 3007 11883
rect 4077 11849 4111 11883
rect 4353 11849 4387 11883
rect 6469 11849 6503 11883
rect 6561 11849 6595 11883
rect 7757 11849 7791 11883
rect 9597 11849 9631 11883
rect 9873 11849 9907 11883
rect 10241 11849 10275 11883
rect 11805 11849 11839 11883
rect 12173 11849 12207 11883
rect 14657 11849 14691 11883
rect 16405 11849 16439 11883
rect 16727 11849 16761 11883
rect 17693 11849 17727 11883
rect 19441 11849 19475 11883
rect 19717 11849 19751 11883
rect 20085 11849 20119 11883
rect 20407 11849 20441 11883
rect 21097 11849 21131 11883
rect 6285 11781 6319 11815
rect 3157 11713 3191 11747
rect 5917 11713 5951 11747
rect 1409 11645 1443 11679
rect 2053 11645 2087 11679
rect 5457 11645 5491 11679
rect 5733 11645 5767 11679
rect 2513 11577 2547 11611
rect 3519 11577 3553 11611
rect 5089 11577 5123 11611
rect 15761 11781 15795 11815
rect 6837 11713 6871 11747
rect 8677 11713 8711 11747
rect 12817 11713 12851 11747
rect 16129 11713 16163 11747
rect 10517 11645 10551 11679
rect 10885 11645 10919 11679
rect 14841 11645 14875 11679
rect 16624 11645 16658 11679
rect 17049 11645 17083 11679
rect 18521 11645 18555 11679
rect 20336 11645 20370 11679
rect 20729 11645 20763 11679
rect 1593 11509 1627 11543
rect 6469 11509 6503 11543
rect 8998 11577 9032 11611
rect 11161 11577 11195 11611
rect 12541 11577 12575 11611
rect 12633 11577 12667 11611
rect 15162 11577 15196 11611
rect 18337 11577 18371 11611
rect 18842 11577 18876 11611
rect 7205 11509 7239 11543
rect 8401 11509 8435 11543
rect 11437 11509 11471 11543
rect 13461 11509 13495 11543
rect 13829 11509 13863 11543
rect 3433 11305 3467 11339
rect 4629 11305 4663 11339
rect 6285 11305 6319 11339
rect 7389 11305 7423 11339
rect 8677 11305 8711 11339
rect 9505 11305 9539 11339
rect 9689 11305 9723 11339
rect 12173 11305 12207 11339
rect 17601 11305 17635 11339
rect 4997 11237 5031 11271
rect 11574 11237 11608 11271
rect 14381 11237 14415 11271
rect 14841 11237 14875 11271
rect 18429 11237 18463 11271
rect 2697 11169 2731 11203
rect 2973 11169 3007 11203
rect 6377 11169 6411 11203
rect 6837 11169 6871 11203
rect 8008 11169 8042 11203
rect 11253 11169 11287 11203
rect 13645 11169 13679 11203
rect 14197 11169 14231 11203
rect 15368 11169 15402 11203
rect 16348 11169 16382 11203
rect 17693 11169 17727 11203
rect 18153 11169 18187 11203
rect 19416 11169 19450 11203
rect 1409 11101 1443 11135
rect 3157 11101 3191 11135
rect 4905 11101 4939 11135
rect 6929 11101 6963 11135
rect 5457 11033 5491 11067
rect 15439 11033 15473 11067
rect 1869 10965 1903 10999
rect 2329 10965 2363 10999
rect 4261 10965 4295 10999
rect 7757 10965 7791 10999
rect 8079 10965 8113 10999
rect 10517 10965 10551 10999
rect 12449 10965 12483 10999
rect 16451 10965 16485 10999
rect 19487 10965 19521 10999
rect 19809 10965 19843 10999
rect 3387 10761 3421 10795
rect 3985 10761 4019 10795
rect 4077 10761 4111 10795
rect 5181 10761 5215 10795
rect 5457 10761 5491 10795
rect 8125 10761 8159 10795
rect 9229 10761 9263 10795
rect 10885 10761 10919 10795
rect 11897 10761 11931 10795
rect 17141 10761 17175 10795
rect 18199 10761 18233 10795
rect 19441 10761 19475 10795
rect 21281 10761 21315 10795
rect 2789 10693 2823 10727
rect 1777 10625 1811 10659
rect 2421 10557 2455 10591
rect 3284 10557 3318 10591
rect 3709 10557 3743 10591
rect 6377 10693 6411 10727
rect 4261 10625 4295 10659
rect 7481 10625 7515 10659
rect 12817 10625 12851 10659
rect 17693 10625 17727 10659
rect 19625 10625 19659 10659
rect 19901 10625 19935 10659
rect 9321 10557 9355 10591
rect 9873 10557 9907 10591
rect 11412 10557 11446 10591
rect 14105 10557 14139 10591
rect 14749 10557 14783 10591
rect 15025 10557 15059 10591
rect 16380 10557 16414 10591
rect 18096 10557 18130 10591
rect 18521 10557 18555 10591
rect 21097 10557 21131 10591
rect 21649 10557 21683 10591
rect 1869 10489 1903 10523
rect 3985 10489 4019 10523
rect 4582 10489 4616 10523
rect 7205 10489 7239 10523
rect 7297 10489 7331 10523
rect 10057 10489 10091 10523
rect 12541 10489 12575 10523
rect 12633 10489 12667 10523
rect 14473 10489 14507 10523
rect 15301 10489 15335 10523
rect 15669 10489 15703 10523
rect 18889 10489 18923 10523
rect 19717 10489 19751 10523
rect 3065 10421 3099 10455
rect 6009 10421 6043 10455
rect 11161 10421 11195 10455
rect 11483 10421 11517 10455
rect 12173 10421 12207 10455
rect 13645 10421 13679 10455
rect 16451 10421 16485 10455
rect 16865 10421 16899 10455
rect 1869 10217 1903 10251
rect 2421 10217 2455 10251
rect 2697 10217 2731 10251
rect 4445 10217 4479 10251
rect 5273 10217 5307 10251
rect 7665 10217 7699 10251
rect 15761 10217 15795 10251
rect 19901 10217 19935 10251
rect 7066 10149 7100 10183
rect 7941 10149 7975 10183
rect 10378 10149 10412 10183
rect 12173 10149 12207 10183
rect 12265 10149 12299 10183
rect 13737 10149 13771 10183
rect 13829 10149 13863 10183
rect 17325 10149 17359 10183
rect 19026 10149 19060 10183
rect 4077 10081 4111 10115
rect 6745 10081 6779 10115
rect 8636 10081 8670 10115
rect 10057 10081 10091 10115
rect 19625 10081 19659 10115
rect 20948 10081 20982 10115
rect 1501 10013 1535 10047
rect 8723 10013 8757 10047
rect 12817 10013 12851 10047
rect 14013 10013 14047 10047
rect 15393 10013 15427 10047
rect 17233 10013 17267 10047
rect 18705 10013 18739 10047
rect 13461 9945 13495 9979
rect 17785 9945 17819 9979
rect 4997 9877 5031 9911
rect 9321 9877 9355 9911
rect 9873 9877 9907 9911
rect 10977 9877 11011 9911
rect 16313 9877 16347 9911
rect 18153 9877 18187 9911
rect 21051 9877 21085 9911
rect 2605 9673 2639 9707
rect 3709 9673 3743 9707
rect 4169 9673 4203 9707
rect 5457 9673 5491 9707
rect 11713 9673 11747 9707
rect 12081 9673 12115 9707
rect 14381 9673 14415 9707
rect 15853 9673 15887 9707
rect 16313 9673 16347 9707
rect 17417 9673 17451 9707
rect 19073 9673 19107 9707
rect 19533 9673 19567 9707
rect 20913 9673 20947 9707
rect 7113 9605 7147 9639
rect 10793 9605 10827 9639
rect 13645 9605 13679 9639
rect 21373 9605 21407 9639
rect 2329 9537 2363 9571
rect 3341 9537 3375 9571
rect 4445 9537 4479 9571
rect 5089 9537 5123 9571
rect 7389 9537 7423 9571
rect 8999 9537 9033 9571
rect 12817 9537 12851 9571
rect 16497 9537 16531 9571
rect 19717 9537 19751 9571
rect 21741 9537 21775 9571
rect 1685 9469 1719 9503
rect 2145 9469 2179 9503
rect 8912 9469 8946 9503
rect 9873 9469 9907 9503
rect 11069 9469 11103 9503
rect 14473 9469 14507 9503
rect 14933 9469 14967 9503
rect 18061 9469 18095 9503
rect 18521 9469 18555 9503
rect 21189 9469 21223 9503
rect 2973 9401 3007 9435
rect 4537 9401 4571 9435
rect 6653 9401 6687 9435
rect 7481 9401 7515 9435
rect 8033 9401 8067 9435
rect 9413 9401 9447 9435
rect 9781 9401 9815 9435
rect 10235 9401 10269 9435
rect 12541 9401 12575 9435
rect 12633 9401 12667 9435
rect 15209 9401 15243 9435
rect 16589 9401 16623 9435
rect 17141 9401 17175 9435
rect 18797 9401 18831 9435
rect 19809 9401 19843 9435
rect 20361 9401 20395 9435
rect 8677 9333 8711 9367
rect 15577 9333 15611 9367
rect 17785 9333 17819 9367
rect 4353 9129 4387 9163
rect 6837 9129 6871 9163
rect 8033 9129 8067 9163
rect 9965 9129 9999 9163
rect 11897 9129 11931 9163
rect 13093 9129 13127 9163
rect 14105 9129 14139 9163
rect 14473 9129 14507 9163
rect 16497 9129 16531 9163
rect 17601 9129 17635 9163
rect 19165 9129 19199 9163
rect 20085 9129 20119 9163
rect 20269 9129 20303 9163
rect 1869 9061 1903 9095
rect 3157 9061 3191 9095
rect 4721 9061 4755 9095
rect 7205 9061 7239 9095
rect 9505 9061 9539 9095
rect 12265 9061 12299 9095
rect 12817 9061 12851 9095
rect 13783 9061 13817 9095
rect 16773 9061 16807 9095
rect 21097 9061 21131 9095
rect 1444 8993 1478 9027
rect 1547 8993 1581 9027
rect 2697 8993 2731 9027
rect 2881 8993 2915 9027
rect 9965 8993 9999 9027
rect 10241 8993 10275 9027
rect 13645 8993 13679 9027
rect 15612 8993 15646 9027
rect 18153 8993 18187 9027
rect 18613 8993 18647 9027
rect 19876 8993 19910 9027
rect 2329 8925 2363 8959
rect 4629 8925 4663 8959
rect 4905 8925 4939 8959
rect 7113 8925 7147 8959
rect 7389 8925 7423 8959
rect 12173 8925 12207 8959
rect 15715 8925 15749 8959
rect 16681 8925 16715 8959
rect 18889 8925 18923 8959
rect 19533 8925 19567 8959
rect 21005 8925 21039 8959
rect 21281 8925 21315 8959
rect 16037 8857 16071 8891
rect 17233 8857 17267 8891
rect 10701 8789 10735 8823
rect 2513 8585 2547 8619
rect 2789 8585 2823 8619
rect 6285 8585 6319 8619
rect 9183 8585 9217 8619
rect 10057 8585 10091 8619
rect 11897 8585 11931 8619
rect 12265 8585 12299 8619
rect 16221 8585 16255 8619
rect 16681 8585 16715 8619
rect 16957 8585 16991 8619
rect 17877 8585 17911 8619
rect 19993 8585 20027 8619
rect 20361 8585 20395 8619
rect 22201 8585 22235 8619
rect 5089 8517 5123 8551
rect 8953 8517 8987 8551
rect 21833 8517 21867 8551
rect 3571 8449 3605 8483
rect 4537 8449 4571 8483
rect 5825 8449 5859 8483
rect 8033 8449 8067 8483
rect 12541 8449 12575 8483
rect 13185 8449 13219 8483
rect 15301 8449 15335 8483
rect 18797 8449 18831 8483
rect 18889 8449 18923 8483
rect 19073 8449 19107 8483
rect 21189 8449 21223 8483
rect 2053 8381 2087 8415
rect 3484 8381 3518 8415
rect 9080 8381 9114 8415
rect 9505 8381 9539 8415
rect 10333 8381 10367 8415
rect 10701 8381 10735 8415
rect 14080 8381 14114 8415
rect 14473 8381 14507 8415
rect 18096 8381 18130 8415
rect 18521 8381 18555 8415
rect 4353 8313 4387 8347
rect 4629 8313 4663 8347
rect 6653 8313 6687 8347
rect 7297 8313 7331 8347
rect 7573 8313 7607 8347
rect 7665 8313 7699 8347
rect 10977 8313 11011 8347
rect 12633 8313 12667 8347
rect 15663 8313 15697 8347
rect 19394 8313 19428 8347
rect 20913 8313 20947 8347
rect 21005 8313 21039 8347
rect 1685 8245 1719 8279
rect 3157 8245 3191 8279
rect 3985 8245 4019 8279
rect 5457 8245 5491 8279
rect 11345 8245 11379 8279
rect 13645 8245 13679 8279
rect 14151 8245 14185 8279
rect 15209 8245 15243 8279
rect 18199 8245 18233 8279
rect 18797 8245 18831 8279
rect 20637 8245 20671 8279
rect 2513 8041 2547 8075
rect 4445 8041 4479 8075
rect 4997 8041 5031 8075
rect 7389 8041 7423 8075
rect 7665 8041 7699 8075
rect 8355 8041 8389 8075
rect 10977 8041 11011 8075
rect 11989 8041 12023 8075
rect 12357 8041 12391 8075
rect 18153 8041 18187 8075
rect 19901 8041 19935 8075
rect 1593 7973 1627 8007
rect 6831 7973 6865 8007
rect 10241 7973 10275 8007
rect 11390 7973 11424 8007
rect 13369 7973 13403 8007
rect 16773 7973 16807 8007
rect 17325 7973 17359 8007
rect 19257 7973 19291 8007
rect 20177 7973 20211 8007
rect 21097 7973 21131 8007
rect 3040 7905 3074 7939
rect 8217 7905 8251 7939
rect 9689 7905 9723 7939
rect 9873 7905 9907 7939
rect 11069 7905 11103 7939
rect 12817 7905 12851 7939
rect 13001 7905 13035 7939
rect 14264 7905 14298 7939
rect 15209 7905 15243 7939
rect 1501 7837 1535 7871
rect 2145 7837 2179 7871
rect 4077 7837 4111 7871
rect 6469 7837 6503 7871
rect 16681 7837 16715 7871
rect 18981 7837 19015 7871
rect 21005 7837 21039 7871
rect 21281 7837 21315 7871
rect 15439 7769 15473 7803
rect 16129 7769 16163 7803
rect 2789 7701 2823 7735
rect 3111 7701 3145 7735
rect 3525 7701 3559 7735
rect 5273 7701 5307 7735
rect 6285 7701 6319 7735
rect 9505 7701 9539 7735
rect 10517 7701 10551 7735
rect 12633 7701 12667 7735
rect 13829 7701 13863 7735
rect 14335 7701 14369 7735
rect 15853 7701 15887 7735
rect 1685 7497 1719 7531
rect 3065 7497 3099 7531
rect 4445 7497 4479 7531
rect 6561 7497 6595 7531
rect 8861 7497 8895 7531
rect 9827 7497 9861 7531
rect 11483 7497 11517 7531
rect 13553 7497 13587 7531
rect 14749 7497 14783 7531
rect 16681 7497 16715 7531
rect 17049 7497 17083 7531
rect 20269 7497 20303 7531
rect 20913 7497 20947 7531
rect 21557 7497 21591 7531
rect 2421 7429 2455 7463
rect 9965 7429 9999 7463
rect 10333 7429 10367 7463
rect 14381 7429 14415 7463
rect 1869 7361 1903 7395
rect 5917 7361 5951 7395
rect 10057 7361 10091 7395
rect 11897 7361 11931 7395
rect 13829 7361 13863 7395
rect 15669 7361 15703 7395
rect 15945 7361 15979 7395
rect 20545 7361 20579 7395
rect 21097 7361 21131 7395
rect 3525 7293 3559 7327
rect 3801 7293 3835 7327
rect 4077 7293 4111 7327
rect 5457 7293 5491 7327
rect 5733 7293 5767 7327
rect 7113 7293 7147 7327
rect 7389 7293 7423 7327
rect 8309 7293 8343 7327
rect 11412 7293 11446 7327
rect 12776 7293 12810 7327
rect 13277 7293 13311 7327
rect 18096 7293 18130 7327
rect 18521 7293 18555 7327
rect 19349 7293 19383 7327
rect 1961 7225 1995 7259
rect 5089 7225 5123 7259
rect 7205 7225 7239 7259
rect 9137 7225 9171 7259
rect 9505 7225 9539 7259
rect 9689 7225 9723 7259
rect 12863 7225 12897 7259
rect 13921 7225 13955 7259
rect 15761 7225 15795 7259
rect 19670 7225 19704 7259
rect 7481 7157 7515 7191
rect 10701 7157 10735 7191
rect 11161 7157 11195 7191
rect 12173 7157 12207 7191
rect 15301 7157 15335 7191
rect 18199 7157 18233 7191
rect 19165 7157 19199 7191
rect 2881 6953 2915 6987
rect 3433 6953 3467 6987
rect 4721 6953 4755 6987
rect 8217 6953 8251 6987
rect 13553 6953 13587 6987
rect 13829 6953 13863 6987
rect 14197 6953 14231 6987
rect 19625 6953 19659 6987
rect 2047 6885 2081 6919
rect 4399 6885 4433 6919
rect 7573 6885 7607 6919
rect 8585 6885 8619 6919
rect 9873 6885 9907 6919
rect 10609 6885 10643 6919
rect 12995 6885 13029 6919
rect 15669 6885 15703 6919
rect 16221 6885 16255 6919
rect 18705 6885 18739 6919
rect 4312 6817 4346 6851
rect 5549 6817 5583 6851
rect 5825 6817 5859 6851
rect 7720 6817 7754 6851
rect 11253 6817 11287 6851
rect 17969 6817 18003 6851
rect 18521 6817 18555 6851
rect 1685 6749 1719 6783
rect 6009 6749 6043 6783
rect 7941 6749 7975 6783
rect 10020 6749 10054 6783
rect 10241 6749 10275 6783
rect 11529 6749 11563 6783
rect 12633 6749 12667 6783
rect 16129 6749 16163 6783
rect 16773 6749 16807 6783
rect 2605 6681 2639 6715
rect 5641 6681 5675 6715
rect 7297 6681 7331 6715
rect 10149 6681 10183 6715
rect 5273 6613 5307 6647
rect 6929 6613 6963 6647
rect 7849 6613 7883 6647
rect 9137 6613 9171 6647
rect 10977 6613 11011 6647
rect 11759 6613 11793 6647
rect 18981 6613 19015 6647
rect 20085 6613 20119 6647
rect 1961 6409 1995 6443
rect 4813 6409 4847 6443
rect 8033 6409 8067 6443
rect 9597 6409 9631 6443
rect 11713 6409 11747 6443
rect 16221 6409 16255 6443
rect 16497 6409 16531 6443
rect 17877 6409 17911 6443
rect 19441 6409 19475 6443
rect 7849 6341 7883 6375
rect 9413 6341 9447 6375
rect 10517 6341 10551 6375
rect 17049 6341 17083 6375
rect 3341 6273 3375 6307
rect 7941 6273 7975 6307
rect 9505 6273 9539 6307
rect 10149 6273 10183 6307
rect 13737 6273 13771 6307
rect 14381 6273 14415 6307
rect 17509 6273 17543 6307
rect 20177 6273 20211 6307
rect 1476 6205 1510 6239
rect 3709 6205 3743 6239
rect 3985 6205 4019 6239
rect 4261 6205 4295 6239
rect 7113 6205 7147 6239
rect 7481 6205 7515 6239
rect 7720 6205 7754 6239
rect 9045 6205 9079 6239
rect 9284 6205 9318 6239
rect 10793 6205 10827 6239
rect 12668 6205 12702 6239
rect 13093 6205 13127 6239
rect 14841 6205 14875 6239
rect 15301 6205 15335 6239
rect 18061 6205 18095 6239
rect 18521 6205 18555 6239
rect 19625 6205 19659 6239
rect 20085 6205 20119 6239
rect 2973 6137 3007 6171
rect 7573 6137 7607 6171
rect 9137 6137 9171 6171
rect 12771 6137 12805 6171
rect 13829 6137 13863 6171
rect 15622 6137 15656 6171
rect 1547 6069 1581 6103
rect 2329 6069 2363 6103
rect 3525 6069 3559 6103
rect 5549 6069 5583 6103
rect 5917 6069 5951 6103
rect 6285 6069 6319 6103
rect 8585 6069 8619 6103
rect 10977 6069 11011 6103
rect 12265 6069 12299 6103
rect 13553 6069 13587 6103
rect 15117 6069 15151 6103
rect 18153 6069 18187 6103
rect 4169 5865 4203 5899
rect 7849 5865 7883 5899
rect 11069 5865 11103 5899
rect 14197 5865 14231 5899
rect 15853 5865 15887 5899
rect 18521 5865 18555 5899
rect 1961 5797 1995 5831
rect 10425 5797 10459 5831
rect 12357 5797 12391 5831
rect 13369 5797 13403 5831
rect 13921 5797 13955 5831
rect 17693 5797 17727 5831
rect 3525 5729 3559 5763
rect 4353 5729 4387 5763
rect 4905 5729 4939 5763
rect 5549 5729 5583 5763
rect 6009 5729 6043 5763
rect 6101 5729 6135 5763
rect 6285 5729 6319 5763
rect 6745 5729 6779 5763
rect 7573 5729 7607 5763
rect 7757 5729 7791 5763
rect 9689 5729 9723 5763
rect 9965 5729 9999 5763
rect 10701 5729 10735 5763
rect 11621 5729 11655 5763
rect 12081 5729 12115 5763
rect 15945 5729 15979 5763
rect 16497 5729 16531 5763
rect 1685 5661 1719 5695
rect 1869 5661 1903 5695
rect 2237 5661 2271 5695
rect 2789 5661 2823 5695
rect 4813 5661 4847 5695
rect 11437 5661 11471 5695
rect 13277 5661 13311 5695
rect 16681 5661 16715 5695
rect 17601 5661 17635 5695
rect 17877 5661 17911 5695
rect 19349 5661 19383 5695
rect 9781 5593 9815 5627
rect 5825 5525 5859 5559
rect 7021 5525 7055 5559
rect 7481 5525 7515 5559
rect 8401 5525 8435 5559
rect 9137 5525 9171 5559
rect 12633 5525 12667 5559
rect 16957 5525 16991 5559
rect 2881 5321 2915 5355
rect 3249 5321 3283 5355
rect 4169 5321 4203 5355
rect 4537 5321 4571 5355
rect 6193 5321 6227 5355
rect 8585 5321 8619 5355
rect 8953 5321 8987 5355
rect 9321 5321 9355 5355
rect 10977 5321 11011 5355
rect 11621 5321 11655 5355
rect 13461 5321 13495 5355
rect 13737 5321 13771 5355
rect 14105 5321 14139 5355
rect 15669 5321 15703 5355
rect 16037 5321 16071 5355
rect 19625 5321 19659 5355
rect 1869 5253 1903 5287
rect 5273 5253 5307 5287
rect 9597 5253 9631 5287
rect 12173 5253 12207 5287
rect 12449 5253 12483 5287
rect 14933 5253 14967 5287
rect 17509 5253 17543 5287
rect 18981 5253 19015 5287
rect 1961 5185 1995 5219
rect 10241 5185 10275 5219
rect 5181 5117 5215 5151
rect 5457 5117 5491 5151
rect 6837 5117 6871 5151
rect 7021 5117 7055 5151
rect 9505 5117 9539 5151
rect 9781 5117 9815 5151
rect 11136 5117 11170 5151
rect 12541 5185 12575 5219
rect 14381 5185 14415 5219
rect 16313 5185 16347 5219
rect 18061 5185 18095 5219
rect 19901 5185 19935 5219
rect 16957 5117 16991 5151
rect 2282 5049 2316 5083
rect 3801 5049 3835 5083
rect 6561 5049 6595 5083
rect 8217 5049 8251 5083
rect 10517 5049 10551 5083
rect 12449 5049 12483 5083
rect 12862 5049 12896 5083
rect 14473 5049 14507 5083
rect 16405 5049 16439 5083
rect 18382 5049 18416 5083
rect 19993 5049 20027 5083
rect 20545 5049 20579 5083
rect 4997 4981 5031 5015
rect 5641 4981 5675 5015
rect 7941 4981 7975 5015
rect 11207 4981 11241 5015
rect 17785 4981 17819 5015
rect 2421 4777 2455 4811
rect 5273 4777 5307 4811
rect 9505 4777 9539 4811
rect 13185 4777 13219 4811
rect 14381 4777 14415 4811
rect 15853 4777 15887 4811
rect 16405 4777 16439 4811
rect 16681 4777 16715 4811
rect 17601 4777 17635 4811
rect 18061 4777 18095 4811
rect 18981 4777 19015 4811
rect 19533 4777 19567 4811
rect 19901 4777 19935 4811
rect 1593 4709 1627 4743
rect 2145 4709 2179 4743
rect 9689 4709 9723 4743
rect 12633 4709 12667 4743
rect 4169 4641 4203 4675
rect 4353 4641 4387 4675
rect 4721 4641 4755 4675
rect 5549 4641 5583 4675
rect 5825 4641 5859 4675
rect 6653 4641 6687 4675
rect 7113 4641 7147 4675
rect 7389 4641 7423 4675
rect 8125 4641 8159 4675
rect 9781 4641 9815 4675
rect 11897 4641 11931 4675
rect 12449 4641 12483 4675
rect 13461 4641 13495 4675
rect 13645 4641 13679 4675
rect 1501 4573 1535 4607
rect 2973 4573 3007 4607
rect 6009 4573 6043 4607
rect 7757 4573 7791 4607
rect 11713 4573 11747 4607
rect 13921 4573 13955 4607
rect 15485 4573 15519 4607
rect 18613 4573 18647 4607
rect 5641 4505 5675 4539
rect 7205 4505 7239 4539
rect 2605 4233 2639 4267
rect 3893 4233 3927 4267
rect 6653 4233 6687 4267
rect 7205 4233 7239 4267
rect 7849 4233 7883 4267
rect 11989 4233 12023 4267
rect 13461 4233 13495 4267
rect 13829 4233 13863 4267
rect 15945 4233 15979 4267
rect 17785 4233 17819 4267
rect 19073 4233 19107 4267
rect 4813 4165 4847 4199
rect 11621 4165 11655 4199
rect 5273 4097 5307 4131
rect 9781 4097 9815 4131
rect 14841 4097 14875 4131
rect 2237 4029 2271 4063
rect 4537 4029 4571 4063
rect 4721 4029 4755 4063
rect 4997 4029 5031 4063
rect 7941 4029 7975 4063
rect 8401 4029 8435 4063
rect 8769 4029 8803 4063
rect 9413 4029 9447 4063
rect 10149 4029 10183 4063
rect 12725 4029 12759 4063
rect 15025 4029 15059 4063
rect 15393 4029 15427 4063
rect 18337 4029 18371 4063
rect 18521 4029 18555 4063
rect 20948 4029 20982 4063
rect 21373 4029 21407 4063
rect 1593 3961 1627 3995
rect 6101 3961 6135 3995
rect 12449 3961 12483 3995
rect 15669 3961 15703 3995
rect 16313 3961 16347 3995
rect 18797 3961 18831 3995
rect 19533 3961 19567 3995
rect 21051 3961 21085 3995
rect 3433 3893 3467 3927
rect 4169 3893 4203 3927
rect 5733 3893 5767 3927
rect 8861 3893 8895 3927
rect 10517 3893 10551 3927
rect 1593 3689 1627 3723
rect 1961 3689 1995 3723
rect 5181 3689 5215 3723
rect 5641 3689 5675 3723
rect 7113 3689 7147 3723
rect 8401 3689 8435 3723
rect 11161 3689 11195 3723
rect 12725 3689 12759 3723
rect 13461 3689 13495 3723
rect 15025 3689 15059 3723
rect 18153 3689 18187 3723
rect 4813 3621 4847 3655
rect 10286 3621 10320 3655
rect 11897 3621 11931 3655
rect 4261 3553 4295 3587
rect 5917 3553 5951 3587
rect 6561 3553 6595 3587
rect 7573 3553 7607 3587
rect 8125 3553 8159 3587
rect 10885 3553 10919 3587
rect 13312 3553 13346 3587
rect 9965 3485 9999 3519
rect 11805 3485 11839 3519
rect 12449 3485 12483 3519
rect 7481 3417 7515 3451
rect 5181 3145 5215 3179
rect 5825 3145 5859 3179
rect 6653 3145 6687 3179
rect 9229 3145 9263 3179
rect 11529 3145 11563 3179
rect 12265 3145 12299 3179
rect 13461 3145 13495 3179
rect 7481 3077 7515 3111
rect 13093 3077 13127 3111
rect 13829 3077 13863 3111
rect 8401 3009 8435 3043
rect 10517 3009 10551 3043
rect 11161 3009 11195 3043
rect 11897 3009 11931 3043
rect 12541 3009 12575 3043
rect 14013 3009 14047 3043
rect 4629 2941 4663 2975
rect 5365 2941 5399 2975
rect 7941 2941 7975 2975
rect 8493 2941 8527 2975
rect 7205 2873 7239 2907
rect 9689 2873 9723 2907
rect 10609 2873 10643 2907
rect 12633 2873 12667 2907
rect 4169 2805 4203 2839
rect 8769 2805 8803 2839
rect 9965 2805 9999 2839
rect 6377 2601 6411 2635
rect 7941 2601 7975 2635
rect 8401 2601 8435 2635
rect 9597 2601 9631 2635
rect 10701 2601 10735 2635
rect 12357 2601 12391 2635
rect 6929 2533 6963 2567
rect 10102 2533 10136 2567
rect 12817 2533 12851 2567
rect 13369 2533 13403 2567
rect 5733 2465 5767 2499
rect 7021 2465 7055 2499
rect 8585 2465 8619 2499
rect 9137 2465 9171 2499
rect 9781 2465 9815 2499
rect 10977 2465 11011 2499
rect 11564 2465 11598 2499
rect 11989 2465 12023 2499
rect 14197 2465 14231 2499
rect 17141 2465 17175 2499
rect 17693 2465 17727 2499
rect 11667 2397 11701 2431
rect 12725 2397 12759 2431
rect 13645 2397 13679 2431
rect 6653 2329 6687 2363
rect 8769 2329 8803 2363
rect 17325 2329 17359 2363
rect 5917 2261 5951 2295
rect 14381 2261 14415 2295
rect 14841 2261 14875 2295
<< metal1 >>
rect 1104 21786 22816 21808
rect 1104 21734 4982 21786
rect 5034 21734 5046 21786
rect 5098 21734 5110 21786
rect 5162 21734 5174 21786
rect 5226 21734 12982 21786
rect 13034 21734 13046 21786
rect 13098 21734 13110 21786
rect 13162 21734 13174 21786
rect 13226 21734 20982 21786
rect 21034 21734 21046 21786
rect 21098 21734 21110 21786
rect 21162 21734 21174 21786
rect 21226 21734 22816 21786
rect 1104 21712 22816 21734
rect 1104 21242 22816 21264
rect 1104 21190 8982 21242
rect 9034 21190 9046 21242
rect 9098 21190 9110 21242
rect 9162 21190 9174 21242
rect 9226 21190 16982 21242
rect 17034 21190 17046 21242
rect 17098 21190 17110 21242
rect 17162 21190 17174 21242
rect 17226 21190 22816 21242
rect 1104 21168 22816 21190
rect 1104 20698 22816 20720
rect 1104 20646 4982 20698
rect 5034 20646 5046 20698
rect 5098 20646 5110 20698
rect 5162 20646 5174 20698
rect 5226 20646 12982 20698
rect 13034 20646 13046 20698
rect 13098 20646 13110 20698
rect 13162 20646 13174 20698
rect 13226 20646 20982 20698
rect 21034 20646 21046 20698
rect 21098 20646 21110 20698
rect 21162 20646 21174 20698
rect 21226 20646 22816 20698
rect 1104 20624 22816 20646
rect 5813 20587 5871 20593
rect 5813 20553 5825 20587
rect 5859 20584 5871 20587
rect 7006 20584 7012 20596
rect 5859 20556 7012 20584
rect 5859 20553 5871 20556
rect 5813 20547 5871 20553
rect 7006 20544 7012 20556
rect 7064 20544 7070 20596
rect 8113 20587 8171 20593
rect 8113 20553 8125 20587
rect 8159 20584 8171 20587
rect 8662 20584 8668 20596
rect 8159 20556 8668 20584
rect 8159 20553 8171 20556
rect 8113 20547 8171 20553
rect 8662 20544 8668 20556
rect 8720 20544 8726 20596
rect 10778 20544 10784 20596
rect 10836 20584 10842 20596
rect 10873 20587 10931 20593
rect 10873 20584 10885 20587
rect 10836 20556 10885 20584
rect 10836 20544 10842 20556
rect 10873 20553 10885 20556
rect 10919 20553 10931 20587
rect 10873 20547 10931 20553
rect 15289 20587 15347 20593
rect 15289 20553 15301 20587
rect 15335 20584 15347 20587
rect 16574 20584 16580 20596
rect 15335 20556 16580 20584
rect 15335 20553 15347 20556
rect 15289 20547 15347 20553
rect 16574 20544 16580 20556
rect 16632 20544 16638 20596
rect 19429 20587 19487 20593
rect 19429 20553 19441 20587
rect 19475 20584 19487 20587
rect 20622 20584 20628 20596
rect 19475 20556 20628 20584
rect 19475 20553 19487 20556
rect 19429 20547 19487 20553
rect 20622 20544 20628 20556
rect 20680 20544 20686 20596
rect 1302 20408 1308 20460
rect 1360 20448 1366 20460
rect 1535 20451 1593 20457
rect 1535 20448 1547 20451
rect 1360 20420 1547 20448
rect 1360 20408 1366 20420
rect 1535 20417 1547 20420
rect 1581 20417 1593 20451
rect 1535 20411 1593 20417
rect 1448 20383 1506 20389
rect 1448 20349 1460 20383
rect 1494 20380 1506 20383
rect 5626 20380 5632 20392
rect 1494 20352 1808 20380
rect 5587 20352 5632 20380
rect 1494 20349 1506 20352
rect 1448 20343 1506 20349
rect 1780 20256 1808 20352
rect 5626 20340 5632 20352
rect 5684 20380 5690 20392
rect 6181 20383 6239 20389
rect 6181 20380 6193 20383
rect 5684 20352 6193 20380
rect 5684 20340 5690 20352
rect 6181 20349 6193 20352
rect 6227 20349 6239 20383
rect 6181 20343 6239 20349
rect 7929 20383 7987 20389
rect 7929 20349 7941 20383
rect 7975 20380 7987 20383
rect 10689 20383 10747 20389
rect 7975 20352 8432 20380
rect 7975 20349 7987 20352
rect 7929 20343 7987 20349
rect 8404 20256 8432 20352
rect 10689 20349 10701 20383
rect 10735 20380 10747 20383
rect 15102 20380 15108 20392
rect 10735 20352 11376 20380
rect 15063 20352 15108 20380
rect 10735 20349 10747 20352
rect 10689 20343 10747 20349
rect 1762 20204 1768 20256
rect 1820 20244 1826 20256
rect 1857 20247 1915 20253
rect 1857 20244 1869 20247
rect 1820 20216 1869 20244
rect 1820 20204 1826 20216
rect 1857 20213 1869 20216
rect 1903 20213 1915 20247
rect 1857 20207 1915 20213
rect 8386 20204 8392 20256
rect 8444 20244 8450 20256
rect 11348 20253 11376 20352
rect 15102 20340 15108 20352
rect 15160 20380 15166 20392
rect 15657 20383 15715 20389
rect 15657 20380 15669 20383
rect 15160 20352 15669 20380
rect 15160 20340 15166 20352
rect 15657 20349 15669 20352
rect 15703 20349 15715 20383
rect 15657 20343 15715 20349
rect 18230 20340 18236 20392
rect 18288 20380 18294 20392
rect 19245 20383 19303 20389
rect 19245 20380 19257 20383
rect 18288 20352 19257 20380
rect 18288 20340 18294 20352
rect 19245 20349 19257 20352
rect 19291 20380 19303 20383
rect 19797 20383 19855 20389
rect 19797 20380 19809 20383
rect 19291 20352 19809 20380
rect 19291 20349 19303 20352
rect 19245 20343 19303 20349
rect 19797 20349 19809 20352
rect 19843 20349 19855 20383
rect 19797 20343 19855 20349
rect 8481 20247 8539 20253
rect 8481 20244 8493 20247
rect 8444 20216 8493 20244
rect 8444 20204 8450 20216
rect 8481 20213 8493 20216
rect 8527 20213 8539 20247
rect 8481 20207 8539 20213
rect 11333 20247 11391 20253
rect 11333 20213 11345 20247
rect 11379 20244 11391 20247
rect 11974 20244 11980 20256
rect 11379 20216 11980 20244
rect 11379 20213 11391 20216
rect 11333 20207 11391 20213
rect 11974 20204 11980 20216
rect 12032 20204 12038 20256
rect 1104 20154 22816 20176
rect 1104 20102 8982 20154
rect 9034 20102 9046 20154
rect 9098 20102 9110 20154
rect 9162 20102 9174 20154
rect 9226 20102 16982 20154
rect 17034 20102 17046 20154
rect 17098 20102 17110 20154
rect 17162 20102 17174 20154
rect 17226 20102 22816 20154
rect 1104 20080 22816 20102
rect 17313 20043 17371 20049
rect 17313 20009 17325 20043
rect 17359 20040 17371 20043
rect 18966 20040 18972 20052
rect 17359 20012 18972 20040
rect 17359 20009 17371 20012
rect 17313 20003 17371 20009
rect 18966 20000 18972 20012
rect 19024 20000 19030 20052
rect 9744 19907 9802 19913
rect 9744 19873 9756 19907
rect 9790 19904 9802 19907
rect 10226 19904 10232 19916
rect 9790 19876 10232 19904
rect 9790 19873 9802 19876
rect 9744 19867 9802 19873
rect 10226 19864 10232 19876
rect 10284 19864 10290 19916
rect 17129 19907 17187 19913
rect 17129 19873 17141 19907
rect 17175 19904 17187 19907
rect 17678 19904 17684 19916
rect 17175 19876 17684 19904
rect 17175 19873 17187 19876
rect 17129 19867 17187 19873
rect 17678 19864 17684 19876
rect 17736 19864 17742 19916
rect 1210 19660 1216 19712
rect 1268 19700 1274 19712
rect 9815 19703 9873 19709
rect 9815 19700 9827 19703
rect 1268 19672 9827 19700
rect 1268 19660 1274 19672
rect 9815 19669 9827 19672
rect 9861 19669 9873 19703
rect 10226 19700 10232 19712
rect 10187 19672 10232 19700
rect 9815 19663 9873 19669
rect 10226 19660 10232 19672
rect 10284 19660 10290 19712
rect 1104 19610 22816 19632
rect 1104 19558 4982 19610
rect 5034 19558 5046 19610
rect 5098 19558 5110 19610
rect 5162 19558 5174 19610
rect 5226 19558 12982 19610
rect 13034 19558 13046 19610
rect 13098 19558 13110 19610
rect 13162 19558 13174 19610
rect 13226 19558 20982 19610
rect 21034 19558 21046 19610
rect 21098 19558 21110 19610
rect 21162 19558 21174 19610
rect 21226 19558 22816 19610
rect 1104 19536 22816 19558
rect 21039 19499 21097 19505
rect 21039 19465 21051 19499
rect 21085 19496 21097 19499
rect 22646 19496 22652 19508
rect 21085 19468 22652 19496
rect 21085 19465 21097 19468
rect 21039 19459 21097 19465
rect 22646 19456 22652 19468
rect 22704 19456 22710 19508
rect 20806 19252 20812 19304
rect 20864 19292 20870 19304
rect 20936 19295 20994 19301
rect 20936 19292 20948 19295
rect 20864 19264 20948 19292
rect 20864 19252 20870 19264
rect 20936 19261 20948 19264
rect 20982 19292 20994 19295
rect 21361 19295 21419 19301
rect 21361 19292 21373 19295
rect 20982 19264 21373 19292
rect 20982 19261 20994 19264
rect 20936 19255 20994 19261
rect 21361 19261 21373 19264
rect 21407 19261 21419 19295
rect 21361 19255 21419 19261
rect 8849 19227 8907 19233
rect 8849 19193 8861 19227
rect 8895 19224 8907 19227
rect 9677 19227 9735 19233
rect 9677 19224 9689 19227
rect 8895 19196 9689 19224
rect 8895 19193 8907 19196
rect 8849 19187 8907 19193
rect 9677 19193 9689 19196
rect 9723 19224 9735 19227
rect 9953 19227 10011 19233
rect 9953 19224 9965 19227
rect 9723 19196 9965 19224
rect 9723 19193 9735 19196
rect 9677 19187 9735 19193
rect 9953 19193 9965 19196
rect 9999 19193 10011 19227
rect 9953 19187 10011 19193
rect 10045 19227 10103 19233
rect 10045 19193 10057 19227
rect 10091 19193 10103 19227
rect 10045 19187 10103 19193
rect 9401 19159 9459 19165
rect 9401 19125 9413 19159
rect 9447 19156 9459 19159
rect 10060 19156 10088 19187
rect 10226 19184 10232 19236
rect 10284 19224 10290 19236
rect 10597 19227 10655 19233
rect 10597 19224 10609 19227
rect 10284 19196 10609 19224
rect 10284 19184 10290 19196
rect 10597 19193 10609 19196
rect 10643 19224 10655 19227
rect 12802 19224 12808 19236
rect 10643 19196 12808 19224
rect 10643 19193 10655 19196
rect 10597 19187 10655 19193
rect 12802 19184 12808 19196
rect 12860 19184 12866 19236
rect 10502 19156 10508 19168
rect 9447 19128 10508 19156
rect 9447 19125 9459 19128
rect 9401 19119 9459 19125
rect 10502 19116 10508 19128
rect 10560 19116 10566 19168
rect 17221 19159 17279 19165
rect 17221 19125 17233 19159
rect 17267 19156 17279 19159
rect 17678 19156 17684 19168
rect 17267 19128 17684 19156
rect 17267 19125 17279 19128
rect 17221 19119 17279 19125
rect 17678 19116 17684 19128
rect 17736 19116 17742 19168
rect 1104 19066 22816 19088
rect 1104 19014 8982 19066
rect 9034 19014 9046 19066
rect 9098 19014 9110 19066
rect 9162 19014 9174 19066
rect 9226 19014 16982 19066
rect 17034 19014 17046 19066
rect 17098 19014 17110 19066
rect 17162 19014 17174 19066
rect 17226 19014 22816 19066
rect 1104 18992 22816 19014
rect 10502 18912 10508 18964
rect 10560 18952 10566 18964
rect 10597 18955 10655 18961
rect 10597 18952 10609 18955
rect 10560 18924 10609 18952
rect 10560 18912 10566 18924
rect 10597 18921 10609 18924
rect 10643 18921 10655 18955
rect 10597 18915 10655 18921
rect 11514 18912 11520 18964
rect 11572 18952 11578 18964
rect 11793 18955 11851 18961
rect 11793 18952 11805 18955
rect 11572 18924 11805 18952
rect 11572 18912 11578 18924
rect 11793 18921 11805 18924
rect 11839 18921 11851 18955
rect 11793 18915 11851 18921
rect 21085 18955 21143 18961
rect 21085 18921 21097 18955
rect 21131 18952 21143 18955
rect 21266 18952 21272 18964
rect 21131 18924 21272 18952
rect 21131 18921 21143 18924
rect 21085 18915 21143 18921
rect 21266 18912 21272 18924
rect 21324 18912 21330 18964
rect 1302 18844 1308 18896
rect 1360 18884 1366 18896
rect 1535 18887 1593 18893
rect 1535 18884 1547 18887
rect 1360 18856 1547 18884
rect 1360 18844 1366 18856
rect 1535 18853 1547 18856
rect 1581 18853 1593 18887
rect 7466 18884 7472 18896
rect 1535 18847 1593 18853
rect 6932 18856 7472 18884
rect 1448 18819 1506 18825
rect 1448 18785 1460 18819
rect 1494 18816 1506 18819
rect 1670 18816 1676 18828
rect 1494 18788 1676 18816
rect 1494 18785 1506 18788
rect 1448 18779 1506 18785
rect 1670 18776 1676 18788
rect 1728 18776 1734 18828
rect 6932 18825 6960 18856
rect 7466 18844 7472 18856
rect 7524 18844 7530 18896
rect 9766 18844 9772 18896
rect 9824 18884 9830 18896
rect 10039 18887 10097 18893
rect 10039 18884 10051 18887
rect 9824 18856 10051 18884
rect 9824 18844 9830 18856
rect 10039 18853 10051 18856
rect 10085 18884 10097 18887
rect 11532 18884 11560 18912
rect 10085 18856 11560 18884
rect 10085 18853 10097 18856
rect 10039 18847 10097 18853
rect 6917 18819 6975 18825
rect 6917 18785 6929 18819
rect 6963 18785 6975 18819
rect 7098 18816 7104 18828
rect 7059 18788 7104 18816
rect 6917 18779 6975 18785
rect 7098 18776 7104 18788
rect 7156 18776 7162 18828
rect 15194 18776 15200 18828
rect 15252 18816 15258 18828
rect 15324 18819 15382 18825
rect 15324 18816 15336 18819
rect 15252 18788 15336 18816
rect 15252 18776 15258 18788
rect 15324 18785 15336 18788
rect 15370 18785 15382 18819
rect 15324 18779 15382 18785
rect 16577 18819 16635 18825
rect 16577 18785 16589 18819
rect 16623 18785 16635 18819
rect 16577 18779 16635 18785
rect 7190 18748 7196 18760
rect 7151 18720 7196 18748
rect 7190 18708 7196 18720
rect 7248 18708 7254 18760
rect 9674 18748 9680 18760
rect 9635 18720 9680 18748
rect 9674 18708 9680 18720
rect 9732 18708 9738 18760
rect 11425 18751 11483 18757
rect 11425 18717 11437 18751
rect 11471 18748 11483 18751
rect 11790 18748 11796 18760
rect 11471 18720 11796 18748
rect 11471 18717 11483 18720
rect 11425 18711 11483 18717
rect 11790 18708 11796 18720
rect 11848 18708 11854 18760
rect 16592 18748 16620 18779
rect 16666 18776 16672 18828
rect 16724 18816 16730 18828
rect 17037 18819 17095 18825
rect 17037 18816 17049 18819
rect 16724 18788 17049 18816
rect 16724 18776 16730 18788
rect 17037 18785 17049 18788
rect 17083 18785 17095 18819
rect 17037 18779 17095 18785
rect 20901 18819 20959 18825
rect 20901 18785 20913 18819
rect 20947 18816 20959 18819
rect 21542 18816 21548 18828
rect 20947 18788 21548 18816
rect 20947 18785 20959 18788
rect 20901 18779 20959 18785
rect 21542 18776 21548 18788
rect 21600 18776 21606 18828
rect 16850 18748 16856 18760
rect 16592 18720 16856 18748
rect 16850 18708 16856 18720
rect 16908 18708 16914 18760
rect 17310 18748 17316 18760
rect 17271 18720 17316 18748
rect 17310 18708 17316 18720
rect 17368 18708 17374 18760
rect 19429 18751 19487 18757
rect 19429 18717 19441 18751
rect 19475 18748 19487 18751
rect 20346 18748 20352 18760
rect 19475 18720 20352 18748
rect 19475 18717 19487 18720
rect 19429 18711 19487 18717
rect 20346 18708 20352 18720
rect 20404 18708 20410 18760
rect 4798 18572 4804 18624
rect 4856 18612 4862 18624
rect 4893 18615 4951 18621
rect 4893 18612 4905 18615
rect 4856 18584 4905 18612
rect 4856 18572 4862 18584
rect 4893 18581 4905 18584
rect 4939 18581 4951 18615
rect 8294 18612 8300 18624
rect 8255 18584 8300 18612
rect 4893 18575 4951 18581
rect 8294 18572 8300 18584
rect 8352 18572 8358 18624
rect 12342 18612 12348 18624
rect 12303 18584 12348 18612
rect 12342 18572 12348 18584
rect 12400 18572 12406 18624
rect 12618 18612 12624 18624
rect 12579 18584 12624 18612
rect 12618 18572 12624 18584
rect 12676 18572 12682 18624
rect 15427 18615 15485 18621
rect 15427 18581 15439 18615
rect 15473 18612 15485 18615
rect 15562 18612 15568 18624
rect 15473 18584 15568 18612
rect 15473 18581 15485 18584
rect 15427 18575 15485 18581
rect 15562 18572 15568 18584
rect 15620 18572 15626 18624
rect 15746 18612 15752 18624
rect 15707 18584 15752 18612
rect 15746 18572 15752 18584
rect 15804 18572 15810 18624
rect 16114 18612 16120 18624
rect 16075 18584 16120 18612
rect 16114 18572 16120 18584
rect 16172 18572 16178 18624
rect 18782 18612 18788 18624
rect 18743 18584 18788 18612
rect 18782 18572 18788 18584
rect 18840 18572 18846 18624
rect 1104 18522 22816 18544
rect 1104 18470 4982 18522
rect 5034 18470 5046 18522
rect 5098 18470 5110 18522
rect 5162 18470 5174 18522
rect 5226 18470 12982 18522
rect 13034 18470 13046 18522
rect 13098 18470 13110 18522
rect 13162 18470 13174 18522
rect 13226 18470 20982 18522
rect 21034 18470 21046 18522
rect 21098 18470 21110 18522
rect 21162 18470 21174 18522
rect 21226 18470 22816 18522
rect 1104 18448 22816 18470
rect 2406 18368 2412 18420
rect 2464 18408 2470 18420
rect 7466 18408 7472 18420
rect 2464 18380 7472 18408
rect 2464 18368 2470 18380
rect 7466 18368 7472 18380
rect 7524 18368 7530 18420
rect 9677 18411 9735 18417
rect 9677 18377 9689 18411
rect 9723 18408 9735 18411
rect 9766 18408 9772 18420
rect 9723 18380 9772 18408
rect 9723 18377 9735 18380
rect 9677 18371 9735 18377
rect 9766 18368 9772 18380
rect 9824 18368 9830 18420
rect 11514 18408 11520 18420
rect 11475 18380 11520 18408
rect 11514 18368 11520 18380
rect 11572 18368 11578 18420
rect 12253 18411 12311 18417
rect 12253 18377 12265 18411
rect 12299 18408 12311 18411
rect 12342 18408 12348 18420
rect 12299 18380 12348 18408
rect 12299 18377 12311 18380
rect 12253 18371 12311 18377
rect 12342 18368 12348 18380
rect 12400 18368 12406 18420
rect 16850 18408 16856 18420
rect 13786 18380 16856 18408
rect 5534 18340 5540 18352
rect 4126 18312 5540 18340
rect 3418 18204 3424 18216
rect 3379 18176 3424 18204
rect 3418 18164 3424 18176
rect 3476 18164 3482 18216
rect 3881 18207 3939 18213
rect 3881 18173 3893 18207
rect 3927 18204 3939 18207
rect 4126 18204 4154 18312
rect 5534 18300 5540 18312
rect 5592 18340 5598 18352
rect 7009 18343 7067 18349
rect 7009 18340 7021 18343
rect 5592 18312 7021 18340
rect 5592 18300 5598 18312
rect 7009 18309 7021 18312
rect 7055 18340 7067 18343
rect 7098 18340 7104 18352
rect 7055 18312 7104 18340
rect 7055 18309 7067 18312
rect 7009 18303 7067 18309
rect 7098 18300 7104 18312
rect 7156 18300 7162 18352
rect 10870 18300 10876 18352
rect 10928 18340 10934 18352
rect 13786 18340 13814 18380
rect 16850 18368 16856 18380
rect 16908 18368 16914 18420
rect 20346 18408 20352 18420
rect 20307 18380 20352 18408
rect 20346 18368 20352 18380
rect 20404 18408 20410 18420
rect 20404 18380 20668 18408
rect 20404 18368 20410 18380
rect 10928 18312 13814 18340
rect 14323 18343 14381 18349
rect 10928 18300 10934 18312
rect 14323 18309 14335 18343
rect 14369 18340 14381 18343
rect 14369 18312 15424 18340
rect 14369 18309 14381 18312
rect 14323 18303 14381 18309
rect 4798 18232 4804 18284
rect 4856 18272 4862 18284
rect 4985 18275 5043 18281
rect 4985 18272 4997 18275
rect 4856 18244 4997 18272
rect 4856 18232 4862 18244
rect 4985 18241 4997 18244
rect 5031 18241 5043 18275
rect 5350 18272 5356 18284
rect 5311 18244 5356 18272
rect 4985 18235 5043 18241
rect 5350 18232 5356 18244
rect 5408 18232 5414 18284
rect 8570 18272 8576 18284
rect 8531 18244 8576 18272
rect 8570 18232 8576 18244
rect 8628 18232 8634 18284
rect 9674 18232 9680 18284
rect 9732 18272 9738 18284
rect 10505 18275 10563 18281
rect 10505 18272 10517 18275
rect 9732 18244 10517 18272
rect 9732 18232 9738 18244
rect 10505 18241 10517 18244
rect 10551 18272 10563 18275
rect 10781 18275 10839 18281
rect 10781 18272 10793 18275
rect 10551 18244 10793 18272
rect 10551 18241 10563 18244
rect 10505 18235 10563 18241
rect 10781 18241 10793 18244
rect 10827 18241 10839 18275
rect 10781 18235 10839 18241
rect 12529 18275 12587 18281
rect 12529 18241 12541 18275
rect 12575 18272 12587 18275
rect 12618 18272 12624 18284
rect 12575 18244 12624 18272
rect 12575 18241 12587 18244
rect 12529 18235 12587 18241
rect 12618 18232 12624 18244
rect 12676 18232 12682 18284
rect 12802 18272 12808 18284
rect 12763 18244 12808 18272
rect 12802 18232 12808 18244
rect 12860 18232 12866 18284
rect 15396 18281 15424 18312
rect 15381 18275 15439 18281
rect 15381 18241 15393 18275
rect 15427 18272 15439 18275
rect 16114 18272 16120 18284
rect 15427 18244 16120 18272
rect 15427 18241 15439 18244
rect 15381 18235 15439 18241
rect 16114 18232 16120 18244
rect 16172 18232 16178 18284
rect 18782 18272 18788 18284
rect 18743 18244 18788 18272
rect 18782 18232 18788 18244
rect 18840 18232 18846 18284
rect 20640 18281 20668 18380
rect 20625 18275 20683 18281
rect 20625 18241 20637 18275
rect 20671 18241 20683 18275
rect 20625 18235 20683 18241
rect 20806 18232 20812 18284
rect 20864 18272 20870 18284
rect 20901 18275 20959 18281
rect 20901 18272 20913 18275
rect 20864 18244 20913 18272
rect 20864 18232 20870 18244
rect 20901 18241 20913 18244
rect 20947 18241 20959 18275
rect 20901 18235 20959 18241
rect 9858 18204 9864 18216
rect 3927 18176 4154 18204
rect 9819 18176 9864 18204
rect 3927 18173 3939 18176
rect 3881 18167 3939 18173
rect 3142 18096 3148 18148
rect 3200 18136 3206 18148
rect 3237 18139 3295 18145
rect 3237 18136 3249 18139
rect 3200 18108 3249 18136
rect 3200 18096 3206 18108
rect 3237 18105 3249 18108
rect 3283 18136 3295 18139
rect 3896 18136 3924 18167
rect 9858 18164 9864 18176
rect 9916 18164 9922 18216
rect 10321 18207 10379 18213
rect 10321 18173 10333 18207
rect 10367 18173 10379 18207
rect 10321 18167 10379 18173
rect 4062 18136 4068 18148
rect 3283 18108 3924 18136
rect 4023 18108 4068 18136
rect 3283 18105 3295 18108
rect 3237 18099 3295 18105
rect 4062 18096 4068 18108
rect 4120 18096 4126 18148
rect 5077 18139 5135 18145
rect 5077 18105 5089 18139
rect 5123 18105 5135 18139
rect 8294 18136 8300 18148
rect 8255 18108 8300 18136
rect 5077 18099 5135 18105
rect 1670 18068 1676 18080
rect 1631 18040 1676 18068
rect 1670 18028 1676 18040
rect 1728 18028 1734 18080
rect 1946 18068 1952 18080
rect 1907 18040 1952 18068
rect 1946 18028 1952 18040
rect 2004 18028 2010 18080
rect 4430 18068 4436 18080
rect 4391 18040 4436 18068
rect 4430 18028 4436 18040
rect 4488 18028 4494 18080
rect 4801 18071 4859 18077
rect 4801 18037 4813 18071
rect 4847 18068 4859 18071
rect 5092 18068 5120 18099
rect 8294 18096 8300 18108
rect 8352 18096 8358 18148
rect 8389 18139 8447 18145
rect 8389 18105 8401 18139
rect 8435 18105 8447 18139
rect 8389 18099 8447 18105
rect 9309 18139 9367 18145
rect 9309 18105 9321 18139
rect 9355 18136 9367 18139
rect 9355 18108 9674 18136
rect 9355 18105 9367 18108
rect 9309 18099 9367 18105
rect 5166 18068 5172 18080
rect 4847 18040 5172 18068
rect 4847 18037 4859 18040
rect 4801 18031 4859 18037
rect 5166 18028 5172 18040
rect 5224 18028 5230 18080
rect 7466 18068 7472 18080
rect 7427 18040 7472 18068
rect 7466 18028 7472 18040
rect 7524 18028 7530 18080
rect 7926 18028 7932 18080
rect 7984 18068 7990 18080
rect 8021 18071 8079 18077
rect 8021 18068 8033 18071
rect 7984 18040 8033 18068
rect 7984 18028 7990 18040
rect 8021 18037 8033 18040
rect 8067 18068 8079 18071
rect 8404 18068 8432 18099
rect 8067 18040 8432 18068
rect 9646 18068 9674 18108
rect 10336 18068 10364 18167
rect 13170 18164 13176 18216
rect 13228 18204 13234 18216
rect 14252 18207 14310 18213
rect 14252 18204 14264 18207
rect 13228 18176 14264 18204
rect 13228 18164 13234 18176
rect 14252 18173 14264 18176
rect 14298 18204 14310 18207
rect 14645 18207 14703 18213
rect 14645 18204 14657 18207
rect 14298 18176 14657 18204
rect 14298 18173 14310 18176
rect 14252 18167 14310 18173
rect 14645 18173 14657 18176
rect 14691 18173 14703 18207
rect 14645 18167 14703 18173
rect 12621 18139 12679 18145
rect 12621 18105 12633 18139
rect 12667 18105 12679 18139
rect 12621 18099 12679 18105
rect 15473 18139 15531 18145
rect 15473 18105 15485 18139
rect 15519 18136 15531 18139
rect 15746 18136 15752 18148
rect 15519 18108 15752 18136
rect 15519 18105 15531 18108
rect 15473 18099 15531 18105
rect 11054 18068 11060 18080
rect 9646 18040 11060 18068
rect 8067 18037 8079 18040
rect 8021 18031 8079 18037
rect 11054 18028 11060 18040
rect 11112 18028 11118 18080
rect 11790 18068 11796 18080
rect 11751 18040 11796 18068
rect 11790 18028 11796 18040
rect 11848 18028 11854 18080
rect 12342 18028 12348 18080
rect 12400 18068 12406 18080
rect 12636 18068 12664 18099
rect 15746 18096 15752 18108
rect 15804 18096 15810 18148
rect 16025 18139 16083 18145
rect 16025 18105 16037 18139
rect 16071 18136 16083 18139
rect 18414 18136 18420 18148
rect 16071 18108 18420 18136
rect 16071 18105 16083 18108
rect 16025 18099 16083 18105
rect 18414 18096 18420 18108
rect 18472 18096 18478 18148
rect 19106 18139 19164 18145
rect 19106 18105 19118 18139
rect 19152 18105 19164 18139
rect 19106 18099 19164 18105
rect 20717 18139 20775 18145
rect 20717 18105 20729 18139
rect 20763 18105 20775 18139
rect 20717 18099 20775 18105
rect 15194 18068 15200 18080
rect 12400 18040 12664 18068
rect 15155 18040 15200 18068
rect 12400 18028 12406 18040
rect 15194 18028 15200 18040
rect 15252 18028 15258 18080
rect 16666 18068 16672 18080
rect 16627 18040 16672 18068
rect 16666 18028 16672 18040
rect 16724 18028 16730 18080
rect 16850 18028 16856 18080
rect 16908 18068 16914 18080
rect 17037 18071 17095 18077
rect 17037 18068 17049 18071
rect 16908 18040 17049 18068
rect 16908 18028 16914 18040
rect 17037 18037 17049 18040
rect 17083 18068 17095 18071
rect 17402 18068 17408 18080
rect 17083 18040 17408 18068
rect 17083 18037 17095 18040
rect 17037 18031 17095 18037
rect 17402 18028 17408 18040
rect 17460 18028 17466 18080
rect 17494 18028 17500 18080
rect 17552 18068 17558 18080
rect 18601 18071 18659 18077
rect 18601 18068 18613 18071
rect 17552 18040 18613 18068
rect 17552 18028 17558 18040
rect 18601 18037 18613 18040
rect 18647 18068 18659 18071
rect 19121 18068 19149 18099
rect 18647 18040 19149 18068
rect 19705 18071 19763 18077
rect 18647 18037 18659 18040
rect 18601 18031 18659 18037
rect 19705 18037 19717 18071
rect 19751 18068 19763 18071
rect 20530 18068 20536 18080
rect 19751 18040 20536 18068
rect 19751 18037 19763 18040
rect 19705 18031 19763 18037
rect 20530 18028 20536 18040
rect 20588 18068 20594 18080
rect 20732 18068 20760 18099
rect 21542 18068 21548 18080
rect 20588 18040 20760 18068
rect 21503 18040 21548 18068
rect 20588 18028 20594 18040
rect 21542 18028 21548 18040
rect 21600 18028 21606 18080
rect 1104 17978 22816 18000
rect 1104 17926 8982 17978
rect 9034 17926 9046 17978
rect 9098 17926 9110 17978
rect 9162 17926 9174 17978
rect 9226 17926 16982 17978
rect 17034 17926 17046 17978
rect 17098 17926 17110 17978
rect 17162 17926 17174 17978
rect 17226 17926 22816 17978
rect 1104 17904 22816 17926
rect 2222 17864 2228 17876
rect 2183 17836 2228 17864
rect 2222 17824 2228 17836
rect 2280 17824 2286 17876
rect 3418 17864 3424 17876
rect 3379 17836 3424 17864
rect 3418 17824 3424 17836
rect 3476 17824 3482 17876
rect 5166 17864 5172 17876
rect 5127 17836 5172 17864
rect 5166 17824 5172 17836
rect 5224 17824 5230 17876
rect 8386 17824 8392 17876
rect 8444 17864 8450 17876
rect 13170 17864 13176 17876
rect 8444 17836 13176 17864
rect 8444 17824 8450 17836
rect 13170 17824 13176 17836
rect 13228 17824 13234 17876
rect 15654 17864 15660 17876
rect 15615 17836 15660 17864
rect 15654 17824 15660 17836
rect 15712 17824 15718 17876
rect 15746 17824 15752 17876
rect 15804 17864 15810 17876
rect 16209 17867 16267 17873
rect 16209 17864 16221 17867
rect 15804 17836 16221 17864
rect 15804 17824 15810 17836
rect 16209 17833 16221 17836
rect 16255 17833 16267 17867
rect 17494 17864 17500 17876
rect 17455 17836 17500 17864
rect 16209 17827 16267 17833
rect 17494 17824 17500 17836
rect 17552 17824 17558 17876
rect 18782 17824 18788 17876
rect 18840 17864 18846 17876
rect 18969 17867 19027 17873
rect 18969 17864 18981 17867
rect 18840 17836 18981 17864
rect 18840 17824 18846 17836
rect 18969 17833 18981 17836
rect 19015 17833 19027 17867
rect 20530 17864 20536 17876
rect 20491 17836 20536 17864
rect 18969 17827 19027 17833
rect 20530 17824 20536 17836
rect 20588 17824 20594 17876
rect 21082 17864 21088 17876
rect 21043 17836 21088 17864
rect 21082 17824 21088 17836
rect 21140 17824 21146 17876
rect 4154 17756 4160 17808
rect 4212 17796 4218 17808
rect 4570 17799 4628 17805
rect 4570 17796 4582 17799
rect 4212 17768 4582 17796
rect 4212 17756 4218 17768
rect 4570 17765 4582 17768
rect 4616 17765 4628 17799
rect 4570 17759 4628 17765
rect 7555 17799 7613 17805
rect 7555 17765 7567 17799
rect 7601 17796 7613 17799
rect 7742 17796 7748 17808
rect 7601 17768 7748 17796
rect 7601 17765 7613 17768
rect 7555 17759 7613 17765
rect 7742 17756 7748 17768
rect 7800 17756 7806 17808
rect 11333 17799 11391 17805
rect 11333 17765 11345 17799
rect 11379 17796 11391 17799
rect 11790 17796 11796 17808
rect 11379 17768 11796 17796
rect 11379 17765 11391 17768
rect 11333 17759 11391 17765
rect 11790 17756 11796 17768
rect 11848 17756 11854 17808
rect 12250 17756 12256 17808
rect 12308 17796 12314 17808
rect 12621 17799 12679 17805
rect 12621 17796 12633 17799
rect 12308 17768 12633 17796
rect 12308 17756 12314 17768
rect 12621 17765 12633 17768
rect 12667 17765 12679 17799
rect 12621 17759 12679 17765
rect 15194 17756 15200 17808
rect 15252 17796 15258 17808
rect 20714 17796 20720 17808
rect 15252 17768 20720 17796
rect 15252 17756 15258 17768
rect 20714 17756 20720 17768
rect 20772 17796 20778 17808
rect 20772 17768 20944 17796
rect 20772 17756 20778 17768
rect 4062 17688 4068 17740
rect 4120 17728 4126 17740
rect 4249 17731 4307 17737
rect 4249 17728 4261 17731
rect 4120 17700 4261 17728
rect 4120 17688 4126 17700
rect 4249 17697 4261 17700
rect 4295 17697 4307 17731
rect 4249 17691 4307 17697
rect 4706 17688 4712 17740
rect 4764 17728 4770 17740
rect 5994 17728 6000 17740
rect 6052 17737 6058 17740
rect 6052 17731 6090 17737
rect 4764 17700 6000 17728
rect 4764 17688 4770 17700
rect 5994 17688 6000 17700
rect 6078 17697 6090 17731
rect 7190 17728 7196 17740
rect 7151 17700 7196 17728
rect 6052 17691 6090 17697
rect 6052 17688 6058 17691
rect 7190 17688 7196 17700
rect 7248 17688 7254 17740
rect 10870 17728 10876 17740
rect 10831 17700 10876 17728
rect 10870 17688 10876 17700
rect 10928 17688 10934 17740
rect 11054 17728 11060 17740
rect 11015 17700 11060 17728
rect 11054 17688 11060 17700
rect 11112 17688 11118 17740
rect 13262 17688 13268 17740
rect 13320 17728 13326 17740
rect 14036 17731 14094 17737
rect 14036 17728 14048 17731
rect 13320 17700 14048 17728
rect 13320 17688 13326 17700
rect 14036 17697 14048 17700
rect 14082 17697 14094 17731
rect 14036 17691 14094 17697
rect 17129 17731 17187 17737
rect 17129 17697 17141 17731
rect 17175 17728 17187 17731
rect 17310 17728 17316 17740
rect 17175 17700 17316 17728
rect 17175 17697 17187 17700
rect 17129 17691 17187 17697
rect 17310 17688 17316 17700
rect 17368 17688 17374 17740
rect 18874 17728 18880 17740
rect 18835 17700 18880 17728
rect 18874 17688 18880 17700
rect 18932 17688 18938 17740
rect 19058 17688 19064 17740
rect 19116 17728 19122 17740
rect 20916 17737 20944 17768
rect 19337 17731 19395 17737
rect 19337 17728 19349 17731
rect 19116 17700 19349 17728
rect 19116 17688 19122 17700
rect 19337 17697 19349 17700
rect 19383 17697 19395 17731
rect 19337 17691 19395 17697
rect 20901 17731 20959 17737
rect 20901 17697 20913 17731
rect 20947 17697 20959 17731
rect 20901 17691 20959 17697
rect 1857 17663 1915 17669
rect 1857 17629 1869 17663
rect 1903 17629 1915 17663
rect 12529 17663 12587 17669
rect 12529 17660 12541 17663
rect 1857 17623 1915 17629
rect 12519 17629 12541 17660
rect 12575 17629 12587 17663
rect 12519 17623 12587 17629
rect 1872 17536 1900 17623
rect 7466 17552 7472 17604
rect 7524 17592 7530 17604
rect 7524 17564 10548 17592
rect 7524 17552 7530 17564
rect 1765 17527 1823 17533
rect 1765 17493 1777 17527
rect 1811 17524 1823 17527
rect 1854 17524 1860 17536
rect 1811 17496 1860 17524
rect 1811 17493 1823 17496
rect 1765 17487 1823 17493
rect 1854 17484 1860 17496
rect 1912 17484 1918 17536
rect 2774 17524 2780 17536
rect 2735 17496 2780 17524
rect 2774 17484 2780 17496
rect 2832 17484 2838 17536
rect 5902 17484 5908 17536
rect 5960 17524 5966 17536
rect 6135 17527 6193 17533
rect 6135 17524 6147 17527
rect 5960 17496 6147 17524
rect 5960 17484 5966 17496
rect 6135 17493 6147 17496
rect 6181 17493 6193 17527
rect 6135 17487 6193 17493
rect 7926 17484 7932 17536
rect 7984 17524 7990 17536
rect 8113 17527 8171 17533
rect 8113 17524 8125 17527
rect 7984 17496 8125 17524
rect 7984 17484 7990 17496
rect 8113 17493 8125 17496
rect 8159 17493 8171 17527
rect 8113 17487 8171 17493
rect 8846 17484 8852 17536
rect 8904 17524 8910 17536
rect 9858 17524 9864 17536
rect 8904 17496 9864 17524
rect 8904 17484 8910 17496
rect 9858 17484 9864 17496
rect 9916 17484 9922 17536
rect 10520 17533 10548 17564
rect 10505 17527 10563 17533
rect 10505 17493 10517 17527
rect 10551 17524 10563 17527
rect 10778 17524 10784 17536
rect 10551 17496 10784 17524
rect 10551 17493 10563 17496
rect 10505 17487 10563 17493
rect 10778 17484 10784 17496
rect 10836 17484 10842 17536
rect 12519 17524 12547 17623
rect 12618 17620 12624 17672
rect 12676 17660 12682 17672
rect 12805 17663 12863 17669
rect 12805 17660 12817 17663
rect 12676 17632 12817 17660
rect 12676 17620 12682 17632
rect 12805 17629 12817 17632
rect 12851 17629 12863 17663
rect 12805 17623 12863 17629
rect 12820 17592 12848 17623
rect 13354 17620 13360 17672
rect 13412 17660 13418 17672
rect 14139 17663 14197 17669
rect 14139 17660 14151 17663
rect 13412 17632 14151 17660
rect 13412 17620 13418 17632
rect 14139 17629 14151 17632
rect 14185 17629 14197 17663
rect 15286 17660 15292 17672
rect 15247 17632 15292 17660
rect 14139 17623 14197 17629
rect 15286 17620 15292 17632
rect 15344 17620 15350 17672
rect 13814 17592 13820 17604
rect 12820 17564 13820 17592
rect 13814 17552 13820 17564
rect 13872 17552 13878 17604
rect 12710 17524 12716 17536
rect 12519 17496 12716 17524
rect 12710 17484 12716 17496
rect 12768 17524 12774 17536
rect 13354 17524 13360 17536
rect 12768 17496 13360 17524
rect 12768 17484 12774 17496
rect 13354 17484 13360 17496
rect 13412 17484 13418 17536
rect 13446 17484 13452 17536
rect 13504 17524 13510 17536
rect 15470 17524 15476 17536
rect 13504 17496 15476 17524
rect 13504 17484 13510 17496
rect 15470 17484 15476 17496
rect 15528 17484 15534 17536
rect 18046 17524 18052 17536
rect 18007 17496 18052 17524
rect 18046 17484 18052 17496
rect 18104 17484 18110 17536
rect 18414 17524 18420 17536
rect 18375 17496 18420 17524
rect 18414 17484 18420 17496
rect 18472 17484 18478 17536
rect 19702 17484 19708 17536
rect 19760 17524 19766 17536
rect 19889 17527 19947 17533
rect 19889 17524 19901 17527
rect 19760 17496 19901 17524
rect 19760 17484 19766 17496
rect 19889 17493 19901 17496
rect 19935 17493 19947 17527
rect 19889 17487 19947 17493
rect 1104 17434 22816 17456
rect 1104 17382 4982 17434
rect 5034 17382 5046 17434
rect 5098 17382 5110 17434
rect 5162 17382 5174 17434
rect 5226 17382 12982 17434
rect 13034 17382 13046 17434
rect 13098 17382 13110 17434
rect 13162 17382 13174 17434
rect 13226 17382 20982 17434
rect 21034 17382 21046 17434
rect 21098 17382 21110 17434
rect 21162 17382 21174 17434
rect 21226 17382 22816 17434
rect 1104 17360 22816 17382
rect 1949 17323 2007 17329
rect 1949 17289 1961 17323
rect 1995 17320 2007 17323
rect 2222 17320 2228 17332
rect 1995 17292 2228 17320
rect 1995 17289 2007 17292
rect 1949 17283 2007 17289
rect 2222 17280 2228 17292
rect 2280 17280 2286 17332
rect 3881 17323 3939 17329
rect 3881 17289 3893 17323
rect 3927 17320 3939 17323
rect 4062 17320 4068 17332
rect 3927 17292 4068 17320
rect 3927 17289 3939 17292
rect 3881 17283 3939 17289
rect 4062 17280 4068 17292
rect 4120 17280 4126 17332
rect 5994 17320 6000 17332
rect 5955 17292 6000 17320
rect 5994 17280 6000 17292
rect 6052 17280 6058 17332
rect 8294 17280 8300 17332
rect 8352 17320 8358 17332
rect 9539 17323 9597 17329
rect 9539 17320 9551 17323
rect 8352 17292 9551 17320
rect 8352 17280 8358 17292
rect 9539 17289 9551 17292
rect 9585 17289 9597 17323
rect 9539 17283 9597 17289
rect 11974 17280 11980 17332
rect 12032 17320 12038 17332
rect 13446 17320 13452 17332
rect 12032 17292 13452 17320
rect 12032 17280 12038 17292
rect 13446 17280 13452 17292
rect 13504 17280 13510 17332
rect 15286 17280 15292 17332
rect 15344 17320 15350 17332
rect 16669 17323 16727 17329
rect 16669 17320 16681 17323
rect 15344 17292 16681 17320
rect 15344 17280 15350 17292
rect 16669 17289 16681 17292
rect 16715 17289 16727 17323
rect 16669 17283 16727 17289
rect 17865 17323 17923 17329
rect 17865 17289 17877 17323
rect 17911 17320 17923 17323
rect 18046 17320 18052 17332
rect 17911 17292 18052 17320
rect 17911 17289 17923 17292
rect 17865 17283 17923 17289
rect 18046 17280 18052 17292
rect 18104 17280 18110 17332
rect 18874 17280 18880 17332
rect 18932 17320 18938 17332
rect 19429 17323 19487 17329
rect 19429 17320 19441 17323
rect 18932 17292 19441 17320
rect 18932 17280 18938 17292
rect 19429 17289 19441 17292
rect 19475 17289 19487 17323
rect 19429 17283 19487 17289
rect 20714 17280 20720 17332
rect 20772 17320 20778 17332
rect 20901 17323 20959 17329
rect 20901 17320 20913 17323
rect 20772 17292 20913 17320
rect 20772 17280 20778 17292
rect 20901 17289 20913 17292
rect 20947 17289 20959 17323
rect 20901 17283 20959 17289
rect 1670 17212 1676 17264
rect 1728 17252 1734 17264
rect 2869 17255 2927 17261
rect 2869 17252 2881 17255
rect 1728 17224 2881 17252
rect 1728 17212 1734 17224
rect 2869 17221 2881 17224
rect 2915 17252 2927 17255
rect 2915 17224 4154 17252
rect 2915 17221 2927 17224
rect 2869 17215 2927 17221
rect 1946 17144 1952 17196
rect 2004 17184 2010 17196
rect 2317 17187 2375 17193
rect 2317 17184 2329 17187
rect 2004 17156 2329 17184
rect 2004 17144 2010 17156
rect 2317 17153 2329 17156
rect 2363 17184 2375 17187
rect 3237 17187 3295 17193
rect 3237 17184 3249 17187
rect 2363 17156 3249 17184
rect 2363 17153 2375 17156
rect 2317 17147 2375 17153
rect 3237 17153 3249 17156
rect 3283 17153 3295 17187
rect 4126 17184 4154 17224
rect 4706 17212 4712 17264
rect 4764 17252 4770 17264
rect 7377 17255 7435 17261
rect 7377 17252 7389 17255
rect 4764 17224 7389 17252
rect 4764 17212 4770 17224
rect 5077 17187 5135 17193
rect 5077 17184 5089 17187
rect 4126 17156 5089 17184
rect 3237 17147 3295 17153
rect 5077 17153 5089 17156
rect 5123 17184 5135 17187
rect 5350 17184 5356 17196
rect 5123 17156 5356 17184
rect 5123 17153 5135 17156
rect 5077 17147 5135 17153
rect 5350 17144 5356 17156
rect 5408 17144 5414 17196
rect 6891 17125 6919 17224
rect 7377 17221 7389 17224
rect 7423 17252 7435 17255
rect 9766 17252 9772 17264
rect 7423 17224 9772 17252
rect 7423 17221 7435 17224
rect 7377 17215 7435 17221
rect 9766 17212 9772 17224
rect 9824 17212 9830 17264
rect 13262 17252 13268 17264
rect 11532 17224 13268 17252
rect 6963 17187 7021 17193
rect 6963 17153 6975 17187
rect 7009 17184 7021 17187
rect 7929 17187 7987 17193
rect 7929 17184 7941 17187
rect 7009 17156 7941 17184
rect 7009 17153 7021 17156
rect 6963 17147 7021 17153
rect 7929 17153 7941 17156
rect 7975 17184 7987 17187
rect 8849 17187 8907 17193
rect 8849 17184 8861 17187
rect 7975 17156 8861 17184
rect 7975 17153 7987 17156
rect 7929 17147 7987 17153
rect 8849 17153 8861 17156
rect 8895 17153 8907 17187
rect 8849 17147 8907 17153
rect 9490 17125 9496 17128
rect 6876 17119 6934 17125
rect 6876 17085 6888 17119
rect 6922 17085 6934 17119
rect 6876 17079 6934 17085
rect 9468 17119 9496 17125
rect 9468 17085 9480 17119
rect 9548 17116 9554 17128
rect 10689 17119 10747 17125
rect 9548 17088 9996 17116
rect 9468 17079 9496 17085
rect 9490 17076 9496 17079
rect 9548 17076 9554 17088
rect 2409 17051 2467 17057
rect 2409 17017 2421 17051
rect 2455 17048 2467 17051
rect 2774 17048 2780 17060
rect 2455 17020 2780 17048
rect 2455 17017 2467 17020
rect 2409 17011 2467 17017
rect 2774 17008 2780 17020
rect 2832 17008 2838 17060
rect 4430 17048 4436 17060
rect 4391 17020 4436 17048
rect 4430 17008 4436 17020
rect 4488 17008 4494 17060
rect 4525 17051 4583 17057
rect 4525 17017 4537 17051
rect 4571 17017 4583 17051
rect 4525 17011 4583 17017
rect 2222 16940 2228 16992
rect 2280 16980 2286 16992
rect 2590 16980 2596 16992
rect 2280 16952 2596 16980
rect 2280 16940 2286 16952
rect 2590 16940 2596 16952
rect 2648 16980 2654 16992
rect 4154 16980 4160 16992
rect 2648 16952 4160 16980
rect 2648 16940 2654 16952
rect 4154 16940 4160 16952
rect 4212 16940 4218 16992
rect 4540 16980 4568 17011
rect 7926 17008 7932 17060
rect 7984 17048 7990 17060
rect 8021 17051 8079 17057
rect 8021 17048 8033 17051
rect 7984 17020 8033 17048
rect 7984 17008 7990 17020
rect 8021 17017 8033 17020
rect 8067 17017 8079 17051
rect 8021 17011 8079 17017
rect 8110 17008 8116 17060
rect 8168 17048 8174 17060
rect 8573 17051 8631 17057
rect 8573 17048 8585 17051
rect 8168 17020 8585 17048
rect 8168 17008 8174 17020
rect 8573 17017 8585 17020
rect 8619 17017 8631 17051
rect 8573 17011 8631 17017
rect 4982 16980 4988 16992
rect 4540 16952 4988 16980
rect 4982 16940 4988 16952
rect 5040 16980 5046 16992
rect 5353 16983 5411 16989
rect 5353 16980 5365 16983
rect 5040 16952 5365 16980
rect 5040 16940 5046 16952
rect 5353 16949 5365 16952
rect 5399 16949 5411 16983
rect 7742 16980 7748 16992
rect 7655 16952 7748 16980
rect 5353 16943 5411 16949
rect 7742 16940 7748 16952
rect 7800 16980 7806 16992
rect 8478 16980 8484 16992
rect 7800 16952 8484 16980
rect 7800 16940 7806 16952
rect 8478 16940 8484 16952
rect 8536 16940 8542 16992
rect 9968 16989 9996 17088
rect 10689 17085 10701 17119
rect 10735 17116 10747 17119
rect 10778 17116 10784 17128
rect 10735 17088 10784 17116
rect 10735 17085 10747 17088
rect 10689 17079 10747 17085
rect 10778 17076 10784 17088
rect 10836 17076 10842 17128
rect 10873 17119 10931 17125
rect 10873 17085 10885 17119
rect 10919 17116 10931 17119
rect 11054 17116 11060 17128
rect 10919 17088 11060 17116
rect 10919 17085 10931 17088
rect 10873 17079 10931 17085
rect 10321 17051 10379 17057
rect 10321 17017 10333 17051
rect 10367 17048 10379 17051
rect 10410 17048 10416 17060
rect 10367 17020 10416 17048
rect 10367 17017 10379 17020
rect 10321 17011 10379 17017
rect 10410 17008 10416 17020
rect 10468 17048 10474 17060
rect 10888 17048 10916 17079
rect 11054 17076 11060 17088
rect 11112 17116 11118 17128
rect 11425 17119 11483 17125
rect 11425 17116 11437 17119
rect 11112 17088 11437 17116
rect 11112 17076 11118 17088
rect 11425 17085 11437 17088
rect 11471 17085 11483 17119
rect 11425 17079 11483 17085
rect 11146 17048 11152 17060
rect 10468 17020 10916 17048
rect 11107 17020 11152 17048
rect 10468 17008 10474 17020
rect 11146 17008 11152 17020
rect 11204 17008 11210 17060
rect 9953 16983 10011 16989
rect 9953 16949 9965 16983
rect 9999 16980 10011 16983
rect 11532 16980 11560 17224
rect 13262 17212 13268 17224
rect 13320 17212 13326 17264
rect 12526 17184 12532 17196
rect 12487 17156 12532 17184
rect 12526 17144 12532 17156
rect 12584 17144 12590 17196
rect 12802 17184 12808 17196
rect 12763 17156 12808 17184
rect 12802 17144 12808 17156
rect 12860 17144 12866 17196
rect 12894 17144 12900 17196
rect 12952 17184 12958 17196
rect 14829 17187 14887 17193
rect 12952 17156 13814 17184
rect 12952 17144 12958 17156
rect 13786 17116 13814 17156
rect 14829 17153 14841 17187
rect 14875 17184 14887 17187
rect 15304 17184 15332 17280
rect 14875 17156 15332 17184
rect 14875 17153 14887 17156
rect 14829 17147 14887 17153
rect 15562 17144 15568 17196
rect 15620 17184 15626 17196
rect 15749 17187 15807 17193
rect 15749 17184 15761 17187
rect 15620 17156 15761 17184
rect 15620 17144 15626 17156
rect 15749 17153 15761 17156
rect 15795 17184 15807 17187
rect 16206 17184 16212 17196
rect 15795 17156 16212 17184
rect 15795 17153 15807 17156
rect 15749 17147 15807 17153
rect 16206 17144 16212 17156
rect 16264 17144 16270 17196
rect 18141 17187 18199 17193
rect 18141 17153 18153 17187
rect 18187 17184 18199 17187
rect 18414 17184 18420 17196
rect 18187 17156 18420 17184
rect 18187 17153 18199 17156
rect 18141 17147 18199 17153
rect 18414 17144 18420 17156
rect 18472 17144 18478 17196
rect 18785 17187 18843 17193
rect 18785 17153 18797 17187
rect 18831 17184 18843 17187
rect 19981 17187 20039 17193
rect 19981 17184 19993 17187
rect 18831 17156 19993 17184
rect 18831 17153 18843 17156
rect 18785 17147 18843 17153
rect 19981 17153 19993 17156
rect 20027 17184 20039 17187
rect 20806 17184 20812 17196
rect 20027 17156 20812 17184
rect 20027 17153 20039 17156
rect 19981 17147 20039 17153
rect 20806 17144 20812 17156
rect 20864 17144 20870 17196
rect 14090 17116 14096 17128
rect 13786 17088 14096 17116
rect 14090 17076 14096 17088
rect 14148 17076 14154 17128
rect 14553 17119 14611 17125
rect 14553 17116 14565 17119
rect 14235 17088 14565 17116
rect 12618 17048 12624 17060
rect 12579 17020 12624 17048
rect 12618 17008 12624 17020
rect 12676 17008 12682 17060
rect 13633 17051 13691 17057
rect 13633 17017 13645 17051
rect 13679 17048 13691 17051
rect 13722 17048 13728 17060
rect 13679 17020 13728 17048
rect 13679 17017 13691 17020
rect 13633 17011 13691 17017
rect 13722 17008 13728 17020
rect 13780 17048 13786 17060
rect 14235 17048 14263 17088
rect 14553 17085 14565 17088
rect 14599 17085 14611 17119
rect 14553 17079 14611 17085
rect 13780 17020 14263 17048
rect 13780 17008 13786 17020
rect 15838 17008 15844 17060
rect 15896 17048 15902 17060
rect 16390 17048 16396 17060
rect 15896 17020 15941 17048
rect 16351 17020 16396 17048
rect 15896 17008 15902 17020
rect 16390 17008 16396 17020
rect 16448 17008 16454 17060
rect 18233 17051 18291 17057
rect 18233 17017 18245 17051
rect 18279 17017 18291 17051
rect 19702 17048 19708 17060
rect 19663 17020 19708 17048
rect 18233 17011 18291 17017
rect 11790 16980 11796 16992
rect 9999 16952 11560 16980
rect 11751 16952 11796 16980
rect 9999 16949 10011 16952
rect 9953 16943 10011 16949
rect 11790 16940 11796 16952
rect 11848 16940 11854 16992
rect 12250 16980 12256 16992
rect 12211 16952 12256 16980
rect 12250 16940 12256 16952
rect 12308 16940 12314 16992
rect 13262 16940 13268 16992
rect 13320 16980 13326 16992
rect 13538 16980 13544 16992
rect 13320 16952 13544 16980
rect 13320 16940 13326 16952
rect 13538 16940 13544 16952
rect 13596 16980 13602 16992
rect 13909 16983 13967 16989
rect 13909 16980 13921 16983
rect 13596 16952 13921 16980
rect 13596 16940 13602 16952
rect 13909 16949 13921 16952
rect 13955 16949 13967 16983
rect 13909 16943 13967 16949
rect 15381 16983 15439 16989
rect 15381 16949 15393 16983
rect 15427 16980 15439 16983
rect 15654 16980 15660 16992
rect 15427 16952 15660 16980
rect 15427 16949 15439 16952
rect 15381 16943 15439 16949
rect 15654 16940 15660 16952
rect 15712 16980 15718 16992
rect 17129 16983 17187 16989
rect 17129 16980 17141 16983
rect 15712 16952 17141 16980
rect 15712 16940 15718 16952
rect 17129 16949 17141 16952
rect 17175 16980 17187 16983
rect 17494 16980 17500 16992
rect 17175 16952 17500 16980
rect 17175 16949 17187 16952
rect 17129 16943 17187 16949
rect 17494 16940 17500 16952
rect 17552 16940 17558 16992
rect 18046 16940 18052 16992
rect 18104 16980 18110 16992
rect 18248 16980 18276 17011
rect 19702 17008 19708 17020
rect 19760 17008 19766 17060
rect 19794 17008 19800 17060
rect 19852 17048 19858 17060
rect 19852 17020 19897 17048
rect 19852 17008 19858 17020
rect 19058 16980 19064 16992
rect 18104 16952 18276 16980
rect 19019 16952 19064 16980
rect 18104 16940 18110 16952
rect 19058 16940 19064 16952
rect 19116 16940 19122 16992
rect 1104 16890 22816 16912
rect 1104 16838 8982 16890
rect 9034 16838 9046 16890
rect 9098 16838 9110 16890
rect 9162 16838 9174 16890
rect 9226 16838 16982 16890
rect 17034 16838 17046 16890
rect 17098 16838 17110 16890
rect 17162 16838 17174 16890
rect 17226 16838 22816 16890
rect 1104 16816 22816 16838
rect 1854 16776 1860 16788
rect 1815 16748 1860 16776
rect 1854 16736 1860 16748
rect 1912 16736 1918 16788
rect 2774 16776 2780 16788
rect 2735 16748 2780 16776
rect 2774 16736 2780 16748
rect 2832 16736 2838 16788
rect 4982 16776 4988 16788
rect 4943 16748 4988 16776
rect 4982 16736 4988 16748
rect 5040 16736 5046 16788
rect 7190 16776 7196 16788
rect 7151 16748 7196 16776
rect 7190 16736 7196 16748
rect 7248 16736 7254 16788
rect 7926 16776 7932 16788
rect 7887 16748 7932 16776
rect 7926 16736 7932 16748
rect 7984 16736 7990 16788
rect 10686 16776 10692 16788
rect 10599 16748 10692 16776
rect 10686 16736 10692 16748
rect 10744 16776 10750 16788
rect 10870 16776 10876 16788
rect 10744 16748 10876 16776
rect 10744 16736 10750 16748
rect 10870 16736 10876 16748
rect 10928 16736 10934 16788
rect 12250 16736 12256 16788
rect 12308 16776 12314 16788
rect 12345 16779 12403 16785
rect 12345 16776 12357 16779
rect 12308 16748 12357 16776
rect 12308 16736 12314 16748
rect 12345 16745 12357 16748
rect 12391 16745 12403 16779
rect 12710 16776 12716 16788
rect 12671 16748 12716 16776
rect 12345 16739 12403 16745
rect 4154 16668 4160 16720
rect 4212 16708 4218 16720
rect 4386 16711 4444 16717
rect 4386 16708 4398 16711
rect 4212 16680 4398 16708
rect 4212 16668 4218 16680
rect 4386 16677 4398 16680
rect 4432 16677 4444 16711
rect 4386 16671 4444 16677
rect 5721 16711 5779 16717
rect 5721 16677 5733 16711
rect 5767 16708 5779 16711
rect 5902 16708 5908 16720
rect 5767 16680 5908 16708
rect 5767 16677 5779 16680
rect 5721 16671 5779 16677
rect 5902 16668 5908 16680
rect 5960 16668 5966 16720
rect 5994 16668 6000 16720
rect 6052 16708 6058 16720
rect 8202 16708 8208 16720
rect 6052 16680 6097 16708
rect 8163 16680 8208 16708
rect 6052 16668 6058 16680
rect 8202 16668 8208 16680
rect 8260 16668 8266 16720
rect 11514 16668 11520 16720
rect 11572 16708 11578 16720
rect 11746 16711 11804 16717
rect 11746 16708 11758 16711
rect 11572 16680 11758 16708
rect 11572 16668 11578 16680
rect 11746 16677 11758 16680
rect 11792 16677 11804 16711
rect 12360 16708 12388 16739
rect 12710 16736 12716 16748
rect 12768 16736 12774 16788
rect 14090 16736 14096 16788
rect 14148 16776 14154 16788
rect 14185 16779 14243 16785
rect 14185 16776 14197 16779
rect 14148 16748 14197 16776
rect 14148 16736 14154 16748
rect 14185 16745 14197 16748
rect 14231 16745 14243 16779
rect 14185 16739 14243 16745
rect 15838 16736 15844 16788
rect 15896 16776 15902 16788
rect 15933 16779 15991 16785
rect 15933 16776 15945 16779
rect 15896 16748 15945 16776
rect 15896 16736 15902 16748
rect 15933 16745 15945 16748
rect 15979 16745 15991 16779
rect 15933 16739 15991 16745
rect 16206 16736 16212 16788
rect 16264 16776 16270 16788
rect 16301 16779 16359 16785
rect 16301 16776 16313 16779
rect 16264 16748 16313 16776
rect 16264 16736 16270 16748
rect 16301 16745 16313 16748
rect 16347 16745 16359 16779
rect 16301 16739 16359 16745
rect 17310 16736 17316 16788
rect 17368 16776 17374 16788
rect 17957 16779 18015 16785
rect 17957 16776 17969 16779
rect 17368 16748 17969 16776
rect 17368 16736 17374 16748
rect 17957 16745 17969 16748
rect 18003 16745 18015 16779
rect 17957 16739 18015 16745
rect 19429 16779 19487 16785
rect 19429 16745 19441 16779
rect 19475 16776 19487 16779
rect 19794 16776 19800 16788
rect 19475 16748 19800 16776
rect 19475 16745 19487 16748
rect 19429 16739 19487 16745
rect 19794 16736 19800 16748
rect 19852 16736 19858 16788
rect 13262 16708 13268 16720
rect 12360 16680 13268 16708
rect 11746 16671 11804 16677
rect 13262 16668 13268 16680
rect 13320 16708 13326 16720
rect 13357 16711 13415 16717
rect 13357 16708 13369 16711
rect 13320 16680 13369 16708
rect 13320 16668 13326 16680
rect 13357 16677 13369 16680
rect 13403 16677 13415 16711
rect 13357 16671 13415 16677
rect 17494 16668 17500 16720
rect 17552 16708 17558 16720
rect 18830 16711 18888 16717
rect 18830 16708 18842 16711
rect 17552 16680 18842 16708
rect 17552 16668 17558 16680
rect 18830 16677 18842 16680
rect 18876 16708 18888 16711
rect 18966 16708 18972 16720
rect 18876 16680 18972 16708
rect 18876 16677 18888 16680
rect 18830 16671 18888 16677
rect 18966 16668 18972 16680
rect 19024 16668 19030 16720
rect 1670 16600 1676 16652
rect 1728 16640 1734 16652
rect 1765 16643 1823 16649
rect 1765 16640 1777 16643
rect 1728 16612 1777 16640
rect 1728 16600 1734 16612
rect 1765 16609 1777 16612
rect 1811 16609 1823 16643
rect 1765 16603 1823 16609
rect 2317 16643 2375 16649
rect 2317 16609 2329 16643
rect 2363 16640 2375 16643
rect 3142 16640 3148 16652
rect 2363 16612 3148 16640
rect 2363 16609 2375 16612
rect 2317 16603 2375 16609
rect 3142 16600 3148 16612
rect 3200 16600 3206 16652
rect 9582 16640 9588 16652
rect 9543 16612 9588 16640
rect 9582 16600 9588 16612
rect 9640 16600 9646 16652
rect 12526 16600 12532 16652
rect 12584 16640 12590 16652
rect 12989 16643 13047 16649
rect 12989 16640 13001 16643
rect 12584 16612 13001 16640
rect 12584 16600 12590 16612
rect 12989 16609 13001 16612
rect 13035 16609 13047 16643
rect 12989 16603 13047 16609
rect 15381 16643 15439 16649
rect 15381 16609 15393 16643
rect 15427 16640 15439 16643
rect 15470 16640 15476 16652
rect 15427 16612 15476 16640
rect 15427 16609 15439 16612
rect 15381 16603 15439 16609
rect 4062 16572 4068 16584
rect 4023 16544 4068 16572
rect 4062 16532 4068 16544
rect 4120 16532 4126 16584
rect 4798 16532 4804 16584
rect 4856 16572 4862 16584
rect 6181 16575 6239 16581
rect 6181 16572 6193 16575
rect 4856 16544 6193 16572
rect 4856 16532 4862 16544
rect 6181 16541 6193 16544
rect 6227 16541 6239 16575
rect 6181 16535 6239 16541
rect 6196 16504 6224 16535
rect 7926 16532 7932 16584
rect 7984 16572 7990 16584
rect 8113 16575 8171 16581
rect 8113 16572 8125 16575
rect 7984 16544 8125 16572
rect 7984 16532 7990 16544
rect 8113 16541 8125 16544
rect 8159 16541 8171 16575
rect 8113 16535 8171 16541
rect 8389 16575 8447 16581
rect 8389 16541 8401 16575
rect 8435 16572 8447 16575
rect 8570 16572 8576 16584
rect 8435 16544 8576 16572
rect 8435 16541 8447 16544
rect 8389 16535 8447 16541
rect 8404 16504 8432 16535
rect 8570 16532 8576 16544
rect 8628 16532 8634 16584
rect 11146 16532 11152 16584
rect 11204 16572 11210 16584
rect 11425 16575 11483 16581
rect 11425 16572 11437 16575
rect 11204 16544 11437 16572
rect 11204 16532 11210 16544
rect 11425 16541 11437 16544
rect 11471 16572 11483 16575
rect 12158 16572 12164 16584
rect 11471 16544 12164 16572
rect 11471 16541 11483 16544
rect 11425 16535 11483 16541
rect 12158 16532 12164 16544
rect 12216 16532 12222 16584
rect 6196 16476 8432 16504
rect 11882 16464 11888 16516
rect 11940 16504 11946 16516
rect 12894 16504 12900 16516
rect 11940 16476 12900 16504
rect 11940 16464 11946 16476
rect 12894 16464 12900 16476
rect 12952 16464 12958 16516
rect 13004 16504 13032 16603
rect 15470 16600 15476 16612
rect 15528 16600 15534 16652
rect 17221 16643 17279 16649
rect 17221 16609 17233 16643
rect 17267 16609 17279 16643
rect 17221 16603 17279 16609
rect 13265 16575 13323 16581
rect 13265 16541 13277 16575
rect 13311 16572 13323 16575
rect 13354 16572 13360 16584
rect 13311 16544 13360 16572
rect 13311 16541 13323 16544
rect 13265 16535 13323 16541
rect 13354 16532 13360 16544
rect 13412 16532 13418 16584
rect 13541 16575 13599 16581
rect 13541 16541 13553 16575
rect 13587 16541 13599 16575
rect 17236 16572 17264 16603
rect 17310 16600 17316 16652
rect 17368 16640 17374 16652
rect 17405 16643 17463 16649
rect 17405 16640 17417 16643
rect 17368 16612 17417 16640
rect 17368 16600 17374 16612
rect 17405 16609 17417 16612
rect 17451 16640 17463 16643
rect 19058 16640 19064 16652
rect 17451 16612 19064 16640
rect 17451 16609 17463 16612
rect 17405 16603 17463 16609
rect 19058 16600 19064 16612
rect 19116 16600 19122 16652
rect 20806 16600 20812 16652
rect 20864 16640 20870 16652
rect 20901 16643 20959 16649
rect 20901 16640 20913 16643
rect 20864 16612 20913 16640
rect 20864 16600 20870 16612
rect 20901 16609 20913 16612
rect 20947 16609 20959 16643
rect 20901 16603 20959 16609
rect 17494 16572 17500 16584
rect 17236 16544 17500 16572
rect 13541 16535 13599 16541
rect 13556 16504 13584 16535
rect 17494 16532 17500 16544
rect 17552 16532 17558 16584
rect 17681 16575 17739 16581
rect 17681 16541 17693 16575
rect 17727 16572 17739 16575
rect 18509 16575 18567 16581
rect 18509 16572 18521 16575
rect 17727 16544 18521 16572
rect 17727 16541 17739 16544
rect 17681 16535 17739 16541
rect 18509 16541 18521 16544
rect 18555 16572 18567 16575
rect 19426 16572 19432 16584
rect 18555 16544 19432 16572
rect 18555 16541 18567 16544
rect 18509 16535 18567 16541
rect 19426 16532 19432 16544
rect 19484 16532 19490 16584
rect 21082 16504 21088 16516
rect 13004 16476 13584 16504
rect 21043 16476 21088 16504
rect 21082 16464 21088 16476
rect 21140 16464 21146 16516
rect 6914 16436 6920 16448
rect 6875 16408 6920 16436
rect 6914 16396 6920 16408
rect 6972 16396 6978 16448
rect 9306 16396 9312 16448
rect 9364 16436 9370 16448
rect 9815 16439 9873 16445
rect 9815 16436 9827 16439
rect 9364 16408 9827 16436
rect 9364 16396 9370 16408
rect 9815 16405 9827 16408
rect 9861 16405 9873 16439
rect 9815 16399 9873 16405
rect 15611 16439 15669 16445
rect 15611 16405 15623 16439
rect 15657 16436 15669 16439
rect 15838 16436 15844 16448
rect 15657 16408 15844 16436
rect 15657 16405 15669 16408
rect 15611 16399 15669 16405
rect 15838 16396 15844 16408
rect 15896 16396 15902 16448
rect 18322 16436 18328 16448
rect 18283 16408 18328 16436
rect 18322 16396 18328 16408
rect 18380 16396 18386 16448
rect 1104 16346 22816 16368
rect 1104 16294 4982 16346
rect 5034 16294 5046 16346
rect 5098 16294 5110 16346
rect 5162 16294 5174 16346
rect 5226 16294 12982 16346
rect 13034 16294 13046 16346
rect 13098 16294 13110 16346
rect 13162 16294 13174 16346
rect 13226 16294 20982 16346
rect 21034 16294 21046 16346
rect 21098 16294 21110 16346
rect 21162 16294 21174 16346
rect 21226 16294 22816 16346
rect 1104 16272 22816 16294
rect 3789 16235 3847 16241
rect 3789 16232 3801 16235
rect 3344 16204 3801 16232
rect 1578 16164 1584 16176
rect 1539 16136 1584 16164
rect 1578 16124 1584 16136
rect 1636 16124 1642 16176
rect 1946 16056 1952 16108
rect 2004 16096 2010 16108
rect 3344 16105 3372 16204
rect 3789 16201 3801 16204
rect 3835 16232 3847 16235
rect 4062 16232 4068 16244
rect 3835 16204 4068 16232
rect 3835 16201 3847 16204
rect 3789 16195 3847 16201
rect 4062 16192 4068 16204
rect 4120 16192 4126 16244
rect 4154 16192 4160 16244
rect 4212 16232 4218 16244
rect 4798 16232 4804 16244
rect 4212 16204 4804 16232
rect 4212 16192 4218 16204
rect 4798 16192 4804 16204
rect 4856 16192 4862 16244
rect 5905 16235 5963 16241
rect 5905 16201 5917 16235
rect 5951 16232 5963 16235
rect 5994 16232 6000 16244
rect 5951 16204 6000 16232
rect 5951 16201 5963 16204
rect 5905 16195 5963 16201
rect 5994 16192 6000 16204
rect 6052 16232 6058 16244
rect 6181 16235 6239 16241
rect 6181 16232 6193 16235
rect 6052 16204 6193 16232
rect 6052 16192 6058 16204
rect 6181 16201 6193 16204
rect 6227 16232 6239 16235
rect 6549 16235 6607 16241
rect 6549 16232 6561 16235
rect 6227 16204 6561 16232
rect 6227 16201 6239 16204
rect 6181 16195 6239 16201
rect 6549 16201 6561 16204
rect 6595 16232 6607 16235
rect 7006 16232 7012 16244
rect 6595 16204 7012 16232
rect 6595 16201 6607 16204
rect 6549 16195 6607 16201
rect 7006 16192 7012 16204
rect 7064 16192 7070 16244
rect 10505 16235 10563 16241
rect 10505 16201 10517 16235
rect 10551 16232 10563 16235
rect 10962 16232 10968 16244
rect 10551 16204 10968 16232
rect 10551 16201 10563 16204
rect 10505 16195 10563 16201
rect 10962 16192 10968 16204
rect 11020 16232 11026 16244
rect 11422 16232 11428 16244
rect 11020 16204 11428 16232
rect 11020 16192 11026 16204
rect 11422 16192 11428 16204
rect 11480 16192 11486 16244
rect 11517 16235 11575 16241
rect 11517 16201 11529 16235
rect 11563 16232 11575 16235
rect 11790 16232 11796 16244
rect 11563 16204 11796 16232
rect 11563 16201 11575 16204
rect 11517 16195 11575 16201
rect 11790 16192 11796 16204
rect 11848 16192 11854 16244
rect 12158 16232 12164 16244
rect 12119 16204 12164 16232
rect 12158 16192 12164 16204
rect 12216 16192 12222 16244
rect 12575 16235 12633 16241
rect 12575 16201 12587 16235
rect 12621 16232 12633 16235
rect 13354 16232 13360 16244
rect 12621 16204 13360 16232
rect 12621 16201 12633 16204
rect 12575 16195 12633 16201
rect 13354 16192 13360 16204
rect 13412 16232 13418 16244
rect 13633 16235 13691 16241
rect 13633 16232 13645 16235
rect 13412 16204 13645 16232
rect 13412 16192 13418 16204
rect 13633 16201 13645 16204
rect 13679 16201 13691 16235
rect 15470 16232 15476 16244
rect 15431 16204 15476 16232
rect 13633 16195 13691 16201
rect 15470 16192 15476 16204
rect 15528 16192 15534 16244
rect 18966 16192 18972 16244
rect 19024 16232 19030 16244
rect 19061 16235 19119 16241
rect 19061 16232 19073 16235
rect 19024 16204 19073 16232
rect 19024 16192 19030 16204
rect 19061 16201 19073 16204
rect 19107 16201 19119 16235
rect 19426 16232 19432 16244
rect 19387 16204 19432 16232
rect 19061 16195 19119 16201
rect 19426 16192 19432 16204
rect 19484 16192 19490 16244
rect 9033 16167 9091 16173
rect 9033 16164 9045 16167
rect 8128 16136 9045 16164
rect 8128 16108 8156 16136
rect 9033 16133 9045 16136
rect 9079 16133 9091 16167
rect 11440 16164 11468 16192
rect 11885 16167 11943 16173
rect 11885 16164 11897 16167
rect 11440 16136 11897 16164
rect 9033 16127 9091 16133
rect 11885 16133 11897 16136
rect 11931 16133 11943 16167
rect 13262 16164 13268 16176
rect 13223 16136 13268 16164
rect 11885 16127 11943 16133
rect 13262 16124 13268 16136
rect 13320 16124 13326 16176
rect 15010 16164 15016 16176
rect 13786 16136 15016 16164
rect 2501 16099 2559 16105
rect 2501 16096 2513 16099
rect 2004 16068 2513 16096
rect 2004 16056 2010 16068
rect 2501 16065 2513 16068
rect 2547 16096 2559 16099
rect 3329 16099 3387 16105
rect 2547 16068 3188 16096
rect 2547 16065 2559 16068
rect 2501 16059 2559 16065
rect 3160 16040 3188 16068
rect 3329 16065 3341 16099
rect 3375 16065 3387 16099
rect 3329 16059 3387 16065
rect 4430 16056 4436 16108
rect 4488 16096 4494 16108
rect 7193 16099 7251 16105
rect 7193 16096 7205 16099
rect 4488 16068 7205 16096
rect 4488 16056 4494 16068
rect 7193 16065 7205 16068
rect 7239 16096 7251 16099
rect 8110 16096 8116 16108
rect 7239 16068 8116 16096
rect 7239 16065 7251 16068
rect 7193 16059 7251 16065
rect 8110 16056 8116 16068
rect 8168 16056 8174 16108
rect 8481 16099 8539 16105
rect 8481 16065 8493 16099
rect 8527 16096 8539 16099
rect 9306 16096 9312 16108
rect 8527 16068 9312 16096
rect 8527 16065 8539 16068
rect 8481 16059 8539 16065
rect 9306 16056 9312 16068
rect 9364 16056 9370 16108
rect 9582 16056 9588 16108
rect 9640 16096 9646 16108
rect 13786 16096 13814 16136
rect 15010 16124 15016 16136
rect 15068 16124 15074 16176
rect 16390 16164 16396 16176
rect 16303 16136 16396 16164
rect 16390 16124 16396 16136
rect 16448 16164 16454 16176
rect 19702 16164 19708 16176
rect 16448 16136 19708 16164
rect 16448 16124 16454 16136
rect 19702 16124 19708 16136
rect 19760 16124 19766 16176
rect 9640 16068 13814 16096
rect 14829 16099 14887 16105
rect 9640 16056 9646 16068
rect 14829 16065 14841 16099
rect 14875 16096 14887 16099
rect 15838 16096 15844 16108
rect 14875 16068 15844 16096
rect 14875 16065 14887 16068
rect 14829 16059 14887 16065
rect 15838 16056 15844 16068
rect 15896 16056 15902 16108
rect 18138 16096 18144 16108
rect 18051 16068 18144 16096
rect 18138 16056 18144 16068
rect 18196 16096 18202 16108
rect 18322 16096 18328 16108
rect 18196 16068 18328 16096
rect 18196 16056 18202 16068
rect 18322 16056 18328 16068
rect 18380 16056 18386 16108
rect 18414 16056 18420 16108
rect 18472 16096 18478 16108
rect 18472 16068 18517 16096
rect 18472 16056 18478 16068
rect 1397 16031 1455 16037
rect 1397 15997 1409 16031
rect 1443 16028 1455 16031
rect 1443 16000 2084 16028
rect 1443 15997 1455 16000
rect 1397 15991 1455 15997
rect 2056 15969 2084 16000
rect 2314 15988 2320 16040
rect 2372 16028 2378 16040
rect 2593 16031 2651 16037
rect 2593 16028 2605 16031
rect 2372 16000 2605 16028
rect 2372 15988 2378 16000
rect 2593 15997 2605 16000
rect 2639 15997 2651 16031
rect 3142 16028 3148 16040
rect 3103 16000 3148 16028
rect 2593 15991 2651 15997
rect 3142 15988 3148 16000
rect 3200 15988 3206 16040
rect 4525 16031 4583 16037
rect 4525 15997 4537 16031
rect 4571 16028 4583 16031
rect 4985 16031 5043 16037
rect 4985 16028 4997 16031
rect 4571 16000 4997 16028
rect 4571 15997 4583 16000
rect 4525 15991 4583 15997
rect 4985 15997 4997 16000
rect 5031 16028 5043 16031
rect 5442 16028 5448 16040
rect 5031 16000 5448 16028
rect 5031 15997 5043 16000
rect 4985 15991 5043 15997
rect 5442 15988 5448 16000
rect 5500 15988 5506 16040
rect 10137 16031 10195 16037
rect 10137 15997 10149 16031
rect 10183 16028 10195 16031
rect 10226 16028 10232 16040
rect 10183 16000 10232 16028
rect 10183 15997 10195 16000
rect 10137 15991 10195 15997
rect 10226 15988 10232 16000
rect 10284 16028 10290 16040
rect 10597 16031 10655 16037
rect 10597 16028 10609 16031
rect 10284 16000 10609 16028
rect 10284 15988 10290 16000
rect 10597 15997 10609 16000
rect 10643 15997 10655 16031
rect 10597 15991 10655 15997
rect 10778 15988 10784 16040
rect 10836 16028 10842 16040
rect 11790 16028 11796 16040
rect 10836 16000 11796 16028
rect 10836 15988 10842 16000
rect 11790 15988 11796 16000
rect 11848 15988 11854 16040
rect 12504 16031 12562 16037
rect 12504 15997 12516 16031
rect 12550 16028 12562 16031
rect 12550 16000 13032 16028
rect 12550 15997 12562 16000
rect 12504 15991 12562 15997
rect 2041 15963 2099 15969
rect 2041 15929 2053 15963
rect 2087 15960 2099 15963
rect 3602 15960 3608 15972
rect 2087 15932 3608 15960
rect 2087 15929 2099 15932
rect 2041 15923 2099 15929
rect 3602 15920 3608 15932
rect 3660 15960 3666 15972
rect 4706 15960 4712 15972
rect 3660 15932 4712 15960
rect 3660 15920 3666 15932
rect 4706 15920 4712 15932
rect 4764 15920 4770 15972
rect 4798 15920 4804 15972
rect 4856 15960 4862 15972
rect 5306 15963 5364 15969
rect 5306 15960 5318 15963
rect 4856 15932 5318 15960
rect 4856 15920 4862 15932
rect 5306 15929 5318 15932
rect 5352 15929 5364 15963
rect 6914 15960 6920 15972
rect 6875 15932 6920 15960
rect 5306 15923 5364 15929
rect 6914 15920 6920 15932
rect 6972 15920 6978 15972
rect 7006 15920 7012 15972
rect 7064 15960 7070 15972
rect 7929 15963 7987 15969
rect 7064 15932 7109 15960
rect 7064 15920 7070 15932
rect 7929 15929 7941 15963
rect 7975 15960 7987 15963
rect 8202 15960 8208 15972
rect 7975 15932 8208 15960
rect 7975 15929 7987 15932
rect 7929 15923 7987 15929
rect 8202 15920 8208 15932
rect 8260 15960 8266 15972
rect 8297 15963 8355 15969
rect 8297 15960 8309 15963
rect 8260 15932 8309 15960
rect 8260 15920 8266 15932
rect 8297 15929 8309 15932
rect 8343 15960 8355 15963
rect 8573 15963 8631 15969
rect 8573 15960 8585 15963
rect 8343 15932 8585 15960
rect 8343 15929 8355 15932
rect 8297 15923 8355 15929
rect 8573 15929 8585 15932
rect 8619 15960 8631 15963
rect 8754 15960 8760 15972
rect 8619 15932 8760 15960
rect 8619 15929 8631 15932
rect 8573 15923 8631 15929
rect 8754 15920 8760 15932
rect 8812 15920 8818 15972
rect 9766 15920 9772 15972
rect 9824 15960 9830 15972
rect 12519 15960 12547 15991
rect 9824 15932 12547 15960
rect 9824 15920 9830 15932
rect 8662 15852 8668 15904
rect 8720 15892 8726 15904
rect 9582 15892 9588 15904
rect 8720 15864 9588 15892
rect 8720 15852 8726 15864
rect 9582 15852 9588 15864
rect 9640 15892 9646 15904
rect 9677 15895 9735 15901
rect 9677 15892 9689 15895
rect 9640 15864 9689 15892
rect 9640 15852 9646 15864
rect 9677 15861 9689 15864
rect 9723 15861 9735 15895
rect 10962 15892 10968 15904
rect 10923 15864 10968 15892
rect 9677 15855 9735 15861
rect 10962 15852 10968 15864
rect 11020 15852 11026 15904
rect 13004 15901 13032 16000
rect 15197 15963 15255 15969
rect 15197 15929 15209 15963
rect 15243 15960 15255 15963
rect 15933 15963 15991 15969
rect 15933 15960 15945 15963
rect 15243 15932 15945 15960
rect 15243 15929 15255 15932
rect 15197 15923 15255 15929
rect 15933 15929 15945 15932
rect 15979 15960 15991 15963
rect 16206 15960 16212 15972
rect 15979 15932 16212 15960
rect 15979 15929 15991 15932
rect 15933 15923 15991 15929
rect 16206 15920 16212 15932
rect 16264 15920 16270 15972
rect 17865 15963 17923 15969
rect 17865 15929 17877 15963
rect 17911 15960 17923 15963
rect 18233 15963 18291 15969
rect 18233 15960 18245 15963
rect 17911 15932 18245 15960
rect 17911 15929 17923 15932
rect 17865 15923 17923 15929
rect 18233 15929 18245 15932
rect 18279 15960 18291 15963
rect 18322 15960 18328 15972
rect 18279 15932 18328 15960
rect 18279 15929 18291 15932
rect 18233 15923 18291 15929
rect 18322 15920 18328 15932
rect 18380 15960 18386 15972
rect 18506 15960 18512 15972
rect 18380 15932 18512 15960
rect 18380 15920 18386 15932
rect 18506 15920 18512 15932
rect 18564 15920 18570 15972
rect 20806 15960 20812 15972
rect 19306 15932 20812 15960
rect 12989 15895 13047 15901
rect 12989 15861 13001 15895
rect 13035 15892 13047 15895
rect 13262 15892 13268 15904
rect 13035 15864 13268 15892
rect 13035 15861 13047 15864
rect 12989 15855 13047 15861
rect 13262 15852 13268 15864
rect 13320 15852 13326 15904
rect 13722 15852 13728 15904
rect 13780 15892 13786 15904
rect 16666 15892 16672 15904
rect 13780 15864 16672 15892
rect 13780 15852 13786 15864
rect 16666 15852 16672 15864
rect 16724 15892 16730 15904
rect 16945 15895 17003 15901
rect 16945 15892 16957 15895
rect 16724 15864 16957 15892
rect 16724 15852 16730 15864
rect 16945 15861 16957 15864
rect 16991 15892 17003 15895
rect 17310 15892 17316 15904
rect 16991 15864 17316 15892
rect 16991 15861 17003 15864
rect 16945 15855 17003 15861
rect 17310 15852 17316 15864
rect 17368 15852 17374 15904
rect 17405 15895 17463 15901
rect 17405 15861 17417 15895
rect 17451 15892 17463 15895
rect 17494 15892 17500 15904
rect 17451 15864 17500 15892
rect 17451 15861 17463 15864
rect 17405 15855 17463 15861
rect 17494 15852 17500 15864
rect 17552 15852 17558 15904
rect 17954 15852 17960 15904
rect 18012 15892 18018 15904
rect 19306 15892 19334 15932
rect 20806 15920 20812 15932
rect 20864 15960 20870 15972
rect 20901 15963 20959 15969
rect 20901 15960 20913 15963
rect 20864 15932 20913 15960
rect 20864 15920 20870 15932
rect 20901 15929 20913 15932
rect 20947 15929 20959 15963
rect 20901 15923 20959 15929
rect 18012 15864 19334 15892
rect 18012 15852 18018 15864
rect 1104 15802 22816 15824
rect 1104 15750 8982 15802
rect 9034 15750 9046 15802
rect 9098 15750 9110 15802
rect 9162 15750 9174 15802
rect 9226 15750 16982 15802
rect 17034 15750 17046 15802
rect 17098 15750 17110 15802
rect 17162 15750 17174 15802
rect 17226 15750 22816 15802
rect 1104 15728 22816 15750
rect 1946 15688 1952 15700
rect 1907 15660 1952 15688
rect 1946 15648 1952 15660
rect 2004 15648 2010 15700
rect 4847 15691 4905 15697
rect 4847 15657 4859 15691
rect 4893 15688 4905 15691
rect 6914 15688 6920 15700
rect 4893 15660 6920 15688
rect 4893 15657 4905 15660
rect 4847 15651 4905 15657
rect 6914 15648 6920 15660
rect 6972 15648 6978 15700
rect 8754 15688 8760 15700
rect 8715 15660 8760 15688
rect 8754 15648 8760 15660
rect 8812 15648 8818 15700
rect 9125 15691 9183 15697
rect 9125 15657 9137 15691
rect 9171 15688 9183 15691
rect 9306 15688 9312 15700
rect 9171 15660 9312 15688
rect 9171 15657 9183 15660
rect 9125 15651 9183 15657
rect 9306 15648 9312 15660
rect 9364 15648 9370 15700
rect 10226 15688 10232 15700
rect 10187 15660 10232 15688
rect 10226 15648 10232 15660
rect 10284 15648 10290 15700
rect 15654 15688 15660 15700
rect 15615 15660 15660 15688
rect 15654 15648 15660 15660
rect 15712 15648 15718 15700
rect 16206 15688 16212 15700
rect 16167 15660 16212 15688
rect 16206 15648 16212 15660
rect 16264 15648 16270 15700
rect 17175 15691 17233 15697
rect 17175 15657 17187 15691
rect 17221 15688 17233 15691
rect 18138 15688 18144 15700
rect 17221 15660 18144 15688
rect 17221 15657 17233 15660
rect 17175 15651 17233 15657
rect 18138 15648 18144 15660
rect 18196 15648 18202 15700
rect 21039 15691 21097 15697
rect 21039 15657 21051 15691
rect 21085 15688 21097 15691
rect 22002 15688 22008 15700
rect 21085 15660 22008 15688
rect 21085 15657 21097 15660
rect 21039 15651 21097 15657
rect 22002 15648 22008 15660
rect 22060 15648 22066 15700
rect 1302 15580 1308 15632
rect 1360 15620 1366 15632
rect 1535 15623 1593 15629
rect 1535 15620 1547 15623
rect 1360 15592 1547 15620
rect 1360 15580 1366 15592
rect 1535 15589 1547 15592
rect 1581 15589 1593 15623
rect 1535 15583 1593 15589
rect 5261 15623 5319 15629
rect 5261 15589 5273 15623
rect 5307 15620 5319 15623
rect 5534 15620 5540 15632
rect 5307 15592 5540 15620
rect 5307 15589 5319 15592
rect 5261 15583 5319 15589
rect 5534 15580 5540 15592
rect 5592 15580 5598 15632
rect 8199 15623 8257 15629
rect 8199 15589 8211 15623
rect 8245 15620 8257 15623
rect 8478 15620 8484 15632
rect 8245 15592 8484 15620
rect 8245 15589 8257 15592
rect 8199 15583 8257 15589
rect 8478 15580 8484 15592
rect 8536 15580 8542 15632
rect 18334 15623 18392 15629
rect 18334 15589 18346 15623
rect 18380 15620 18392 15623
rect 18506 15620 18512 15632
rect 18380 15592 18512 15620
rect 18380 15589 18392 15592
rect 18334 15583 18392 15589
rect 18506 15580 18512 15592
rect 18564 15580 18570 15632
rect 18877 15623 18935 15629
rect 18877 15589 18889 15623
rect 18923 15620 18935 15623
rect 19702 15620 19708 15632
rect 18923 15592 19708 15620
rect 18923 15589 18935 15592
rect 18877 15583 18935 15589
rect 19702 15580 19708 15592
rect 19760 15580 19766 15632
rect 1448 15555 1506 15561
rect 1448 15521 1460 15555
rect 1494 15552 1506 15555
rect 2130 15552 2136 15564
rect 1494 15524 2136 15552
rect 1494 15521 1506 15524
rect 1448 15515 1506 15521
rect 2130 15512 2136 15524
rect 2188 15552 2194 15564
rect 3050 15552 3056 15564
rect 2188 15524 3056 15552
rect 2188 15512 2194 15524
rect 3050 15512 3056 15524
rect 3108 15512 3114 15564
rect 4617 15555 4675 15561
rect 4617 15521 4629 15555
rect 4663 15552 4675 15555
rect 4798 15552 4804 15564
rect 4663 15524 4804 15552
rect 4663 15521 4675 15524
rect 4617 15515 4675 15521
rect 4798 15512 4804 15524
rect 4856 15512 4862 15564
rect 5994 15552 6000 15564
rect 5955 15524 6000 15552
rect 5994 15512 6000 15524
rect 6052 15512 6058 15564
rect 6178 15552 6184 15564
rect 6139 15524 6184 15552
rect 6178 15512 6184 15524
rect 6236 15512 6242 15564
rect 10229 15555 10287 15561
rect 10229 15521 10241 15555
rect 10275 15521 10287 15555
rect 10410 15552 10416 15564
rect 10371 15524 10416 15552
rect 10229 15515 10287 15521
rect 6454 15484 6460 15496
rect 6415 15456 6460 15484
rect 6454 15444 6460 15456
rect 6512 15444 6518 15496
rect 7834 15484 7840 15496
rect 7795 15456 7840 15484
rect 7834 15444 7840 15456
rect 7892 15444 7898 15496
rect 10244 15484 10272 15515
rect 10410 15512 10416 15524
rect 10468 15512 10474 15564
rect 11952 15555 12010 15561
rect 11952 15521 11964 15555
rect 11998 15552 12010 15555
rect 12066 15552 12072 15564
rect 11998 15524 12072 15552
rect 11998 15521 12010 15524
rect 11952 15515 12010 15521
rect 12066 15512 12072 15524
rect 12124 15512 12130 15564
rect 13357 15555 13415 15561
rect 13357 15521 13369 15555
rect 13403 15552 13415 15555
rect 13538 15552 13544 15564
rect 13403 15524 13544 15552
rect 13403 15521 13415 15524
rect 13357 15515 13415 15521
rect 13538 15512 13544 15524
rect 13596 15512 13602 15564
rect 17126 15561 17132 15564
rect 17104 15555 17132 15561
rect 17104 15521 17116 15555
rect 17184 15552 17190 15564
rect 17954 15552 17960 15564
rect 17184 15524 17960 15552
rect 17104 15515 17132 15521
rect 17126 15512 17132 15515
rect 17184 15512 17190 15524
rect 17954 15512 17960 15524
rect 18012 15512 18018 15564
rect 20806 15512 20812 15564
rect 20864 15552 20870 15564
rect 20936 15555 20994 15561
rect 20936 15552 20948 15555
rect 20864 15524 20948 15552
rect 20864 15512 20870 15524
rect 20936 15521 20948 15524
rect 20982 15521 20994 15555
rect 20936 15515 20994 15521
rect 10594 15484 10600 15496
rect 10244 15456 10600 15484
rect 10594 15444 10600 15456
rect 10652 15444 10658 15496
rect 12529 15487 12587 15493
rect 12529 15453 12541 15487
rect 12575 15484 12587 15487
rect 12618 15484 12624 15496
rect 12575 15456 12624 15484
rect 12575 15453 12587 15456
rect 12529 15447 12587 15453
rect 12618 15444 12624 15456
rect 12676 15444 12682 15496
rect 14734 15444 14740 15496
rect 14792 15484 14798 15496
rect 15289 15487 15347 15493
rect 15289 15484 15301 15487
rect 14792 15456 15301 15484
rect 14792 15444 14798 15456
rect 15289 15453 15301 15456
rect 15335 15453 15347 15487
rect 15289 15447 15347 15453
rect 18233 15487 18291 15493
rect 18233 15453 18245 15487
rect 18279 15484 18291 15487
rect 18690 15484 18696 15496
rect 18279 15456 18696 15484
rect 18279 15453 18291 15456
rect 18233 15447 18291 15453
rect 18690 15444 18696 15456
rect 18748 15444 18754 15496
rect 1670 15376 1676 15428
rect 1728 15416 1734 15428
rect 2225 15419 2283 15425
rect 2225 15416 2237 15419
rect 1728 15388 2237 15416
rect 1728 15376 1734 15388
rect 2225 15385 2237 15388
rect 2271 15385 2283 15419
rect 2225 15379 2283 15385
rect 7193 15419 7251 15425
rect 7193 15385 7205 15419
rect 7239 15416 7251 15419
rect 7926 15416 7932 15428
rect 7239 15388 7932 15416
rect 7239 15385 7251 15388
rect 7193 15379 7251 15385
rect 7926 15376 7932 15388
rect 7984 15376 7990 15428
rect 12023 15419 12081 15425
rect 12023 15385 12035 15419
rect 12069 15416 12081 15419
rect 13587 15419 13645 15425
rect 12069 15388 12572 15416
rect 12069 15385 12081 15388
rect 12023 15379 12081 15385
rect 12544 15360 12572 15388
rect 13587 15385 13599 15419
rect 13633 15416 13645 15419
rect 16114 15416 16120 15428
rect 13633 15388 16120 15416
rect 13633 15385 13645 15388
rect 13587 15379 13645 15385
rect 16114 15376 16120 15388
rect 16172 15376 16178 15428
rect 2314 15308 2320 15360
rect 2372 15348 2378 15360
rect 2593 15351 2651 15357
rect 2593 15348 2605 15351
rect 2372 15320 2605 15348
rect 2372 15308 2378 15320
rect 2593 15317 2605 15320
rect 2639 15317 2651 15351
rect 2593 15311 2651 15317
rect 7561 15351 7619 15357
rect 7561 15317 7573 15351
rect 7607 15348 7619 15351
rect 7650 15348 7656 15360
rect 7607 15320 7656 15348
rect 7607 15317 7619 15320
rect 7561 15311 7619 15317
rect 7650 15308 7656 15320
rect 7708 15308 7714 15360
rect 12526 15308 12532 15360
rect 12584 15348 12590 15360
rect 12805 15351 12863 15357
rect 12805 15348 12817 15351
rect 12584 15320 12817 15348
rect 12584 15308 12590 15320
rect 12805 15317 12817 15320
rect 12851 15317 12863 15351
rect 13998 15348 14004 15360
rect 13959 15320 14004 15348
rect 12805 15311 12863 15317
rect 13998 15308 14004 15320
rect 14056 15308 14062 15360
rect 16482 15348 16488 15360
rect 16443 15320 16488 15348
rect 16482 15308 16488 15320
rect 16540 15308 16546 15360
rect 19518 15348 19524 15360
rect 19479 15320 19524 15348
rect 19518 15308 19524 15320
rect 19576 15308 19582 15360
rect 1104 15258 22816 15280
rect 1104 15206 4982 15258
rect 5034 15206 5046 15258
rect 5098 15206 5110 15258
rect 5162 15206 5174 15258
rect 5226 15206 12982 15258
rect 13034 15206 13046 15258
rect 13098 15206 13110 15258
rect 13162 15206 13174 15258
rect 13226 15206 20982 15258
rect 21034 15206 21046 15258
rect 21098 15206 21110 15258
rect 21162 15206 21174 15258
rect 21226 15206 22816 15258
rect 1104 15184 22816 15206
rect 3050 15144 3056 15156
rect 3011 15116 3056 15144
rect 3050 15104 3056 15116
rect 3108 15104 3114 15156
rect 5534 15104 5540 15156
rect 5592 15144 5598 15156
rect 5902 15144 5908 15156
rect 5592 15116 5908 15144
rect 5592 15104 5598 15116
rect 5902 15104 5908 15116
rect 5960 15144 5966 15156
rect 7285 15147 7343 15153
rect 7285 15144 7297 15147
rect 5960 15116 7297 15144
rect 5960 15104 5966 15116
rect 7285 15113 7297 15116
rect 7331 15113 7343 15147
rect 7285 15107 7343 15113
rect 9401 15147 9459 15153
rect 9401 15113 9413 15147
rect 9447 15144 9459 15147
rect 9766 15144 9772 15156
rect 9447 15116 9772 15144
rect 9447 15113 9459 15116
rect 9401 15107 9459 15113
rect 6178 15008 6184 15020
rect 4172 14980 6184 15008
rect 2314 14940 2320 14952
rect 2275 14912 2320 14940
rect 2314 14900 2320 14912
rect 2372 14900 2378 14952
rect 2593 14943 2651 14949
rect 2593 14909 2605 14943
rect 2639 14909 2651 14943
rect 2593 14903 2651 14909
rect 1946 14804 1952 14816
rect 1907 14776 1952 14804
rect 1946 14764 1952 14776
rect 2004 14804 2010 14816
rect 2608 14804 2636 14903
rect 3418 14900 3424 14952
rect 3476 14940 3482 14952
rect 4172 14949 4200 14980
rect 6178 14968 6184 14980
rect 6236 14968 6242 15020
rect 7300 15008 7328 15107
rect 9766 15104 9772 15116
rect 9824 15104 9830 15156
rect 13538 15144 13544 15156
rect 13499 15116 13544 15144
rect 13538 15104 13544 15116
rect 13596 15104 13602 15156
rect 16945 15147 17003 15153
rect 16945 15113 16957 15147
rect 16991 15144 17003 15147
rect 18233 15147 18291 15153
rect 18233 15144 18245 15147
rect 16991 15116 18245 15144
rect 16991 15113 17003 15116
rect 16945 15107 17003 15113
rect 18233 15113 18245 15116
rect 18279 15144 18291 15147
rect 18322 15144 18328 15156
rect 18279 15116 18328 15144
rect 18279 15113 18291 15116
rect 18233 15107 18291 15113
rect 18322 15104 18328 15116
rect 18380 15104 18386 15156
rect 20806 15104 20812 15156
rect 20864 15144 20870 15156
rect 20901 15147 20959 15153
rect 20901 15144 20913 15147
rect 20864 15116 20913 15144
rect 20864 15104 20870 15116
rect 20901 15113 20913 15116
rect 20947 15113 20959 15147
rect 20901 15107 20959 15113
rect 8202 15036 8208 15088
rect 8260 15076 8266 15088
rect 9490 15076 9496 15088
rect 8260 15048 9496 15076
rect 8260 15036 8266 15048
rect 9490 15036 9496 15048
rect 9548 15036 9554 15088
rect 7300 14980 7788 15008
rect 3605 14943 3663 14949
rect 3605 14940 3617 14943
rect 3476 14912 3617 14940
rect 3476 14900 3482 14912
rect 3605 14909 3617 14912
rect 3651 14909 3663 14943
rect 3605 14903 3663 14909
rect 4157 14943 4215 14949
rect 4157 14909 4169 14943
rect 4203 14909 4215 14943
rect 4157 14903 4215 14909
rect 5445 14943 5503 14949
rect 5445 14909 5457 14943
rect 5491 14909 5503 14943
rect 5445 14903 5503 14909
rect 2774 14872 2780 14884
rect 2735 14844 2780 14872
rect 2774 14832 2780 14844
rect 2832 14832 2838 14884
rect 4172 14872 4200 14903
rect 3436 14844 4200 14872
rect 3436 14813 3464 14844
rect 5350 14832 5356 14884
rect 5408 14872 5414 14884
rect 5460 14872 5488 14903
rect 5534 14900 5540 14952
rect 5592 14940 5598 14952
rect 5629 14943 5687 14949
rect 5629 14940 5641 14943
rect 5592 14912 5641 14940
rect 5592 14900 5598 14912
rect 5629 14909 5641 14912
rect 5675 14909 5687 14943
rect 7650 14940 7656 14952
rect 7611 14912 7656 14940
rect 5629 14903 5687 14909
rect 7650 14900 7656 14912
rect 7708 14900 7714 14952
rect 7760 14940 7788 14980
rect 7834 14968 7840 15020
rect 7892 15008 7898 15020
rect 8021 15011 8079 15017
rect 8021 15008 8033 15011
rect 7892 14980 8033 15008
rect 7892 14968 7898 14980
rect 8021 14977 8033 14980
rect 8067 14977 8079 15011
rect 12526 15008 12532 15020
rect 12487 14980 12532 15008
rect 8021 14971 8079 14977
rect 12526 14968 12532 14980
rect 12584 14968 12590 15020
rect 7929 14943 7987 14949
rect 7929 14940 7941 14943
rect 7760 14912 7941 14940
rect 7929 14909 7941 14912
rect 7975 14909 7987 14943
rect 7929 14903 7987 14909
rect 9033 14943 9091 14949
rect 9033 14909 9045 14943
rect 9079 14940 9091 14943
rect 9490 14940 9496 14952
rect 9079 14912 9496 14940
rect 9079 14909 9091 14912
rect 9033 14903 9091 14909
rect 5994 14872 6000 14884
rect 5408 14844 6000 14872
rect 5408 14832 5414 14844
rect 5994 14832 6000 14844
rect 6052 14872 6058 14884
rect 6641 14875 6699 14881
rect 6641 14872 6653 14875
rect 6052 14844 6653 14872
rect 6052 14832 6058 14844
rect 6641 14841 6653 14844
rect 6687 14872 6699 14875
rect 9048 14872 9076 14903
rect 9490 14900 9496 14912
rect 9548 14900 9554 14952
rect 9766 14900 9772 14952
rect 9824 14940 9830 14952
rect 9953 14943 10011 14949
rect 9953 14940 9965 14943
rect 9824 14912 9965 14940
rect 9824 14900 9830 14912
rect 9953 14909 9965 14912
rect 9999 14940 10011 14943
rect 10410 14940 10416 14952
rect 9999 14912 10416 14940
rect 9999 14909 10011 14912
rect 9953 14903 10011 14909
rect 10410 14900 10416 14912
rect 10468 14940 10474 14952
rect 10505 14943 10563 14949
rect 10505 14940 10517 14943
rect 10468 14912 10517 14940
rect 10468 14900 10474 14912
rect 10505 14909 10517 14912
rect 10551 14909 10563 14943
rect 11238 14940 11244 14952
rect 11199 14912 11244 14940
rect 10505 14903 10563 14909
rect 11238 14900 11244 14912
rect 11296 14940 11302 14952
rect 11368 14943 11426 14949
rect 11368 14940 11380 14943
rect 11296 14912 11380 14940
rect 11296 14900 11302 14912
rect 11368 14909 11380 14912
rect 11414 14909 11426 14943
rect 13998 14940 14004 14952
rect 13959 14912 14004 14940
rect 11368 14903 11426 14909
rect 13998 14900 14004 14912
rect 14056 14900 14062 14952
rect 14550 14940 14556 14952
rect 14511 14912 14556 14940
rect 14550 14900 14556 14912
rect 14608 14900 14614 14952
rect 15470 14900 15476 14952
rect 15528 14940 15534 14952
rect 16025 14943 16083 14949
rect 16025 14940 16037 14943
rect 15528 14912 16037 14940
rect 15528 14900 15534 14912
rect 16025 14909 16037 14912
rect 16071 14940 16083 14943
rect 16482 14940 16488 14952
rect 16071 14912 16488 14940
rect 16071 14909 16083 14912
rect 16025 14903 16083 14909
rect 16482 14900 16488 14912
rect 16540 14900 16546 14952
rect 18598 14900 18604 14952
rect 18656 14940 18662 14952
rect 19518 14940 19524 14952
rect 18656 14912 19524 14940
rect 18656 14900 18662 14912
rect 19518 14900 19524 14912
rect 19576 14900 19582 14952
rect 10226 14872 10232 14884
rect 6687 14844 9076 14872
rect 10187 14844 10232 14872
rect 6687 14841 6699 14844
rect 6641 14835 6699 14841
rect 10226 14832 10232 14844
rect 10284 14832 10290 14884
rect 12618 14872 12624 14884
rect 12579 14844 12624 14872
rect 12618 14832 12624 14844
rect 12676 14832 12682 14884
rect 13173 14875 13231 14881
rect 13173 14841 13185 14875
rect 13219 14872 13231 14875
rect 13814 14872 13820 14884
rect 13219 14844 13820 14872
rect 13219 14841 13231 14844
rect 13173 14835 13231 14841
rect 13814 14832 13820 14844
rect 13872 14832 13878 14884
rect 13909 14875 13967 14881
rect 13909 14841 13921 14875
rect 13955 14872 13967 14875
rect 14568 14872 14596 14900
rect 14734 14872 14740 14884
rect 13955 14844 14596 14872
rect 14695 14844 14740 14872
rect 13955 14841 13967 14844
rect 13909 14835 13967 14841
rect 3421 14807 3479 14813
rect 3421 14804 3433 14807
rect 2004 14776 3433 14804
rect 2004 14764 2010 14776
rect 3421 14773 3433 14776
rect 3467 14773 3479 14807
rect 3878 14804 3884 14816
rect 3839 14776 3884 14804
rect 3421 14767 3479 14773
rect 3878 14764 3884 14776
rect 3936 14764 3942 14816
rect 4798 14804 4804 14816
rect 4759 14776 4804 14804
rect 4798 14764 4804 14776
rect 4856 14764 4862 14816
rect 5442 14804 5448 14816
rect 5403 14776 5448 14804
rect 5442 14764 5448 14776
rect 5500 14764 5506 14816
rect 8478 14764 8484 14816
rect 8536 14804 8542 14816
rect 8573 14807 8631 14813
rect 8573 14804 8585 14807
rect 8536 14776 8585 14804
rect 8536 14764 8542 14776
rect 8573 14773 8585 14776
rect 8619 14804 8631 14807
rect 10962 14804 10968 14816
rect 8619 14776 10968 14804
rect 8619 14773 8631 14776
rect 8573 14767 8631 14773
rect 10962 14764 10968 14776
rect 11020 14764 11026 14816
rect 11471 14807 11529 14813
rect 11471 14773 11483 14807
rect 11517 14804 11529 14807
rect 11882 14804 11888 14816
rect 11517 14776 11888 14804
rect 11517 14773 11529 14776
rect 11471 14767 11529 14773
rect 11882 14764 11888 14776
rect 11940 14764 11946 14816
rect 11977 14807 12035 14813
rect 11977 14773 11989 14807
rect 12023 14804 12035 14807
rect 12066 14804 12072 14816
rect 12023 14776 12072 14804
rect 12023 14773 12035 14776
rect 11977 14767 12035 14773
rect 12066 14764 12072 14776
rect 12124 14764 12130 14816
rect 13722 14764 13728 14816
rect 13780 14804 13786 14816
rect 13924 14804 13952 14835
rect 14734 14832 14740 14844
rect 14792 14832 14798 14884
rect 16346 14875 16404 14881
rect 16346 14872 16358 14875
rect 15856 14844 16358 14872
rect 13780 14776 13952 14804
rect 13780 14764 13786 14776
rect 14642 14764 14648 14816
rect 14700 14804 14706 14816
rect 15289 14807 15347 14813
rect 15289 14804 15301 14807
rect 14700 14776 15301 14804
rect 14700 14764 14706 14776
rect 15289 14773 15301 14776
rect 15335 14804 15347 14807
rect 15654 14804 15660 14816
rect 15335 14776 15660 14804
rect 15335 14773 15347 14776
rect 15289 14767 15347 14773
rect 15654 14764 15660 14776
rect 15712 14804 15718 14816
rect 15856 14813 15884 14844
rect 16346 14841 16358 14844
rect 16392 14841 16404 14875
rect 16346 14835 16404 14841
rect 16574 14832 16580 14884
rect 16632 14872 16638 14884
rect 17126 14872 17132 14884
rect 16632 14844 17132 14872
rect 16632 14832 16638 14844
rect 17126 14832 17132 14844
rect 17184 14872 17190 14884
rect 17221 14875 17279 14881
rect 17221 14872 17233 14875
rect 17184 14844 17233 14872
rect 17184 14832 17190 14844
rect 17221 14841 17233 14844
rect 17267 14841 17279 14875
rect 17221 14835 17279 14841
rect 15841 14807 15899 14813
rect 15841 14804 15853 14807
rect 15712 14776 15853 14804
rect 15712 14764 15718 14776
rect 15841 14773 15853 14776
rect 15887 14773 15899 14807
rect 18690 14804 18696 14816
rect 18651 14776 18696 14804
rect 15841 14767 15899 14773
rect 18690 14764 18696 14776
rect 18748 14764 18754 14816
rect 19426 14804 19432 14816
rect 19339 14776 19432 14804
rect 19426 14764 19432 14776
rect 19484 14804 19490 14816
rect 19889 14807 19947 14813
rect 19889 14804 19901 14807
rect 19484 14776 19901 14804
rect 19484 14764 19490 14776
rect 19889 14773 19901 14776
rect 19935 14773 19947 14807
rect 20438 14804 20444 14816
rect 20399 14776 20444 14804
rect 19889 14767 19947 14773
rect 20438 14764 20444 14776
rect 20496 14764 20502 14816
rect 20990 14764 20996 14816
rect 21048 14804 21054 14816
rect 21269 14807 21327 14813
rect 21269 14804 21281 14807
rect 21048 14776 21281 14804
rect 21048 14764 21054 14776
rect 21269 14773 21281 14776
rect 21315 14773 21327 14807
rect 21269 14767 21327 14773
rect 1104 14714 22816 14736
rect 1104 14662 8982 14714
rect 9034 14662 9046 14714
rect 9098 14662 9110 14714
rect 9162 14662 9174 14714
rect 9226 14662 16982 14714
rect 17034 14662 17046 14714
rect 17098 14662 17110 14714
rect 17162 14662 17174 14714
rect 17226 14662 22816 14714
rect 1104 14640 22816 14662
rect 2590 14600 2596 14612
rect 2551 14572 2596 14600
rect 2590 14560 2596 14572
rect 2648 14560 2654 14612
rect 3418 14560 3424 14612
rect 3476 14600 3482 14612
rect 3605 14603 3663 14609
rect 3605 14600 3617 14603
rect 3476 14572 3617 14600
rect 3476 14560 3482 14572
rect 3605 14569 3617 14572
rect 3651 14600 3663 14603
rect 3694 14600 3700 14612
rect 3651 14572 3700 14600
rect 3651 14569 3663 14572
rect 3605 14563 3663 14569
rect 3694 14560 3700 14572
rect 3752 14560 3758 14612
rect 4154 14560 4160 14612
rect 4212 14600 4218 14612
rect 4433 14603 4491 14609
rect 4433 14600 4445 14603
rect 4212 14572 4445 14600
rect 4212 14560 4218 14572
rect 4433 14569 4445 14572
rect 4479 14569 4491 14603
rect 5350 14600 5356 14612
rect 5311 14572 5356 14600
rect 4433 14563 4491 14569
rect 5350 14560 5356 14572
rect 5408 14560 5414 14612
rect 7834 14600 7840 14612
rect 6891 14572 7696 14600
rect 7795 14572 7840 14600
rect 2133 14535 2191 14541
rect 2133 14501 2145 14535
rect 2179 14532 2191 14535
rect 2314 14532 2320 14544
rect 2179 14504 2320 14532
rect 2179 14501 2191 14504
rect 2133 14495 2191 14501
rect 2314 14492 2320 14504
rect 2372 14532 2378 14544
rect 6891 14532 6919 14572
rect 7006 14532 7012 14544
rect 2372 14504 6919 14532
rect 6967 14504 7012 14532
rect 2372 14492 2378 14504
rect 7006 14492 7012 14504
rect 7064 14492 7070 14544
rect 7668 14532 7696 14572
rect 7834 14560 7840 14572
rect 7892 14560 7898 14612
rect 7926 14560 7932 14612
rect 7984 14600 7990 14612
rect 8711 14603 8769 14609
rect 8711 14600 8723 14603
rect 7984 14572 8723 14600
rect 7984 14560 7990 14572
rect 8711 14569 8723 14572
rect 8757 14569 8769 14603
rect 12802 14600 12808 14612
rect 8711 14563 8769 14569
rect 12176 14572 12808 14600
rect 10591 14535 10649 14541
rect 7668 14504 9674 14532
rect 3878 14424 3884 14476
rect 3936 14464 3942 14476
rect 4065 14467 4123 14473
rect 4065 14464 4077 14467
rect 3936 14436 4077 14464
rect 3936 14424 3942 14436
rect 4065 14433 4077 14436
rect 4111 14433 4123 14467
rect 4065 14427 4123 14433
rect 8640 14467 8698 14473
rect 8640 14433 8652 14467
rect 8686 14464 8698 14467
rect 8754 14464 8760 14476
rect 8686 14436 8760 14464
rect 8686 14433 8698 14436
rect 8640 14427 8698 14433
rect 8754 14424 8760 14436
rect 8812 14424 8818 14476
rect 2225 14399 2283 14405
rect 2225 14365 2237 14399
rect 2271 14396 2283 14399
rect 2774 14396 2780 14408
rect 2271 14368 2780 14396
rect 2271 14365 2283 14368
rect 2225 14359 2283 14365
rect 2774 14356 2780 14368
rect 2832 14356 2838 14408
rect 6917 14399 6975 14405
rect 6917 14365 6929 14399
rect 6963 14365 6975 14399
rect 6917 14359 6975 14365
rect 3145 14331 3203 14337
rect 3145 14297 3157 14331
rect 3191 14328 3203 14331
rect 3786 14328 3792 14340
rect 3191 14300 3792 14328
rect 3191 14297 3203 14300
rect 3145 14291 3203 14297
rect 3786 14288 3792 14300
rect 3844 14288 3850 14340
rect 1578 14260 1584 14272
rect 1539 14232 1584 14260
rect 1578 14220 1584 14232
rect 1636 14220 1642 14272
rect 4522 14220 4528 14272
rect 4580 14260 4586 14272
rect 4985 14263 5043 14269
rect 4985 14260 4997 14263
rect 4580 14232 4997 14260
rect 4580 14220 4586 14232
rect 4985 14229 4997 14232
rect 5031 14229 5043 14263
rect 4985 14223 5043 14229
rect 6362 14220 6368 14272
rect 6420 14260 6426 14272
rect 6641 14263 6699 14269
rect 6641 14260 6653 14263
rect 6420 14232 6653 14260
rect 6420 14220 6426 14232
rect 6641 14229 6653 14232
rect 6687 14260 6699 14263
rect 6932 14260 6960 14359
rect 7466 14328 7472 14340
rect 7427 14300 7472 14328
rect 7466 14288 7472 14300
rect 7524 14288 7530 14340
rect 6687 14232 6960 14260
rect 9646 14260 9674 14504
rect 10591 14501 10603 14535
rect 10637 14532 10649 14535
rect 10962 14532 10968 14544
rect 10637 14504 10968 14532
rect 10637 14501 10649 14504
rect 10591 14495 10649 14501
rect 10962 14492 10968 14504
rect 11020 14492 11026 14544
rect 11882 14492 11888 14544
rect 11940 14532 11946 14544
rect 12176 14541 12204 14572
rect 12802 14560 12808 14572
rect 12860 14560 12866 14612
rect 14734 14560 14740 14612
rect 14792 14600 14798 14612
rect 15473 14603 15531 14609
rect 15473 14600 15485 14603
rect 14792 14572 15485 14600
rect 14792 14560 14798 14572
rect 15473 14569 15485 14572
rect 15519 14569 15531 14603
rect 15473 14563 15531 14569
rect 17402 14560 17408 14612
rect 17460 14600 17466 14612
rect 18506 14600 18512 14612
rect 17460 14572 18512 14600
rect 17460 14560 17466 14572
rect 18506 14560 18512 14572
rect 18564 14560 18570 14612
rect 18690 14560 18696 14612
rect 18748 14600 18754 14612
rect 19567 14603 19625 14609
rect 19567 14600 19579 14603
rect 18748 14572 19579 14600
rect 18748 14560 18754 14572
rect 19567 14569 19579 14572
rect 19613 14569 19625 14603
rect 19567 14563 19625 14569
rect 20438 14560 20444 14612
rect 20496 14600 20502 14612
rect 20496 14572 21128 14600
rect 20496 14560 20502 14572
rect 12161 14535 12219 14541
rect 12161 14532 12173 14535
rect 11940 14504 12173 14532
rect 11940 14492 11946 14504
rect 12161 14501 12173 14504
rect 12207 14501 12219 14535
rect 12161 14495 12219 14501
rect 12250 14492 12256 14544
rect 12308 14532 12314 14544
rect 12618 14532 12624 14544
rect 12308 14504 12624 14532
rect 12308 14492 12314 14504
rect 12618 14492 12624 14504
rect 12676 14492 12682 14544
rect 13814 14492 13820 14544
rect 13872 14532 13878 14544
rect 15838 14532 15844 14544
rect 13872 14504 13917 14532
rect 15751 14504 15844 14532
rect 13872 14492 13878 14504
rect 15838 14492 15844 14504
rect 15896 14532 15902 14544
rect 16206 14532 16212 14544
rect 15896 14504 16212 14532
rect 15896 14492 15902 14504
rect 16206 14492 16212 14504
rect 16264 14492 16270 14544
rect 16393 14535 16451 14541
rect 16393 14501 16405 14535
rect 16439 14532 16451 14535
rect 18414 14532 18420 14544
rect 16439 14504 18420 14532
rect 16439 14501 16451 14504
rect 16393 14495 16451 14501
rect 18414 14492 18420 14504
rect 18472 14492 18478 14544
rect 18598 14532 18604 14544
rect 18559 14504 18604 14532
rect 18598 14492 18604 14504
rect 18656 14492 18662 14544
rect 20714 14492 20720 14544
rect 20772 14532 20778 14544
rect 20990 14532 20996 14544
rect 20772 14504 20996 14532
rect 20772 14492 20778 14504
rect 20990 14492 20996 14504
rect 21048 14492 21054 14544
rect 21100 14541 21128 14572
rect 21085 14535 21143 14541
rect 21085 14501 21097 14535
rect 21131 14532 21143 14535
rect 22186 14532 22192 14544
rect 21131 14504 22192 14532
rect 21131 14501 21143 14504
rect 21085 14495 21143 14501
rect 22186 14492 22192 14504
rect 22244 14492 22250 14544
rect 10226 14464 10232 14476
rect 10187 14436 10232 14464
rect 10226 14424 10232 14436
rect 10284 14424 10290 14476
rect 17862 14464 17868 14476
rect 17823 14436 17868 14464
rect 17862 14424 17868 14436
rect 17920 14424 17926 14476
rect 18325 14467 18383 14473
rect 18325 14433 18337 14467
rect 18371 14433 18383 14467
rect 18325 14427 18383 14433
rect 19496 14467 19554 14473
rect 19496 14433 19508 14467
rect 19542 14464 19554 14467
rect 20346 14464 20352 14476
rect 19542 14436 20352 14464
rect 19542 14433 19554 14436
rect 19496 14427 19554 14433
rect 12434 14396 12440 14408
rect 12395 14368 12440 14396
rect 12434 14356 12440 14368
rect 12492 14356 12498 14408
rect 13722 14396 13728 14408
rect 13683 14368 13728 14396
rect 13722 14356 13728 14368
rect 13780 14356 13786 14408
rect 13906 14356 13912 14408
rect 13964 14396 13970 14408
rect 14001 14399 14059 14405
rect 14001 14396 14013 14399
rect 13964 14368 14013 14396
rect 13964 14356 13970 14368
rect 14001 14365 14013 14368
rect 14047 14365 14059 14399
rect 15746 14396 15752 14408
rect 15707 14368 15752 14396
rect 14001 14359 14059 14365
rect 15746 14356 15752 14368
rect 15804 14356 15810 14408
rect 17494 14356 17500 14408
rect 17552 14396 17558 14408
rect 18340 14396 18368 14427
rect 20346 14424 20352 14436
rect 20404 14424 20410 14476
rect 17552 14368 18368 14396
rect 17552 14356 17558 14368
rect 20806 14356 20812 14408
rect 20864 14396 20870 14408
rect 21266 14396 21272 14408
rect 20864 14368 21272 14396
rect 20864 14356 20870 14368
rect 21266 14356 21272 14368
rect 21324 14356 21330 14408
rect 11149 14331 11207 14337
rect 11149 14297 11161 14331
rect 11195 14328 11207 14331
rect 12250 14328 12256 14340
rect 11195 14300 12256 14328
rect 11195 14297 11207 14300
rect 11149 14291 11207 14297
rect 12250 14288 12256 14300
rect 12308 14288 12314 14340
rect 10045 14263 10103 14269
rect 10045 14260 10057 14263
rect 9646 14232 10057 14260
rect 6687 14229 6699 14232
rect 6641 14223 6699 14229
rect 10045 14229 10057 14232
rect 10091 14260 10103 14263
rect 10594 14260 10600 14272
rect 10091 14232 10600 14260
rect 10091 14229 10103 14232
rect 10045 14223 10103 14229
rect 10594 14220 10600 14232
rect 10652 14220 10658 14272
rect 19058 14260 19064 14272
rect 19019 14232 19064 14260
rect 19058 14220 19064 14232
rect 19116 14220 19122 14272
rect 1104 14170 22816 14192
rect 1104 14118 4982 14170
rect 5034 14118 5046 14170
rect 5098 14118 5110 14170
rect 5162 14118 5174 14170
rect 5226 14118 12982 14170
rect 13034 14118 13046 14170
rect 13098 14118 13110 14170
rect 13162 14118 13174 14170
rect 13226 14118 20982 14170
rect 21034 14118 21046 14170
rect 21098 14118 21110 14170
rect 21162 14118 21174 14170
rect 21226 14118 22816 14170
rect 1104 14096 22816 14118
rect 2590 14056 2596 14068
rect 2551 14028 2596 14056
rect 2590 14016 2596 14028
rect 2648 14016 2654 14068
rect 2774 14016 2780 14068
rect 2832 14056 2838 14068
rect 2869 14059 2927 14065
rect 2869 14056 2881 14059
rect 2832 14028 2881 14056
rect 2832 14016 2838 14028
rect 2869 14025 2881 14028
rect 2915 14025 2927 14059
rect 2869 14019 2927 14025
rect 3605 14059 3663 14065
rect 3605 14025 3617 14059
rect 3651 14056 3663 14059
rect 3878 14056 3884 14068
rect 3651 14028 3884 14056
rect 3651 14025 3663 14028
rect 3605 14019 3663 14025
rect 3878 14016 3884 14028
rect 3936 14016 3942 14068
rect 4154 14016 4160 14068
rect 4212 14056 4218 14068
rect 4709 14059 4767 14065
rect 4709 14056 4721 14059
rect 4212 14028 4721 14056
rect 4212 14016 4218 14028
rect 4709 14025 4721 14028
rect 4755 14056 4767 14059
rect 6457 14059 6515 14065
rect 6457 14056 6469 14059
rect 4755 14028 6469 14056
rect 4755 14025 4767 14028
rect 4709 14019 4767 14025
rect 6457 14025 6469 14028
rect 6503 14056 6515 14059
rect 6549 14059 6607 14065
rect 6549 14056 6561 14059
rect 6503 14028 6561 14056
rect 6503 14025 6515 14028
rect 6457 14019 6515 14025
rect 6549 14025 6561 14028
rect 6595 14025 6607 14059
rect 6549 14019 6607 14025
rect 9585 14059 9643 14065
rect 9585 14025 9597 14059
rect 9631 14056 9643 14059
rect 10226 14056 10232 14068
rect 9631 14028 10232 14056
rect 9631 14025 9643 14028
rect 9585 14019 9643 14025
rect 10226 14016 10232 14028
rect 10284 14016 10290 14068
rect 10318 14016 10324 14068
rect 10376 14056 10382 14068
rect 10962 14056 10968 14068
rect 10376 14028 10968 14056
rect 10376 14016 10382 14028
rect 10962 14016 10968 14028
rect 11020 14016 11026 14068
rect 11885 14059 11943 14065
rect 11885 14025 11897 14059
rect 11931 14056 11943 14059
rect 12250 14056 12256 14068
rect 11931 14028 12256 14056
rect 11931 14025 11943 14028
rect 11885 14019 11943 14025
rect 12250 14016 12256 14028
rect 12308 14016 12314 14068
rect 15746 14016 15752 14068
rect 15804 14056 15810 14068
rect 16117 14059 16175 14065
rect 16117 14056 16129 14059
rect 15804 14028 16129 14056
rect 15804 14016 15810 14028
rect 16117 14025 16129 14028
rect 16163 14056 16175 14059
rect 16439 14059 16497 14065
rect 16439 14056 16451 14059
rect 16163 14028 16451 14056
rect 16163 14025 16175 14028
rect 16117 14019 16175 14025
rect 16439 14025 16451 14028
rect 16485 14025 16497 14059
rect 17862 14056 17868 14068
rect 17823 14028 17868 14056
rect 16439 14019 16497 14025
rect 17862 14016 17868 14028
rect 17920 14056 17926 14068
rect 19150 14056 19156 14068
rect 17920 14028 19156 14056
rect 17920 14016 17926 14028
rect 19150 14016 19156 14028
rect 19208 14016 19214 14068
rect 20714 14056 20720 14068
rect 20675 14028 20720 14056
rect 20714 14016 20720 14028
rect 20772 14016 20778 14068
rect 22186 14056 22192 14068
rect 22147 14028 22192 14056
rect 22186 14016 22192 14028
rect 22244 14016 22250 14068
rect 2130 13988 2136 14000
rect 2091 13960 2136 13988
rect 2130 13948 2136 13960
rect 2188 13988 2194 14000
rect 4246 13988 4252 14000
rect 2188 13960 4252 13988
rect 2188 13948 2194 13960
rect 4246 13948 4252 13960
rect 4304 13948 4310 14000
rect 4614 13988 4620 14000
rect 4401 13960 4620 13988
rect 1578 13920 1584 13932
rect 1539 13892 1584 13920
rect 1578 13880 1584 13892
rect 1636 13880 1642 13932
rect 3789 13923 3847 13929
rect 3789 13889 3801 13923
rect 3835 13920 3847 13923
rect 4401 13920 4429 13960
rect 4614 13948 4620 13960
rect 4672 13988 4678 14000
rect 5077 13991 5135 13997
rect 5077 13988 5089 13991
rect 4672 13960 5089 13988
rect 4672 13948 4678 13960
rect 5077 13957 5089 13960
rect 5123 13957 5135 13991
rect 5077 13951 5135 13957
rect 6273 13991 6331 13997
rect 6273 13957 6285 13991
rect 6319 13988 6331 13991
rect 11238 13988 11244 14000
rect 6319 13960 11244 13988
rect 6319 13957 6331 13960
rect 6273 13951 6331 13957
rect 3835 13892 4429 13920
rect 3835 13889 3847 13892
rect 3789 13883 3847 13889
rect 4890 13812 4896 13864
rect 4948 13852 4954 13864
rect 5788 13855 5846 13861
rect 5788 13852 5800 13855
rect 4948 13824 5800 13852
rect 4948 13812 4954 13824
rect 5788 13821 5800 13824
rect 5834 13852 5846 13855
rect 6288 13852 6316 13951
rect 11238 13948 11244 13960
rect 11296 13948 11302 14000
rect 11333 13991 11391 13997
rect 11333 13957 11345 13991
rect 11379 13988 11391 13991
rect 12161 13991 12219 13997
rect 12161 13988 12173 13991
rect 11379 13960 12173 13988
rect 11379 13957 11391 13960
rect 11333 13951 11391 13957
rect 12161 13957 12173 13960
rect 12207 13988 12219 13991
rect 12618 13988 12624 14000
rect 12207 13960 12624 13988
rect 12207 13957 12219 13960
rect 12161 13951 12219 13957
rect 12618 13948 12624 13960
rect 12676 13988 12682 14000
rect 13633 13991 13691 13997
rect 13633 13988 13645 13991
rect 12676 13960 13645 13988
rect 12676 13948 12682 13960
rect 13633 13957 13645 13960
rect 13679 13988 13691 13991
rect 13814 13988 13820 14000
rect 13679 13960 13820 13988
rect 13679 13957 13691 13960
rect 13633 13951 13691 13957
rect 13814 13948 13820 13960
rect 13872 13948 13878 14000
rect 15838 13988 15844 14000
rect 15799 13960 15844 13988
rect 15838 13948 15844 13960
rect 15896 13948 15902 14000
rect 6454 13880 6460 13932
rect 6512 13920 6518 13932
rect 6825 13923 6883 13929
rect 6825 13920 6837 13923
rect 6512 13892 6837 13920
rect 6512 13880 6518 13892
rect 6825 13889 6837 13892
rect 6871 13889 6883 13923
rect 9950 13920 9956 13932
rect 9863 13892 9956 13920
rect 6825 13883 6883 13889
rect 9950 13880 9956 13892
rect 10008 13920 10014 13932
rect 10318 13920 10324 13932
rect 10008 13892 10324 13920
rect 10008 13880 10014 13892
rect 10318 13880 10324 13892
rect 10376 13880 10382 13932
rect 12526 13880 12532 13932
rect 12584 13920 12590 13932
rect 12805 13923 12863 13929
rect 12805 13920 12817 13923
rect 12584 13892 12817 13920
rect 12584 13880 12590 13892
rect 12805 13889 12817 13892
rect 12851 13889 12863 13923
rect 15470 13920 15476 13932
rect 15431 13892 15476 13920
rect 12805 13883 12863 13889
rect 15470 13880 15476 13892
rect 15528 13880 15534 13932
rect 18782 13880 18788 13932
rect 18840 13920 18846 13932
rect 19058 13920 19064 13932
rect 18840 13892 19064 13920
rect 18840 13880 18846 13892
rect 19058 13880 19064 13892
rect 19116 13880 19122 13932
rect 20346 13920 20352 13932
rect 20307 13892 20352 13920
rect 20346 13880 20352 13892
rect 20404 13880 20410 13932
rect 21266 13920 21272 13932
rect 21227 13892 21272 13920
rect 21266 13880 21272 13892
rect 21324 13880 21330 13932
rect 10410 13852 10416 13864
rect 5834 13824 6316 13852
rect 10371 13824 10416 13852
rect 5834 13821 5846 13824
rect 5788 13815 5846 13821
rect 10410 13812 10416 13824
rect 10468 13812 10474 13864
rect 14734 13852 14740 13864
rect 14695 13824 14740 13852
rect 14734 13812 14740 13824
rect 14792 13812 14798 13864
rect 15197 13855 15255 13861
rect 15197 13821 15209 13855
rect 15243 13821 15255 13855
rect 15197 13815 15255 13821
rect 16368 13855 16426 13861
rect 16368 13821 16380 13855
rect 16414 13852 16426 13855
rect 16853 13855 16911 13861
rect 16853 13852 16865 13855
rect 16414 13824 16865 13852
rect 16414 13821 16426 13824
rect 16368 13815 16426 13821
rect 16853 13821 16865 13824
rect 16899 13852 16911 13855
rect 18046 13852 18052 13864
rect 18104 13861 18110 13864
rect 18104 13855 18142 13861
rect 16899 13824 18052 13852
rect 16899 13821 16911 13824
rect 16853 13815 16911 13821
rect 1673 13787 1731 13793
rect 1673 13753 1685 13787
rect 1719 13784 1731 13787
rect 2038 13784 2044 13796
rect 1719 13756 2044 13784
rect 1719 13753 1731 13756
rect 1673 13747 1731 13753
rect 2038 13744 2044 13756
rect 2096 13744 2102 13796
rect 3878 13784 3884 13796
rect 3839 13756 3884 13784
rect 3878 13744 3884 13756
rect 3936 13744 3942 13796
rect 4246 13744 4252 13796
rect 4304 13784 4310 13796
rect 4433 13787 4491 13793
rect 4433 13784 4445 13787
rect 4304 13756 4445 13784
rect 4304 13744 4310 13756
rect 4433 13753 4445 13756
rect 4479 13753 4491 13787
rect 4433 13747 4491 13753
rect 6457 13787 6515 13793
rect 6457 13753 6469 13787
rect 6503 13784 6515 13787
rect 7146 13787 7204 13793
rect 7146 13784 7158 13787
rect 6503 13756 7158 13784
rect 6503 13753 6515 13756
rect 6457 13747 6515 13753
rect 7146 13753 7158 13756
rect 7192 13753 7204 13787
rect 7146 13747 7204 13753
rect 10775 13787 10833 13793
rect 10775 13753 10787 13787
rect 10821 13784 10833 13787
rect 11330 13784 11336 13796
rect 10821 13756 11336 13784
rect 10821 13753 10833 13756
rect 10775 13747 10833 13753
rect 11330 13744 11336 13756
rect 11388 13744 11394 13796
rect 12529 13787 12587 13793
rect 12529 13753 12541 13787
rect 12575 13753 12587 13787
rect 12529 13747 12587 13753
rect 5859 13719 5917 13725
rect 5859 13685 5871 13719
rect 5905 13716 5917 13719
rect 6270 13716 6276 13728
rect 5905 13688 6276 13716
rect 5905 13685 5917 13688
rect 5859 13679 5917 13685
rect 6270 13676 6276 13688
rect 6328 13676 6334 13728
rect 7745 13719 7803 13725
rect 7745 13685 7757 13719
rect 7791 13716 7803 13719
rect 7834 13716 7840 13728
rect 7791 13688 7840 13716
rect 7791 13685 7803 13688
rect 7745 13679 7803 13685
rect 7834 13676 7840 13688
rect 7892 13716 7898 13728
rect 8021 13719 8079 13725
rect 8021 13716 8033 13719
rect 7892 13688 8033 13716
rect 7892 13676 7898 13688
rect 8021 13685 8033 13688
rect 8067 13685 8079 13719
rect 8662 13716 8668 13728
rect 8575 13688 8668 13716
rect 8021 13679 8079 13685
rect 8662 13676 8668 13688
rect 8720 13716 8726 13728
rect 10134 13716 10140 13728
rect 8720 13688 10140 13716
rect 8720 13676 8726 13688
rect 10134 13676 10140 13688
rect 10192 13676 10198 13728
rect 12434 13676 12440 13728
rect 12492 13716 12498 13728
rect 12544 13716 12572 13747
rect 12618 13744 12624 13796
rect 12676 13784 12682 13796
rect 12676 13756 12721 13784
rect 12676 13744 12682 13756
rect 12492 13688 12572 13716
rect 12492 13676 12498 13688
rect 13170 13676 13176 13728
rect 13228 13716 13234 13728
rect 13722 13716 13728 13728
rect 13228 13688 13728 13716
rect 13228 13676 13234 13688
rect 13722 13676 13728 13688
rect 13780 13716 13786 13728
rect 14001 13719 14059 13725
rect 14001 13716 14013 13719
rect 13780 13688 14013 13716
rect 13780 13676 13786 13688
rect 14001 13685 14013 13688
rect 14047 13685 14059 13719
rect 14550 13716 14556 13728
rect 14511 13688 14556 13716
rect 14001 13679 14059 13685
rect 14550 13676 14556 13688
rect 14608 13716 14614 13728
rect 15212 13716 15240 13815
rect 18046 13812 18052 13824
rect 18130 13852 18142 13855
rect 18509 13855 18567 13861
rect 18509 13852 18521 13855
rect 18130 13824 18521 13852
rect 18130 13821 18142 13824
rect 18104 13815 18142 13821
rect 18509 13821 18521 13824
rect 18555 13821 18567 13855
rect 19426 13852 19432 13864
rect 18509 13815 18567 13821
rect 19260 13824 19432 13852
rect 18104 13812 18110 13815
rect 17494 13716 17500 13728
rect 14608 13688 15240 13716
rect 17455 13688 17500 13716
rect 14608 13676 14614 13688
rect 17494 13676 17500 13688
rect 17552 13676 17558 13728
rect 17586 13676 17592 13728
rect 17644 13716 17650 13728
rect 18187 13719 18245 13725
rect 18187 13716 18199 13719
rect 17644 13688 18199 13716
rect 17644 13676 17650 13688
rect 18187 13685 18199 13688
rect 18233 13685 18245 13719
rect 18874 13716 18880 13728
rect 18835 13688 18880 13716
rect 18187 13679 18245 13685
rect 18874 13676 18880 13688
rect 18932 13716 18938 13728
rect 19260 13716 19288 13824
rect 18932 13688 19288 13716
rect 19352 13716 19380 13824
rect 19426 13812 19432 13824
rect 19484 13812 19490 13864
rect 20622 13744 20628 13796
rect 20680 13784 20686 13796
rect 20901 13787 20959 13793
rect 20901 13784 20913 13787
rect 20680 13756 20913 13784
rect 20680 13744 20686 13756
rect 20901 13753 20913 13756
rect 20947 13753 20959 13787
rect 20901 13747 20959 13753
rect 20990 13744 20996 13796
rect 21048 13784 21054 13796
rect 21821 13787 21879 13793
rect 21821 13784 21833 13787
rect 21048 13756 21833 13784
rect 21048 13744 21054 13756
rect 21821 13753 21833 13756
rect 21867 13753 21879 13787
rect 21821 13747 21879 13753
rect 19429 13719 19487 13725
rect 19429 13716 19441 13719
rect 19352 13688 19441 13716
rect 18932 13676 18938 13688
rect 19429 13685 19441 13688
rect 19475 13685 19487 13719
rect 19429 13679 19487 13685
rect 19981 13719 20039 13725
rect 19981 13685 19993 13719
rect 20027 13716 20039 13719
rect 20806 13716 20812 13728
rect 20027 13688 20812 13716
rect 20027 13685 20039 13688
rect 19981 13679 20039 13685
rect 20806 13676 20812 13688
rect 20864 13716 20870 13728
rect 21082 13716 21088 13728
rect 20864 13688 21088 13716
rect 20864 13676 20870 13688
rect 21082 13676 21088 13688
rect 21140 13676 21146 13728
rect 1104 13626 22816 13648
rect 1104 13574 8982 13626
rect 9034 13574 9046 13626
rect 9098 13574 9110 13626
rect 9162 13574 9174 13626
rect 9226 13574 16982 13626
rect 17034 13574 17046 13626
rect 17098 13574 17110 13626
rect 17162 13574 17174 13626
rect 17226 13574 22816 13626
rect 1104 13552 22816 13574
rect 2038 13472 2044 13524
rect 2096 13512 2102 13524
rect 2317 13515 2375 13521
rect 2317 13512 2329 13515
rect 2096 13484 2329 13512
rect 2096 13472 2102 13484
rect 2317 13481 2329 13484
rect 2363 13512 2375 13515
rect 2593 13515 2651 13521
rect 2593 13512 2605 13515
rect 2363 13484 2605 13512
rect 2363 13481 2375 13484
rect 2317 13475 2375 13481
rect 2593 13481 2605 13484
rect 2639 13481 2651 13515
rect 2593 13475 2651 13481
rect 3789 13515 3847 13521
rect 3789 13481 3801 13515
rect 3835 13512 3847 13515
rect 3878 13512 3884 13524
rect 3835 13484 3884 13512
rect 3835 13481 3847 13484
rect 3789 13475 3847 13481
rect 3878 13472 3884 13484
rect 3936 13472 3942 13524
rect 6043 13515 6101 13521
rect 6043 13481 6055 13515
rect 6089 13512 6101 13515
rect 6362 13512 6368 13524
rect 6089 13484 6368 13512
rect 6089 13481 6101 13484
rect 6043 13475 6101 13481
rect 6362 13472 6368 13484
rect 6420 13472 6426 13524
rect 6454 13472 6460 13524
rect 6512 13512 6518 13524
rect 6733 13515 6791 13521
rect 6733 13512 6745 13515
rect 6512 13484 6745 13512
rect 6512 13472 6518 13484
rect 6733 13481 6745 13484
rect 6779 13481 6791 13515
rect 6733 13475 6791 13481
rect 9950 13472 9956 13524
rect 10008 13512 10014 13524
rect 11330 13512 11336 13524
rect 10008 13484 11336 13512
rect 10008 13472 10014 13484
rect 11330 13472 11336 13484
rect 11388 13472 11394 13524
rect 12802 13512 12808 13524
rect 12763 13484 12808 13512
rect 12802 13472 12808 13484
rect 12860 13472 12866 13524
rect 14734 13512 14740 13524
rect 14695 13484 14740 13512
rect 14734 13472 14740 13484
rect 14792 13472 14798 13524
rect 17678 13512 17684 13524
rect 15764 13484 17684 13512
rect 1759 13447 1817 13453
rect 1759 13413 1771 13447
rect 1805 13444 1817 13447
rect 1854 13444 1860 13456
rect 1805 13416 1860 13444
rect 1805 13413 1817 13416
rect 1759 13407 1817 13413
rect 1854 13404 1860 13416
rect 1912 13444 1918 13456
rect 2498 13444 2504 13456
rect 1912 13416 2504 13444
rect 1912 13404 1918 13416
rect 2498 13404 2504 13416
rect 2556 13404 2562 13456
rect 4522 13444 4528 13456
rect 4483 13416 4528 13444
rect 4522 13404 4528 13416
rect 4580 13404 4586 13456
rect 7006 13404 7012 13456
rect 7064 13444 7070 13456
rect 7101 13447 7159 13453
rect 7101 13444 7113 13447
rect 7064 13416 7113 13444
rect 7064 13404 7070 13416
rect 7101 13413 7113 13416
rect 7147 13444 7159 13447
rect 7834 13444 7840 13456
rect 7147 13416 7840 13444
rect 7147 13413 7159 13416
rect 7101 13407 7159 13413
rect 7834 13404 7840 13416
rect 7892 13404 7898 13456
rect 10410 13444 10416 13456
rect 10323 13416 10416 13444
rect 10410 13404 10416 13416
rect 10468 13444 10474 13456
rect 10689 13447 10747 13453
rect 10689 13444 10701 13447
rect 10468 13416 10701 13444
rect 10468 13404 10474 13416
rect 10689 13413 10701 13416
rect 10735 13413 10747 13447
rect 10689 13407 10747 13413
rect 12023 13447 12081 13453
rect 12023 13413 12035 13447
rect 12069 13444 12081 13447
rect 13170 13444 13176 13456
rect 12069 13416 13176 13444
rect 12069 13413 12081 13416
rect 12023 13407 12081 13413
rect 13170 13404 13176 13416
rect 13228 13404 13234 13456
rect 5972 13379 6030 13385
rect 5972 13345 5984 13379
rect 6018 13376 6030 13379
rect 6178 13376 6184 13388
rect 6018 13348 6184 13376
rect 6018 13345 6030 13348
rect 5972 13339 6030 13345
rect 6178 13336 6184 13348
rect 6236 13336 6242 13388
rect 7650 13336 7656 13388
rect 7708 13376 7714 13388
rect 9582 13376 9588 13388
rect 7708 13348 9588 13376
rect 7708 13336 7714 13348
rect 9582 13336 9588 13348
rect 9640 13376 9646 13388
rect 9677 13379 9735 13385
rect 9677 13376 9689 13379
rect 9640 13348 9689 13376
rect 9640 13336 9646 13348
rect 9677 13345 9689 13348
rect 9723 13345 9735 13379
rect 9677 13339 9735 13345
rect 9766 13336 9772 13388
rect 9824 13376 9830 13388
rect 10137 13379 10195 13385
rect 10137 13376 10149 13379
rect 9824 13348 10149 13376
rect 9824 13336 9830 13348
rect 10137 13345 10149 13348
rect 10183 13345 10195 13379
rect 11882 13376 11888 13388
rect 11843 13348 11888 13376
rect 10137 13339 10195 13345
rect 11882 13336 11888 13348
rect 11940 13336 11946 13388
rect 13722 13376 13728 13388
rect 13683 13348 13728 13376
rect 13722 13336 13728 13348
rect 13780 13336 13786 13388
rect 14182 13376 14188 13388
rect 14095 13348 14188 13376
rect 14182 13336 14188 13348
rect 14240 13376 14246 13388
rect 14752 13376 14780 13472
rect 14240 13348 14780 13376
rect 14240 13336 14246 13348
rect 1397 13311 1455 13317
rect 1397 13277 1409 13311
rect 1443 13308 1455 13311
rect 2130 13308 2136 13320
rect 1443 13280 2136 13308
rect 1443 13277 1455 13280
rect 1397 13271 1455 13277
rect 2130 13268 2136 13280
rect 2188 13268 2194 13320
rect 4430 13308 4436 13320
rect 4391 13280 4436 13308
rect 4430 13268 4436 13280
rect 4488 13268 4494 13320
rect 4709 13311 4767 13317
rect 4709 13277 4721 13311
rect 4755 13277 4767 13311
rect 4709 13271 4767 13277
rect 4246 13200 4252 13252
rect 4304 13240 4310 13252
rect 4724 13240 4752 13271
rect 6270 13268 6276 13320
rect 6328 13308 6334 13320
rect 7009 13311 7067 13317
rect 7009 13308 7021 13311
rect 6328 13280 7021 13308
rect 6328 13268 6334 13280
rect 7009 13277 7021 13280
rect 7055 13277 7067 13311
rect 7282 13308 7288 13320
rect 7243 13280 7288 13308
rect 7009 13271 7067 13277
rect 7282 13268 7288 13280
rect 7340 13268 7346 13320
rect 14274 13308 14280 13320
rect 14235 13280 14280 13308
rect 14274 13268 14280 13280
rect 14332 13268 14338 13320
rect 4304 13212 4752 13240
rect 4304 13200 4310 13212
rect 11882 13200 11888 13252
rect 11940 13240 11946 13252
rect 15764 13240 15792 13484
rect 17678 13472 17684 13484
rect 17736 13472 17742 13524
rect 18506 13512 18512 13524
rect 18467 13484 18512 13512
rect 18506 13472 18512 13484
rect 18564 13472 18570 13524
rect 19334 13472 19340 13524
rect 19392 13512 19398 13524
rect 19429 13515 19487 13521
rect 19429 13512 19441 13515
rect 19392 13484 19441 13512
rect 19392 13472 19398 13484
rect 19429 13481 19441 13484
rect 19475 13481 19487 13515
rect 19429 13475 19487 13481
rect 19981 13515 20039 13521
rect 19981 13481 19993 13515
rect 20027 13512 20039 13515
rect 20990 13512 20996 13524
rect 20027 13484 20996 13512
rect 20027 13481 20039 13484
rect 19981 13475 20039 13481
rect 20990 13472 20996 13484
rect 21048 13472 21054 13524
rect 16022 13444 16028 13456
rect 15983 13416 16028 13444
rect 16022 13404 16028 13416
rect 16080 13404 16086 13456
rect 21082 13444 21088 13456
rect 21043 13416 21088 13444
rect 21082 13404 21088 13416
rect 21140 13404 21146 13456
rect 17494 13376 17500 13388
rect 17455 13348 17500 13376
rect 17494 13336 17500 13348
rect 17552 13336 17558 13388
rect 18049 13379 18107 13385
rect 18049 13345 18061 13379
rect 18095 13345 18107 13379
rect 18049 13339 18107 13345
rect 15930 13308 15936 13320
rect 15843 13280 15936 13308
rect 15930 13268 15936 13280
rect 15988 13308 15994 13320
rect 17586 13308 17592 13320
rect 15988 13280 17592 13308
rect 15988 13268 15994 13280
rect 17586 13268 17592 13280
rect 17644 13268 17650 13320
rect 11940 13212 15792 13240
rect 16485 13243 16543 13249
rect 11940 13200 11946 13212
rect 16485 13209 16497 13243
rect 16531 13240 16543 13243
rect 17954 13240 17960 13252
rect 16531 13212 17960 13240
rect 16531 13209 16543 13212
rect 16485 13203 16543 13209
rect 17954 13200 17960 13212
rect 18012 13200 18018 13252
rect 6454 13172 6460 13184
rect 6415 13144 6460 13172
rect 6454 13132 6460 13144
rect 6512 13132 6518 13184
rect 8662 13172 8668 13184
rect 8623 13144 8668 13172
rect 8662 13132 8668 13144
rect 8720 13132 8726 13184
rect 12434 13172 12440 13184
rect 12395 13144 12440 13172
rect 12434 13132 12440 13144
rect 12492 13132 12498 13184
rect 16114 13132 16120 13184
rect 16172 13172 16178 13184
rect 16853 13175 16911 13181
rect 16853 13172 16865 13175
rect 16172 13144 16865 13172
rect 16172 13132 16178 13144
rect 16853 13141 16865 13144
rect 16899 13141 16911 13175
rect 16853 13135 16911 13141
rect 17402 13132 17408 13184
rect 17460 13172 17466 13184
rect 18064 13172 18092 13339
rect 18233 13311 18291 13317
rect 18233 13277 18245 13311
rect 18279 13308 18291 13311
rect 19058 13308 19064 13320
rect 18279 13280 19064 13308
rect 18279 13277 18291 13280
rect 18233 13271 18291 13277
rect 19058 13268 19064 13280
rect 19116 13268 19122 13320
rect 20993 13311 21051 13317
rect 20993 13277 21005 13311
rect 21039 13277 21051 13311
rect 21266 13308 21272 13320
rect 21227 13280 21272 13308
rect 20993 13271 21051 13277
rect 21008 13240 21036 13271
rect 21266 13268 21272 13280
rect 21324 13268 21330 13320
rect 21358 13240 21364 13252
rect 21008 13212 21364 13240
rect 21358 13200 21364 13212
rect 21416 13200 21422 13252
rect 20622 13172 20628 13184
rect 17460 13144 18092 13172
rect 20583 13144 20628 13172
rect 17460 13132 17466 13144
rect 20622 13132 20628 13144
rect 20680 13132 20686 13184
rect 1104 13082 22816 13104
rect 1104 13030 4982 13082
rect 5034 13030 5046 13082
rect 5098 13030 5110 13082
rect 5162 13030 5174 13082
rect 5226 13030 12982 13082
rect 13034 13030 13046 13082
rect 13098 13030 13110 13082
rect 13162 13030 13174 13082
rect 13226 13030 20982 13082
rect 21034 13030 21046 13082
rect 21098 13030 21110 13082
rect 21162 13030 21174 13082
rect 21226 13030 22816 13082
rect 1104 13008 22816 13030
rect 3602 12968 3608 12980
rect 3563 12940 3608 12968
rect 3602 12928 3608 12940
rect 3660 12928 3666 12980
rect 4522 12928 4528 12980
rect 4580 12968 4586 12980
rect 5077 12971 5135 12977
rect 5077 12968 5089 12971
rect 4580 12940 5089 12968
rect 4580 12928 4586 12940
rect 5077 12937 5089 12940
rect 5123 12937 5135 12971
rect 5077 12931 5135 12937
rect 5626 12928 5632 12980
rect 5684 12968 5690 12980
rect 6457 12971 6515 12977
rect 6457 12968 6469 12971
rect 5684 12940 6469 12968
rect 5684 12928 5690 12940
rect 6457 12937 6469 12940
rect 6503 12937 6515 12971
rect 6457 12931 6515 12937
rect 9582 12928 9588 12980
rect 9640 12968 9646 12980
rect 11333 12971 11391 12977
rect 11333 12968 11345 12971
rect 9640 12940 11345 12968
rect 9640 12928 9646 12940
rect 11333 12937 11345 12940
rect 11379 12968 11391 12971
rect 11379 12940 12020 12968
rect 11379 12937 11391 12940
rect 11333 12931 11391 12937
rect 4430 12860 4436 12912
rect 4488 12900 4494 12912
rect 4709 12903 4767 12909
rect 4709 12900 4721 12903
rect 4488 12872 4721 12900
rect 4488 12860 4494 12872
rect 4709 12869 4721 12872
rect 4755 12900 4767 12903
rect 7466 12900 7472 12912
rect 4755 12872 7472 12900
rect 4755 12869 4767 12872
rect 4709 12863 4767 12869
rect 7466 12860 7472 12872
rect 7524 12860 7530 12912
rect 10134 12860 10140 12912
rect 10192 12900 10198 12912
rect 11882 12900 11888 12912
rect 10192 12872 11888 12900
rect 10192 12860 10198 12872
rect 11882 12860 11888 12872
rect 11940 12860 11946 12912
rect 11992 12900 12020 12940
rect 12434 12928 12440 12980
rect 12492 12968 12498 12980
rect 12575 12971 12633 12977
rect 12575 12968 12587 12971
rect 12492 12940 12587 12968
rect 12492 12928 12498 12940
rect 12575 12937 12587 12940
rect 12621 12937 12633 12971
rect 12575 12931 12633 12937
rect 13722 12928 13728 12980
rect 13780 12968 13786 12980
rect 15197 12971 15255 12977
rect 13780 12940 15148 12968
rect 13780 12928 13786 12940
rect 13265 12903 13323 12909
rect 13265 12900 13277 12903
rect 11992 12872 13277 12900
rect 13265 12869 13277 12872
rect 13311 12900 13323 12903
rect 14182 12900 14188 12912
rect 13311 12872 14188 12900
rect 13311 12869 13323 12872
rect 13265 12863 13323 12869
rect 14182 12860 14188 12872
rect 14240 12860 14246 12912
rect 15120 12900 15148 12940
rect 15197 12937 15209 12971
rect 15243 12968 15255 12971
rect 15565 12971 15623 12977
rect 15565 12968 15577 12971
rect 15243 12940 15577 12968
rect 15243 12937 15255 12940
rect 15197 12931 15255 12937
rect 15565 12937 15577 12940
rect 15611 12968 15623 12971
rect 15933 12971 15991 12977
rect 15933 12968 15945 12971
rect 15611 12940 15945 12968
rect 15611 12937 15623 12940
rect 15565 12931 15623 12937
rect 15933 12937 15945 12940
rect 15979 12968 15991 12971
rect 16022 12968 16028 12980
rect 15979 12940 16028 12968
rect 15979 12937 15991 12940
rect 15933 12931 15991 12937
rect 16022 12928 16028 12940
rect 16080 12928 16086 12980
rect 19306 12940 20484 12968
rect 17405 12903 17463 12909
rect 17405 12900 17417 12903
rect 15120 12872 17417 12900
rect 17405 12869 17417 12872
rect 17451 12900 17463 12903
rect 17494 12900 17500 12912
rect 17451 12872 17500 12900
rect 17451 12869 17463 12872
rect 17405 12863 17463 12869
rect 17494 12860 17500 12872
rect 17552 12900 17558 12912
rect 17773 12903 17831 12909
rect 17773 12900 17785 12903
rect 17552 12872 17785 12900
rect 17552 12860 17558 12872
rect 17773 12869 17785 12872
rect 17819 12869 17831 12903
rect 17773 12863 17831 12869
rect 2130 12832 2136 12844
rect 2043 12804 2136 12832
rect 2130 12792 2136 12804
rect 2188 12832 2194 12844
rect 2777 12835 2835 12841
rect 2777 12832 2789 12835
rect 2188 12804 2789 12832
rect 2188 12792 2194 12804
rect 2777 12801 2789 12804
rect 2823 12801 2835 12835
rect 2777 12795 2835 12801
rect 4157 12835 4215 12841
rect 4157 12801 4169 12835
rect 4203 12832 4215 12835
rect 5445 12835 5503 12841
rect 5445 12832 5457 12835
rect 4203 12804 5457 12832
rect 4203 12801 4215 12804
rect 4157 12795 4215 12801
rect 5445 12801 5457 12804
rect 5491 12832 5503 12835
rect 5767 12835 5825 12841
rect 5767 12832 5779 12835
rect 5491 12804 5779 12832
rect 5491 12801 5503 12804
rect 5445 12795 5503 12801
rect 5767 12801 5779 12804
rect 5813 12801 5825 12835
rect 5767 12795 5825 12801
rect 6454 12792 6460 12844
rect 6512 12832 6518 12844
rect 6917 12835 6975 12841
rect 6917 12832 6929 12835
rect 6512 12804 6929 12832
rect 6512 12792 6518 12804
rect 6917 12801 6929 12804
rect 6963 12832 6975 12835
rect 7926 12832 7932 12844
rect 6963 12804 7932 12832
rect 6963 12801 6975 12804
rect 6917 12795 6975 12801
rect 7926 12792 7932 12804
rect 7984 12792 7990 12844
rect 8481 12835 8539 12841
rect 8481 12801 8493 12835
rect 8527 12832 8539 12835
rect 14274 12832 14280 12844
rect 8527 12804 9076 12832
rect 14235 12804 14280 12832
rect 8527 12801 8539 12804
rect 8481 12795 8539 12801
rect 1670 12764 1676 12776
rect 1631 12736 1676 12764
rect 1670 12724 1676 12736
rect 1728 12724 1734 12776
rect 1946 12764 1952 12776
rect 1859 12736 1952 12764
rect 1946 12724 1952 12736
rect 2004 12764 2010 12776
rect 3120 12767 3178 12773
rect 2004 12736 2544 12764
rect 2004 12724 2010 12736
rect 2516 12637 2544 12736
rect 3120 12733 3132 12767
rect 3166 12764 3178 12767
rect 3602 12764 3608 12776
rect 3166 12736 3608 12764
rect 3166 12733 3178 12736
rect 3120 12727 3178 12733
rect 3602 12724 3608 12736
rect 3660 12724 3666 12776
rect 4798 12724 4804 12776
rect 4856 12764 4862 12776
rect 5626 12764 5632 12776
rect 4856 12736 5632 12764
rect 4856 12724 4862 12736
rect 5626 12724 5632 12736
rect 5684 12724 5690 12776
rect 8662 12764 8668 12776
rect 8623 12736 8668 12764
rect 8662 12724 8668 12736
rect 8720 12724 8726 12776
rect 9048 12773 9076 12804
rect 14274 12792 14280 12804
rect 14332 12792 14338 12844
rect 16114 12832 16120 12844
rect 16075 12804 16120 12832
rect 16114 12792 16120 12804
rect 16172 12792 16178 12844
rect 9033 12767 9091 12773
rect 9033 12733 9045 12767
rect 9079 12764 9091 12767
rect 10137 12767 10195 12773
rect 10137 12764 10149 12767
rect 9079 12736 10149 12764
rect 9079 12733 9091 12736
rect 9033 12727 9091 12733
rect 10137 12733 10149 12736
rect 10183 12733 10195 12767
rect 10594 12764 10600 12776
rect 10555 12736 10600 12764
rect 10137 12727 10195 12733
rect 3973 12699 4031 12705
rect 3973 12665 3985 12699
rect 4019 12696 4031 12699
rect 4246 12696 4252 12708
rect 4019 12668 4252 12696
rect 4019 12665 4031 12668
rect 3973 12659 4031 12665
rect 4246 12656 4252 12668
rect 4304 12656 4310 12708
rect 7006 12696 7012 12708
rect 6967 12668 7012 12696
rect 7006 12656 7012 12668
rect 7064 12656 7070 12708
rect 10152 12696 10180 12727
rect 10594 12724 10600 12736
rect 10652 12724 10658 12776
rect 10781 12767 10839 12773
rect 10781 12733 10793 12767
rect 10827 12733 10839 12767
rect 10781 12727 10839 12733
rect 10226 12696 10232 12708
rect 10139 12668 10232 12696
rect 10226 12656 10232 12668
rect 10284 12696 10290 12708
rect 10796 12696 10824 12727
rect 12342 12724 12348 12776
rect 12400 12764 12406 12776
rect 12472 12767 12530 12773
rect 12472 12764 12484 12767
rect 12400 12736 12484 12764
rect 12400 12724 12406 12736
rect 12472 12733 12484 12736
rect 12518 12764 12530 12767
rect 12897 12767 12955 12773
rect 12897 12764 12909 12767
rect 12518 12736 12909 12764
rect 12518 12733 12530 12736
rect 12472 12727 12530 12733
rect 12897 12733 12909 12736
rect 12943 12764 12955 12767
rect 15838 12764 15844 12776
rect 12943 12736 15844 12764
rect 12943 12733 12955 12736
rect 12897 12727 12955 12733
rect 15838 12724 15844 12736
rect 15896 12724 15902 12776
rect 17788 12764 17816 12863
rect 17954 12860 17960 12912
rect 18012 12900 18018 12912
rect 19306 12900 19334 12940
rect 18012 12872 19334 12900
rect 18012 12860 18018 12872
rect 18782 12832 18788 12844
rect 18743 12804 18788 12832
rect 18782 12792 18788 12804
rect 18840 12792 18846 12844
rect 18049 12767 18107 12773
rect 18049 12764 18061 12767
rect 17788 12736 18061 12764
rect 18049 12733 18061 12736
rect 18095 12733 18107 12767
rect 18506 12764 18512 12776
rect 18467 12736 18512 12764
rect 18049 12727 18107 12733
rect 18506 12724 18512 12736
rect 18564 12724 18570 12776
rect 10284 12668 10824 12696
rect 11057 12699 11115 12705
rect 10284 12656 10290 12668
rect 11057 12665 11069 12699
rect 11103 12696 11115 12699
rect 11238 12696 11244 12708
rect 11103 12668 11244 12696
rect 11103 12665 11115 12668
rect 11057 12659 11115 12665
rect 11238 12656 11244 12668
rect 11296 12656 11302 12708
rect 11330 12656 11336 12708
rect 11388 12696 11394 12708
rect 16209 12699 16267 12705
rect 11388 12668 14228 12696
rect 11388 12656 11394 12668
rect 2501 12631 2559 12637
rect 2501 12597 2513 12631
rect 2547 12628 2559 12631
rect 2866 12628 2872 12640
rect 2547 12600 2872 12628
rect 2547 12597 2559 12600
rect 2501 12591 2559 12597
rect 2866 12588 2872 12600
rect 2924 12588 2930 12640
rect 3191 12631 3249 12637
rect 3191 12597 3203 12631
rect 3237 12628 3249 12631
rect 3418 12628 3424 12640
rect 3237 12600 3424 12628
rect 3237 12597 3249 12600
rect 3191 12591 3249 12597
rect 3418 12588 3424 12600
rect 3476 12588 3482 12640
rect 6178 12628 6184 12640
rect 6139 12600 6184 12628
rect 6178 12588 6184 12600
rect 6236 12588 6242 12640
rect 7190 12588 7196 12640
rect 7248 12628 7254 12640
rect 7837 12631 7895 12637
rect 7837 12628 7849 12631
rect 7248 12600 7849 12628
rect 7248 12588 7254 12600
rect 7837 12597 7849 12600
rect 7883 12597 7895 12631
rect 8846 12628 8852 12640
rect 8807 12600 8852 12628
rect 7837 12591 7895 12597
rect 8846 12588 8852 12600
rect 8904 12588 8910 12640
rect 9674 12588 9680 12640
rect 9732 12628 9738 12640
rect 13722 12628 13728 12640
rect 9732 12600 9777 12628
rect 13683 12600 13728 12628
rect 9732 12588 9738 12600
rect 13722 12588 13728 12600
rect 13780 12588 13786 12640
rect 14200 12637 14228 12668
rect 16209 12665 16221 12699
rect 16255 12665 16267 12699
rect 16758 12696 16764 12708
rect 16719 12668 16764 12696
rect 16209 12659 16267 12665
rect 14185 12631 14243 12637
rect 14185 12597 14197 12631
rect 14231 12628 14243 12631
rect 14642 12628 14648 12640
rect 14231 12600 14648 12628
rect 14231 12597 14243 12600
rect 14185 12591 14243 12597
rect 14642 12588 14648 12600
rect 14700 12588 14706 12640
rect 16022 12588 16028 12640
rect 16080 12628 16086 12640
rect 16224 12628 16252 12659
rect 16758 12656 16764 12668
rect 16816 12656 16822 12708
rect 19794 12696 19800 12708
rect 19755 12668 19800 12696
rect 19794 12656 19800 12668
rect 19852 12656 19858 12708
rect 20456 12705 20484 12940
rect 20806 12928 20812 12980
rect 20864 12968 20870 12980
rect 20901 12971 20959 12977
rect 20901 12968 20913 12971
rect 20864 12940 20913 12968
rect 20864 12928 20870 12940
rect 20901 12937 20913 12940
rect 20947 12937 20959 12971
rect 21910 12968 21916 12980
rect 21871 12940 21916 12968
rect 20901 12931 20959 12937
rect 21910 12928 21916 12940
rect 21968 12928 21974 12980
rect 21453 12903 21511 12909
rect 21453 12869 21465 12903
rect 21499 12900 21511 12903
rect 23566 12900 23572 12912
rect 21499 12872 23572 12900
rect 21499 12869 21511 12872
rect 21453 12863 21511 12869
rect 23566 12860 23572 12872
rect 23624 12860 23630 12912
rect 21269 12767 21327 12773
rect 21269 12733 21281 12767
rect 21315 12764 21327 12767
rect 21910 12764 21916 12776
rect 21315 12736 21916 12764
rect 21315 12733 21327 12736
rect 21269 12727 21327 12733
rect 21910 12724 21916 12736
rect 21968 12724 21974 12776
rect 19889 12699 19947 12705
rect 19889 12665 19901 12699
rect 19935 12665 19947 12699
rect 19889 12659 19947 12665
rect 20441 12699 20499 12705
rect 20441 12665 20453 12699
rect 20487 12696 20499 12699
rect 21358 12696 21364 12708
rect 20487 12668 21364 12696
rect 20487 12665 20499 12668
rect 20441 12659 20499 12665
rect 16080 12600 16252 12628
rect 17129 12631 17187 12637
rect 16080 12588 16086 12600
rect 17129 12597 17141 12631
rect 17175 12628 17187 12631
rect 17402 12628 17408 12640
rect 17175 12600 17408 12628
rect 17175 12597 17187 12600
rect 17129 12591 17187 12597
rect 17402 12588 17408 12600
rect 17460 12588 17466 12640
rect 18874 12588 18880 12640
rect 18932 12628 18938 12640
rect 19061 12631 19119 12637
rect 19061 12628 19073 12631
rect 18932 12600 19073 12628
rect 18932 12588 18938 12600
rect 19061 12597 19073 12600
rect 19107 12597 19119 12631
rect 19061 12591 19119 12597
rect 19426 12588 19432 12640
rect 19484 12628 19490 12640
rect 19613 12631 19671 12637
rect 19613 12628 19625 12631
rect 19484 12600 19625 12628
rect 19484 12588 19490 12600
rect 19613 12597 19625 12600
rect 19659 12628 19671 12631
rect 19904 12628 19932 12659
rect 21358 12656 21364 12668
rect 21416 12656 21422 12708
rect 19659 12600 19932 12628
rect 19659 12597 19671 12600
rect 19613 12591 19671 12597
rect 1104 12538 22816 12560
rect 1104 12486 8982 12538
rect 9034 12486 9046 12538
rect 9098 12486 9110 12538
rect 9162 12486 9174 12538
rect 9226 12486 16982 12538
rect 17034 12486 17046 12538
rect 17098 12486 17110 12538
rect 17162 12486 17174 12538
rect 17226 12486 22816 12538
rect 1104 12464 22816 12486
rect 1397 12427 1455 12433
rect 1397 12393 1409 12427
rect 1443 12424 1455 12427
rect 1578 12424 1584 12436
rect 1443 12396 1584 12424
rect 1443 12393 1455 12396
rect 1397 12387 1455 12393
rect 1578 12384 1584 12396
rect 1636 12384 1642 12436
rect 1670 12384 1676 12436
rect 1728 12424 1734 12436
rect 2225 12427 2283 12433
rect 2225 12424 2237 12427
rect 1728 12396 2237 12424
rect 1728 12384 1734 12396
rect 2225 12393 2237 12396
rect 2271 12393 2283 12427
rect 2225 12387 2283 12393
rect 3881 12427 3939 12433
rect 3881 12393 3893 12427
rect 3927 12424 3939 12427
rect 4430 12424 4436 12436
rect 3927 12396 4436 12424
rect 3927 12393 3939 12396
rect 3881 12387 3939 12393
rect 4430 12384 4436 12396
rect 4488 12384 4494 12436
rect 6270 12424 6276 12436
rect 6231 12396 6276 12424
rect 6270 12384 6276 12396
rect 6328 12384 6334 12436
rect 7834 12424 7840 12436
rect 7795 12396 7840 12424
rect 7834 12384 7840 12396
rect 7892 12384 7898 12436
rect 7926 12384 7932 12436
rect 7984 12424 7990 12436
rect 8435 12427 8493 12433
rect 8435 12424 8447 12427
rect 7984 12396 8447 12424
rect 7984 12384 7990 12396
rect 8435 12393 8447 12396
rect 8481 12393 8493 12427
rect 8846 12424 8852 12436
rect 8807 12396 8852 12424
rect 8435 12387 8493 12393
rect 8846 12384 8852 12396
rect 8904 12384 8910 12436
rect 10594 12384 10600 12436
rect 10652 12424 10658 12436
rect 10781 12427 10839 12433
rect 10781 12424 10793 12427
rect 10652 12396 10793 12424
rect 10652 12384 10658 12396
rect 10781 12393 10793 12396
rect 10827 12424 10839 12427
rect 14274 12424 14280 12436
rect 10827 12396 13768 12424
rect 14235 12396 14280 12424
rect 10827 12393 10839 12396
rect 10781 12387 10839 12393
rect 1854 12356 1860 12368
rect 1815 12328 1860 12356
rect 1854 12316 1860 12328
rect 1912 12316 1918 12368
rect 4246 12356 4252 12368
rect 4207 12328 4252 12356
rect 4246 12316 4252 12328
rect 4304 12316 4310 12368
rect 6917 12359 6975 12365
rect 6917 12325 6929 12359
rect 6963 12356 6975 12359
rect 7190 12356 7196 12368
rect 6963 12328 7196 12356
rect 6963 12325 6975 12328
rect 6917 12319 6975 12325
rect 7190 12316 7196 12328
rect 7248 12316 7254 12368
rect 9582 12316 9588 12368
rect 9640 12356 9646 12368
rect 9861 12359 9919 12365
rect 9861 12356 9873 12359
rect 9640 12328 9873 12356
rect 9640 12316 9646 12328
rect 9861 12325 9873 12328
rect 9907 12325 9919 12359
rect 9861 12319 9919 12325
rect 11330 12316 11336 12368
rect 11388 12356 11394 12368
rect 11562 12359 11620 12365
rect 11562 12356 11574 12359
rect 11388 12328 11574 12356
rect 11388 12316 11394 12328
rect 11562 12325 11574 12328
rect 11608 12325 11620 12359
rect 11562 12319 11620 12325
rect 13173 12359 13231 12365
rect 13173 12325 13185 12359
rect 13219 12356 13231 12359
rect 13446 12356 13452 12368
rect 13219 12328 13452 12356
rect 13219 12325 13231 12328
rect 13173 12319 13231 12325
rect 13446 12316 13452 12328
rect 13504 12316 13510 12368
rect 13740 12356 13768 12396
rect 14274 12384 14280 12396
rect 14332 12384 14338 12436
rect 15930 12424 15936 12436
rect 15891 12396 15936 12424
rect 15930 12384 15936 12396
rect 15988 12384 15994 12436
rect 17402 12424 17408 12436
rect 16040 12396 17408 12424
rect 16040 12356 16068 12396
rect 17402 12384 17408 12396
rect 17460 12384 17466 12436
rect 19058 12424 19064 12436
rect 19019 12396 19064 12424
rect 19058 12384 19064 12396
rect 19116 12384 19122 12436
rect 19794 12384 19800 12436
rect 19852 12424 19858 12436
rect 20257 12427 20315 12433
rect 20257 12424 20269 12427
rect 19852 12396 20269 12424
rect 19852 12384 19858 12396
rect 20257 12393 20269 12396
rect 20303 12424 20315 12427
rect 21039 12427 21097 12433
rect 21039 12424 21051 12427
rect 20303 12396 21051 12424
rect 20303 12393 20315 12396
rect 20257 12387 20315 12393
rect 21039 12393 21051 12396
rect 21085 12393 21097 12427
rect 21358 12424 21364 12436
rect 21319 12396 21364 12424
rect 21039 12387 21097 12393
rect 21358 12384 21364 12396
rect 21416 12384 21422 12436
rect 16206 12356 16212 12368
rect 13740 12328 16068 12356
rect 16119 12328 16212 12356
rect 16206 12316 16212 12328
rect 16264 12356 16270 12368
rect 17770 12356 17776 12368
rect 16264 12328 17776 12356
rect 16264 12316 16270 12328
rect 17770 12316 17776 12328
rect 17828 12316 17834 12368
rect 19426 12356 19432 12368
rect 19387 12328 19432 12356
rect 19426 12316 19432 12328
rect 19484 12316 19490 12368
rect 2409 12291 2467 12297
rect 2409 12257 2421 12291
rect 2455 12257 2467 12291
rect 2866 12288 2872 12300
rect 2827 12260 2872 12288
rect 2409 12251 2467 12257
rect 2424 12220 2452 12251
rect 2866 12248 2872 12260
rect 2924 12248 2930 12300
rect 5772 12291 5830 12297
rect 5772 12257 5784 12291
rect 5818 12288 5830 12291
rect 5994 12288 6000 12300
rect 5818 12260 6000 12288
rect 5818 12257 5830 12260
rect 5772 12251 5830 12257
rect 5994 12248 6000 12260
rect 6052 12248 6058 12300
rect 8297 12291 8355 12297
rect 8297 12257 8309 12291
rect 8343 12288 8355 12291
rect 8386 12288 8392 12300
rect 8343 12260 8392 12288
rect 8343 12257 8355 12260
rect 8297 12251 8355 12257
rect 8386 12248 8392 12260
rect 8444 12248 8450 12300
rect 10410 12248 10416 12300
rect 10468 12288 10474 12300
rect 10468 12260 10513 12288
rect 10468 12248 10474 12260
rect 16758 12248 16764 12300
rect 16816 12288 16822 12300
rect 16816 12260 16861 12288
rect 16816 12248 16822 12260
rect 20346 12248 20352 12300
rect 20404 12288 20410 12300
rect 20806 12288 20812 12300
rect 20404 12260 20812 12288
rect 20404 12248 20410 12260
rect 20806 12248 20812 12260
rect 20864 12288 20870 12300
rect 20936 12291 20994 12297
rect 20936 12288 20948 12291
rect 20864 12260 20948 12288
rect 20864 12248 20870 12260
rect 20936 12257 20948 12260
rect 20982 12257 20994 12291
rect 20936 12251 20994 12257
rect 2590 12220 2596 12232
rect 2424 12192 2596 12220
rect 2590 12180 2596 12192
rect 2648 12180 2654 12232
rect 3142 12220 3148 12232
rect 3103 12192 3148 12220
rect 3142 12180 3148 12192
rect 3200 12180 3206 12232
rect 3418 12180 3424 12232
rect 3476 12220 3482 12232
rect 4154 12220 4160 12232
rect 3476 12192 4160 12220
rect 3476 12180 3482 12192
rect 4154 12180 4160 12192
rect 4212 12220 4218 12232
rect 4614 12220 4620 12232
rect 4212 12192 4257 12220
rect 4575 12192 4620 12220
rect 4212 12180 4218 12192
rect 4614 12180 4620 12192
rect 4672 12180 4678 12232
rect 5859 12223 5917 12229
rect 5859 12189 5871 12223
rect 5905 12220 5917 12223
rect 6270 12220 6276 12232
rect 5905 12192 6276 12220
rect 5905 12189 5917 12192
rect 5859 12183 5917 12189
rect 6270 12180 6276 12192
rect 6328 12220 6334 12232
rect 6825 12223 6883 12229
rect 6825 12220 6837 12223
rect 6328 12192 6837 12220
rect 6328 12180 6334 12192
rect 6825 12189 6837 12192
rect 6871 12189 6883 12223
rect 6825 12183 6883 12189
rect 7101 12223 7159 12229
rect 7101 12189 7113 12223
rect 7147 12220 7159 12223
rect 7282 12220 7288 12232
rect 7147 12192 7288 12220
rect 7147 12189 7159 12192
rect 7101 12183 7159 12189
rect 4632 12152 4660 12180
rect 7116 12152 7144 12183
rect 7282 12180 7288 12192
rect 7340 12180 7346 12232
rect 9766 12220 9772 12232
rect 9727 12192 9772 12220
rect 9766 12180 9772 12192
rect 9824 12180 9830 12232
rect 11238 12220 11244 12232
rect 11199 12192 11244 12220
rect 11238 12180 11244 12192
rect 11296 12180 11302 12232
rect 13081 12223 13139 12229
rect 13081 12189 13093 12223
rect 13127 12220 13139 12223
rect 13814 12220 13820 12232
rect 13127 12192 13820 12220
rect 13127 12189 13139 12192
rect 13081 12183 13139 12189
rect 13814 12180 13820 12192
rect 13872 12180 13878 12232
rect 16114 12220 16120 12232
rect 16075 12192 16120 12220
rect 16114 12180 16120 12192
rect 16172 12180 16178 12232
rect 13630 12152 13636 12164
rect 4632 12124 7144 12152
rect 13591 12124 13636 12152
rect 13630 12112 13636 12124
rect 13688 12112 13694 12164
rect 16776 12152 16804 12248
rect 17678 12220 17684 12232
rect 17639 12192 17684 12220
rect 17678 12180 17684 12192
rect 17736 12180 17742 12232
rect 17954 12220 17960 12232
rect 17915 12192 17960 12220
rect 17954 12180 17960 12192
rect 18012 12180 18018 12232
rect 19337 12223 19395 12229
rect 19337 12189 19349 12223
rect 19383 12220 19395 12223
rect 20070 12220 20076 12232
rect 19383 12192 20076 12220
rect 19383 12189 19395 12192
rect 19337 12183 19395 12189
rect 20070 12180 20076 12192
rect 20128 12180 20134 12232
rect 19889 12155 19947 12161
rect 19889 12152 19901 12155
rect 16776 12124 19901 12152
rect 19889 12121 19901 12124
rect 19935 12152 19947 12155
rect 20622 12152 20628 12164
rect 19935 12124 20628 12152
rect 19935 12121 19947 12124
rect 19889 12115 19947 12121
rect 20622 12112 20628 12124
rect 20680 12112 20686 12164
rect 5261 12087 5319 12093
rect 5261 12053 5273 12087
rect 5307 12084 5319 12087
rect 5534 12084 5540 12096
rect 5307 12056 5540 12084
rect 5307 12053 5319 12056
rect 5261 12047 5319 12053
rect 5534 12044 5540 12056
rect 5592 12044 5598 12096
rect 6546 12084 6552 12096
rect 6507 12056 6552 12084
rect 6546 12044 6552 12056
rect 6604 12044 6610 12096
rect 12158 12084 12164 12096
rect 12119 12056 12164 12084
rect 12158 12044 12164 12056
rect 12216 12044 12222 12096
rect 12526 12084 12532 12096
rect 12487 12056 12532 12084
rect 12526 12044 12532 12056
rect 12584 12044 12590 12096
rect 13354 12044 13360 12096
rect 13412 12084 13418 12096
rect 14550 12084 14556 12096
rect 13412 12056 14556 12084
rect 13412 12044 13418 12056
rect 14550 12044 14556 12056
rect 14608 12044 14614 12096
rect 18414 12044 18420 12096
rect 18472 12084 18478 12096
rect 18601 12087 18659 12093
rect 18601 12084 18613 12087
rect 18472 12056 18613 12084
rect 18472 12044 18478 12056
rect 18601 12053 18613 12056
rect 18647 12053 18659 12087
rect 18601 12047 18659 12053
rect 1104 11994 22816 12016
rect 1104 11942 4982 11994
rect 5034 11942 5046 11994
rect 5098 11942 5110 11994
rect 5162 11942 5174 11994
rect 5226 11942 12982 11994
rect 13034 11942 13046 11994
rect 13098 11942 13110 11994
rect 13162 11942 13174 11994
rect 13226 11942 20982 11994
rect 21034 11942 21046 11994
rect 21098 11942 21110 11994
rect 21162 11942 21174 11994
rect 21226 11942 22816 11994
rect 1104 11920 22816 11942
rect 1854 11840 1860 11892
rect 1912 11880 1918 11892
rect 2961 11883 3019 11889
rect 2961 11880 2973 11883
rect 1912 11852 2973 11880
rect 1912 11840 1918 11852
rect 2961 11849 2973 11852
rect 3007 11880 3019 11883
rect 3510 11880 3516 11892
rect 3007 11852 3516 11880
rect 3007 11849 3019 11852
rect 2961 11843 3019 11849
rect 3510 11840 3516 11852
rect 3568 11840 3574 11892
rect 4065 11883 4123 11889
rect 4065 11849 4077 11883
rect 4111 11880 4123 11883
rect 4246 11880 4252 11892
rect 4111 11852 4252 11880
rect 4111 11849 4123 11852
rect 4065 11843 4123 11849
rect 4246 11840 4252 11852
rect 4304 11880 4310 11892
rect 4341 11883 4399 11889
rect 4341 11880 4353 11883
rect 4304 11852 4353 11880
rect 4304 11840 4310 11852
rect 4341 11849 4353 11852
rect 4387 11849 4399 11883
rect 6457 11883 6515 11889
rect 6457 11880 6469 11883
rect 4341 11843 4399 11849
rect 4724 11852 6469 11880
rect 3528 11812 3556 11840
rect 4724 11812 4752 11852
rect 6457 11849 6469 11852
rect 6503 11880 6515 11883
rect 6549 11883 6607 11889
rect 6549 11880 6561 11883
rect 6503 11852 6561 11880
rect 6503 11849 6515 11852
rect 6457 11843 6515 11849
rect 6549 11849 6561 11852
rect 6595 11849 6607 11883
rect 6549 11843 6607 11849
rect 7190 11840 7196 11892
rect 7248 11880 7254 11892
rect 7745 11883 7803 11889
rect 7745 11880 7757 11883
rect 7248 11852 7757 11880
rect 7248 11840 7254 11852
rect 7745 11849 7757 11852
rect 7791 11849 7803 11883
rect 9582 11880 9588 11892
rect 9543 11852 9588 11880
rect 7745 11843 7803 11849
rect 9582 11840 9588 11852
rect 9640 11840 9646 11892
rect 9766 11840 9772 11892
rect 9824 11880 9830 11892
rect 9861 11883 9919 11889
rect 9861 11880 9873 11883
rect 9824 11852 9873 11880
rect 9824 11840 9830 11852
rect 9861 11849 9873 11852
rect 9907 11849 9919 11883
rect 10226 11880 10232 11892
rect 10187 11852 10232 11880
rect 9861 11843 9919 11849
rect 10226 11840 10232 11852
rect 10284 11840 10290 11892
rect 11238 11840 11244 11892
rect 11296 11880 11302 11892
rect 11793 11883 11851 11889
rect 11793 11880 11805 11883
rect 11296 11852 11805 11880
rect 11296 11840 11302 11852
rect 11793 11849 11805 11852
rect 11839 11849 11851 11883
rect 12158 11880 12164 11892
rect 12119 11852 12164 11880
rect 11793 11843 11851 11849
rect 12158 11840 12164 11852
rect 12216 11840 12222 11892
rect 14642 11880 14648 11892
rect 14603 11852 14648 11880
rect 14642 11840 14648 11852
rect 14700 11840 14706 11892
rect 16114 11840 16120 11892
rect 16172 11880 16178 11892
rect 16393 11883 16451 11889
rect 16393 11880 16405 11883
rect 16172 11852 16405 11880
rect 16172 11840 16178 11852
rect 16393 11849 16405 11852
rect 16439 11880 16451 11883
rect 16715 11883 16773 11889
rect 16715 11880 16727 11883
rect 16439 11852 16727 11880
rect 16439 11849 16451 11852
rect 16393 11843 16451 11849
rect 16715 11849 16727 11852
rect 16761 11849 16773 11883
rect 16715 11843 16773 11849
rect 17681 11883 17739 11889
rect 17681 11849 17693 11883
rect 17727 11880 17739 11883
rect 17770 11880 17776 11892
rect 17727 11852 17776 11880
rect 17727 11849 17739 11852
rect 17681 11843 17739 11849
rect 17770 11840 17776 11852
rect 17828 11840 17834 11892
rect 19426 11880 19432 11892
rect 19387 11852 19432 11880
rect 19426 11840 19432 11852
rect 19484 11880 19490 11892
rect 19705 11883 19763 11889
rect 19705 11880 19717 11883
rect 19484 11852 19717 11880
rect 19484 11840 19490 11852
rect 19705 11849 19717 11852
rect 19751 11849 19763 11883
rect 20070 11880 20076 11892
rect 20031 11852 20076 11880
rect 19705 11843 19763 11849
rect 20070 11840 20076 11852
rect 20128 11880 20134 11892
rect 20395 11883 20453 11889
rect 20395 11880 20407 11883
rect 20128 11852 20407 11880
rect 20128 11840 20134 11852
rect 20395 11849 20407 11852
rect 20441 11849 20453 11883
rect 20395 11843 20453 11849
rect 20806 11840 20812 11892
rect 20864 11880 20870 11892
rect 21085 11883 21143 11889
rect 21085 11880 21097 11883
rect 20864 11852 21097 11880
rect 20864 11840 20870 11852
rect 21085 11849 21097 11852
rect 21131 11849 21143 11883
rect 21085 11843 21143 11849
rect 5994 11812 6000 11824
rect 3528 11784 4752 11812
rect 5092 11784 6000 11812
rect 3142 11744 3148 11756
rect 3103 11716 3148 11744
rect 3142 11704 3148 11716
rect 3200 11704 3206 11756
rect 1397 11679 1455 11685
rect 1397 11645 1409 11679
rect 1443 11676 1455 11679
rect 2041 11679 2099 11685
rect 2041 11676 2053 11679
rect 1443 11648 2053 11676
rect 1443 11645 1455 11648
rect 1397 11639 1455 11645
rect 2041 11645 2053 11648
rect 2087 11676 2099 11679
rect 5092 11676 5120 11784
rect 5994 11772 6000 11784
rect 6052 11812 6058 11824
rect 6273 11815 6331 11821
rect 6273 11812 6285 11815
rect 6052 11784 6285 11812
rect 6052 11772 6058 11784
rect 6273 11781 6285 11784
rect 6319 11812 6331 11815
rect 8570 11812 8576 11824
rect 6319 11784 8576 11812
rect 6319 11781 6331 11784
rect 6273 11775 6331 11781
rect 8570 11772 8576 11784
rect 8628 11772 8634 11824
rect 5905 11747 5963 11753
rect 5905 11713 5917 11747
rect 5951 11744 5963 11747
rect 6546 11744 6552 11756
rect 5951 11716 6552 11744
rect 5951 11713 5963 11716
rect 5905 11707 5963 11713
rect 6546 11704 6552 11716
rect 6604 11744 6610 11756
rect 6825 11747 6883 11753
rect 6825 11744 6837 11747
rect 6604 11716 6837 11744
rect 6604 11704 6610 11716
rect 6825 11713 6837 11716
rect 6871 11713 6883 11747
rect 6825 11707 6883 11713
rect 8665 11747 8723 11753
rect 8665 11713 8677 11747
rect 8711 11744 8723 11747
rect 8846 11744 8852 11756
rect 8711 11716 8852 11744
rect 8711 11713 8723 11716
rect 8665 11707 8723 11713
rect 8846 11704 8852 11716
rect 8904 11704 8910 11756
rect 10244 11744 10272 11840
rect 10410 11772 10416 11824
rect 10468 11812 10474 11824
rect 13630 11812 13636 11824
rect 10468 11784 13636 11812
rect 10468 11772 10474 11784
rect 12820 11753 12848 11784
rect 13630 11772 13636 11784
rect 13688 11772 13694 11824
rect 15749 11815 15807 11821
rect 15749 11781 15761 11815
rect 15795 11781 15807 11815
rect 15749 11775 15807 11781
rect 12805 11747 12863 11753
rect 10244 11716 10916 11744
rect 2087 11648 5120 11676
rect 5445 11679 5503 11685
rect 2087 11645 2099 11648
rect 2041 11639 2099 11645
rect 5445 11645 5457 11679
rect 5491 11676 5503 11679
rect 5534 11676 5540 11688
rect 5491 11648 5540 11676
rect 5491 11645 5503 11648
rect 5445 11639 5503 11645
rect 5534 11636 5540 11648
rect 5592 11636 5598 11688
rect 5718 11676 5724 11688
rect 5679 11648 5724 11676
rect 5718 11636 5724 11648
rect 5776 11636 5782 11688
rect 10502 11676 10508 11688
rect 10463 11648 10508 11676
rect 10502 11636 10508 11648
rect 10560 11636 10566 11688
rect 10888 11685 10916 11716
rect 12805 11713 12817 11747
rect 12851 11713 12863 11747
rect 15764 11744 15792 11775
rect 16117 11747 16175 11753
rect 16117 11744 16129 11747
rect 15764 11716 16129 11744
rect 12805 11707 12863 11713
rect 16117 11713 16129 11716
rect 16163 11744 16175 11747
rect 16206 11744 16212 11756
rect 16163 11716 16212 11744
rect 16163 11713 16175 11716
rect 16117 11707 16175 11713
rect 16206 11704 16212 11716
rect 16264 11704 16270 11756
rect 10873 11679 10931 11685
rect 10873 11645 10885 11679
rect 10919 11645 10931 11679
rect 14826 11676 14832 11688
rect 14787 11648 14832 11676
rect 10873 11639 10931 11645
rect 14826 11636 14832 11648
rect 14884 11636 14890 11688
rect 15838 11636 15844 11688
rect 15896 11676 15902 11688
rect 16612 11679 16670 11685
rect 16612 11676 16624 11679
rect 15896 11648 16624 11676
rect 15896 11636 15902 11648
rect 16612 11645 16624 11648
rect 16658 11676 16670 11679
rect 16850 11676 16856 11688
rect 16658 11648 16856 11676
rect 16658 11645 16670 11648
rect 16612 11639 16670 11645
rect 16850 11636 16856 11648
rect 16908 11676 16914 11688
rect 17037 11679 17095 11685
rect 17037 11676 17049 11679
rect 16908 11648 17049 11676
rect 16908 11636 16914 11648
rect 17037 11645 17049 11648
rect 17083 11645 17095 11679
rect 17037 11639 17095 11645
rect 18414 11636 18420 11688
rect 18472 11676 18478 11688
rect 18509 11679 18567 11685
rect 18509 11676 18521 11679
rect 18472 11648 18521 11676
rect 18472 11636 18478 11648
rect 18509 11645 18521 11648
rect 18555 11645 18567 11679
rect 18509 11639 18567 11645
rect 20324 11679 20382 11685
rect 20324 11645 20336 11679
rect 20370 11676 20382 11679
rect 20714 11676 20720 11688
rect 20370 11648 20720 11676
rect 20370 11645 20382 11648
rect 20324 11639 20382 11645
rect 20714 11636 20720 11648
rect 20772 11676 20778 11688
rect 21542 11676 21548 11688
rect 20772 11648 21548 11676
rect 20772 11636 20778 11648
rect 21542 11636 21548 11648
rect 21600 11636 21606 11688
rect 2501 11611 2559 11617
rect 2501 11577 2513 11611
rect 2547 11608 2559 11611
rect 2866 11608 2872 11620
rect 2547 11580 2872 11608
rect 2547 11577 2559 11580
rect 2501 11571 2559 11577
rect 2866 11568 2872 11580
rect 2924 11608 2930 11620
rect 3510 11617 3516 11620
rect 3507 11608 3516 11617
rect 2924 11580 3418 11608
rect 3471 11580 3516 11608
rect 2924 11568 2930 11580
rect 106 11500 112 11552
rect 164 11540 170 11552
rect 1581 11543 1639 11549
rect 1581 11540 1593 11543
rect 164 11512 1593 11540
rect 164 11500 170 11512
rect 1581 11509 1593 11512
rect 1627 11509 1639 11543
rect 3390 11540 3418 11580
rect 3507 11571 3516 11580
rect 3510 11568 3516 11571
rect 3568 11568 3574 11620
rect 5077 11611 5135 11617
rect 5077 11577 5089 11611
rect 5123 11608 5135 11611
rect 5736 11608 5764 11636
rect 8986 11611 9044 11617
rect 8986 11608 8998 11611
rect 5123 11580 5764 11608
rect 8128 11580 8998 11608
rect 5123 11577 5135 11580
rect 5077 11571 5135 11577
rect 5092 11540 5120 11571
rect 8128 11552 8156 11580
rect 8986 11577 8998 11580
rect 9032 11608 9044 11611
rect 11146 11608 11152 11620
rect 9032 11580 9674 11608
rect 11107 11580 11152 11608
rect 9032 11577 9044 11580
rect 8986 11571 9044 11577
rect 3390 11512 5120 11540
rect 6457 11543 6515 11549
rect 1581 11503 1639 11509
rect 6457 11509 6469 11543
rect 6503 11540 6515 11543
rect 7193 11543 7251 11549
rect 7193 11540 7205 11543
rect 6503 11512 7205 11540
rect 6503 11509 6515 11512
rect 6457 11503 6515 11509
rect 7193 11509 7205 11512
rect 7239 11540 7251 11543
rect 8110 11540 8116 11552
rect 7239 11512 8116 11540
rect 7239 11509 7251 11512
rect 7193 11503 7251 11509
rect 8110 11500 8116 11512
rect 8168 11500 8174 11552
rect 8386 11540 8392 11552
rect 8347 11512 8392 11540
rect 8386 11500 8392 11512
rect 8444 11500 8450 11552
rect 9646 11540 9674 11580
rect 11146 11568 11152 11580
rect 11204 11568 11210 11620
rect 12526 11608 12532 11620
rect 12487 11580 12532 11608
rect 12526 11568 12532 11580
rect 12584 11568 12590 11620
rect 12621 11611 12679 11617
rect 12621 11577 12633 11611
rect 12667 11577 12679 11611
rect 12621 11571 12679 11577
rect 11238 11540 11244 11552
rect 9646 11512 11244 11540
rect 11238 11500 11244 11512
rect 11296 11540 11302 11552
rect 11425 11543 11483 11549
rect 11425 11540 11437 11543
rect 11296 11512 11437 11540
rect 11296 11500 11302 11512
rect 11425 11509 11437 11512
rect 11471 11509 11483 11543
rect 11425 11503 11483 11509
rect 12158 11500 12164 11552
rect 12216 11540 12222 11552
rect 12636 11540 12664 11571
rect 14642 11568 14648 11620
rect 14700 11608 14706 11620
rect 15150 11611 15208 11617
rect 15150 11608 15162 11611
rect 14700 11580 15162 11608
rect 14700 11568 14706 11580
rect 15150 11577 15162 11580
rect 15196 11608 15208 11611
rect 15746 11608 15752 11620
rect 15196 11580 15752 11608
rect 15196 11577 15208 11580
rect 15150 11571 15208 11577
rect 15746 11568 15752 11580
rect 15804 11608 15810 11620
rect 18874 11617 18880 11620
rect 18325 11611 18383 11617
rect 18325 11608 18337 11611
rect 15804 11580 18337 11608
rect 15804 11568 15810 11580
rect 18325 11577 18337 11580
rect 18371 11608 18383 11611
rect 18830 11611 18880 11617
rect 18830 11608 18842 11611
rect 18371 11580 18842 11608
rect 18371 11577 18383 11580
rect 18325 11571 18383 11577
rect 18830 11577 18842 11580
rect 18876 11577 18880 11611
rect 18830 11571 18880 11577
rect 18874 11568 18880 11571
rect 18932 11568 18938 11620
rect 13446 11540 13452 11552
rect 12216 11512 12664 11540
rect 13407 11512 13452 11540
rect 12216 11500 12222 11512
rect 13446 11500 13452 11512
rect 13504 11500 13510 11552
rect 13814 11500 13820 11552
rect 13872 11540 13878 11552
rect 13872 11512 13917 11540
rect 13872 11500 13878 11512
rect 1104 11450 22816 11472
rect 1104 11398 8982 11450
rect 9034 11398 9046 11450
rect 9098 11398 9110 11450
rect 9162 11398 9174 11450
rect 9226 11398 16982 11450
rect 17034 11398 17046 11450
rect 17098 11398 17110 11450
rect 17162 11398 17174 11450
rect 17226 11398 22816 11450
rect 1104 11376 22816 11398
rect 3142 11296 3148 11348
rect 3200 11336 3206 11348
rect 3421 11339 3479 11345
rect 3421 11336 3433 11339
rect 3200 11308 3433 11336
rect 3200 11296 3206 11308
rect 3421 11305 3433 11308
rect 3467 11305 3479 11339
rect 3421 11299 3479 11305
rect 4154 11296 4160 11348
rect 4212 11336 4218 11348
rect 4617 11339 4675 11345
rect 4617 11336 4629 11339
rect 4212 11308 4629 11336
rect 4212 11296 4218 11308
rect 4617 11305 4629 11308
rect 4663 11305 4675 11339
rect 6270 11336 6276 11348
rect 6231 11308 6276 11336
rect 4617 11299 4675 11305
rect 6270 11296 6276 11308
rect 6328 11296 6334 11348
rect 7190 11296 7196 11348
rect 7248 11336 7254 11348
rect 7377 11339 7435 11345
rect 7377 11336 7389 11339
rect 7248 11308 7389 11336
rect 7248 11296 7254 11308
rect 7377 11305 7389 11308
rect 7423 11305 7435 11339
rect 7377 11299 7435 11305
rect 8110 11296 8116 11348
rect 8168 11336 8174 11348
rect 8665 11339 8723 11345
rect 8665 11336 8677 11339
rect 8168 11308 8677 11336
rect 8168 11296 8174 11308
rect 8665 11305 8677 11308
rect 8711 11305 8723 11339
rect 8665 11299 8723 11305
rect 9493 11339 9551 11345
rect 9493 11305 9505 11339
rect 9539 11336 9551 11339
rect 9582 11336 9588 11348
rect 9539 11308 9588 11336
rect 9539 11305 9551 11308
rect 9493 11299 9551 11305
rect 9582 11296 9588 11308
rect 9640 11296 9646 11348
rect 9677 11339 9735 11345
rect 9677 11305 9689 11339
rect 9723 11336 9735 11339
rect 9766 11336 9772 11348
rect 9723 11308 9772 11336
rect 9723 11305 9735 11308
rect 9677 11299 9735 11305
rect 9766 11296 9772 11308
rect 9824 11296 9830 11348
rect 12161 11339 12219 11345
rect 12161 11305 12173 11339
rect 12207 11336 12219 11339
rect 13446 11336 13452 11348
rect 12207 11308 13452 11336
rect 12207 11305 12219 11308
rect 12161 11299 12219 11305
rect 13446 11296 13452 11308
rect 13504 11296 13510 11348
rect 17589 11339 17647 11345
rect 17589 11305 17601 11339
rect 17635 11336 17647 11339
rect 17678 11336 17684 11348
rect 17635 11308 17684 11336
rect 17635 11305 17647 11308
rect 17589 11299 17647 11305
rect 17678 11296 17684 11308
rect 17736 11296 17742 11348
rect 2314 11228 2320 11280
rect 2372 11268 2378 11280
rect 3050 11268 3056 11280
rect 2372 11240 3056 11268
rect 2372 11228 2378 11240
rect 2700 11209 2728 11240
rect 3050 11228 3056 11240
rect 3108 11228 3114 11280
rect 4985 11271 5043 11277
rect 4985 11237 4997 11271
rect 5031 11268 5043 11271
rect 5350 11268 5356 11280
rect 5031 11240 5356 11268
rect 5031 11237 5043 11240
rect 4985 11231 5043 11237
rect 5350 11228 5356 11240
rect 5408 11228 5414 11280
rect 7650 11268 7656 11280
rect 6380 11240 7656 11268
rect 2685 11203 2743 11209
rect 2685 11169 2697 11203
rect 2731 11169 2743 11203
rect 2685 11163 2743 11169
rect 2774 11160 2780 11212
rect 2832 11200 2838 11212
rect 2961 11203 3019 11209
rect 2961 11200 2973 11203
rect 2832 11172 2973 11200
rect 2832 11160 2838 11172
rect 2961 11169 2973 11172
rect 3007 11200 3019 11203
rect 4706 11200 4712 11212
rect 3007 11172 4712 11200
rect 3007 11169 3019 11172
rect 2961 11163 3019 11169
rect 4706 11160 4712 11172
rect 4764 11160 4770 11212
rect 5534 11160 5540 11212
rect 5592 11200 5598 11212
rect 5994 11200 6000 11212
rect 5592 11172 6000 11200
rect 5592 11160 5598 11172
rect 5994 11160 6000 11172
rect 6052 11200 6058 11212
rect 6380 11209 6408 11240
rect 7650 11228 7656 11240
rect 7708 11228 7714 11280
rect 11330 11228 11336 11280
rect 11388 11268 11394 11280
rect 11562 11271 11620 11277
rect 11562 11268 11574 11271
rect 11388 11240 11574 11268
rect 11388 11228 11394 11240
rect 11562 11237 11574 11240
rect 11608 11237 11620 11271
rect 11562 11231 11620 11237
rect 14369 11271 14427 11277
rect 14369 11237 14381 11271
rect 14415 11268 14427 11271
rect 14826 11268 14832 11280
rect 14415 11240 14832 11268
rect 14415 11237 14427 11240
rect 14369 11231 14427 11237
rect 14826 11228 14832 11240
rect 14884 11228 14890 11280
rect 18414 11268 18420 11280
rect 18375 11240 18420 11268
rect 18414 11228 18420 11240
rect 18472 11228 18478 11280
rect 6365 11203 6423 11209
rect 6365 11200 6377 11203
rect 6052 11172 6377 11200
rect 6052 11160 6058 11172
rect 6365 11169 6377 11172
rect 6411 11169 6423 11203
rect 6822 11200 6828 11212
rect 6783 11172 6828 11200
rect 6365 11163 6423 11169
rect 6822 11160 6828 11172
rect 6880 11160 6886 11212
rect 7996 11203 8054 11209
rect 7996 11169 8008 11203
rect 8042 11200 8054 11203
rect 8110 11200 8116 11212
rect 8042 11172 8116 11200
rect 8042 11169 8054 11172
rect 7996 11163 8054 11169
rect 8110 11160 8116 11172
rect 8168 11200 8174 11212
rect 8570 11200 8576 11212
rect 8168 11172 8576 11200
rect 8168 11160 8174 11172
rect 8570 11160 8576 11172
rect 8628 11160 8634 11212
rect 11146 11160 11152 11212
rect 11204 11200 11210 11212
rect 11241 11203 11299 11209
rect 11241 11200 11253 11203
rect 11204 11172 11253 11200
rect 11204 11160 11210 11172
rect 11241 11169 11253 11172
rect 11287 11169 11299 11203
rect 13630 11200 13636 11212
rect 13591 11172 13636 11200
rect 11241 11163 11299 11169
rect 13630 11160 13636 11172
rect 13688 11160 13694 11212
rect 14182 11200 14188 11212
rect 14143 11172 14188 11200
rect 14182 11160 14188 11172
rect 14240 11160 14246 11212
rect 15194 11160 15200 11212
rect 15252 11200 15258 11212
rect 15356 11203 15414 11209
rect 15356 11200 15368 11203
rect 15252 11172 15368 11200
rect 15252 11160 15258 11172
rect 15356 11169 15368 11172
rect 15402 11200 15414 11203
rect 16206 11200 16212 11212
rect 15402 11172 16212 11200
rect 15402 11169 15414 11172
rect 15356 11163 15414 11169
rect 16206 11160 16212 11172
rect 16264 11200 16270 11212
rect 16336 11203 16394 11209
rect 16336 11200 16348 11203
rect 16264 11172 16348 11200
rect 16264 11160 16270 11172
rect 16336 11169 16348 11172
rect 16382 11169 16394 11203
rect 16336 11163 16394 11169
rect 17494 11160 17500 11212
rect 17552 11200 17558 11212
rect 17681 11203 17739 11209
rect 17681 11200 17693 11203
rect 17552 11172 17693 11200
rect 17552 11160 17558 11172
rect 17681 11169 17693 11172
rect 17727 11169 17739 11203
rect 18138 11200 18144 11212
rect 18099 11172 18144 11200
rect 17681 11163 17739 11169
rect 18138 11160 18144 11172
rect 18196 11160 18202 11212
rect 19426 11209 19432 11212
rect 19404 11203 19432 11209
rect 19404 11200 19416 11203
rect 19339 11172 19416 11200
rect 19404 11169 19416 11172
rect 19484 11200 19490 11212
rect 20346 11200 20352 11212
rect 19484 11172 20352 11200
rect 19404 11163 19432 11169
rect 19426 11160 19432 11163
rect 19484 11160 19490 11172
rect 20346 11160 20352 11172
rect 20404 11160 20410 11212
rect 1397 11135 1455 11141
rect 1397 11101 1409 11135
rect 1443 11132 1455 11135
rect 3142 11132 3148 11144
rect 1443 11104 1808 11132
rect 3103 11104 3148 11132
rect 1443 11101 1455 11104
rect 1397 11095 1455 11101
rect 1780 11008 1808 11104
rect 3142 11092 3148 11104
rect 3200 11092 3206 11144
rect 4893 11135 4951 11141
rect 4893 11132 4905 11135
rect 4816 11104 4905 11132
rect 4816 11076 4844 11104
rect 4893 11101 4905 11104
rect 4939 11101 4951 11135
rect 6914 11132 6920 11144
rect 6875 11104 6920 11132
rect 4893 11095 4951 11101
rect 6914 11092 6920 11104
rect 6972 11092 6978 11144
rect 4798 11024 4804 11076
rect 4856 11024 4862 11076
rect 5442 11064 5448 11076
rect 5403 11036 5448 11064
rect 5442 11024 5448 11036
rect 5500 11024 5506 11076
rect 15427 11067 15485 11073
rect 15427 11064 15439 11067
rect 14292 11036 15439 11064
rect 1762 10956 1768 11008
rect 1820 10996 1826 11008
rect 1857 10999 1915 11005
rect 1857 10996 1869 10999
rect 1820 10968 1869 10996
rect 1820 10956 1826 10968
rect 1857 10965 1869 10968
rect 1903 10965 1915 10999
rect 1857 10959 1915 10965
rect 2317 10999 2375 11005
rect 2317 10965 2329 10999
rect 2363 10996 2375 10999
rect 2590 10996 2596 11008
rect 2363 10968 2596 10996
rect 2363 10965 2375 10968
rect 2317 10959 2375 10965
rect 2590 10956 2596 10968
rect 2648 10996 2654 11008
rect 3510 10996 3516 11008
rect 2648 10968 3516 10996
rect 2648 10956 2654 10968
rect 3510 10956 3516 10968
rect 3568 10956 3574 11008
rect 4246 10996 4252 11008
rect 4207 10968 4252 10996
rect 4246 10956 4252 10968
rect 4304 10956 4310 11008
rect 7742 10996 7748 11008
rect 7703 10968 7748 10996
rect 7742 10956 7748 10968
rect 7800 10956 7806 11008
rect 7926 10956 7932 11008
rect 7984 10996 7990 11008
rect 8067 10999 8125 11005
rect 8067 10996 8079 10999
rect 7984 10968 8079 10996
rect 7984 10956 7990 10968
rect 8067 10965 8079 10968
rect 8113 10965 8125 10999
rect 10502 10996 10508 11008
rect 10463 10968 10508 10996
rect 8067 10959 8125 10965
rect 10502 10956 10508 10968
rect 10560 10956 10566 11008
rect 12342 10956 12348 11008
rect 12400 10996 12406 11008
rect 12437 10999 12495 11005
rect 12437 10996 12449 10999
rect 12400 10968 12449 10996
rect 12400 10956 12406 10968
rect 12437 10965 12449 10968
rect 12483 10965 12495 10999
rect 12437 10959 12495 10965
rect 13722 10956 13728 11008
rect 13780 10996 13786 11008
rect 14292 10996 14320 11036
rect 15427 11033 15439 11036
rect 15473 11033 15485 11067
rect 15427 11027 15485 11033
rect 13780 10968 14320 10996
rect 16439 10999 16497 11005
rect 13780 10956 13786 10968
rect 16439 10965 16451 10999
rect 16485 10996 16497 10999
rect 16574 10996 16580 11008
rect 16485 10968 16580 10996
rect 16485 10965 16497 10968
rect 16439 10959 16497 10965
rect 16574 10956 16580 10968
rect 16632 10956 16638 11008
rect 19475 10999 19533 11005
rect 19475 10965 19487 10999
rect 19521 10996 19533 10999
rect 19610 10996 19616 11008
rect 19521 10968 19616 10996
rect 19521 10965 19533 10968
rect 19475 10959 19533 10965
rect 19610 10956 19616 10968
rect 19668 10956 19674 11008
rect 19794 10996 19800 11008
rect 19755 10968 19800 10996
rect 19794 10956 19800 10968
rect 19852 10956 19858 11008
rect 1104 10906 22816 10928
rect 1104 10854 4982 10906
rect 5034 10854 5046 10906
rect 5098 10854 5110 10906
rect 5162 10854 5174 10906
rect 5226 10854 12982 10906
rect 13034 10854 13046 10906
rect 13098 10854 13110 10906
rect 13162 10854 13174 10906
rect 13226 10854 20982 10906
rect 21034 10854 21046 10906
rect 21098 10854 21110 10906
rect 21162 10854 21174 10906
rect 21226 10854 22816 10906
rect 1104 10832 22816 10854
rect 2222 10752 2228 10804
rect 2280 10792 2286 10804
rect 3375 10795 3433 10801
rect 3375 10792 3387 10795
rect 2280 10764 3387 10792
rect 2280 10752 2286 10764
rect 3375 10761 3387 10764
rect 3421 10761 3433 10795
rect 3375 10755 3433 10761
rect 3602 10752 3608 10804
rect 3660 10792 3666 10804
rect 3973 10795 4031 10801
rect 3973 10792 3985 10795
rect 3660 10764 3985 10792
rect 3660 10752 3666 10764
rect 3973 10761 3985 10764
rect 4019 10792 4031 10795
rect 4065 10795 4123 10801
rect 4065 10792 4077 10795
rect 4019 10764 4077 10792
rect 4019 10761 4031 10764
rect 3973 10755 4031 10761
rect 4065 10761 4077 10764
rect 4111 10761 4123 10795
rect 4065 10755 4123 10761
rect 5169 10795 5227 10801
rect 5169 10761 5181 10795
rect 5215 10792 5227 10795
rect 5350 10792 5356 10804
rect 5215 10764 5356 10792
rect 5215 10761 5227 10764
rect 5169 10755 5227 10761
rect 5350 10752 5356 10764
rect 5408 10792 5414 10804
rect 5445 10795 5503 10801
rect 5445 10792 5457 10795
rect 5408 10764 5457 10792
rect 5408 10752 5414 10764
rect 5445 10761 5457 10764
rect 5491 10761 5503 10795
rect 8110 10792 8116 10804
rect 8071 10764 8116 10792
rect 5445 10755 5503 10761
rect 8110 10752 8116 10764
rect 8168 10752 8174 10804
rect 9217 10795 9275 10801
rect 9217 10761 9229 10795
rect 9263 10792 9275 10795
rect 10226 10792 10232 10804
rect 9263 10764 10232 10792
rect 9263 10761 9275 10764
rect 9217 10755 9275 10761
rect 2774 10724 2780 10736
rect 2735 10696 2780 10724
rect 2774 10684 2780 10696
rect 2832 10684 2838 10736
rect 4706 10684 4712 10736
rect 4764 10724 4770 10736
rect 6365 10727 6423 10733
rect 6365 10724 6377 10727
rect 4764 10696 6377 10724
rect 4764 10684 4770 10696
rect 6365 10693 6377 10696
rect 6411 10724 6423 10727
rect 6822 10724 6828 10736
rect 6411 10696 6828 10724
rect 6411 10693 6423 10696
rect 6365 10687 6423 10693
rect 6822 10684 6828 10696
rect 6880 10684 6886 10736
rect 1762 10656 1768 10668
rect 1723 10628 1768 10656
rect 1762 10616 1768 10628
rect 1820 10616 1826 10668
rect 3602 10616 3608 10668
rect 3660 10656 3666 10668
rect 4246 10656 4252 10668
rect 3660 10628 4252 10656
rect 3660 10616 3666 10628
rect 4246 10616 4252 10628
rect 4304 10616 4310 10668
rect 7466 10656 7472 10668
rect 7427 10628 7472 10656
rect 7466 10616 7472 10628
rect 7524 10616 7530 10668
rect 2409 10591 2467 10597
rect 2409 10557 2421 10591
rect 2455 10588 2467 10591
rect 3272 10591 3330 10597
rect 3272 10588 3284 10591
rect 2455 10560 3284 10588
rect 2455 10557 2467 10560
rect 2409 10551 2467 10557
rect 3272 10557 3284 10560
rect 3318 10588 3330 10591
rect 3697 10591 3755 10597
rect 3697 10588 3709 10591
rect 3318 10560 3709 10588
rect 3318 10557 3330 10560
rect 3272 10551 3330 10557
rect 3697 10557 3709 10560
rect 3743 10588 3755 10591
rect 5442 10588 5448 10600
rect 3743 10560 5448 10588
rect 3743 10557 3755 10560
rect 3697 10551 3755 10557
rect 5442 10548 5448 10560
rect 5500 10548 5506 10600
rect 9306 10588 9312 10600
rect 9267 10560 9312 10588
rect 9306 10548 9312 10560
rect 9364 10548 9370 10600
rect 9876 10597 9904 10764
rect 10226 10752 10232 10764
rect 10284 10752 10290 10804
rect 10873 10795 10931 10801
rect 10873 10761 10885 10795
rect 10919 10792 10931 10795
rect 11146 10792 11152 10804
rect 10919 10764 11152 10792
rect 10919 10761 10931 10764
rect 10873 10755 10931 10761
rect 11146 10752 11152 10764
rect 11204 10752 11210 10804
rect 11885 10795 11943 10801
rect 11885 10761 11897 10795
rect 11931 10792 11943 10795
rect 11974 10792 11980 10804
rect 11931 10764 11980 10792
rect 11931 10761 11943 10764
rect 11885 10755 11943 10761
rect 9861 10591 9919 10597
rect 9861 10557 9873 10591
rect 9907 10557 9919 10591
rect 9861 10551 9919 10557
rect 11400 10591 11458 10597
rect 11400 10557 11412 10591
rect 11446 10588 11458 10591
rect 11900 10588 11928 10755
rect 11974 10752 11980 10764
rect 12032 10792 12038 10804
rect 13446 10792 13452 10804
rect 12032 10764 13452 10792
rect 12032 10752 12038 10764
rect 13446 10752 13452 10764
rect 13504 10752 13510 10804
rect 16850 10752 16856 10804
rect 16908 10792 16914 10804
rect 17129 10795 17187 10801
rect 17129 10792 17141 10795
rect 16908 10764 17141 10792
rect 16908 10752 16914 10764
rect 17129 10761 17141 10764
rect 17175 10761 17187 10795
rect 17129 10755 17187 10761
rect 17144 10724 17172 10755
rect 17678 10752 17684 10804
rect 17736 10792 17742 10804
rect 18187 10795 18245 10801
rect 18187 10792 18199 10795
rect 17736 10764 18199 10792
rect 17736 10752 17742 10764
rect 18187 10761 18199 10764
rect 18233 10761 18245 10795
rect 19426 10792 19432 10804
rect 19387 10764 19432 10792
rect 18187 10755 18245 10761
rect 19426 10752 19432 10764
rect 19484 10752 19490 10804
rect 21266 10792 21272 10804
rect 21227 10764 21272 10792
rect 21266 10752 21272 10764
rect 21324 10752 21330 10804
rect 17144 10696 20300 10724
rect 12802 10656 12808 10668
rect 12763 10628 12808 10656
rect 12802 10616 12808 10628
rect 12860 10656 12866 10668
rect 13814 10656 13820 10668
rect 12860 10628 13820 10656
rect 12860 10616 12866 10628
rect 13814 10616 13820 10628
rect 13872 10616 13878 10668
rect 16758 10656 16764 10668
rect 14752 10628 16764 10656
rect 14093 10591 14151 10597
rect 14093 10588 14105 10591
rect 11446 10560 11928 10588
rect 13786 10560 14105 10588
rect 11446 10557 11458 10560
rect 11400 10551 11458 10557
rect 1857 10523 1915 10529
rect 1857 10489 1869 10523
rect 1903 10520 1915 10523
rect 2222 10520 2228 10532
rect 1903 10492 2228 10520
rect 1903 10489 1915 10492
rect 1857 10483 1915 10489
rect 2222 10480 2228 10492
rect 2280 10480 2286 10532
rect 3973 10523 4031 10529
rect 3973 10489 3985 10523
rect 4019 10520 4031 10523
rect 4430 10520 4436 10532
rect 4019 10492 4436 10520
rect 4019 10489 4031 10492
rect 3973 10483 4031 10489
rect 4430 10480 4436 10492
rect 4488 10520 4494 10532
rect 4570 10523 4628 10529
rect 4570 10520 4582 10523
rect 4488 10492 4582 10520
rect 4488 10480 4494 10492
rect 4570 10489 4582 10492
rect 4616 10489 4628 10523
rect 7190 10520 7196 10532
rect 7151 10492 7196 10520
rect 4570 10483 4628 10489
rect 7190 10480 7196 10492
rect 7248 10480 7254 10532
rect 7285 10523 7343 10529
rect 7285 10489 7297 10523
rect 7331 10520 7343 10523
rect 7650 10520 7656 10532
rect 7331 10492 7656 10520
rect 7331 10489 7343 10492
rect 7285 10483 7343 10489
rect 7650 10480 7656 10492
rect 7708 10480 7714 10532
rect 10042 10520 10048 10532
rect 10003 10492 10048 10520
rect 10042 10480 10048 10492
rect 10100 10480 10106 10532
rect 12342 10480 12348 10532
rect 12400 10520 12406 10532
rect 12529 10523 12587 10529
rect 12529 10520 12541 10523
rect 12400 10492 12541 10520
rect 12400 10480 12406 10492
rect 12529 10489 12541 10492
rect 12575 10489 12587 10523
rect 12529 10483 12587 10489
rect 12621 10523 12679 10529
rect 12621 10489 12633 10523
rect 12667 10489 12679 10523
rect 12621 10483 12679 10489
rect 3050 10452 3056 10464
rect 3011 10424 3056 10452
rect 3050 10412 3056 10424
rect 3108 10412 3114 10464
rect 5994 10452 6000 10464
rect 5955 10424 6000 10452
rect 5994 10412 6000 10424
rect 6052 10412 6058 10464
rect 11146 10452 11152 10464
rect 11107 10424 11152 10452
rect 11146 10412 11152 10424
rect 11204 10412 11210 10464
rect 11471 10455 11529 10461
rect 11471 10421 11483 10455
rect 11517 10452 11529 10455
rect 11698 10452 11704 10464
rect 11517 10424 11704 10452
rect 11517 10421 11529 10424
rect 11471 10415 11529 10421
rect 11698 10412 11704 10424
rect 11756 10412 11762 10464
rect 12158 10452 12164 10464
rect 12119 10424 12164 10452
rect 12158 10412 12164 10424
rect 12216 10452 12222 10464
rect 12636 10452 12664 10483
rect 13170 10480 13176 10532
rect 13228 10520 13234 10532
rect 13786 10520 13814 10560
rect 14093 10557 14105 10560
rect 14139 10588 14151 10591
rect 14182 10588 14188 10600
rect 14139 10560 14188 10588
rect 14139 10557 14151 10560
rect 14093 10551 14151 10557
rect 14182 10548 14188 10560
rect 14240 10588 14246 10600
rect 14752 10597 14780 10628
rect 16758 10616 16764 10628
rect 16816 10616 16822 10668
rect 17494 10616 17500 10668
rect 17552 10656 17558 10668
rect 17681 10659 17739 10665
rect 17681 10656 17693 10659
rect 17552 10628 17693 10656
rect 17552 10616 17558 10628
rect 17681 10625 17693 10628
rect 17727 10625 17739 10659
rect 19610 10656 19616 10668
rect 19571 10628 19616 10656
rect 17681 10619 17739 10625
rect 19610 10616 19616 10628
rect 19668 10616 19674 10668
rect 19886 10656 19892 10668
rect 19847 10628 19892 10656
rect 19886 10616 19892 10628
rect 19944 10616 19950 10668
rect 14737 10591 14795 10597
rect 14737 10588 14749 10591
rect 14240 10560 14749 10588
rect 14240 10548 14246 10560
rect 14737 10557 14749 10560
rect 14783 10557 14795 10591
rect 15013 10591 15071 10597
rect 15013 10588 15025 10591
rect 14737 10551 14795 10557
rect 14844 10560 15025 10588
rect 13228 10492 13814 10520
rect 13228 10480 13234 10492
rect 14366 10480 14372 10532
rect 14424 10520 14430 10532
rect 14461 10523 14519 10529
rect 14461 10520 14473 10523
rect 14424 10492 14473 10520
rect 14424 10480 14430 10492
rect 14461 10489 14473 10492
rect 14507 10520 14519 10523
rect 14844 10520 14872 10560
rect 15013 10557 15025 10560
rect 15059 10557 15071 10591
rect 15013 10551 15071 10557
rect 16368 10591 16426 10597
rect 16368 10557 16380 10591
rect 16414 10588 16426 10591
rect 16850 10588 16856 10600
rect 16414 10560 16856 10588
rect 16414 10557 16426 10560
rect 16368 10551 16426 10557
rect 16850 10548 16856 10560
rect 16908 10548 16914 10600
rect 17862 10548 17868 10600
rect 17920 10588 17926 10600
rect 18084 10591 18142 10597
rect 18084 10588 18096 10591
rect 17920 10560 18096 10588
rect 17920 10548 17926 10560
rect 18084 10557 18096 10560
rect 18130 10588 18142 10591
rect 18509 10591 18567 10597
rect 18509 10588 18521 10591
rect 18130 10560 18521 10588
rect 18130 10557 18142 10560
rect 18084 10551 18142 10557
rect 18509 10557 18521 10560
rect 18555 10557 18567 10591
rect 20272 10588 20300 10696
rect 21085 10591 21143 10597
rect 21085 10588 21097 10591
rect 20272 10560 21097 10588
rect 18509 10551 18567 10557
rect 21085 10557 21097 10560
rect 21131 10588 21143 10591
rect 21637 10591 21695 10597
rect 21637 10588 21649 10591
rect 21131 10560 21649 10588
rect 21131 10557 21143 10560
rect 21085 10551 21143 10557
rect 21637 10557 21649 10560
rect 21683 10557 21695 10591
rect 21637 10551 21695 10557
rect 14507 10492 14872 10520
rect 15289 10523 15347 10529
rect 14507 10489 14519 10492
rect 14461 10483 14519 10489
rect 15289 10489 15301 10523
rect 15335 10520 15347 10523
rect 15378 10520 15384 10532
rect 15335 10492 15384 10520
rect 15335 10489 15347 10492
rect 15289 10483 15347 10489
rect 15378 10480 15384 10492
rect 15436 10480 15442 10532
rect 15657 10523 15715 10529
rect 15657 10489 15669 10523
rect 15703 10520 15715 10523
rect 16206 10520 16212 10532
rect 15703 10492 16212 10520
rect 15703 10489 15715 10492
rect 15657 10483 15715 10489
rect 16206 10480 16212 10492
rect 16264 10520 16270 10532
rect 18877 10523 18935 10529
rect 18877 10520 18889 10523
rect 16264 10492 16896 10520
rect 16264 10480 16270 10492
rect 12216 10424 12664 10452
rect 12216 10412 12222 10424
rect 12710 10412 12716 10464
rect 12768 10452 12774 10464
rect 13630 10452 13636 10464
rect 12768 10424 13636 10452
rect 12768 10412 12774 10424
rect 13630 10412 13636 10424
rect 13688 10412 13694 10464
rect 16439 10455 16497 10461
rect 16439 10421 16451 10455
rect 16485 10452 16497 10455
rect 16666 10452 16672 10464
rect 16485 10424 16672 10452
rect 16485 10421 16497 10424
rect 16439 10415 16497 10421
rect 16666 10412 16672 10424
rect 16724 10412 16730 10464
rect 16868 10461 16896 10492
rect 18385 10492 18889 10520
rect 16853 10455 16911 10461
rect 16853 10421 16865 10455
rect 16899 10452 16911 10455
rect 17494 10452 17500 10464
rect 16899 10424 17500 10452
rect 16899 10421 16911 10424
rect 16853 10415 16911 10421
rect 17494 10412 17500 10424
rect 17552 10412 17558 10464
rect 18138 10412 18144 10464
rect 18196 10452 18202 10464
rect 18385 10452 18413 10492
rect 18877 10489 18889 10492
rect 18923 10489 18935 10523
rect 18877 10483 18935 10489
rect 19705 10523 19763 10529
rect 19705 10489 19717 10523
rect 19751 10520 19763 10523
rect 19794 10520 19800 10532
rect 19751 10492 19800 10520
rect 19751 10489 19763 10492
rect 19705 10483 19763 10489
rect 19794 10480 19800 10492
rect 19852 10480 19858 10532
rect 18196 10424 18413 10452
rect 18196 10412 18202 10424
rect 1104 10362 22816 10384
rect 1104 10310 8982 10362
rect 9034 10310 9046 10362
rect 9098 10310 9110 10362
rect 9162 10310 9174 10362
rect 9226 10310 16982 10362
rect 17034 10310 17046 10362
rect 17098 10310 17110 10362
rect 17162 10310 17174 10362
rect 17226 10310 22816 10362
rect 1104 10288 22816 10310
rect 1857 10251 1915 10257
rect 1857 10217 1869 10251
rect 1903 10248 1915 10251
rect 1946 10248 1952 10260
rect 1903 10220 1952 10248
rect 1903 10217 1915 10220
rect 1857 10211 1915 10217
rect 1946 10208 1952 10220
rect 2004 10208 2010 10260
rect 2222 10208 2228 10260
rect 2280 10248 2286 10260
rect 2409 10251 2467 10257
rect 2409 10248 2421 10251
rect 2280 10220 2421 10248
rect 2280 10208 2286 10220
rect 2409 10217 2421 10220
rect 2455 10248 2467 10251
rect 2685 10251 2743 10257
rect 2685 10248 2697 10251
rect 2455 10220 2697 10248
rect 2455 10217 2467 10220
rect 2409 10211 2467 10217
rect 2685 10217 2697 10220
rect 2731 10217 2743 10251
rect 4430 10248 4436 10260
rect 4391 10220 4436 10248
rect 2685 10211 2743 10217
rect 4430 10208 4436 10220
rect 4488 10208 4494 10260
rect 4798 10208 4804 10260
rect 4856 10248 4862 10260
rect 5261 10251 5319 10257
rect 5261 10248 5273 10251
rect 4856 10220 5273 10248
rect 4856 10208 4862 10220
rect 5261 10217 5273 10220
rect 5307 10217 5319 10251
rect 5261 10211 5319 10217
rect 7653 10251 7711 10257
rect 7653 10217 7665 10251
rect 7699 10248 7711 10251
rect 7742 10248 7748 10260
rect 7699 10220 7748 10248
rect 7699 10217 7711 10220
rect 7653 10211 7711 10217
rect 7742 10208 7748 10220
rect 7800 10208 7806 10260
rect 13538 10208 13544 10260
rect 13596 10248 13602 10260
rect 15746 10248 15752 10260
rect 13596 10220 13860 10248
rect 15707 10220 15752 10248
rect 13596 10208 13602 10220
rect 4448 10180 4476 10208
rect 7098 10189 7104 10192
rect 7054 10183 7104 10189
rect 7054 10180 7066 10183
rect 4448 10152 7066 10180
rect 7054 10149 7066 10152
rect 7100 10149 7104 10183
rect 7054 10143 7104 10149
rect 7098 10140 7104 10143
rect 7156 10140 7162 10192
rect 7190 10140 7196 10192
rect 7248 10180 7254 10192
rect 7929 10183 7987 10189
rect 7929 10180 7941 10183
rect 7248 10152 7941 10180
rect 7248 10140 7254 10152
rect 7929 10149 7941 10152
rect 7975 10180 7987 10183
rect 8754 10180 8760 10192
rect 7975 10152 8760 10180
rect 7975 10149 7987 10152
rect 7929 10143 7987 10149
rect 8754 10140 8760 10152
rect 8812 10140 8818 10192
rect 9766 10140 9772 10192
rect 9824 10180 9830 10192
rect 10366 10183 10424 10189
rect 10366 10180 10378 10183
rect 9824 10152 10378 10180
rect 9824 10140 9830 10152
rect 10366 10149 10378 10152
rect 10412 10149 10424 10183
rect 10366 10143 10424 10149
rect 11698 10140 11704 10192
rect 11756 10180 11762 10192
rect 12161 10183 12219 10189
rect 12161 10180 12173 10183
rect 11756 10152 12173 10180
rect 11756 10140 11762 10152
rect 12161 10149 12173 10152
rect 12207 10149 12219 10183
rect 12161 10143 12219 10149
rect 12250 10140 12256 10192
rect 12308 10180 12314 10192
rect 13722 10180 13728 10192
rect 12308 10152 12353 10180
rect 13683 10152 13728 10180
rect 12308 10140 12314 10152
rect 13722 10140 13728 10152
rect 13780 10140 13786 10192
rect 13832 10189 13860 10220
rect 15746 10208 15752 10220
rect 15804 10208 15810 10260
rect 19610 10208 19616 10260
rect 19668 10248 19674 10260
rect 19889 10251 19947 10257
rect 19889 10248 19901 10251
rect 19668 10220 19901 10248
rect 19668 10208 19674 10220
rect 19889 10217 19901 10220
rect 19935 10217 19947 10251
rect 19889 10211 19947 10217
rect 13817 10183 13875 10189
rect 13817 10149 13829 10183
rect 13863 10149 13875 10183
rect 17310 10180 17316 10192
rect 17271 10152 17316 10180
rect 13817 10143 13875 10149
rect 17310 10140 17316 10152
rect 17368 10140 17374 10192
rect 18874 10140 18880 10192
rect 18932 10180 18938 10192
rect 19014 10183 19072 10189
rect 19014 10180 19026 10183
rect 18932 10152 19026 10180
rect 18932 10140 18938 10152
rect 19014 10149 19026 10152
rect 19060 10149 19072 10183
rect 19014 10143 19072 10149
rect 3142 10072 3148 10124
rect 3200 10112 3206 10124
rect 3694 10112 3700 10124
rect 3200 10084 3700 10112
rect 3200 10072 3206 10084
rect 3694 10072 3700 10084
rect 3752 10112 3758 10124
rect 4065 10115 4123 10121
rect 4065 10112 4077 10115
rect 3752 10084 4077 10112
rect 3752 10072 3758 10084
rect 4065 10081 4077 10084
rect 4111 10081 4123 10115
rect 4065 10075 4123 10081
rect 6733 10115 6791 10121
rect 6733 10081 6745 10115
rect 6779 10112 6791 10115
rect 6914 10112 6920 10124
rect 6779 10084 6920 10112
rect 6779 10081 6791 10084
rect 6733 10075 6791 10081
rect 6914 10072 6920 10084
rect 6972 10072 6978 10124
rect 8478 10072 8484 10124
rect 8536 10112 8542 10124
rect 8624 10115 8682 10121
rect 8624 10112 8636 10115
rect 8536 10084 8636 10112
rect 8536 10072 8542 10084
rect 8624 10081 8636 10084
rect 8670 10112 8682 10115
rect 8846 10112 8852 10124
rect 8670 10084 8852 10112
rect 8670 10081 8682 10084
rect 8624 10075 8682 10081
rect 8846 10072 8852 10084
rect 8904 10072 8910 10124
rect 10042 10112 10048 10124
rect 10003 10084 10048 10112
rect 10042 10072 10048 10084
rect 10100 10072 10106 10124
rect 19613 10115 19671 10121
rect 19613 10081 19625 10115
rect 19659 10112 19671 10115
rect 19794 10112 19800 10124
rect 19659 10084 19800 10112
rect 19659 10081 19671 10084
rect 19613 10075 19671 10081
rect 19794 10072 19800 10084
rect 19852 10072 19858 10124
rect 20714 10072 20720 10124
rect 20772 10112 20778 10124
rect 20936 10115 20994 10121
rect 20936 10112 20948 10115
rect 20772 10084 20948 10112
rect 20772 10072 20778 10084
rect 20936 10081 20948 10084
rect 20982 10081 20994 10115
rect 20936 10075 20994 10081
rect 1486 10044 1492 10056
rect 1447 10016 1492 10044
rect 1486 10004 1492 10016
rect 1544 10004 1550 10056
rect 8711 10047 8769 10053
rect 8711 10013 8723 10047
rect 8757 10044 8769 10047
rect 12342 10044 12348 10056
rect 8757 10016 12348 10044
rect 8757 10013 8769 10016
rect 8711 10007 8769 10013
rect 12342 10004 12348 10016
rect 12400 10004 12406 10056
rect 12526 10004 12532 10056
rect 12584 10044 12590 10056
rect 12805 10047 12863 10053
rect 12805 10044 12817 10047
rect 12584 10016 12817 10044
rect 12584 10004 12590 10016
rect 12805 10013 12817 10016
rect 12851 10044 12863 10047
rect 13906 10044 13912 10056
rect 12851 10016 13912 10044
rect 12851 10013 12863 10016
rect 12805 10007 12863 10013
rect 13906 10004 13912 10016
rect 13964 10044 13970 10056
rect 14001 10047 14059 10053
rect 14001 10044 14013 10047
rect 13964 10016 14013 10044
rect 13964 10004 13970 10016
rect 14001 10013 14013 10016
rect 14047 10013 14059 10047
rect 15378 10044 15384 10056
rect 15339 10016 15384 10044
rect 14001 10007 14059 10013
rect 15378 10004 15384 10016
rect 15436 10004 15442 10056
rect 16666 10004 16672 10056
rect 16724 10044 16730 10056
rect 17221 10047 17279 10053
rect 17221 10044 17233 10047
rect 16724 10016 17233 10044
rect 16724 10004 16730 10016
rect 17221 10013 17233 10016
rect 17267 10044 17279 10047
rect 17586 10044 17592 10056
rect 17267 10016 17592 10044
rect 17267 10013 17279 10016
rect 17221 10007 17279 10013
rect 17586 10004 17592 10016
rect 17644 10004 17650 10056
rect 18693 10047 18751 10053
rect 18693 10013 18705 10047
rect 18739 10044 18751 10047
rect 18782 10044 18788 10056
rect 18739 10016 18788 10044
rect 18739 10013 18751 10016
rect 18693 10007 18751 10013
rect 18782 10004 18788 10016
rect 18840 10004 18846 10056
rect 13170 9976 13176 9988
rect 9324 9948 13176 9976
rect 9324 9920 9352 9948
rect 13170 9936 13176 9948
rect 13228 9976 13234 9988
rect 13449 9979 13507 9985
rect 13449 9976 13461 9979
rect 13228 9948 13461 9976
rect 13228 9936 13234 9948
rect 13449 9945 13461 9948
rect 13495 9945 13507 9979
rect 17770 9976 17776 9988
rect 17731 9948 17776 9976
rect 13449 9939 13507 9945
rect 17770 9936 17776 9948
rect 17828 9936 17834 9988
rect 4062 9868 4068 9920
rect 4120 9908 4126 9920
rect 4985 9911 5043 9917
rect 4985 9908 4997 9911
rect 4120 9880 4997 9908
rect 4120 9868 4126 9880
rect 4985 9877 4997 9880
rect 5031 9877 5043 9911
rect 4985 9871 5043 9877
rect 5534 9868 5540 9920
rect 5592 9908 5598 9920
rect 9306 9908 9312 9920
rect 5592 9880 9312 9908
rect 5592 9868 5598 9880
rect 9306 9868 9312 9880
rect 9364 9868 9370 9920
rect 9766 9868 9772 9920
rect 9824 9908 9830 9920
rect 9861 9911 9919 9917
rect 9861 9908 9873 9911
rect 9824 9880 9873 9908
rect 9824 9868 9830 9880
rect 9861 9877 9873 9880
rect 9907 9877 9919 9911
rect 10962 9908 10968 9920
rect 10923 9880 10968 9908
rect 9861 9871 9919 9877
rect 10962 9868 10968 9880
rect 11020 9868 11026 9920
rect 16298 9908 16304 9920
rect 16259 9880 16304 9908
rect 16298 9868 16304 9880
rect 16356 9868 16362 9920
rect 18138 9908 18144 9920
rect 18099 9880 18144 9908
rect 18138 9868 18144 9880
rect 18196 9868 18202 9920
rect 20254 9868 20260 9920
rect 20312 9908 20318 9920
rect 21039 9911 21097 9917
rect 21039 9908 21051 9911
rect 20312 9880 21051 9908
rect 20312 9868 20318 9880
rect 21039 9877 21051 9880
rect 21085 9877 21097 9911
rect 21039 9871 21097 9877
rect 1104 9818 22816 9840
rect 1104 9766 4982 9818
rect 5034 9766 5046 9818
rect 5098 9766 5110 9818
rect 5162 9766 5174 9818
rect 5226 9766 12982 9818
rect 13034 9766 13046 9818
rect 13098 9766 13110 9818
rect 13162 9766 13174 9818
rect 13226 9766 20982 9818
rect 21034 9766 21046 9818
rect 21098 9766 21110 9818
rect 21162 9766 21174 9818
rect 21226 9766 22816 9818
rect 1104 9744 22816 9766
rect 1946 9664 1952 9716
rect 2004 9704 2010 9716
rect 2593 9707 2651 9713
rect 2593 9704 2605 9707
rect 2004 9676 2605 9704
rect 2004 9664 2010 9676
rect 2593 9673 2605 9676
rect 2639 9673 2651 9707
rect 3694 9704 3700 9716
rect 3655 9676 3700 9704
rect 2593 9667 2651 9673
rect 3694 9664 3700 9676
rect 3752 9664 3758 9716
rect 4157 9707 4215 9713
rect 4157 9673 4169 9707
rect 4203 9704 4215 9707
rect 4430 9704 4436 9716
rect 4203 9676 4436 9704
rect 4203 9673 4215 9676
rect 4157 9667 4215 9673
rect 4430 9664 4436 9676
rect 4488 9664 4494 9716
rect 5350 9664 5356 9716
rect 5408 9704 5414 9716
rect 5445 9707 5503 9713
rect 5445 9704 5457 9707
rect 5408 9676 5457 9704
rect 5408 9664 5414 9676
rect 5445 9673 5457 9676
rect 5491 9704 5503 9707
rect 8018 9704 8024 9716
rect 5491 9676 8024 9704
rect 5491 9673 5503 9676
rect 5445 9667 5503 9673
rect 8018 9664 8024 9676
rect 8076 9664 8082 9716
rect 10962 9664 10968 9716
rect 11020 9704 11026 9716
rect 11701 9707 11759 9713
rect 11701 9704 11713 9707
rect 11020 9676 11713 9704
rect 11020 9664 11026 9676
rect 11701 9673 11713 9676
rect 11747 9704 11759 9707
rect 12069 9707 12127 9713
rect 12069 9704 12081 9707
rect 11747 9676 12081 9704
rect 11747 9673 11759 9676
rect 11701 9667 11759 9673
rect 12069 9673 12081 9676
rect 12115 9704 12127 9707
rect 12250 9704 12256 9716
rect 12115 9676 12256 9704
rect 12115 9673 12127 9676
rect 12069 9667 12127 9673
rect 12250 9664 12256 9676
rect 12308 9664 12314 9716
rect 13814 9664 13820 9716
rect 13872 9704 13878 9716
rect 14366 9704 14372 9716
rect 13872 9676 14372 9704
rect 13872 9664 13878 9676
rect 14366 9664 14372 9676
rect 14424 9664 14430 9716
rect 15378 9664 15384 9716
rect 15436 9704 15442 9716
rect 15841 9707 15899 9713
rect 15841 9704 15853 9707
rect 15436 9676 15853 9704
rect 15436 9664 15442 9676
rect 15841 9673 15853 9676
rect 15887 9673 15899 9707
rect 16298 9704 16304 9716
rect 16211 9676 16304 9704
rect 15841 9667 15899 9673
rect 16298 9664 16304 9676
rect 16356 9704 16362 9716
rect 17310 9704 17316 9716
rect 16356 9676 17316 9704
rect 16356 9664 16362 9676
rect 17310 9664 17316 9676
rect 17368 9704 17374 9716
rect 17405 9707 17463 9713
rect 17405 9704 17417 9707
rect 17368 9676 17417 9704
rect 17368 9664 17374 9676
rect 17405 9673 17417 9676
rect 17451 9673 17463 9707
rect 17405 9667 17463 9673
rect 18874 9664 18880 9716
rect 18932 9704 18938 9716
rect 19061 9707 19119 9713
rect 19061 9704 19073 9707
rect 18932 9676 19073 9704
rect 18932 9664 18938 9676
rect 19061 9673 19073 9676
rect 19107 9673 19119 9707
rect 19061 9667 19119 9673
rect 19521 9707 19579 9713
rect 19521 9673 19533 9707
rect 19567 9704 19579 9707
rect 19794 9704 19800 9716
rect 19567 9676 19800 9704
rect 19567 9673 19579 9676
rect 19521 9667 19579 9673
rect 19794 9664 19800 9676
rect 19852 9664 19858 9716
rect 20714 9664 20720 9716
rect 20772 9704 20778 9716
rect 20901 9707 20959 9713
rect 20901 9704 20913 9707
rect 20772 9676 20913 9704
rect 20772 9664 20778 9676
rect 20901 9673 20913 9676
rect 20947 9673 20959 9707
rect 20901 9667 20959 9673
rect 5368 9636 5396 9664
rect 7098 9636 7104 9648
rect 4448 9608 5396 9636
rect 7059 9608 7104 9636
rect 1486 9528 1492 9580
rect 1544 9568 1550 9580
rect 4448 9577 4476 9608
rect 7098 9596 7104 9608
rect 7156 9596 7162 9648
rect 10781 9639 10839 9645
rect 10781 9605 10793 9639
rect 10827 9636 10839 9639
rect 12158 9636 12164 9648
rect 10827 9608 12164 9636
rect 10827 9605 10839 9608
rect 10781 9599 10839 9605
rect 12158 9596 12164 9608
rect 12216 9636 12222 9648
rect 13538 9636 13544 9648
rect 12216 9608 13544 9636
rect 12216 9596 12222 9608
rect 13538 9596 13544 9608
rect 13596 9636 13602 9648
rect 13633 9639 13691 9645
rect 13633 9636 13645 9639
rect 13596 9608 13645 9636
rect 13596 9596 13602 9608
rect 13633 9605 13645 9608
rect 13679 9605 13691 9639
rect 13633 9599 13691 9605
rect 13998 9596 14004 9648
rect 14056 9636 14062 9648
rect 18138 9636 18144 9648
rect 14056 9608 18144 9636
rect 14056 9596 14062 9608
rect 2317 9571 2375 9577
rect 2317 9568 2329 9571
rect 1544 9540 2329 9568
rect 1544 9528 1550 9540
rect 2317 9537 2329 9540
rect 2363 9568 2375 9571
rect 3329 9571 3387 9577
rect 3329 9568 3341 9571
rect 2363 9540 3341 9568
rect 2363 9537 2375 9540
rect 2317 9531 2375 9537
rect 3329 9537 3341 9540
rect 3375 9537 3387 9571
rect 3329 9531 3387 9537
rect 4433 9571 4491 9577
rect 4433 9537 4445 9571
rect 4479 9537 4491 9571
rect 4433 9531 4491 9537
rect 5077 9571 5135 9577
rect 5077 9537 5089 9571
rect 5123 9568 5135 9571
rect 5442 9568 5448 9580
rect 5123 9540 5448 9568
rect 5123 9537 5135 9540
rect 5077 9531 5135 9537
rect 5442 9528 5448 9540
rect 5500 9528 5506 9580
rect 7377 9571 7435 9577
rect 7377 9537 7389 9571
rect 7423 9568 7435 9571
rect 7834 9568 7840 9580
rect 7423 9540 7840 9568
rect 7423 9537 7435 9540
rect 7377 9531 7435 9537
rect 7834 9528 7840 9540
rect 7892 9528 7898 9580
rect 8754 9528 8760 9580
rect 8812 9568 8818 9580
rect 8987 9571 9045 9577
rect 8987 9568 8999 9571
rect 8812 9540 8999 9568
rect 8812 9528 8818 9540
rect 8987 9537 8999 9540
rect 9033 9537 9045 9571
rect 12802 9568 12808 9580
rect 12763 9540 12808 9568
rect 8987 9531 9045 9537
rect 12802 9528 12808 9540
rect 12860 9528 12866 9580
rect 13446 9528 13452 9580
rect 13504 9568 13510 9580
rect 13722 9568 13728 9580
rect 13504 9540 13728 9568
rect 13504 9528 13510 9540
rect 13722 9528 13728 9540
rect 13780 9568 13786 9580
rect 16485 9571 16543 9577
rect 13780 9540 14964 9568
rect 13780 9528 13786 9540
rect 1670 9500 1676 9512
rect 1631 9472 1676 9500
rect 1670 9460 1676 9472
rect 1728 9460 1734 9512
rect 2133 9503 2191 9509
rect 2133 9469 2145 9503
rect 2179 9500 2191 9503
rect 2866 9500 2872 9512
rect 2179 9472 2872 9500
rect 2179 9469 2191 9472
rect 2133 9463 2191 9469
rect 2866 9460 2872 9472
rect 2924 9460 2930 9512
rect 8386 9460 8392 9512
rect 8444 9500 8450 9512
rect 8900 9503 8958 9509
rect 8900 9500 8912 9503
rect 8444 9472 8912 9500
rect 8444 9460 8450 9472
rect 8900 9469 8912 9472
rect 8946 9500 8958 9503
rect 9861 9503 9919 9509
rect 8946 9472 9444 9500
rect 8946 9469 8958 9472
rect 8900 9463 8958 9469
rect 1688 9432 1716 9460
rect 9416 9444 9444 9472
rect 9861 9469 9873 9503
rect 9907 9500 9919 9503
rect 9950 9500 9956 9512
rect 9907 9472 9956 9500
rect 9907 9469 9919 9472
rect 9861 9463 9919 9469
rect 9950 9460 9956 9472
rect 10008 9500 10014 9512
rect 11057 9503 11115 9509
rect 11057 9500 11069 9503
rect 10008 9472 11069 9500
rect 10008 9460 10014 9472
rect 11057 9469 11069 9472
rect 11103 9469 11115 9503
rect 14458 9500 14464 9512
rect 14419 9472 14464 9500
rect 11057 9463 11115 9469
rect 14458 9460 14464 9472
rect 14516 9460 14522 9512
rect 14936 9509 14964 9540
rect 16485 9537 16497 9571
rect 16531 9568 16543 9571
rect 16574 9568 16580 9580
rect 16531 9540 16580 9568
rect 16531 9537 16543 9540
rect 16485 9531 16543 9537
rect 16574 9528 16580 9540
rect 16632 9528 16638 9580
rect 18064 9509 18092 9608
rect 18138 9596 18144 9608
rect 18196 9596 18202 9648
rect 21358 9636 21364 9648
rect 21319 9608 21364 9636
rect 21358 9596 21364 9608
rect 21416 9596 21422 9648
rect 19705 9571 19763 9577
rect 19705 9537 19717 9571
rect 19751 9568 19763 9571
rect 20162 9568 20168 9580
rect 19751 9540 20168 9568
rect 19751 9537 19763 9540
rect 19705 9531 19763 9537
rect 20162 9528 20168 9540
rect 20220 9528 20226 9580
rect 20346 9528 20352 9580
rect 20404 9568 20410 9580
rect 21729 9571 21787 9577
rect 21729 9568 21741 9571
rect 20404 9540 21741 9568
rect 20404 9528 20410 9540
rect 21192 9509 21220 9540
rect 21729 9537 21741 9540
rect 21775 9537 21787 9571
rect 21729 9531 21787 9537
rect 14921 9503 14979 9509
rect 14921 9469 14933 9503
rect 14967 9500 14979 9503
rect 18049 9503 18107 9509
rect 14967 9472 16252 9500
rect 14967 9469 14979 9472
rect 14921 9463 14979 9469
rect 2958 9432 2964 9444
rect 1688 9404 2964 9432
rect 2958 9392 2964 9404
rect 3016 9392 3022 9444
rect 4525 9435 4583 9441
rect 4126 9404 4292 9432
rect 4126 9376 4154 9404
rect 4062 9324 4068 9376
rect 4120 9336 4154 9376
rect 4264 9364 4292 9404
rect 4525 9401 4537 9435
rect 4571 9401 4583 9435
rect 4525 9395 4583 9401
rect 6641 9435 6699 9441
rect 6641 9401 6653 9435
rect 6687 9432 6699 9435
rect 7469 9435 7527 9441
rect 7469 9432 7481 9435
rect 6687 9404 7481 9432
rect 6687 9401 6699 9404
rect 6641 9395 6699 9401
rect 7469 9401 7481 9404
rect 7515 9432 7527 9435
rect 7742 9432 7748 9444
rect 7515 9404 7748 9432
rect 7515 9401 7527 9404
rect 7469 9395 7527 9401
rect 4540 9364 4568 9395
rect 7742 9392 7748 9404
rect 7800 9392 7806 9444
rect 8018 9432 8024 9444
rect 7979 9404 8024 9432
rect 8018 9392 8024 9404
rect 8076 9392 8082 9444
rect 9398 9432 9404 9444
rect 9359 9404 9404 9432
rect 9398 9392 9404 9404
rect 9456 9392 9462 9444
rect 9766 9432 9772 9444
rect 9679 9404 9772 9432
rect 9766 9392 9772 9404
rect 9824 9432 9830 9444
rect 10223 9435 10281 9441
rect 10223 9432 10235 9435
rect 9824 9404 10235 9432
rect 9824 9392 9830 9404
rect 10223 9401 10235 9404
rect 10269 9432 10281 9435
rect 11146 9432 11152 9444
rect 10269 9404 11152 9432
rect 10269 9401 10281 9404
rect 10223 9395 10281 9401
rect 11146 9392 11152 9404
rect 11204 9392 11210 9444
rect 12526 9432 12532 9444
rect 12487 9404 12532 9432
rect 12526 9392 12532 9404
rect 12584 9392 12590 9444
rect 12621 9435 12679 9441
rect 12621 9401 12633 9435
rect 12667 9401 12679 9435
rect 15194 9432 15200 9444
rect 15155 9404 15200 9432
rect 12621 9395 12679 9401
rect 4264 9336 4568 9364
rect 8665 9367 8723 9373
rect 4120 9324 4126 9336
rect 8665 9333 8677 9367
rect 8711 9364 8723 9367
rect 8754 9364 8760 9376
rect 8711 9336 8760 9364
rect 8711 9333 8723 9336
rect 8665 9327 8723 9333
rect 8754 9324 8760 9336
rect 8812 9324 8818 9376
rect 12250 9324 12256 9376
rect 12308 9364 12314 9376
rect 12636 9364 12664 9395
rect 15194 9392 15200 9404
rect 15252 9392 15258 9444
rect 12308 9336 12664 9364
rect 15565 9367 15623 9373
rect 12308 9324 12314 9336
rect 15565 9333 15577 9367
rect 15611 9364 15623 9367
rect 15838 9364 15844 9376
rect 15611 9336 15844 9364
rect 15611 9333 15623 9336
rect 15565 9327 15623 9333
rect 15838 9324 15844 9336
rect 15896 9324 15902 9376
rect 16224 9364 16252 9472
rect 18049 9469 18061 9503
rect 18095 9469 18107 9503
rect 18049 9463 18107 9469
rect 18509 9503 18567 9509
rect 18509 9469 18521 9503
rect 18555 9469 18567 9503
rect 18509 9463 18567 9469
rect 21177 9503 21235 9509
rect 21177 9469 21189 9503
rect 21223 9469 21235 9503
rect 21177 9463 21235 9469
rect 16298 9392 16304 9444
rect 16356 9432 16362 9444
rect 16577 9435 16635 9441
rect 16577 9432 16589 9435
rect 16356 9404 16589 9432
rect 16356 9392 16362 9404
rect 16577 9401 16589 9404
rect 16623 9401 16635 9435
rect 16577 9395 16635 9401
rect 17129 9435 17187 9441
rect 17129 9401 17141 9435
rect 17175 9432 17187 9435
rect 17310 9432 17316 9444
rect 17175 9404 17316 9432
rect 17175 9401 17187 9404
rect 17129 9395 17187 9401
rect 17310 9392 17316 9404
rect 17368 9392 17374 9444
rect 18524 9432 18552 9463
rect 18598 9432 18604 9444
rect 17788 9404 18604 9432
rect 17788 9373 17816 9404
rect 18598 9392 18604 9404
rect 18656 9392 18662 9444
rect 18782 9432 18788 9444
rect 18743 9404 18788 9432
rect 18782 9392 18788 9404
rect 18840 9392 18846 9444
rect 19794 9392 19800 9444
rect 19852 9432 19858 9444
rect 20349 9435 20407 9441
rect 19852 9404 19897 9432
rect 19852 9392 19858 9404
rect 20349 9401 20361 9435
rect 20395 9432 20407 9435
rect 20438 9432 20444 9444
rect 20395 9404 20444 9432
rect 20395 9401 20407 9404
rect 20349 9395 20407 9401
rect 20438 9392 20444 9404
rect 20496 9392 20502 9444
rect 17773 9367 17831 9373
rect 17773 9364 17785 9367
rect 16224 9336 17785 9364
rect 17773 9333 17785 9336
rect 17819 9333 17831 9367
rect 17773 9327 17831 9333
rect 1104 9274 22816 9296
rect 1104 9222 8982 9274
rect 9034 9222 9046 9274
rect 9098 9222 9110 9274
rect 9162 9222 9174 9274
rect 9226 9222 16982 9274
rect 17034 9222 17046 9274
rect 17098 9222 17110 9274
rect 17162 9222 17174 9274
rect 17226 9222 22816 9274
rect 1104 9200 22816 9222
rect 3786 9160 3792 9172
rect 2700 9132 3792 9160
rect 1854 9092 1860 9104
rect 1479 9064 1860 9092
rect 14 8984 20 9036
rect 72 9024 78 9036
rect 1479 9033 1507 9064
rect 1854 9052 1860 9064
rect 1912 9052 1918 9104
rect 2700 9036 2728 9132
rect 3786 9120 3792 9132
rect 3844 9120 3850 9172
rect 4062 9120 4068 9172
rect 4120 9160 4126 9172
rect 4341 9163 4399 9169
rect 4341 9160 4353 9163
rect 4120 9132 4353 9160
rect 4120 9120 4126 9132
rect 4341 9129 4353 9132
rect 4387 9129 4399 9163
rect 4341 9123 4399 9129
rect 6825 9163 6883 9169
rect 6825 9129 6837 9163
rect 6871 9160 6883 9163
rect 6914 9160 6920 9172
rect 6871 9132 6920 9160
rect 6871 9129 6883 9132
rect 6825 9123 6883 9129
rect 6914 9120 6920 9132
rect 6972 9120 6978 9172
rect 7926 9120 7932 9172
rect 7984 9160 7990 9172
rect 8021 9163 8079 9169
rect 8021 9160 8033 9163
rect 7984 9132 8033 9160
rect 7984 9120 7990 9132
rect 8021 9129 8033 9132
rect 8067 9129 8079 9163
rect 9950 9160 9956 9172
rect 9911 9132 9956 9160
rect 8021 9123 8079 9129
rect 9950 9120 9956 9132
rect 10008 9120 10014 9172
rect 11698 9120 11704 9172
rect 11756 9160 11762 9172
rect 11885 9163 11943 9169
rect 11885 9160 11897 9163
rect 11756 9132 11897 9160
rect 11756 9120 11762 9132
rect 11885 9129 11897 9132
rect 11931 9129 11943 9163
rect 11885 9123 11943 9129
rect 12526 9120 12532 9172
rect 12584 9160 12590 9172
rect 13081 9163 13139 9169
rect 13081 9160 13093 9163
rect 12584 9132 13093 9160
rect 12584 9120 12590 9132
rect 13081 9129 13093 9132
rect 13127 9129 13139 9163
rect 13081 9123 13139 9129
rect 3145 9095 3203 9101
rect 3145 9061 3157 9095
rect 3191 9092 3203 9095
rect 3602 9092 3608 9104
rect 3191 9064 3608 9092
rect 3191 9061 3203 9064
rect 3145 9055 3203 9061
rect 3602 9052 3608 9064
rect 3660 9052 3666 9104
rect 4706 9092 4712 9104
rect 4667 9064 4712 9092
rect 4706 9052 4712 9064
rect 4764 9052 4770 9104
rect 7193 9095 7251 9101
rect 7193 9061 7205 9095
rect 7239 9092 7251 9095
rect 7374 9092 7380 9104
rect 7239 9064 7380 9092
rect 7239 9061 7251 9064
rect 7193 9055 7251 9061
rect 7374 9052 7380 9064
rect 7432 9052 7438 9104
rect 9493 9095 9551 9101
rect 9493 9061 9505 9095
rect 9539 9092 9551 9095
rect 10042 9092 10048 9104
rect 9539 9064 10048 9092
rect 9539 9061 9551 9064
rect 9493 9055 9551 9061
rect 10042 9052 10048 9064
rect 10100 9052 10106 9104
rect 12250 9092 12256 9104
rect 12211 9064 12256 9092
rect 12250 9052 12256 9064
rect 12308 9052 12314 9104
rect 12802 9092 12808 9104
rect 12763 9064 12808 9092
rect 12802 9052 12808 9064
rect 12860 9052 12866 9104
rect 13096 9092 13124 9123
rect 13630 9120 13636 9172
rect 13688 9160 13694 9172
rect 14093 9163 14151 9169
rect 14093 9160 14105 9163
rect 13688 9132 14105 9160
rect 13688 9120 13694 9132
rect 14093 9129 14105 9132
rect 14139 9129 14151 9163
rect 14458 9160 14464 9172
rect 14419 9132 14464 9160
rect 14093 9123 14151 9129
rect 14458 9120 14464 9132
rect 14516 9120 14522 9172
rect 16485 9163 16543 9169
rect 16485 9129 16497 9163
rect 16531 9160 16543 9163
rect 16574 9160 16580 9172
rect 16531 9132 16580 9160
rect 16531 9129 16543 9132
rect 16485 9123 16543 9129
rect 16574 9120 16580 9132
rect 16632 9120 16638 9172
rect 17586 9160 17592 9172
rect 17547 9132 17592 9160
rect 17586 9120 17592 9132
rect 17644 9120 17650 9172
rect 18782 9120 18788 9172
rect 18840 9160 18846 9172
rect 19153 9163 19211 9169
rect 19153 9160 19165 9163
rect 18840 9132 19165 9160
rect 18840 9120 18846 9132
rect 19153 9129 19165 9132
rect 19199 9129 19211 9163
rect 19153 9123 19211 9129
rect 19978 9120 19984 9172
rect 20036 9160 20042 9172
rect 20073 9163 20131 9169
rect 20073 9160 20085 9163
rect 20036 9132 20085 9160
rect 20036 9120 20042 9132
rect 20073 9129 20085 9132
rect 20119 9129 20131 9163
rect 20254 9160 20260 9172
rect 20215 9132 20260 9160
rect 20073 9123 20131 9129
rect 20254 9120 20260 9132
rect 20312 9120 20318 9172
rect 13771 9095 13829 9101
rect 13771 9092 13783 9095
rect 13096 9064 13783 9092
rect 13771 9061 13783 9064
rect 13817 9061 13829 9095
rect 16758 9092 16764 9104
rect 16719 9064 16764 9092
rect 13771 9055 13829 9061
rect 16758 9052 16764 9064
rect 16816 9052 16822 9104
rect 20346 9052 20352 9104
rect 20404 9092 20410 9104
rect 21085 9095 21143 9101
rect 21085 9092 21097 9095
rect 20404 9064 21097 9092
rect 20404 9052 20410 9064
rect 21085 9061 21097 9064
rect 21131 9061 21143 9095
rect 21085 9055 21143 9061
rect 1432 9027 1507 9033
rect 1432 9024 1444 9027
rect 72 8996 1444 9024
rect 72 8984 78 8996
rect 1432 8993 1444 8996
rect 1478 8996 1507 9027
rect 1535 9027 1593 9033
rect 1478 8993 1490 8996
rect 1432 8987 1490 8993
rect 1535 8993 1547 9027
rect 1581 8993 1593 9027
rect 2682 9024 2688 9036
rect 2595 8996 2688 9024
rect 1535 8987 1593 8993
rect 1550 8900 1578 8987
rect 2682 8984 2688 8996
rect 2740 8984 2746 9036
rect 2866 9024 2872 9036
rect 2827 8996 2872 9024
rect 2866 8984 2872 8996
rect 2924 8984 2930 9036
rect 9953 9027 10011 9033
rect 9953 8993 9965 9027
rect 9999 8993 10011 9027
rect 10226 9024 10232 9036
rect 10187 8996 10232 9024
rect 9953 8987 10011 8993
rect 2317 8959 2375 8965
rect 2317 8925 2329 8959
rect 2363 8956 2375 8959
rect 2498 8956 2504 8968
rect 2363 8928 2504 8956
rect 2363 8925 2375 8928
rect 2317 8919 2375 8925
rect 2498 8916 2504 8928
rect 2556 8956 2562 8968
rect 2884 8956 2912 8984
rect 2556 8928 2912 8956
rect 4617 8959 4675 8965
rect 2556 8916 2562 8928
rect 4617 8925 4629 8959
rect 4663 8956 4675 8959
rect 4798 8956 4804 8968
rect 4663 8928 4804 8956
rect 4663 8925 4675 8928
rect 4617 8919 4675 8925
rect 4798 8916 4804 8928
rect 4856 8916 4862 8968
rect 4890 8916 4896 8968
rect 4948 8956 4954 8968
rect 7098 8956 7104 8968
rect 4948 8928 4993 8956
rect 7059 8928 7104 8956
rect 4948 8916 4954 8928
rect 7098 8916 7104 8928
rect 7156 8916 7162 8968
rect 7377 8959 7435 8965
rect 7377 8925 7389 8959
rect 7423 8956 7435 8959
rect 7466 8956 7472 8968
rect 7423 8928 7472 8956
rect 7423 8925 7435 8928
rect 7377 8919 7435 8925
rect 1486 8848 1492 8900
rect 1544 8860 1578 8900
rect 4908 8888 4936 8916
rect 7392 8888 7420 8919
rect 7466 8916 7472 8928
rect 7524 8916 7530 8968
rect 9968 8956 9996 8987
rect 10226 8984 10232 8996
rect 10284 8984 10290 9036
rect 13538 8984 13544 9036
rect 13596 9024 13602 9036
rect 13633 9027 13691 9033
rect 13633 9024 13645 9027
rect 13596 8996 13645 9024
rect 13596 8984 13602 8996
rect 13633 8993 13645 8996
rect 13679 8993 13691 9027
rect 13633 8987 13691 8993
rect 15470 8984 15476 9036
rect 15528 9024 15534 9036
rect 15600 9027 15658 9033
rect 15600 9024 15612 9027
rect 15528 8996 15612 9024
rect 15528 8984 15534 8996
rect 15600 8993 15612 8996
rect 15646 8993 15658 9027
rect 15600 8987 15658 8993
rect 17402 8984 17408 9036
rect 17460 9024 17466 9036
rect 18138 9024 18144 9036
rect 17460 8996 18144 9024
rect 17460 8984 17466 8996
rect 18138 8984 18144 8996
rect 18196 8984 18202 9036
rect 18598 9024 18604 9036
rect 18559 8996 18604 9024
rect 18598 8984 18604 8996
rect 18656 8984 18662 9036
rect 19864 9027 19922 9033
rect 19864 8993 19876 9027
rect 19910 9024 19922 9027
rect 20162 9024 20168 9036
rect 19910 8996 20168 9024
rect 19910 8993 19922 8996
rect 19864 8987 19922 8993
rect 20162 8984 20168 8996
rect 20220 8984 20226 9036
rect 11330 8956 11336 8968
rect 9968 8928 11336 8956
rect 11330 8916 11336 8928
rect 11388 8916 11394 8968
rect 12161 8959 12219 8965
rect 12161 8925 12173 8959
rect 12207 8956 12219 8959
rect 12342 8956 12348 8968
rect 12207 8928 12348 8956
rect 12207 8925 12219 8928
rect 12161 8919 12219 8925
rect 12342 8916 12348 8928
rect 12400 8916 12406 8968
rect 15703 8959 15761 8965
rect 15703 8925 15715 8959
rect 15749 8956 15761 8959
rect 16669 8959 16727 8965
rect 16669 8956 16681 8959
rect 15749 8928 16681 8956
rect 15749 8925 15761 8928
rect 15703 8919 15761 8925
rect 16669 8925 16681 8928
rect 16715 8956 16727 8959
rect 16942 8956 16948 8968
rect 16715 8928 16948 8956
rect 16715 8925 16727 8928
rect 16669 8919 16727 8925
rect 16942 8916 16948 8928
rect 17000 8916 17006 8968
rect 18877 8959 18935 8965
rect 18877 8925 18889 8959
rect 18923 8956 18935 8959
rect 19058 8956 19064 8968
rect 18923 8928 19064 8956
rect 18923 8925 18935 8928
rect 18877 8919 18935 8925
rect 19058 8916 19064 8928
rect 19116 8956 19122 8968
rect 19521 8959 19579 8965
rect 19521 8956 19533 8959
rect 19116 8928 19533 8956
rect 19116 8916 19122 8928
rect 19521 8925 19533 8928
rect 19567 8925 19579 8959
rect 19521 8919 19579 8925
rect 20438 8916 20444 8968
rect 20496 8956 20502 8968
rect 20993 8959 21051 8965
rect 20993 8956 21005 8959
rect 20496 8928 21005 8956
rect 20496 8916 20502 8928
rect 20993 8925 21005 8928
rect 21039 8925 21051 8959
rect 21266 8956 21272 8968
rect 21227 8928 21272 8956
rect 20993 8919 21051 8925
rect 4908 8860 7420 8888
rect 1544 8848 1550 8860
rect 15194 8848 15200 8900
rect 15252 8888 15258 8900
rect 16025 8891 16083 8897
rect 16025 8888 16037 8891
rect 15252 8860 16037 8888
rect 15252 8848 15258 8860
rect 16025 8857 16037 8860
rect 16071 8857 16083 8891
rect 16025 8851 16083 8857
rect 17221 8891 17279 8897
rect 17221 8857 17233 8891
rect 17267 8888 17279 8891
rect 17770 8888 17776 8900
rect 17267 8860 17776 8888
rect 17267 8857 17279 8860
rect 17221 8851 17279 8857
rect 17770 8848 17776 8860
rect 17828 8888 17834 8900
rect 20456 8888 20484 8916
rect 17828 8860 20484 8888
rect 21008 8888 21036 8919
rect 21266 8916 21272 8928
rect 21324 8916 21330 8968
rect 22186 8888 22192 8900
rect 21008 8860 22192 8888
rect 17828 8848 17834 8860
rect 22186 8848 22192 8860
rect 22244 8848 22250 8900
rect 5994 8780 6000 8832
rect 6052 8820 6058 8832
rect 10318 8820 10324 8832
rect 6052 8792 10324 8820
rect 6052 8780 6058 8792
rect 10318 8780 10324 8792
rect 10376 8820 10382 8832
rect 10689 8823 10747 8829
rect 10689 8820 10701 8823
rect 10376 8792 10701 8820
rect 10376 8780 10382 8792
rect 10689 8789 10701 8792
rect 10735 8820 10747 8823
rect 14458 8820 14464 8832
rect 10735 8792 14464 8820
rect 10735 8789 10747 8792
rect 10689 8783 10747 8789
rect 14458 8780 14464 8792
rect 14516 8780 14522 8832
rect 1104 8730 22816 8752
rect 1104 8678 4982 8730
rect 5034 8678 5046 8730
rect 5098 8678 5110 8730
rect 5162 8678 5174 8730
rect 5226 8678 12982 8730
rect 13034 8678 13046 8730
rect 13098 8678 13110 8730
rect 13162 8678 13174 8730
rect 13226 8678 20982 8730
rect 21034 8678 21046 8730
rect 21098 8678 21110 8730
rect 21162 8678 21174 8730
rect 21226 8678 22816 8730
rect 1104 8656 22816 8678
rect 2498 8616 2504 8628
rect 2459 8588 2504 8616
rect 2498 8576 2504 8588
rect 2556 8576 2562 8628
rect 2682 8576 2688 8628
rect 2740 8616 2746 8628
rect 2777 8619 2835 8625
rect 2777 8616 2789 8619
rect 2740 8588 2789 8616
rect 2740 8576 2746 8588
rect 2777 8585 2789 8588
rect 2823 8585 2835 8619
rect 2777 8579 2835 8585
rect 6273 8619 6331 8625
rect 6273 8585 6285 8619
rect 6319 8616 6331 8619
rect 7098 8616 7104 8628
rect 6319 8588 7104 8616
rect 6319 8585 6331 8588
rect 6273 8579 6331 8585
rect 7098 8576 7104 8588
rect 7156 8616 7162 8628
rect 9171 8619 9229 8625
rect 9171 8616 9183 8619
rect 7156 8588 9183 8616
rect 7156 8576 7162 8588
rect 9171 8585 9183 8588
rect 9217 8585 9229 8619
rect 9171 8579 9229 8585
rect 10045 8619 10103 8625
rect 10045 8585 10057 8619
rect 10091 8616 10103 8619
rect 10226 8616 10232 8628
rect 10091 8588 10232 8616
rect 10091 8585 10103 8588
rect 10045 8579 10103 8585
rect 5077 8551 5135 8557
rect 5077 8517 5089 8551
rect 5123 8548 5135 8551
rect 5350 8548 5356 8560
rect 5123 8520 5356 8548
rect 5123 8517 5135 8520
rect 5077 8511 5135 8517
rect 5350 8508 5356 8520
rect 5408 8508 5414 8560
rect 6178 8508 6184 8560
rect 6236 8548 6242 8560
rect 6546 8548 6552 8560
rect 6236 8520 6552 8548
rect 6236 8508 6242 8520
rect 6546 8508 6552 8520
rect 6604 8548 6610 8560
rect 8941 8551 8999 8557
rect 6604 8520 8248 8548
rect 6604 8508 6610 8520
rect 3559 8483 3617 8489
rect 3559 8449 3571 8483
rect 3605 8480 3617 8483
rect 4525 8483 4583 8489
rect 4525 8480 4537 8483
rect 3605 8452 4537 8480
rect 3605 8449 3617 8452
rect 3559 8443 3617 8449
rect 4525 8449 4537 8452
rect 4571 8480 4583 8483
rect 5813 8483 5871 8489
rect 5813 8480 5825 8483
rect 4571 8452 5825 8480
rect 4571 8449 4583 8452
rect 4525 8443 4583 8449
rect 5813 8449 5825 8452
rect 5859 8449 5871 8483
rect 8018 8480 8024 8492
rect 7979 8452 8024 8480
rect 5813 8443 5871 8449
rect 8018 8440 8024 8452
rect 8076 8440 8082 8492
rect 1946 8372 1952 8424
rect 2004 8412 2010 8424
rect 2041 8415 2099 8421
rect 2041 8412 2053 8415
rect 2004 8384 2053 8412
rect 2004 8372 2010 8384
rect 2041 8381 2053 8384
rect 2087 8412 2099 8415
rect 3472 8415 3530 8421
rect 2087 8384 3188 8412
rect 2087 8381 2099 8384
rect 2041 8375 2099 8381
rect 3160 8288 3188 8384
rect 3472 8381 3484 8415
rect 3518 8412 3530 8415
rect 8220 8412 8248 8520
rect 8941 8517 8953 8551
rect 8987 8548 8999 8551
rect 10060 8548 10088 8579
rect 10226 8576 10232 8588
rect 10284 8576 10290 8628
rect 11885 8619 11943 8625
rect 11885 8585 11897 8619
rect 11931 8616 11943 8619
rect 12250 8616 12256 8628
rect 11931 8588 12256 8616
rect 11931 8585 11943 8588
rect 11885 8579 11943 8585
rect 12250 8576 12256 8588
rect 12308 8576 12314 8628
rect 16209 8619 16267 8625
rect 16209 8585 16221 8619
rect 16255 8616 16267 8619
rect 16669 8619 16727 8625
rect 16669 8616 16681 8619
rect 16255 8588 16681 8616
rect 16255 8585 16267 8588
rect 16209 8579 16267 8585
rect 16669 8585 16681 8588
rect 16715 8616 16727 8619
rect 16758 8616 16764 8628
rect 16715 8588 16764 8616
rect 16715 8585 16727 8588
rect 16669 8579 16727 8585
rect 16758 8576 16764 8588
rect 16816 8576 16822 8628
rect 16942 8616 16948 8628
rect 16903 8588 16948 8616
rect 16942 8576 16948 8588
rect 17000 8576 17006 8628
rect 17865 8619 17923 8625
rect 17865 8585 17877 8619
rect 17911 8616 17923 8619
rect 18598 8616 18604 8628
rect 17911 8588 18604 8616
rect 17911 8585 17923 8588
rect 17865 8579 17923 8585
rect 18598 8576 18604 8588
rect 18656 8576 18662 8628
rect 19981 8619 20039 8625
rect 19981 8585 19993 8619
rect 20027 8616 20039 8619
rect 20346 8616 20352 8628
rect 20027 8588 20352 8616
rect 20027 8585 20039 8588
rect 19981 8579 20039 8585
rect 20346 8576 20352 8588
rect 20404 8576 20410 8628
rect 22186 8616 22192 8628
rect 22147 8588 22192 8616
rect 22186 8576 22192 8588
rect 22244 8576 22250 8628
rect 8987 8520 10088 8548
rect 8987 8517 8999 8520
rect 8941 8511 8999 8517
rect 10060 8480 10088 8520
rect 20898 8508 20904 8560
rect 20956 8548 20962 8560
rect 21821 8551 21879 8557
rect 21821 8548 21833 8551
rect 20956 8520 21833 8548
rect 20956 8508 20962 8520
rect 21821 8517 21833 8520
rect 21867 8517 21879 8551
rect 21821 8511 21879 8517
rect 12529 8483 12587 8489
rect 10060 8452 10732 8480
rect 9068 8415 9126 8421
rect 9068 8412 9080 8415
rect 3518 8384 4016 8412
rect 8220 8384 9080 8412
rect 3518 8381 3530 8384
rect 3472 8375 3530 8381
rect 3988 8288 4016 8384
rect 9068 8381 9080 8384
rect 9114 8412 9126 8415
rect 9493 8415 9551 8421
rect 9493 8412 9505 8415
rect 9114 8384 9505 8412
rect 9114 8381 9126 8384
rect 9068 8375 9126 8381
rect 9493 8381 9505 8384
rect 9539 8381 9551 8415
rect 10318 8412 10324 8424
rect 10279 8384 10324 8412
rect 9493 8375 9551 8381
rect 10318 8372 10324 8384
rect 10376 8372 10382 8424
rect 10704 8421 10732 8452
rect 12529 8449 12541 8483
rect 12575 8480 12587 8483
rect 12618 8480 12624 8492
rect 12575 8452 12624 8480
rect 12575 8449 12587 8452
rect 12529 8443 12587 8449
rect 12618 8440 12624 8452
rect 12676 8440 12682 8492
rect 13173 8483 13231 8489
rect 13173 8449 13185 8483
rect 13219 8480 13231 8483
rect 13906 8480 13912 8492
rect 13219 8452 13912 8480
rect 13219 8449 13231 8452
rect 13173 8443 13231 8449
rect 13906 8440 13912 8452
rect 13964 8440 13970 8492
rect 15194 8440 15200 8492
rect 15252 8480 15258 8492
rect 15289 8483 15347 8489
rect 15289 8480 15301 8483
rect 15252 8452 15301 8480
rect 15252 8440 15258 8452
rect 15289 8449 15301 8452
rect 15335 8449 15347 8483
rect 15289 8443 15347 8449
rect 15838 8440 15844 8492
rect 15896 8480 15902 8492
rect 18785 8483 18843 8489
rect 18785 8480 18797 8483
rect 15896 8452 18797 8480
rect 15896 8440 15902 8452
rect 18785 8449 18797 8452
rect 18831 8480 18843 8483
rect 18877 8483 18935 8489
rect 18877 8480 18889 8483
rect 18831 8452 18889 8480
rect 18831 8449 18843 8452
rect 18785 8443 18843 8449
rect 18877 8449 18889 8452
rect 18923 8449 18935 8483
rect 19058 8480 19064 8492
rect 19019 8452 19064 8480
rect 18877 8443 18935 8449
rect 19058 8440 19064 8452
rect 19116 8440 19122 8492
rect 20162 8440 20168 8492
rect 20220 8480 20226 8492
rect 21177 8483 21235 8489
rect 21177 8480 21189 8483
rect 20220 8452 21189 8480
rect 20220 8440 20226 8452
rect 21177 8449 21189 8452
rect 21223 8480 21235 8483
rect 21266 8480 21272 8492
rect 21223 8452 21272 8480
rect 21223 8449 21235 8452
rect 21177 8443 21235 8449
rect 21266 8440 21272 8452
rect 21324 8440 21330 8492
rect 10689 8415 10747 8421
rect 10689 8381 10701 8415
rect 10735 8381 10747 8415
rect 10689 8375 10747 8381
rect 14068 8415 14126 8421
rect 14068 8381 14080 8415
rect 14114 8412 14126 8415
rect 14458 8412 14464 8424
rect 14114 8384 14464 8412
rect 14114 8381 14126 8384
rect 14068 8375 14126 8381
rect 14458 8372 14464 8384
rect 14516 8372 14522 8424
rect 18046 8412 18052 8424
rect 18104 8421 18110 8424
rect 18104 8415 18142 8421
rect 17994 8384 18052 8412
rect 18046 8372 18052 8384
rect 18130 8412 18142 8415
rect 18509 8415 18567 8421
rect 18509 8412 18521 8415
rect 18130 8384 18521 8412
rect 18130 8381 18142 8384
rect 18104 8375 18142 8381
rect 18509 8381 18521 8384
rect 18555 8381 18567 8415
rect 18509 8375 18567 8381
rect 19029 8384 19518 8412
rect 18104 8372 18110 8375
rect 4341 8347 4399 8353
rect 4341 8313 4353 8347
rect 4387 8344 4399 8347
rect 4617 8347 4675 8353
rect 4617 8344 4629 8347
rect 4387 8316 4629 8344
rect 4387 8313 4399 8316
rect 4341 8307 4399 8313
rect 4617 8313 4629 8316
rect 4663 8313 4675 8347
rect 4617 8307 4675 8313
rect 6641 8347 6699 8353
rect 6641 8313 6653 8347
rect 6687 8344 6699 8347
rect 7285 8347 7343 8353
rect 7285 8344 7297 8347
rect 6687 8316 7297 8344
rect 6687 8313 6699 8316
rect 6641 8307 6699 8313
rect 7285 8313 7297 8316
rect 7331 8344 7343 8347
rect 7374 8344 7380 8356
rect 7331 8316 7380 8344
rect 7331 8313 7343 8316
rect 7285 8307 7343 8313
rect 1670 8276 1676 8288
rect 1631 8248 1676 8276
rect 1670 8236 1676 8248
rect 1728 8236 1734 8288
rect 3142 8276 3148 8288
rect 3103 8248 3148 8276
rect 3142 8236 3148 8248
rect 3200 8236 3206 8288
rect 3970 8276 3976 8288
rect 3931 8248 3976 8276
rect 3970 8236 3976 8248
rect 4028 8236 4034 8288
rect 4632 8276 4660 8307
rect 7374 8304 7380 8316
rect 7432 8304 7438 8356
rect 7558 8344 7564 8356
rect 7519 8316 7564 8344
rect 7558 8304 7564 8316
rect 7616 8304 7622 8356
rect 7653 8347 7711 8353
rect 7653 8313 7665 8347
rect 7699 8313 7711 8347
rect 10962 8344 10968 8356
rect 10923 8316 10968 8344
rect 7653 8307 7711 8313
rect 4706 8276 4712 8288
rect 4619 8248 4712 8276
rect 4706 8236 4712 8248
rect 4764 8276 4770 8288
rect 4982 8276 4988 8288
rect 4764 8248 4988 8276
rect 4764 8236 4770 8248
rect 4982 8236 4988 8248
rect 5040 8276 5046 8288
rect 5445 8279 5503 8285
rect 5445 8276 5457 8279
rect 5040 8248 5457 8276
rect 5040 8236 5046 8248
rect 5445 8245 5457 8248
rect 5491 8245 5503 8279
rect 7392 8276 7420 8304
rect 7668 8276 7696 8307
rect 10962 8304 10968 8316
rect 11020 8304 11026 8356
rect 12621 8347 12679 8353
rect 12621 8313 12633 8347
rect 12667 8313 12679 8347
rect 12621 8307 12679 8313
rect 15651 8347 15709 8353
rect 15651 8313 15663 8347
rect 15697 8344 15709 8347
rect 15838 8344 15844 8356
rect 15697 8316 15844 8344
rect 15697 8313 15709 8316
rect 15651 8307 15709 8313
rect 11330 8276 11336 8288
rect 7392 8248 7696 8276
rect 11291 8248 11336 8276
rect 5445 8239 5503 8245
rect 11330 8236 11336 8248
rect 11388 8236 11394 8288
rect 12250 8236 12256 8288
rect 12308 8276 12314 8288
rect 12636 8276 12664 8307
rect 15838 8304 15844 8316
rect 15896 8304 15902 8356
rect 17310 8304 17316 8356
rect 17368 8344 17374 8356
rect 19029 8344 19057 8384
rect 17368 8316 19057 8344
rect 19382 8347 19440 8353
rect 17368 8304 17374 8316
rect 19382 8313 19394 8347
rect 19428 8313 19440 8347
rect 19490 8344 19518 8384
rect 19886 8344 19892 8356
rect 19490 8316 19892 8344
rect 19382 8307 19440 8313
rect 12308 8248 12664 8276
rect 12308 8236 12314 8248
rect 13538 8236 13544 8288
rect 13596 8276 13602 8288
rect 13633 8279 13691 8285
rect 13633 8276 13645 8279
rect 13596 8248 13645 8276
rect 13596 8236 13602 8248
rect 13633 8245 13645 8248
rect 13679 8245 13691 8279
rect 13633 8239 13691 8245
rect 13722 8236 13728 8288
rect 13780 8276 13786 8288
rect 14139 8279 14197 8285
rect 14139 8276 14151 8279
rect 13780 8248 14151 8276
rect 13780 8236 13786 8248
rect 14139 8245 14151 8248
rect 14185 8245 14197 8279
rect 14139 8239 14197 8245
rect 15197 8279 15255 8285
rect 15197 8245 15209 8279
rect 15243 8276 15255 8279
rect 15470 8276 15476 8288
rect 15243 8248 15476 8276
rect 15243 8245 15255 8248
rect 15197 8239 15255 8245
rect 15470 8236 15476 8248
rect 15528 8276 15534 8288
rect 17402 8276 17408 8288
rect 15528 8248 17408 8276
rect 15528 8236 15534 8248
rect 17402 8236 17408 8248
rect 17460 8236 17466 8288
rect 17862 8236 17868 8288
rect 17920 8276 17926 8288
rect 18187 8279 18245 8285
rect 18187 8276 18199 8279
rect 17920 8248 18199 8276
rect 17920 8236 17926 8248
rect 18187 8245 18199 8248
rect 18233 8245 18245 8279
rect 18187 8239 18245 8245
rect 18785 8279 18843 8285
rect 18785 8245 18797 8279
rect 18831 8276 18843 8279
rect 19242 8276 19248 8288
rect 18831 8248 19248 8276
rect 18831 8245 18843 8248
rect 18785 8239 18843 8245
rect 19242 8236 19248 8248
rect 19300 8276 19306 8288
rect 19397 8276 19425 8307
rect 19886 8304 19892 8316
rect 19944 8344 19950 8356
rect 20898 8344 20904 8356
rect 19944 8316 20904 8344
rect 19944 8304 19950 8316
rect 20898 8304 20904 8316
rect 20956 8304 20962 8356
rect 20993 8347 21051 8353
rect 20993 8313 21005 8347
rect 21039 8313 21051 8347
rect 20993 8307 21051 8313
rect 20622 8276 20628 8288
rect 19300 8248 19425 8276
rect 20583 8248 20628 8276
rect 19300 8236 19306 8248
rect 20622 8236 20628 8248
rect 20680 8276 20686 8288
rect 21008 8276 21036 8307
rect 20680 8248 21036 8276
rect 20680 8236 20686 8248
rect 1104 8186 22816 8208
rect 1104 8134 8982 8186
rect 9034 8134 9046 8186
rect 9098 8134 9110 8186
rect 9162 8134 9174 8186
rect 9226 8134 16982 8186
rect 17034 8134 17046 8186
rect 17098 8134 17110 8186
rect 17162 8134 17174 8186
rect 17226 8134 22816 8186
rect 1104 8112 22816 8134
rect 2501 8075 2559 8081
rect 2501 8041 2513 8075
rect 2547 8072 2559 8075
rect 3142 8072 3148 8084
rect 2547 8044 3148 8072
rect 2547 8041 2559 8044
rect 2501 8035 2559 8041
rect 3142 8032 3148 8044
rect 3200 8032 3206 8084
rect 4430 8072 4436 8084
rect 4391 8044 4436 8072
rect 4430 8032 4436 8044
rect 4488 8032 4494 8084
rect 4982 8072 4988 8084
rect 4943 8044 4988 8072
rect 4982 8032 4988 8044
rect 5040 8032 5046 8084
rect 7374 8072 7380 8084
rect 7335 8044 7380 8072
rect 7374 8032 7380 8044
rect 7432 8032 7438 8084
rect 7558 8032 7564 8084
rect 7616 8072 7622 8084
rect 7653 8075 7711 8081
rect 7653 8072 7665 8075
rect 7616 8044 7665 8072
rect 7616 8032 7622 8044
rect 7653 8041 7665 8044
rect 7699 8072 7711 8075
rect 8343 8075 8401 8081
rect 8343 8072 8355 8075
rect 7699 8044 8355 8072
rect 7699 8041 7711 8044
rect 7653 8035 7711 8041
rect 8343 8041 8355 8044
rect 8389 8041 8401 8075
rect 10962 8072 10968 8084
rect 10923 8044 10968 8072
rect 8343 8035 8401 8041
rect 10962 8032 10968 8044
rect 11020 8072 11026 8084
rect 11977 8075 12035 8081
rect 11020 8044 11100 8072
rect 11020 8032 11026 8044
rect 1581 8007 1639 8013
rect 1581 7973 1593 8007
rect 1627 8004 1639 8007
rect 1670 8004 1676 8016
rect 1627 7976 1676 8004
rect 1627 7973 1639 7976
rect 1581 7967 1639 7973
rect 1670 7964 1676 7976
rect 1728 7964 1734 8016
rect 6819 8007 6877 8013
rect 6819 7973 6831 8007
rect 6865 8004 6877 8007
rect 7006 8004 7012 8016
rect 6865 7976 7012 8004
rect 6865 7973 6877 7976
rect 6819 7967 6877 7973
rect 7006 7964 7012 7976
rect 7064 7964 7070 8016
rect 10226 8004 10232 8016
rect 10187 7976 10232 8004
rect 10226 7964 10232 7976
rect 10284 7964 10290 8016
rect 3028 7939 3086 7945
rect 3028 7905 3040 7939
rect 3074 7936 3086 7939
rect 3142 7936 3148 7948
rect 3074 7908 3148 7936
rect 3074 7905 3086 7908
rect 3028 7899 3086 7905
rect 3142 7896 3148 7908
rect 3200 7896 3206 7948
rect 5902 7896 5908 7948
rect 5960 7936 5966 7948
rect 8018 7936 8024 7948
rect 5960 7908 8024 7936
rect 5960 7896 5966 7908
rect 8018 7896 8024 7908
rect 8076 7896 8082 7948
rect 8205 7939 8263 7945
rect 8205 7905 8217 7939
rect 8251 7936 8263 7939
rect 8294 7936 8300 7948
rect 8251 7908 8300 7936
rect 8251 7905 8263 7908
rect 8205 7899 8263 7905
rect 8294 7896 8300 7908
rect 8352 7896 8358 7948
rect 9677 7939 9735 7945
rect 9677 7905 9689 7939
rect 9723 7905 9735 7939
rect 9858 7936 9864 7948
rect 9819 7908 9864 7936
rect 9677 7899 9735 7905
rect 1486 7868 1492 7880
rect 1447 7840 1492 7868
rect 1486 7828 1492 7840
rect 1544 7828 1550 7880
rect 2130 7868 2136 7880
rect 2091 7840 2136 7868
rect 2130 7828 2136 7840
rect 2188 7828 2194 7880
rect 4062 7868 4068 7880
rect 4023 7840 4068 7868
rect 4062 7828 4068 7840
rect 4120 7828 4126 7880
rect 6457 7871 6515 7877
rect 6457 7837 6469 7871
rect 6503 7837 6515 7871
rect 6457 7831 6515 7837
rect 2774 7732 2780 7744
rect 2735 7704 2780 7732
rect 2774 7692 2780 7704
rect 2832 7732 2838 7744
rect 3099 7735 3157 7741
rect 3099 7732 3111 7735
rect 2832 7704 3111 7732
rect 2832 7692 2838 7704
rect 3099 7701 3111 7704
rect 3145 7701 3157 7735
rect 3510 7732 3516 7744
rect 3471 7704 3516 7732
rect 3099 7695 3157 7701
rect 3510 7692 3516 7704
rect 3568 7692 3574 7744
rect 4798 7692 4804 7744
rect 4856 7732 4862 7744
rect 5261 7735 5319 7741
rect 5261 7732 5273 7735
rect 4856 7704 5273 7732
rect 4856 7692 4862 7704
rect 5261 7701 5273 7704
rect 5307 7701 5319 7735
rect 5261 7695 5319 7701
rect 5902 7692 5908 7744
rect 5960 7732 5966 7744
rect 6273 7735 6331 7741
rect 6273 7732 6285 7735
rect 5960 7704 6285 7732
rect 5960 7692 5966 7704
rect 6273 7701 6285 7704
rect 6319 7732 6331 7735
rect 6472 7732 6500 7831
rect 8846 7828 8852 7880
rect 8904 7868 8910 7880
rect 9692 7868 9720 7899
rect 9858 7896 9864 7908
rect 9916 7896 9922 7948
rect 11072 7945 11100 8044
rect 11977 8041 11989 8075
rect 12023 8072 12035 8075
rect 12250 8072 12256 8084
rect 12023 8044 12256 8072
rect 12023 8041 12035 8044
rect 11977 8035 12035 8041
rect 12250 8032 12256 8044
rect 12308 8032 12314 8084
rect 12342 8032 12348 8084
rect 12400 8072 12406 8084
rect 13722 8072 13728 8084
rect 12400 8044 13728 8072
rect 12400 8032 12406 8044
rect 13722 8032 13728 8044
rect 13780 8032 13786 8084
rect 15010 8032 15016 8084
rect 15068 8072 15074 8084
rect 18138 8072 18144 8084
rect 15068 8044 18144 8072
rect 15068 8032 15074 8044
rect 18138 8032 18144 8044
rect 18196 8032 18202 8084
rect 19889 8075 19947 8081
rect 19889 8041 19901 8075
rect 19935 8072 19947 8075
rect 20622 8072 20628 8084
rect 19935 8044 20628 8072
rect 19935 8041 19947 8044
rect 19889 8035 19947 8041
rect 20622 8032 20628 8044
rect 20680 8032 20686 8084
rect 11146 7964 11152 8016
rect 11204 8004 11210 8016
rect 11378 8007 11436 8013
rect 11378 8004 11390 8007
rect 11204 7976 11390 8004
rect 11204 7964 11210 7976
rect 11378 7973 11390 7976
rect 11424 7973 11436 8007
rect 11378 7967 11436 7973
rect 12526 7964 12532 8016
rect 12584 8004 12590 8016
rect 13354 8004 13360 8016
rect 12584 7976 13032 8004
rect 13315 7976 13360 8004
rect 12584 7964 12590 7976
rect 11057 7939 11115 7945
rect 11057 7905 11069 7939
rect 11103 7905 11115 7939
rect 12802 7936 12808 7948
rect 12763 7908 12808 7936
rect 11057 7899 11115 7905
rect 12802 7896 12808 7908
rect 12860 7896 12866 7948
rect 13004 7945 13032 7976
rect 13354 7964 13360 7976
rect 13412 7964 13418 8016
rect 16758 8004 16764 8016
rect 16719 7976 16764 8004
rect 16758 7964 16764 7976
rect 16816 7964 16822 8016
rect 17310 8004 17316 8016
rect 17271 7976 17316 8004
rect 17310 7964 17316 7976
rect 17368 7964 17374 8016
rect 19242 8004 19248 8016
rect 19203 7976 19248 8004
rect 19242 7964 19248 7976
rect 19300 7964 19306 8016
rect 20162 8004 20168 8016
rect 20123 7976 20168 8004
rect 20162 7964 20168 7976
rect 20220 7964 20226 8016
rect 20254 7964 20260 8016
rect 20312 8004 20318 8016
rect 21085 8007 21143 8013
rect 21085 8004 21097 8007
rect 20312 7976 21097 8004
rect 20312 7964 20318 7976
rect 21085 7973 21097 7976
rect 21131 8004 21143 8007
rect 21450 8004 21456 8016
rect 21131 7976 21456 8004
rect 21131 7973 21143 7976
rect 21085 7967 21143 7973
rect 21450 7964 21456 7976
rect 21508 7964 21514 8016
rect 12989 7939 13047 7945
rect 12989 7905 13001 7939
rect 13035 7905 13047 7939
rect 12989 7899 13047 7905
rect 14252 7939 14310 7945
rect 14252 7905 14264 7939
rect 14298 7936 14310 7939
rect 14734 7936 14740 7948
rect 14298 7908 14740 7936
rect 14298 7905 14310 7908
rect 14252 7899 14310 7905
rect 14734 7896 14740 7908
rect 14792 7896 14798 7948
rect 15197 7939 15255 7945
rect 15197 7905 15209 7939
rect 15243 7936 15255 7939
rect 15286 7936 15292 7948
rect 15243 7908 15292 7936
rect 15243 7905 15255 7908
rect 15197 7899 15255 7905
rect 15286 7896 15292 7908
rect 15344 7896 15350 7948
rect 10410 7868 10416 7880
rect 8904 7840 10416 7868
rect 8904 7828 8910 7840
rect 10410 7828 10416 7840
rect 10468 7868 10474 7880
rect 12820 7868 12848 7896
rect 10468 7840 12848 7868
rect 16669 7871 16727 7877
rect 10468 7828 10474 7840
rect 16669 7837 16681 7871
rect 16715 7868 16727 7871
rect 17034 7868 17040 7880
rect 16715 7840 17040 7868
rect 16715 7837 16727 7840
rect 16669 7831 16727 7837
rect 17034 7828 17040 7840
rect 17092 7868 17098 7880
rect 17862 7868 17868 7880
rect 17092 7840 17868 7868
rect 17092 7828 17098 7840
rect 17862 7828 17868 7840
rect 17920 7828 17926 7880
rect 18966 7868 18972 7880
rect 18927 7840 18972 7868
rect 18966 7828 18972 7840
rect 19024 7828 19030 7880
rect 20806 7828 20812 7880
rect 20864 7868 20870 7880
rect 20993 7871 21051 7877
rect 20993 7868 21005 7871
rect 20864 7840 21005 7868
rect 20864 7828 20870 7840
rect 20993 7837 21005 7840
rect 21039 7837 21051 7871
rect 21266 7868 21272 7880
rect 21227 7840 21272 7868
rect 20993 7831 21051 7837
rect 21266 7828 21272 7840
rect 21324 7828 21330 7880
rect 15427 7803 15485 7809
rect 15427 7769 15439 7803
rect 15473 7800 15485 7803
rect 15654 7800 15660 7812
rect 15473 7772 15660 7800
rect 15473 7769 15485 7772
rect 15427 7763 15485 7769
rect 15654 7760 15660 7772
rect 15712 7800 15718 7812
rect 16117 7803 16175 7809
rect 16117 7800 16129 7803
rect 15712 7772 16129 7800
rect 15712 7760 15718 7772
rect 16117 7769 16129 7772
rect 16163 7769 16175 7803
rect 16117 7763 16175 7769
rect 9490 7732 9496 7744
rect 6319 7704 6500 7732
rect 9451 7704 9496 7732
rect 6319 7701 6331 7704
rect 6273 7695 6331 7701
rect 9490 7692 9496 7704
rect 9548 7692 9554 7744
rect 10134 7692 10140 7744
rect 10192 7732 10198 7744
rect 10505 7735 10563 7741
rect 10505 7732 10517 7735
rect 10192 7704 10517 7732
rect 10192 7692 10198 7704
rect 10505 7701 10517 7704
rect 10551 7701 10563 7735
rect 12618 7732 12624 7744
rect 12579 7704 12624 7732
rect 10505 7695 10563 7701
rect 12618 7692 12624 7704
rect 12676 7692 12682 7744
rect 13814 7692 13820 7744
rect 13872 7732 13878 7744
rect 13872 7704 13917 7732
rect 13872 7692 13878 7704
rect 14182 7692 14188 7744
rect 14240 7732 14246 7744
rect 14323 7735 14381 7741
rect 14323 7732 14335 7735
rect 14240 7704 14335 7732
rect 14240 7692 14246 7704
rect 14323 7701 14335 7704
rect 14369 7701 14381 7735
rect 15838 7732 15844 7744
rect 15799 7704 15844 7732
rect 14323 7695 14381 7701
rect 15838 7692 15844 7704
rect 15896 7692 15902 7744
rect 1104 7642 22816 7664
rect 1104 7590 4982 7642
rect 5034 7590 5046 7642
rect 5098 7590 5110 7642
rect 5162 7590 5174 7642
rect 5226 7590 12982 7642
rect 13034 7590 13046 7642
rect 13098 7590 13110 7642
rect 13162 7590 13174 7642
rect 13226 7590 20982 7642
rect 21034 7590 21046 7642
rect 21098 7590 21110 7642
rect 21162 7590 21174 7642
rect 21226 7590 22816 7642
rect 1104 7568 22816 7590
rect 1670 7528 1676 7540
rect 1631 7500 1676 7528
rect 1670 7488 1676 7500
rect 1728 7488 1734 7540
rect 3053 7531 3111 7537
rect 3053 7497 3065 7531
rect 3099 7528 3111 7531
rect 3142 7528 3148 7540
rect 3099 7500 3148 7528
rect 3099 7497 3111 7500
rect 3053 7491 3111 7497
rect 3142 7488 3148 7500
rect 3200 7488 3206 7540
rect 4430 7528 4436 7540
rect 4343 7500 4436 7528
rect 4430 7488 4436 7500
rect 4488 7528 4494 7540
rect 6549 7531 6607 7537
rect 6549 7528 6561 7531
rect 4488 7500 6561 7528
rect 4488 7488 4494 7500
rect 6549 7497 6561 7500
rect 6595 7528 6607 7531
rect 7006 7528 7012 7540
rect 6595 7500 7012 7528
rect 6595 7497 6607 7500
rect 6549 7491 6607 7497
rect 7006 7488 7012 7500
rect 7064 7488 7070 7540
rect 8846 7528 8852 7540
rect 8807 7500 8852 7528
rect 8846 7488 8852 7500
rect 8904 7488 8910 7540
rect 9490 7488 9496 7540
rect 9548 7528 9554 7540
rect 9815 7531 9873 7537
rect 9815 7528 9827 7531
rect 9548 7500 9827 7528
rect 9548 7488 9554 7500
rect 9815 7497 9827 7500
rect 9861 7497 9873 7531
rect 9815 7491 9873 7497
rect 11471 7531 11529 7537
rect 11471 7497 11483 7531
rect 11517 7528 11529 7531
rect 12618 7528 12624 7540
rect 11517 7500 12624 7528
rect 11517 7497 11529 7500
rect 11471 7491 11529 7497
rect 12618 7488 12624 7500
rect 12676 7488 12682 7540
rect 12802 7488 12808 7540
rect 12860 7528 12866 7540
rect 13541 7531 13599 7537
rect 13541 7528 13553 7531
rect 12860 7500 13553 7528
rect 12860 7488 12866 7500
rect 13541 7497 13553 7500
rect 13587 7497 13599 7531
rect 14734 7528 14740 7540
rect 14695 7500 14740 7528
rect 13541 7491 13599 7497
rect 14734 7488 14740 7500
rect 14792 7488 14798 7540
rect 16669 7531 16727 7537
rect 16669 7497 16681 7531
rect 16715 7528 16727 7531
rect 16758 7528 16764 7540
rect 16715 7500 16764 7528
rect 16715 7497 16727 7500
rect 16669 7491 16727 7497
rect 16758 7488 16764 7500
rect 16816 7488 16822 7540
rect 17034 7528 17040 7540
rect 16995 7500 17040 7528
rect 17034 7488 17040 7500
rect 17092 7488 17098 7540
rect 20254 7528 20260 7540
rect 20215 7500 20260 7528
rect 20254 7488 20260 7500
rect 20312 7488 20318 7540
rect 20806 7488 20812 7540
rect 20864 7528 20870 7540
rect 20901 7531 20959 7537
rect 20901 7528 20913 7531
rect 20864 7500 20913 7528
rect 20864 7488 20870 7500
rect 20901 7497 20913 7500
rect 20947 7497 20959 7531
rect 20901 7491 20959 7497
rect 2130 7420 2136 7472
rect 2188 7460 2194 7472
rect 2409 7463 2467 7469
rect 2409 7460 2421 7463
rect 2188 7432 2421 7460
rect 2188 7420 2194 7432
rect 2409 7429 2421 7432
rect 2455 7429 2467 7463
rect 2409 7423 2467 7429
rect 9953 7463 10011 7469
rect 9953 7429 9965 7463
rect 9999 7460 10011 7463
rect 10134 7460 10140 7472
rect 9999 7432 10140 7460
rect 9999 7429 10011 7432
rect 9953 7423 10011 7429
rect 10134 7420 10140 7432
rect 10192 7420 10198 7472
rect 10321 7463 10379 7469
rect 10321 7429 10333 7463
rect 10367 7460 10379 7463
rect 13446 7460 13452 7472
rect 10367 7432 13452 7460
rect 10367 7429 10379 7432
rect 10321 7423 10379 7429
rect 13446 7420 13452 7432
rect 13504 7420 13510 7472
rect 14369 7463 14427 7469
rect 14369 7429 14381 7463
rect 14415 7460 14427 7463
rect 14918 7460 14924 7472
rect 14415 7432 14924 7460
rect 14415 7429 14427 7432
rect 14369 7423 14427 7429
rect 14918 7420 14924 7432
rect 14976 7460 14982 7472
rect 14976 7432 15976 7460
rect 14976 7420 14982 7432
rect 1857 7395 1915 7401
rect 1857 7361 1869 7395
rect 1903 7392 1915 7395
rect 2774 7392 2780 7404
rect 1903 7364 2780 7392
rect 1903 7361 1915 7364
rect 1857 7355 1915 7361
rect 2774 7352 2780 7364
rect 2832 7352 2838 7404
rect 2866 7352 2872 7404
rect 2924 7392 2930 7404
rect 3418 7392 3424 7404
rect 2924 7364 3424 7392
rect 2924 7352 2930 7364
rect 3418 7352 3424 7364
rect 3476 7392 3482 7404
rect 5902 7392 5908 7404
rect 3476 7364 5120 7392
rect 5863 7364 5908 7392
rect 3476 7352 3482 7364
rect 3510 7324 3516 7336
rect 3471 7296 3516 7324
rect 3510 7284 3516 7296
rect 3568 7284 3574 7336
rect 3804 7333 3832 7364
rect 3789 7327 3847 7333
rect 3789 7324 3801 7327
rect 3767 7296 3801 7324
rect 3789 7293 3801 7296
rect 3835 7293 3847 7327
rect 4062 7324 4068 7336
rect 4023 7296 4068 7324
rect 3789 7287 3847 7293
rect 4062 7284 4068 7296
rect 4120 7284 4126 7336
rect 1946 7256 1952 7268
rect 1907 7228 1952 7256
rect 1946 7216 1952 7228
rect 2004 7216 2010 7268
rect 5092 7265 5120 7364
rect 5902 7352 5908 7364
rect 5960 7352 5966 7404
rect 10045 7395 10103 7401
rect 10045 7361 10057 7395
rect 10091 7392 10103 7395
rect 10226 7392 10232 7404
rect 10091 7364 10232 7392
rect 10091 7361 10103 7364
rect 10045 7355 10103 7361
rect 10226 7352 10232 7364
rect 10284 7352 10290 7404
rect 11885 7395 11943 7401
rect 11885 7392 11897 7395
rect 11415 7364 11897 7392
rect 5442 7324 5448 7336
rect 5403 7296 5448 7324
rect 5442 7284 5448 7296
rect 5500 7284 5506 7336
rect 5721 7327 5779 7333
rect 5721 7293 5733 7327
rect 5767 7293 5779 7327
rect 5721 7287 5779 7293
rect 7101 7327 7159 7333
rect 7101 7293 7113 7327
rect 7147 7324 7159 7327
rect 7377 7327 7435 7333
rect 7377 7324 7389 7327
rect 7147 7296 7389 7324
rect 7147 7293 7159 7296
rect 7101 7287 7159 7293
rect 7377 7293 7389 7296
rect 7423 7324 7435 7327
rect 7466 7324 7472 7336
rect 7423 7296 7472 7324
rect 7423 7293 7435 7296
rect 7377 7287 7435 7293
rect 5077 7259 5135 7265
rect 5077 7225 5089 7259
rect 5123 7256 5135 7259
rect 5736 7256 5764 7287
rect 7466 7284 7472 7296
rect 7524 7284 7530 7336
rect 8294 7324 8300 7336
rect 8207 7296 8300 7324
rect 8294 7284 8300 7296
rect 8352 7324 8358 7336
rect 11415 7333 11443 7364
rect 11885 7361 11897 7364
rect 11931 7392 11943 7395
rect 13817 7395 13875 7401
rect 11931 7364 13676 7392
rect 11931 7361 11943 7364
rect 11885 7355 11943 7361
rect 11400 7327 11458 7333
rect 11400 7324 11412 7327
rect 8352 7296 11412 7324
rect 8352 7284 8358 7296
rect 11400 7293 11412 7296
rect 11446 7293 11458 7327
rect 11400 7287 11458 7293
rect 12764 7327 12822 7333
rect 12764 7293 12776 7327
rect 12810 7324 12822 7327
rect 13265 7327 13323 7333
rect 13265 7324 13277 7327
rect 12810 7296 13277 7324
rect 12810 7293 12822 7296
rect 12764 7287 12822 7293
rect 13265 7293 13277 7296
rect 13311 7324 13323 7327
rect 13354 7324 13360 7336
rect 13311 7296 13360 7324
rect 13311 7293 13323 7296
rect 13265 7287 13323 7293
rect 13354 7284 13360 7296
rect 13412 7284 13418 7336
rect 5123 7228 7138 7256
rect 5123 7225 5135 7228
rect 5077 7219 5135 7225
rect 3142 7148 3148 7200
rect 3200 7188 3206 7200
rect 4430 7188 4436 7200
rect 3200 7160 4436 7188
rect 3200 7148 3206 7160
rect 4430 7148 4436 7160
rect 4488 7148 4494 7200
rect 7110 7188 7138 7228
rect 7190 7216 7196 7268
rect 7248 7256 7254 7268
rect 7484 7256 7512 7284
rect 9125 7259 9183 7265
rect 9125 7256 9137 7259
rect 7248 7228 7293 7256
rect 7484 7228 9137 7256
rect 7248 7216 7254 7228
rect 9125 7225 9137 7228
rect 9171 7256 9183 7259
rect 9493 7259 9551 7265
rect 9493 7256 9505 7259
rect 9171 7228 9505 7256
rect 9171 7225 9183 7228
rect 9125 7219 9183 7225
rect 9493 7225 9505 7228
rect 9539 7256 9551 7259
rect 9677 7259 9735 7265
rect 9677 7256 9689 7259
rect 9539 7228 9689 7256
rect 9539 7225 9551 7228
rect 9493 7219 9551 7225
rect 9677 7225 9689 7228
rect 9723 7256 9735 7259
rect 9858 7256 9864 7268
rect 9723 7228 9864 7256
rect 9723 7225 9735 7228
rect 9677 7219 9735 7225
rect 9858 7216 9864 7228
rect 9916 7216 9922 7268
rect 12851 7259 12909 7265
rect 12851 7225 12863 7259
rect 12897 7256 12909 7259
rect 13446 7256 13452 7268
rect 12897 7228 13452 7256
rect 12897 7225 12909 7228
rect 12851 7219 12909 7225
rect 13446 7216 13452 7228
rect 13504 7216 13510 7268
rect 7469 7191 7527 7197
rect 7469 7188 7481 7191
rect 7110 7160 7481 7188
rect 7469 7157 7481 7160
rect 7515 7157 7527 7191
rect 7469 7151 7527 7157
rect 10226 7148 10232 7200
rect 10284 7188 10290 7200
rect 10689 7191 10747 7197
rect 10689 7188 10701 7191
rect 10284 7160 10701 7188
rect 10284 7148 10290 7160
rect 10689 7157 10701 7160
rect 10735 7157 10747 7191
rect 11146 7188 11152 7200
rect 11107 7160 11152 7188
rect 10689 7151 10747 7157
rect 11146 7148 11152 7160
rect 11204 7148 11210 7200
rect 11238 7148 11244 7200
rect 11296 7188 11302 7200
rect 12161 7191 12219 7197
rect 12161 7188 12173 7191
rect 11296 7160 12173 7188
rect 11296 7148 11302 7160
rect 12161 7157 12173 7160
rect 12207 7188 12219 7191
rect 12618 7188 12624 7200
rect 12207 7160 12624 7188
rect 12207 7157 12219 7160
rect 12161 7151 12219 7157
rect 12618 7148 12624 7160
rect 12676 7148 12682 7200
rect 13648 7188 13676 7364
rect 13817 7361 13829 7395
rect 13863 7392 13875 7395
rect 14182 7392 14188 7404
rect 13863 7364 14188 7392
rect 13863 7361 13875 7364
rect 13817 7355 13875 7361
rect 14182 7352 14188 7364
rect 14240 7352 14246 7404
rect 15654 7392 15660 7404
rect 15615 7364 15660 7392
rect 15654 7352 15660 7364
rect 15712 7352 15718 7404
rect 15948 7401 15976 7432
rect 15933 7395 15991 7401
rect 15933 7361 15945 7395
rect 15979 7361 15991 7395
rect 15933 7355 15991 7361
rect 18966 7352 18972 7404
rect 19024 7392 19030 7404
rect 20533 7395 20591 7401
rect 20533 7392 20545 7395
rect 19024 7364 20545 7392
rect 19024 7352 19030 7364
rect 20533 7361 20545 7364
rect 20579 7361 20591 7395
rect 20916 7392 20944 7491
rect 21450 7488 21456 7540
rect 21508 7528 21514 7540
rect 21545 7531 21603 7537
rect 21545 7528 21557 7531
rect 21508 7500 21557 7528
rect 21508 7488 21514 7500
rect 21545 7497 21557 7500
rect 21591 7497 21603 7531
rect 21545 7491 21603 7497
rect 21085 7395 21143 7401
rect 21085 7392 21097 7395
rect 20916 7364 21097 7392
rect 20533 7355 20591 7361
rect 21085 7361 21097 7364
rect 21131 7361 21143 7395
rect 21085 7355 21143 7361
rect 17954 7284 17960 7336
rect 18012 7324 18018 7336
rect 18084 7327 18142 7333
rect 18084 7324 18096 7327
rect 18012 7296 18096 7324
rect 18012 7284 18018 7296
rect 18084 7293 18096 7296
rect 18130 7324 18142 7327
rect 18509 7327 18567 7333
rect 18509 7324 18521 7327
rect 18130 7296 18521 7324
rect 18130 7293 18142 7296
rect 18084 7287 18142 7293
rect 18509 7293 18521 7296
rect 18555 7293 18567 7327
rect 18509 7287 18567 7293
rect 19337 7327 19395 7333
rect 19337 7293 19349 7327
rect 19383 7324 19395 7327
rect 20162 7324 20168 7336
rect 19383 7296 20168 7324
rect 19383 7293 19395 7296
rect 19337 7287 19395 7293
rect 20162 7284 20168 7296
rect 20220 7284 20226 7336
rect 13814 7216 13820 7268
rect 13872 7256 13878 7268
rect 13909 7259 13967 7265
rect 13909 7256 13921 7259
rect 13872 7228 13921 7256
rect 13872 7216 13878 7228
rect 13909 7225 13921 7228
rect 13955 7225 13967 7259
rect 15746 7256 15752 7268
rect 15707 7228 15752 7256
rect 13909 7219 13967 7225
rect 15746 7216 15752 7228
rect 15804 7216 15810 7268
rect 19658 7259 19716 7265
rect 19658 7256 19670 7259
rect 19306 7228 19670 7256
rect 15286 7188 15292 7200
rect 13648 7160 15292 7188
rect 15286 7148 15292 7160
rect 15344 7148 15350 7200
rect 16114 7148 16120 7200
rect 16172 7188 16178 7200
rect 18187 7191 18245 7197
rect 18187 7188 18199 7191
rect 16172 7160 18199 7188
rect 16172 7148 16178 7160
rect 18187 7157 18199 7160
rect 18233 7157 18245 7191
rect 18187 7151 18245 7157
rect 19058 7148 19064 7200
rect 19116 7188 19122 7200
rect 19153 7191 19211 7197
rect 19153 7188 19165 7191
rect 19116 7160 19165 7188
rect 19116 7148 19122 7160
rect 19153 7157 19165 7160
rect 19199 7188 19211 7191
rect 19306 7188 19334 7228
rect 19658 7225 19670 7228
rect 19704 7225 19716 7259
rect 19658 7219 19716 7225
rect 19199 7160 19334 7188
rect 19199 7157 19211 7160
rect 19153 7151 19211 7157
rect 1104 7098 22816 7120
rect 1104 7046 8982 7098
rect 9034 7046 9046 7098
rect 9098 7046 9110 7098
rect 9162 7046 9174 7098
rect 9226 7046 16982 7098
rect 17034 7046 17046 7098
rect 17098 7046 17110 7098
rect 17162 7046 17174 7098
rect 17226 7046 22816 7098
rect 1104 7024 22816 7046
rect 1486 6944 1492 6996
rect 1544 6984 1550 6996
rect 2869 6987 2927 6993
rect 2869 6984 2881 6987
rect 1544 6956 2881 6984
rect 1544 6944 1550 6956
rect 2869 6953 2881 6956
rect 2915 6953 2927 6987
rect 3418 6984 3424 6996
rect 3379 6956 3424 6984
rect 2869 6947 2927 6953
rect 3418 6944 3424 6956
rect 3476 6944 3482 6996
rect 4062 6944 4068 6996
rect 4120 6984 4126 6996
rect 4709 6987 4767 6993
rect 4709 6984 4721 6987
rect 4120 6956 4721 6984
rect 4120 6944 4126 6956
rect 4709 6953 4721 6956
rect 4755 6953 4767 6987
rect 4709 6947 4767 6953
rect 5718 6944 5724 6996
rect 5776 6984 5782 6996
rect 8205 6987 8263 6993
rect 8205 6984 8217 6987
rect 5776 6956 8217 6984
rect 5776 6944 5782 6956
rect 8205 6953 8217 6956
rect 8251 6953 8263 6987
rect 8205 6947 8263 6953
rect 11146 6944 11152 6996
rect 11204 6984 11210 6996
rect 13541 6987 13599 6993
rect 11204 6956 13026 6984
rect 11204 6944 11210 6956
rect 2038 6925 2044 6928
rect 2035 6916 2044 6925
rect 1951 6888 2044 6916
rect 2035 6879 2044 6888
rect 2096 6916 2102 6928
rect 3142 6916 3148 6928
rect 2096 6888 3148 6916
rect 2038 6876 2044 6879
rect 2096 6876 2102 6888
rect 3142 6876 3148 6888
rect 3200 6876 3206 6928
rect 4387 6919 4445 6925
rect 4387 6885 4399 6919
rect 4433 6916 4445 6919
rect 4798 6916 4804 6928
rect 4433 6888 4804 6916
rect 4433 6885 4445 6888
rect 4387 6879 4445 6885
rect 4798 6876 4804 6888
rect 4856 6876 4862 6928
rect 5350 6876 5356 6928
rect 5408 6916 5414 6928
rect 7561 6919 7619 6925
rect 7561 6916 7573 6919
rect 5408 6888 7573 6916
rect 5408 6876 5414 6888
rect 7561 6885 7573 6888
rect 7607 6916 7619 6919
rect 8573 6919 8631 6925
rect 8573 6916 8585 6919
rect 7607 6888 8585 6916
rect 7607 6885 7619 6888
rect 7561 6879 7619 6885
rect 8573 6885 8585 6888
rect 8619 6916 8631 6919
rect 9861 6919 9919 6925
rect 9861 6916 9873 6919
rect 8619 6888 9873 6916
rect 8619 6885 8631 6888
rect 8573 6879 8631 6885
rect 9861 6885 9873 6888
rect 9907 6885 9919 6919
rect 9861 6879 9919 6885
rect 10597 6919 10655 6925
rect 10597 6885 10609 6919
rect 10643 6916 10655 6919
rect 12710 6916 12716 6928
rect 10643 6888 12716 6916
rect 10643 6885 10655 6888
rect 10597 6879 10655 6885
rect 4300 6851 4358 6857
rect 4300 6817 4312 6851
rect 4346 6848 4358 6851
rect 4614 6848 4620 6860
rect 4346 6820 4620 6848
rect 4346 6817 4358 6820
rect 4300 6811 4358 6817
rect 4614 6808 4620 6820
rect 4672 6808 4678 6860
rect 5534 6848 5540 6860
rect 5495 6820 5540 6848
rect 5534 6808 5540 6820
rect 5592 6808 5598 6860
rect 5813 6851 5871 6857
rect 5813 6817 5825 6851
rect 5859 6848 5871 6851
rect 5902 6848 5908 6860
rect 5859 6820 5908 6848
rect 5859 6817 5871 6820
rect 5813 6811 5871 6817
rect 5902 6808 5908 6820
rect 5960 6808 5966 6860
rect 7650 6808 7656 6860
rect 7708 6857 7714 6860
rect 7708 6851 7766 6857
rect 7708 6817 7720 6851
rect 7754 6817 7766 6851
rect 9876 6848 9904 6879
rect 12710 6876 12716 6888
rect 12768 6876 12774 6928
rect 12998 6925 13026 6956
rect 13541 6953 13553 6987
rect 13587 6984 13599 6987
rect 13814 6984 13820 6996
rect 13587 6956 13820 6984
rect 13587 6953 13599 6956
rect 13541 6947 13599 6953
rect 13814 6944 13820 6956
rect 13872 6984 13878 6996
rect 14182 6984 14188 6996
rect 13872 6956 13917 6984
rect 14143 6956 14188 6984
rect 13872 6944 13878 6956
rect 14182 6944 14188 6956
rect 14240 6944 14246 6996
rect 19150 6944 19156 6996
rect 19208 6984 19214 6996
rect 19610 6984 19616 6996
rect 19208 6956 19616 6984
rect 19208 6944 19214 6956
rect 19610 6944 19616 6956
rect 19668 6944 19674 6996
rect 12983 6919 13041 6925
rect 12983 6885 12995 6919
rect 13029 6885 13041 6919
rect 12983 6879 13041 6885
rect 15657 6919 15715 6925
rect 15657 6885 15669 6919
rect 15703 6916 15715 6919
rect 15746 6916 15752 6928
rect 15703 6888 15752 6916
rect 15703 6885 15715 6888
rect 15657 6879 15715 6885
rect 15746 6876 15752 6888
rect 15804 6916 15810 6928
rect 16206 6916 16212 6928
rect 15804 6888 16212 6916
rect 15804 6876 15810 6888
rect 16206 6876 16212 6888
rect 16264 6876 16270 6928
rect 18693 6919 18751 6925
rect 18693 6885 18705 6919
rect 18739 6916 18751 6919
rect 18966 6916 18972 6928
rect 18739 6888 18972 6916
rect 18739 6885 18751 6888
rect 18693 6879 18751 6885
rect 18966 6876 18972 6888
rect 19024 6876 19030 6928
rect 11238 6848 11244 6860
rect 9876 6820 11244 6848
rect 7708 6811 7766 6817
rect 7708 6808 7714 6811
rect 11238 6808 11244 6820
rect 11296 6808 11302 6860
rect 17954 6848 17960 6860
rect 17915 6820 17960 6848
rect 17954 6808 17960 6820
rect 18012 6808 18018 6860
rect 18509 6851 18567 6857
rect 18509 6817 18521 6851
rect 18555 6848 18567 6851
rect 18598 6848 18604 6860
rect 18555 6820 18604 6848
rect 18555 6817 18567 6820
rect 18509 6811 18567 6817
rect 18598 6808 18604 6820
rect 18656 6808 18662 6860
rect 1673 6783 1731 6789
rect 1673 6749 1685 6783
rect 1719 6780 1731 6783
rect 2314 6780 2320 6792
rect 1719 6752 2320 6780
rect 1719 6749 1731 6752
rect 1673 6743 1731 6749
rect 2314 6740 2320 6752
rect 2372 6740 2378 6792
rect 5994 6780 6000 6792
rect 5955 6752 6000 6780
rect 5994 6740 6000 6752
rect 6052 6740 6058 6792
rect 7926 6780 7932 6792
rect 7024 6752 7932 6780
rect 1946 6672 1952 6724
rect 2004 6712 2010 6724
rect 2593 6715 2651 6721
rect 2593 6712 2605 6715
rect 2004 6684 2605 6712
rect 2004 6672 2010 6684
rect 2593 6681 2605 6684
rect 2639 6681 2651 6715
rect 2593 6675 2651 6681
rect 5629 6715 5687 6721
rect 5629 6681 5641 6715
rect 5675 6712 5687 6715
rect 6086 6712 6092 6724
rect 5675 6684 6092 6712
rect 5675 6681 5687 6684
rect 5629 6675 5687 6681
rect 6086 6672 6092 6684
rect 6144 6672 6150 6724
rect 7024 6656 7052 6752
rect 7926 6740 7932 6752
rect 7984 6740 7990 6792
rect 9490 6740 9496 6792
rect 9548 6780 9554 6792
rect 10008 6783 10066 6789
rect 10008 6780 10020 6783
rect 9548 6752 10020 6780
rect 9548 6740 9554 6752
rect 10008 6749 10020 6752
rect 10054 6749 10066 6783
rect 10226 6780 10232 6792
rect 10187 6752 10232 6780
rect 10008 6743 10066 6749
rect 10226 6740 10232 6752
rect 10284 6740 10290 6792
rect 11517 6783 11575 6789
rect 11517 6749 11529 6783
rect 11563 6780 11575 6783
rect 11698 6780 11704 6792
rect 11563 6752 11704 6780
rect 11563 6749 11575 6752
rect 11517 6743 11575 6749
rect 11698 6740 11704 6752
rect 11756 6740 11762 6792
rect 12342 6740 12348 6792
rect 12400 6780 12406 6792
rect 12621 6783 12679 6789
rect 12621 6780 12633 6783
rect 12400 6752 12633 6780
rect 12400 6740 12406 6752
rect 12621 6749 12633 6752
rect 12667 6749 12679 6783
rect 16114 6780 16120 6792
rect 16075 6752 16120 6780
rect 12621 6743 12679 6749
rect 16114 6740 16120 6752
rect 16172 6740 16178 6792
rect 16298 6740 16304 6792
rect 16356 6780 16362 6792
rect 16761 6783 16819 6789
rect 16761 6780 16773 6783
rect 16356 6752 16773 6780
rect 16356 6740 16362 6752
rect 16761 6749 16773 6752
rect 16807 6780 16819 6783
rect 17586 6780 17592 6792
rect 16807 6752 17592 6780
rect 16807 6749 16819 6752
rect 16761 6743 16819 6749
rect 17586 6740 17592 6752
rect 17644 6740 17650 6792
rect 7190 6672 7196 6724
rect 7248 6712 7254 6724
rect 7285 6715 7343 6721
rect 7285 6712 7297 6715
rect 7248 6684 7297 6712
rect 7248 6672 7254 6684
rect 7285 6681 7297 6684
rect 7331 6712 7343 6715
rect 7742 6712 7748 6724
rect 7331 6684 7748 6712
rect 7331 6681 7343 6684
rect 7285 6675 7343 6681
rect 7742 6672 7748 6684
rect 7800 6672 7806 6724
rect 10134 6712 10140 6724
rect 10047 6684 10140 6712
rect 10134 6672 10140 6684
rect 10192 6712 10198 6724
rect 10192 6684 11008 6712
rect 10192 6672 10198 6684
rect 10980 6656 11008 6684
rect 5261 6647 5319 6653
rect 5261 6613 5273 6647
rect 5307 6644 5319 6647
rect 5442 6644 5448 6656
rect 5307 6616 5448 6644
rect 5307 6613 5319 6616
rect 5261 6607 5319 6613
rect 5442 6604 5448 6616
rect 5500 6644 5506 6656
rect 5718 6644 5724 6656
rect 5500 6616 5724 6644
rect 5500 6604 5506 6616
rect 5718 6604 5724 6616
rect 5776 6604 5782 6656
rect 6917 6647 6975 6653
rect 6917 6613 6929 6647
rect 6963 6644 6975 6647
rect 7006 6644 7012 6656
rect 6963 6616 7012 6644
rect 6963 6613 6975 6616
rect 6917 6607 6975 6613
rect 7006 6604 7012 6616
rect 7064 6604 7070 6656
rect 7834 6644 7840 6656
rect 7795 6616 7840 6644
rect 7834 6604 7840 6616
rect 7892 6604 7898 6656
rect 9122 6644 9128 6656
rect 9083 6616 9128 6644
rect 9122 6604 9128 6616
rect 9180 6604 9186 6656
rect 10962 6644 10968 6656
rect 10923 6616 10968 6644
rect 10962 6604 10968 6616
rect 11020 6604 11026 6656
rect 11747 6647 11805 6653
rect 11747 6613 11759 6647
rect 11793 6644 11805 6647
rect 12802 6644 12808 6656
rect 11793 6616 12808 6644
rect 11793 6613 11805 6616
rect 11747 6607 11805 6613
rect 12802 6604 12808 6616
rect 12860 6604 12866 6656
rect 18966 6644 18972 6656
rect 18927 6616 18972 6644
rect 18966 6604 18972 6616
rect 19024 6604 19030 6656
rect 20073 6647 20131 6653
rect 20073 6613 20085 6647
rect 20119 6644 20131 6647
rect 20162 6644 20168 6656
rect 20119 6616 20168 6644
rect 20119 6613 20131 6616
rect 20073 6607 20131 6613
rect 20162 6604 20168 6616
rect 20220 6604 20226 6656
rect 1104 6554 22816 6576
rect 1104 6502 4982 6554
rect 5034 6502 5046 6554
rect 5098 6502 5110 6554
rect 5162 6502 5174 6554
rect 5226 6502 12982 6554
rect 13034 6502 13046 6554
rect 13098 6502 13110 6554
rect 13162 6502 13174 6554
rect 13226 6502 20982 6554
rect 21034 6502 21046 6554
rect 21098 6502 21110 6554
rect 21162 6502 21174 6554
rect 21226 6502 22816 6554
rect 1104 6480 22816 6502
rect 1949 6443 2007 6449
rect 1949 6409 1961 6443
rect 1995 6440 2007 6443
rect 2038 6440 2044 6452
rect 1995 6412 2044 6440
rect 1995 6409 2007 6412
rect 1949 6403 2007 6409
rect 2038 6400 2044 6412
rect 2096 6400 2102 6452
rect 4614 6400 4620 6452
rect 4672 6440 4678 6452
rect 4801 6443 4859 6449
rect 4801 6440 4813 6443
rect 4672 6412 4813 6440
rect 4672 6400 4678 6412
rect 4801 6409 4813 6412
rect 4847 6409 4859 6443
rect 8018 6440 8024 6452
rect 7979 6412 8024 6440
rect 4801 6403 4859 6409
rect 8018 6400 8024 6412
rect 8076 6400 8082 6452
rect 9585 6443 9643 6449
rect 9585 6409 9597 6443
rect 9631 6440 9643 6443
rect 9674 6440 9680 6452
rect 9631 6412 9680 6440
rect 9631 6409 9643 6412
rect 9585 6403 9643 6409
rect 9674 6400 9680 6412
rect 9732 6400 9738 6452
rect 11698 6440 11704 6452
rect 11659 6412 11704 6440
rect 11698 6400 11704 6412
rect 11756 6400 11762 6452
rect 16206 6440 16212 6452
rect 16119 6412 16212 6440
rect 16206 6400 16212 6412
rect 16264 6440 16270 6452
rect 16485 6443 16543 6449
rect 16485 6440 16497 6443
rect 16264 6412 16497 6440
rect 16264 6400 16270 6412
rect 16485 6409 16497 6412
rect 16531 6409 16543 6443
rect 16485 6403 16543 6409
rect 17865 6443 17923 6449
rect 17865 6409 17877 6443
rect 17911 6440 17923 6443
rect 18598 6440 18604 6452
rect 17911 6412 18604 6440
rect 17911 6409 17923 6412
rect 17865 6403 17923 6409
rect 18598 6400 18604 6412
rect 18656 6440 18662 6452
rect 19429 6443 19487 6449
rect 19429 6440 19441 6443
rect 18656 6412 19441 6440
rect 18656 6400 18662 6412
rect 19429 6409 19441 6412
rect 19475 6409 19487 6443
rect 19429 6403 19487 6409
rect 7834 6332 7840 6384
rect 7892 6372 7898 6384
rect 8294 6372 8300 6384
rect 7892 6344 8300 6372
rect 7892 6332 7898 6344
rect 8294 6332 8300 6344
rect 8352 6332 8358 6384
rect 9398 6372 9404 6384
rect 9359 6344 9404 6372
rect 9398 6332 9404 6344
rect 9456 6372 9462 6384
rect 10505 6375 10563 6381
rect 10505 6372 10517 6375
rect 9456 6344 10517 6372
rect 9456 6332 9462 6344
rect 10505 6341 10517 6344
rect 10551 6341 10563 6375
rect 10505 6335 10563 6341
rect 3329 6307 3387 6313
rect 3329 6273 3341 6307
rect 3375 6304 3387 6307
rect 7926 6304 7932 6316
rect 3375 6276 4154 6304
rect 7887 6276 7932 6304
rect 3375 6273 3387 6276
rect 3329 6267 3387 6273
rect 1464 6239 1522 6245
rect 1464 6205 1476 6239
rect 1510 6236 1522 6239
rect 2222 6236 2228 6248
rect 1510 6208 2228 6236
rect 1510 6205 1522 6208
rect 1464 6199 1522 6205
rect 2222 6196 2228 6208
rect 2280 6196 2286 6248
rect 3694 6236 3700 6248
rect 3655 6208 3700 6236
rect 3694 6196 3700 6208
rect 3752 6196 3758 6248
rect 3973 6239 4031 6245
rect 3973 6205 3985 6239
rect 4019 6205 4031 6239
rect 4126 6236 4154 6276
rect 7926 6264 7932 6276
rect 7984 6304 7990 6316
rect 9493 6307 9551 6313
rect 9493 6304 9505 6307
rect 7984 6276 9505 6304
rect 7984 6264 7990 6276
rect 9493 6273 9505 6276
rect 9539 6304 9551 6307
rect 9950 6304 9956 6316
rect 9539 6276 9956 6304
rect 9539 6273 9551 6276
rect 9493 6267 9551 6273
rect 9950 6264 9956 6276
rect 10008 6304 10014 6316
rect 10137 6307 10195 6313
rect 10137 6304 10149 6307
rect 10008 6276 10149 6304
rect 10008 6264 10014 6276
rect 10137 6273 10149 6276
rect 10183 6304 10195 6307
rect 10226 6304 10232 6316
rect 10183 6276 10232 6304
rect 10183 6273 10195 6276
rect 10137 6267 10195 6273
rect 10226 6264 10232 6276
rect 10284 6264 10290 6316
rect 4249 6239 4307 6245
rect 4249 6236 4261 6239
rect 4126 6208 4261 6236
rect 3973 6199 4031 6205
rect 4249 6205 4261 6208
rect 4295 6236 4307 6239
rect 5534 6236 5540 6248
rect 4295 6208 5540 6236
rect 4295 6205 4307 6208
rect 4249 6199 4307 6205
rect 2961 6171 3019 6177
rect 2961 6137 2973 6171
rect 3007 6168 3019 6171
rect 3007 6140 3832 6168
rect 3007 6137 3019 6140
rect 2961 6131 3019 6137
rect 106 6060 112 6112
rect 164 6100 170 6112
rect 1535 6103 1593 6109
rect 1535 6100 1547 6103
rect 164 6072 1547 6100
rect 164 6060 170 6072
rect 1535 6069 1547 6072
rect 1581 6069 1593 6103
rect 2314 6100 2320 6112
rect 2227 6072 2320 6100
rect 1535 6063 1593 6069
rect 2314 6060 2320 6072
rect 2372 6100 2378 6112
rect 3513 6103 3571 6109
rect 3513 6100 3525 6103
rect 2372 6072 3525 6100
rect 2372 6060 2378 6072
rect 3513 6069 3525 6072
rect 3559 6069 3571 6103
rect 3804 6100 3832 6140
rect 3988 6100 4016 6199
rect 5534 6196 5540 6208
rect 5592 6196 5598 6248
rect 7101 6239 7159 6245
rect 7101 6205 7113 6239
rect 7147 6236 7159 6239
rect 7469 6239 7527 6245
rect 7469 6236 7481 6239
rect 7147 6208 7481 6236
rect 7147 6205 7159 6208
rect 7101 6199 7159 6205
rect 7469 6205 7481 6208
rect 7515 6236 7527 6239
rect 7650 6236 7656 6248
rect 7515 6208 7656 6236
rect 7515 6205 7527 6208
rect 7469 6199 7527 6205
rect 7650 6196 7656 6208
rect 7708 6245 7714 6248
rect 7708 6239 7766 6245
rect 7708 6205 7720 6239
rect 7754 6236 7766 6239
rect 9033 6239 9091 6245
rect 9033 6236 9045 6239
rect 7754 6208 9045 6236
rect 7754 6205 7766 6208
rect 7708 6199 7766 6205
rect 9033 6205 9045 6208
rect 9079 6236 9091 6239
rect 9272 6239 9330 6245
rect 9272 6236 9284 6239
rect 9079 6208 9284 6236
rect 9079 6205 9091 6208
rect 9033 6199 9091 6205
rect 9272 6205 9284 6208
rect 9318 6236 9330 6239
rect 9766 6236 9772 6248
rect 9318 6208 9772 6236
rect 9318 6205 9330 6208
rect 9272 6199 9330 6205
rect 7708 6196 7714 6199
rect 9766 6196 9772 6208
rect 9824 6196 9830 6248
rect 10520 6236 10548 6335
rect 15930 6332 15936 6384
rect 15988 6372 15994 6384
rect 17037 6375 17095 6381
rect 17037 6372 17049 6375
rect 15988 6344 17049 6372
rect 15988 6332 15994 6344
rect 17037 6341 17049 6344
rect 17083 6372 17095 6375
rect 17954 6372 17960 6384
rect 17083 6344 17960 6372
rect 17083 6341 17095 6344
rect 17037 6335 17095 6341
rect 17954 6332 17960 6344
rect 18012 6332 18018 6384
rect 13446 6264 13452 6316
rect 13504 6304 13510 6316
rect 13725 6307 13783 6313
rect 13725 6304 13737 6307
rect 13504 6276 13737 6304
rect 13504 6264 13510 6276
rect 13725 6273 13737 6276
rect 13771 6273 13783 6307
rect 13725 6267 13783 6273
rect 13906 6264 13912 6316
rect 13964 6304 13970 6316
rect 14369 6307 14427 6313
rect 14369 6304 14381 6307
rect 13964 6276 14381 6304
rect 13964 6264 13970 6276
rect 14369 6273 14381 6276
rect 14415 6304 14427 6307
rect 16298 6304 16304 6316
rect 14415 6276 16304 6304
rect 14415 6273 14427 6276
rect 14369 6267 14427 6273
rect 16298 6264 16304 6276
rect 16356 6264 16362 6316
rect 16482 6264 16488 6316
rect 16540 6304 16546 6316
rect 17497 6307 17555 6313
rect 17497 6304 17509 6307
rect 16540 6276 17509 6304
rect 16540 6264 16546 6276
rect 17497 6273 17509 6276
rect 17543 6304 17555 6307
rect 19444 6304 19472 6403
rect 20162 6304 20168 6316
rect 17543 6276 18184 6304
rect 19444 6276 19748 6304
rect 20123 6276 20168 6304
rect 17543 6273 17555 6276
rect 17497 6267 17555 6273
rect 10781 6239 10839 6245
rect 10781 6236 10793 6239
rect 10520 6208 10793 6236
rect 10781 6205 10793 6208
rect 10827 6205 10839 6239
rect 10781 6199 10839 6205
rect 12526 6196 12532 6248
rect 12584 6236 12590 6248
rect 12656 6239 12714 6245
rect 12656 6236 12668 6239
rect 12584 6208 12668 6236
rect 12584 6196 12590 6208
rect 12656 6205 12668 6208
rect 12702 6236 12714 6239
rect 13081 6239 13139 6245
rect 13081 6236 13093 6239
rect 12702 6208 13093 6236
rect 12702 6205 12714 6208
rect 12656 6199 12714 6205
rect 13081 6205 13093 6208
rect 13127 6236 13139 6239
rect 13538 6236 13544 6248
rect 13127 6208 13544 6236
rect 13127 6205 13139 6208
rect 13081 6199 13139 6205
rect 13538 6196 13544 6208
rect 13596 6196 13602 6248
rect 14829 6239 14887 6245
rect 14829 6205 14841 6239
rect 14875 6236 14887 6239
rect 15289 6239 15347 6245
rect 15289 6236 15301 6239
rect 14875 6208 15301 6236
rect 14875 6205 14887 6208
rect 14829 6199 14887 6205
rect 15289 6205 15301 6208
rect 15335 6236 15347 6239
rect 15335 6208 16068 6236
rect 15335 6205 15347 6208
rect 15289 6199 15347 6205
rect 7561 6171 7619 6177
rect 7561 6137 7573 6171
rect 7607 6137 7619 6171
rect 7561 6131 7619 6137
rect 4798 6100 4804 6112
rect 3804 6072 4804 6100
rect 3513 6063 3571 6069
rect 4798 6060 4804 6072
rect 4856 6060 4862 6112
rect 5534 6100 5540 6112
rect 5495 6072 5540 6100
rect 5534 6060 5540 6072
rect 5592 6060 5598 6112
rect 5902 6100 5908 6112
rect 5863 6072 5908 6100
rect 5902 6060 5908 6072
rect 5960 6060 5966 6112
rect 6086 6060 6092 6112
rect 6144 6100 6150 6112
rect 6273 6103 6331 6109
rect 6273 6100 6285 6103
rect 6144 6072 6285 6100
rect 6144 6060 6150 6072
rect 6273 6069 6285 6072
rect 6319 6069 6331 6103
rect 6273 6063 6331 6069
rect 7466 6060 7472 6112
rect 7524 6100 7530 6112
rect 7576 6100 7604 6131
rect 8018 6128 8024 6180
rect 8076 6168 8082 6180
rect 9122 6168 9128 6180
rect 8076 6140 9128 6168
rect 8076 6128 8082 6140
rect 9122 6128 9128 6140
rect 9180 6128 9186 6180
rect 12759 6171 12817 6177
rect 12759 6137 12771 6171
rect 12805 6168 12817 6171
rect 13262 6168 13268 6180
rect 12805 6140 13268 6168
rect 12805 6137 12817 6140
rect 12759 6131 12817 6137
rect 13262 6128 13268 6140
rect 13320 6128 13326 6180
rect 13814 6128 13820 6180
rect 13872 6168 13878 6180
rect 15610 6171 15668 6177
rect 15610 6168 15622 6171
rect 13872 6140 13917 6168
rect 15120 6140 15622 6168
rect 13872 6128 13878 6140
rect 7524 6072 7604 6100
rect 7524 6060 7530 6072
rect 8294 6060 8300 6112
rect 8352 6100 8358 6112
rect 8573 6103 8631 6109
rect 8573 6100 8585 6103
rect 8352 6072 8585 6100
rect 8352 6060 8358 6072
rect 8573 6069 8585 6072
rect 8619 6069 8631 6103
rect 10962 6100 10968 6112
rect 10923 6072 10968 6100
rect 8573 6063 8631 6069
rect 10962 6060 10968 6072
rect 11020 6060 11026 6112
rect 12253 6103 12311 6109
rect 12253 6069 12265 6103
rect 12299 6100 12311 6103
rect 12342 6100 12348 6112
rect 12299 6072 12348 6100
rect 12299 6069 12311 6072
rect 12253 6063 12311 6069
rect 12342 6060 12348 6072
rect 12400 6060 12406 6112
rect 13538 6100 13544 6112
rect 13499 6072 13544 6100
rect 13538 6060 13544 6072
rect 13596 6100 13602 6112
rect 15120 6109 15148 6140
rect 15610 6137 15622 6140
rect 15656 6168 15668 6171
rect 15838 6168 15844 6180
rect 15656 6140 15844 6168
rect 15656 6137 15668 6140
rect 15610 6131 15668 6137
rect 15838 6128 15844 6140
rect 15896 6128 15902 6180
rect 16040 6168 16068 6208
rect 16850 6196 16856 6248
rect 16908 6236 16914 6248
rect 17862 6236 17868 6248
rect 16908 6208 17868 6236
rect 16908 6196 16914 6208
rect 17862 6196 17868 6208
rect 17920 6236 17926 6248
rect 18049 6239 18107 6245
rect 18049 6236 18061 6239
rect 17920 6208 18061 6236
rect 17920 6196 17926 6208
rect 18049 6205 18061 6208
rect 18095 6205 18107 6239
rect 18156 6236 18184 6276
rect 18509 6239 18567 6245
rect 18509 6236 18521 6239
rect 18156 6208 18521 6236
rect 18049 6199 18107 6205
rect 18509 6205 18521 6208
rect 18555 6205 18567 6239
rect 19610 6236 19616 6248
rect 19571 6208 19616 6236
rect 18509 6199 18567 6205
rect 19610 6196 19616 6208
rect 19668 6196 19674 6248
rect 19720 6236 19748 6276
rect 20162 6264 20168 6276
rect 20220 6264 20226 6316
rect 20073 6239 20131 6245
rect 20073 6236 20085 6239
rect 19720 6208 20085 6236
rect 20073 6205 20085 6208
rect 20119 6205 20131 6239
rect 20073 6199 20131 6205
rect 16040 6140 18092 6168
rect 15105 6103 15163 6109
rect 15105 6100 15117 6103
rect 13596 6072 15117 6100
rect 13596 6060 13602 6072
rect 15105 6069 15117 6072
rect 15151 6069 15163 6103
rect 18064 6100 18092 6140
rect 18141 6103 18199 6109
rect 18141 6100 18153 6103
rect 18064 6072 18153 6100
rect 15105 6063 15163 6069
rect 18141 6069 18153 6072
rect 18187 6069 18199 6103
rect 18141 6063 18199 6069
rect 1104 6010 22816 6032
rect 1104 5958 8982 6010
rect 9034 5958 9046 6010
rect 9098 5958 9110 6010
rect 9162 5958 9174 6010
rect 9226 5958 16982 6010
rect 17034 5958 17046 6010
rect 17098 5958 17110 6010
rect 17162 5958 17174 6010
rect 17226 5958 22816 6010
rect 1104 5936 22816 5958
rect 3234 5856 3240 5908
rect 3292 5896 3298 5908
rect 4157 5899 4215 5905
rect 4157 5896 4169 5899
rect 3292 5868 4169 5896
rect 3292 5856 3298 5868
rect 4157 5865 4169 5868
rect 4203 5865 4215 5899
rect 4157 5859 4215 5865
rect 4724 5868 4936 5896
rect 1946 5828 1952 5840
rect 1907 5800 1952 5828
rect 1946 5788 1952 5800
rect 2004 5788 2010 5840
rect 3513 5763 3571 5769
rect 3513 5729 3525 5763
rect 3559 5760 3571 5763
rect 3694 5760 3700 5772
rect 3559 5732 3700 5760
rect 3559 5729 3571 5732
rect 3513 5723 3571 5729
rect 3694 5720 3700 5732
rect 3752 5760 3758 5772
rect 4154 5760 4160 5772
rect 3752 5732 4160 5760
rect 3752 5720 3758 5732
rect 4154 5720 4160 5732
rect 4212 5760 4218 5772
rect 4341 5763 4399 5769
rect 4341 5760 4353 5763
rect 4212 5732 4353 5760
rect 4212 5720 4218 5732
rect 4341 5729 4353 5732
rect 4387 5760 4399 5763
rect 4724 5760 4752 5868
rect 4908 5828 4936 5868
rect 4982 5856 4988 5908
rect 5040 5896 5046 5908
rect 7837 5899 7895 5905
rect 7837 5896 7849 5899
rect 5040 5868 7849 5896
rect 5040 5856 5046 5868
rect 7837 5865 7849 5868
rect 7883 5896 7895 5899
rect 8018 5896 8024 5908
rect 7883 5868 8024 5896
rect 7883 5865 7895 5868
rect 7837 5859 7895 5865
rect 8018 5856 8024 5868
rect 8076 5856 8082 5908
rect 9490 5856 9496 5908
rect 9548 5896 9554 5908
rect 11057 5899 11115 5905
rect 11057 5896 11069 5899
rect 9548 5868 11069 5896
rect 9548 5856 9554 5868
rect 11057 5865 11069 5868
rect 11103 5865 11115 5899
rect 11057 5859 11115 5865
rect 13446 5856 13452 5908
rect 13504 5896 13510 5908
rect 14185 5899 14243 5905
rect 14185 5896 14197 5899
rect 13504 5868 14197 5896
rect 13504 5856 13510 5868
rect 14185 5865 14197 5868
rect 14231 5865 14243 5899
rect 14185 5859 14243 5865
rect 15841 5899 15899 5905
rect 15841 5865 15853 5899
rect 15887 5896 15899 5899
rect 16114 5896 16120 5908
rect 15887 5868 16120 5896
rect 15887 5865 15899 5868
rect 15841 5859 15899 5865
rect 16114 5856 16120 5868
rect 16172 5856 16178 5908
rect 17862 5856 17868 5908
rect 17920 5896 17926 5908
rect 18509 5899 18567 5905
rect 18509 5896 18521 5899
rect 17920 5868 18521 5896
rect 17920 5856 17926 5868
rect 18509 5865 18521 5868
rect 18555 5865 18567 5899
rect 18509 5859 18567 5865
rect 10410 5828 10416 5840
rect 4908 5800 10416 5828
rect 10410 5788 10416 5800
rect 10468 5788 10474 5840
rect 12342 5828 12348 5840
rect 12303 5800 12348 5828
rect 12342 5788 12348 5800
rect 12400 5788 12406 5840
rect 13354 5828 13360 5840
rect 13315 5800 13360 5828
rect 13354 5788 13360 5800
rect 13412 5788 13418 5840
rect 13906 5828 13912 5840
rect 13867 5800 13912 5828
rect 13906 5788 13912 5800
rect 13964 5788 13970 5840
rect 17678 5828 17684 5840
rect 17639 5800 17684 5828
rect 17678 5788 17684 5800
rect 17736 5788 17742 5840
rect 4387 5732 4752 5760
rect 4893 5763 4951 5769
rect 4387 5729 4399 5732
rect 4341 5723 4399 5729
rect 4893 5729 4905 5763
rect 4939 5760 4951 5763
rect 5537 5763 5595 5769
rect 5537 5760 5549 5763
rect 4939 5732 5549 5760
rect 4939 5729 4951 5732
rect 4893 5723 4951 5729
rect 5537 5729 5549 5732
rect 5583 5760 5595 5763
rect 5994 5760 6000 5772
rect 5583 5732 6000 5760
rect 5583 5729 5595 5732
rect 5537 5723 5595 5729
rect 5994 5720 6000 5732
rect 6052 5720 6058 5772
rect 6086 5720 6092 5772
rect 6144 5760 6150 5772
rect 6273 5763 6331 5769
rect 6144 5732 6189 5760
rect 6144 5720 6150 5732
rect 6273 5729 6285 5763
rect 6319 5729 6331 5763
rect 6730 5760 6736 5772
rect 6691 5732 6736 5760
rect 6273 5723 6331 5729
rect 1673 5695 1731 5701
rect 1673 5661 1685 5695
rect 1719 5692 1731 5695
rect 1857 5695 1915 5701
rect 1857 5692 1869 5695
rect 1719 5664 1869 5692
rect 1719 5661 1731 5664
rect 1673 5655 1731 5661
rect 1857 5661 1869 5664
rect 1903 5692 1915 5695
rect 2130 5692 2136 5704
rect 1903 5664 2136 5692
rect 1903 5661 1915 5664
rect 1857 5655 1915 5661
rect 2130 5652 2136 5664
rect 2188 5652 2194 5704
rect 2222 5652 2228 5704
rect 2280 5692 2286 5704
rect 2777 5695 2835 5701
rect 2777 5692 2789 5695
rect 2280 5664 2789 5692
rect 2280 5652 2286 5664
rect 2777 5661 2789 5664
rect 2823 5661 2835 5695
rect 4798 5692 4804 5704
rect 4759 5664 4804 5692
rect 2777 5655 2835 5661
rect 4798 5652 4804 5664
rect 4856 5652 4862 5704
rect 6288 5692 6316 5723
rect 6730 5720 6736 5732
rect 6788 5720 6794 5772
rect 7558 5760 7564 5772
rect 7519 5732 7564 5760
rect 7558 5720 7564 5732
rect 7616 5720 7622 5772
rect 7745 5763 7803 5769
rect 7745 5729 7757 5763
rect 7791 5760 7803 5763
rect 8110 5760 8116 5772
rect 7791 5732 8116 5760
rect 7791 5729 7803 5732
rect 7745 5723 7803 5729
rect 8110 5720 8116 5732
rect 8168 5720 8174 5772
rect 9677 5763 9735 5769
rect 9677 5729 9689 5763
rect 9723 5760 9735 5763
rect 9766 5760 9772 5772
rect 9723 5732 9772 5760
rect 9723 5729 9735 5732
rect 9677 5723 9735 5729
rect 9766 5720 9772 5732
rect 9824 5720 9830 5772
rect 9950 5760 9956 5772
rect 9911 5732 9956 5760
rect 9950 5720 9956 5732
rect 10008 5760 10014 5772
rect 10689 5763 10747 5769
rect 10689 5760 10701 5763
rect 10008 5732 10701 5760
rect 10008 5720 10014 5732
rect 10689 5729 10701 5732
rect 10735 5729 10747 5763
rect 10689 5723 10747 5729
rect 11609 5763 11667 5769
rect 11609 5729 11621 5763
rect 11655 5729 11667 5763
rect 11609 5723 11667 5729
rect 5828 5664 6316 5692
rect 5626 5516 5632 5568
rect 5684 5556 5690 5568
rect 5828 5565 5856 5664
rect 10318 5652 10324 5704
rect 10376 5692 10382 5704
rect 11425 5695 11483 5701
rect 11425 5692 11437 5695
rect 10376 5664 11437 5692
rect 10376 5652 10382 5664
rect 11425 5661 11437 5664
rect 11471 5692 11483 5695
rect 11624 5692 11652 5723
rect 11974 5720 11980 5772
rect 12032 5760 12038 5772
rect 12069 5763 12127 5769
rect 12069 5760 12081 5763
rect 12032 5732 12081 5760
rect 12032 5720 12038 5732
rect 12069 5729 12081 5732
rect 12115 5729 12127 5763
rect 15930 5760 15936 5772
rect 15891 5732 15936 5760
rect 12069 5723 12127 5729
rect 15930 5720 15936 5732
rect 15988 5720 15994 5772
rect 16482 5760 16488 5772
rect 16443 5732 16488 5760
rect 16482 5720 16488 5732
rect 16540 5720 16546 5772
rect 11471 5664 11652 5692
rect 11471 5661 11483 5664
rect 11425 5655 11483 5661
rect 12802 5652 12808 5704
rect 12860 5692 12866 5704
rect 13265 5695 13323 5701
rect 13265 5692 13277 5695
rect 12860 5664 13277 5692
rect 12860 5652 12866 5664
rect 13265 5661 13277 5664
rect 13311 5661 13323 5695
rect 16666 5692 16672 5704
rect 16627 5664 16672 5692
rect 13265 5655 13323 5661
rect 16666 5652 16672 5664
rect 16724 5652 16730 5704
rect 17586 5692 17592 5704
rect 17547 5664 17592 5692
rect 17586 5652 17592 5664
rect 17644 5652 17650 5704
rect 17862 5692 17868 5704
rect 17823 5664 17868 5692
rect 17862 5652 17868 5664
rect 17920 5652 17926 5704
rect 19334 5692 19340 5704
rect 19295 5664 19340 5692
rect 19334 5652 19340 5664
rect 19392 5652 19398 5704
rect 9769 5627 9827 5633
rect 9769 5593 9781 5627
rect 9815 5624 9827 5627
rect 10962 5624 10968 5636
rect 9815 5596 10968 5624
rect 9815 5593 9827 5596
rect 9769 5587 9827 5593
rect 10962 5584 10968 5596
rect 11020 5584 11026 5636
rect 5813 5559 5871 5565
rect 5813 5556 5825 5559
rect 5684 5528 5825 5556
rect 5684 5516 5690 5528
rect 5813 5525 5825 5528
rect 5859 5525 5871 5559
rect 7006 5556 7012 5568
rect 6967 5528 7012 5556
rect 5813 5519 5871 5525
rect 7006 5516 7012 5528
rect 7064 5516 7070 5568
rect 7466 5556 7472 5568
rect 7427 5528 7472 5556
rect 7466 5516 7472 5528
rect 7524 5516 7530 5568
rect 8294 5516 8300 5568
rect 8352 5556 8358 5568
rect 8389 5559 8447 5565
rect 8389 5556 8401 5559
rect 8352 5528 8401 5556
rect 8352 5516 8358 5528
rect 8389 5525 8401 5528
rect 8435 5556 8447 5559
rect 9125 5559 9183 5565
rect 9125 5556 9137 5559
rect 8435 5528 9137 5556
rect 8435 5525 8447 5528
rect 8389 5519 8447 5525
rect 9125 5525 9137 5528
rect 9171 5556 9183 5559
rect 9306 5556 9312 5568
rect 9171 5528 9312 5556
rect 9171 5525 9183 5528
rect 9125 5519 9183 5525
rect 9306 5516 9312 5528
rect 9364 5516 9370 5568
rect 12618 5556 12624 5568
rect 12579 5528 12624 5556
rect 12618 5516 12624 5528
rect 12676 5516 12682 5568
rect 16942 5556 16948 5568
rect 16903 5528 16948 5556
rect 16942 5516 16948 5528
rect 17000 5516 17006 5568
rect 1104 5466 22816 5488
rect 1104 5414 4982 5466
rect 5034 5414 5046 5466
rect 5098 5414 5110 5466
rect 5162 5414 5174 5466
rect 5226 5414 12982 5466
rect 13034 5414 13046 5466
rect 13098 5414 13110 5466
rect 13162 5414 13174 5466
rect 13226 5414 20982 5466
rect 21034 5414 21046 5466
rect 21098 5414 21110 5466
rect 21162 5414 21174 5466
rect 21226 5414 22816 5466
rect 1104 5392 22816 5414
rect 1946 5312 1952 5364
rect 2004 5352 2010 5364
rect 2406 5352 2412 5364
rect 2004 5324 2412 5352
rect 2004 5312 2010 5324
rect 2406 5312 2412 5324
rect 2464 5352 2470 5364
rect 2869 5355 2927 5361
rect 2869 5352 2881 5355
rect 2464 5324 2881 5352
rect 2464 5312 2470 5324
rect 2869 5321 2881 5324
rect 2915 5321 2927 5355
rect 3234 5352 3240 5364
rect 3195 5324 3240 5352
rect 2869 5315 2927 5321
rect 3234 5312 3240 5324
rect 3292 5312 3298 5364
rect 4154 5352 4160 5364
rect 4115 5324 4160 5352
rect 4154 5312 4160 5324
rect 4212 5312 4218 5364
rect 4525 5355 4583 5361
rect 4525 5321 4537 5355
rect 4571 5352 4583 5355
rect 4798 5352 4804 5364
rect 4571 5324 4804 5352
rect 4571 5321 4583 5324
rect 4525 5315 4583 5321
rect 4798 5312 4804 5324
rect 4856 5312 4862 5364
rect 6086 5352 6092 5364
rect 5276 5324 6092 5352
rect 1857 5287 1915 5293
rect 1857 5253 1869 5287
rect 1903 5284 1915 5287
rect 2038 5284 2044 5296
rect 1903 5256 2044 5284
rect 1903 5253 1915 5256
rect 1857 5247 1915 5253
rect 2038 5244 2044 5256
rect 2096 5244 2102 5296
rect 1949 5219 2007 5225
rect 1949 5185 1961 5219
rect 1995 5216 2007 5219
rect 3252 5216 3280 5312
rect 5276 5296 5304 5324
rect 6086 5312 6092 5324
rect 6144 5352 6150 5364
rect 6181 5355 6239 5361
rect 6181 5352 6193 5355
rect 6144 5324 6193 5352
rect 6144 5312 6150 5324
rect 6181 5321 6193 5324
rect 6227 5321 6239 5355
rect 6181 5315 6239 5321
rect 7006 5312 7012 5364
rect 7064 5352 7070 5364
rect 8573 5355 8631 5361
rect 8573 5352 8585 5355
rect 7064 5324 8585 5352
rect 7064 5312 7070 5324
rect 8573 5321 8585 5324
rect 8619 5352 8631 5355
rect 8941 5355 8999 5361
rect 8941 5352 8953 5355
rect 8619 5324 8953 5352
rect 8619 5321 8631 5324
rect 8573 5315 8631 5321
rect 8941 5321 8953 5324
rect 8987 5321 8999 5355
rect 9306 5352 9312 5364
rect 9267 5324 9312 5352
rect 8941 5315 8999 5321
rect 5258 5284 5264 5296
rect 5171 5256 5264 5284
rect 5258 5244 5264 5256
rect 5316 5244 5322 5296
rect 5994 5216 6000 5228
rect 1995 5188 3280 5216
rect 5184 5188 6000 5216
rect 1995 5185 2007 5188
rect 1949 5179 2007 5185
rect 4798 5148 4804 5160
rect 4126 5120 4804 5148
rect 2038 5040 2044 5092
rect 2096 5080 2102 5092
rect 2270 5083 2328 5089
rect 2270 5080 2282 5083
rect 2096 5052 2282 5080
rect 2096 5040 2102 5052
rect 2270 5049 2282 5052
rect 2316 5080 2328 5083
rect 2866 5080 2872 5092
rect 2316 5052 2872 5080
rect 2316 5049 2328 5052
rect 2270 5043 2328 5049
rect 2866 5040 2872 5052
rect 2924 5040 2930 5092
rect 3789 5083 3847 5089
rect 3789 5049 3801 5083
rect 3835 5080 3847 5083
rect 4126 5080 4154 5120
rect 4798 5108 4804 5120
rect 4856 5148 4862 5160
rect 5184 5157 5212 5188
rect 5994 5176 6000 5188
rect 6052 5176 6058 5228
rect 8956 5216 8984 5315
rect 9306 5312 9312 5324
rect 9364 5352 9370 5364
rect 10962 5352 10968 5364
rect 9364 5324 9628 5352
rect 10923 5324 10968 5352
rect 9364 5312 9370 5324
rect 9600 5293 9628 5324
rect 10962 5312 10968 5324
rect 11020 5312 11026 5364
rect 11609 5355 11667 5361
rect 11609 5321 11621 5355
rect 11655 5352 11667 5355
rect 11698 5352 11704 5364
rect 11655 5324 11704 5352
rect 11655 5321 11667 5324
rect 11609 5315 11667 5321
rect 11698 5312 11704 5324
rect 11756 5312 11762 5364
rect 13354 5312 13360 5364
rect 13412 5352 13418 5364
rect 13449 5355 13507 5361
rect 13449 5352 13461 5355
rect 13412 5324 13461 5352
rect 13412 5312 13418 5324
rect 13449 5321 13461 5324
rect 13495 5352 13507 5355
rect 13725 5355 13783 5361
rect 13725 5352 13737 5355
rect 13495 5324 13737 5352
rect 13495 5321 13507 5324
rect 13449 5315 13507 5321
rect 13725 5321 13737 5324
rect 13771 5352 13783 5355
rect 14093 5355 14151 5361
rect 14093 5352 14105 5355
rect 13771 5324 14105 5352
rect 13771 5321 13783 5324
rect 13725 5315 13783 5321
rect 14093 5321 14105 5324
rect 14139 5352 14151 5355
rect 14458 5352 14464 5364
rect 14139 5324 14464 5352
rect 14139 5321 14151 5324
rect 14093 5315 14151 5321
rect 14458 5312 14464 5324
rect 14516 5312 14522 5364
rect 15657 5355 15715 5361
rect 15657 5321 15669 5355
rect 15703 5352 15715 5355
rect 15930 5352 15936 5364
rect 15703 5324 15936 5352
rect 15703 5321 15715 5324
rect 15657 5315 15715 5321
rect 15930 5312 15936 5324
rect 15988 5312 15994 5364
rect 16025 5355 16083 5361
rect 16025 5321 16037 5355
rect 16071 5352 16083 5355
rect 16482 5352 16488 5364
rect 16071 5324 16488 5352
rect 16071 5321 16083 5324
rect 16025 5315 16083 5321
rect 16482 5312 16488 5324
rect 16540 5312 16546 5364
rect 19334 5312 19340 5364
rect 19392 5352 19398 5364
rect 19613 5355 19671 5361
rect 19613 5352 19625 5355
rect 19392 5324 19625 5352
rect 19392 5312 19398 5324
rect 19613 5321 19625 5324
rect 19659 5321 19671 5355
rect 19613 5315 19671 5321
rect 9585 5287 9643 5293
rect 9585 5253 9597 5287
rect 9631 5253 9643 5287
rect 9585 5247 9643 5253
rect 9950 5244 9956 5296
rect 10008 5284 10014 5296
rect 12161 5287 12219 5293
rect 12161 5284 12173 5287
rect 10008 5256 12173 5284
rect 10008 5244 10014 5256
rect 12161 5253 12173 5256
rect 12207 5284 12219 5287
rect 12437 5287 12495 5293
rect 12437 5284 12449 5287
rect 12207 5256 12449 5284
rect 12207 5253 12219 5256
rect 12161 5247 12219 5253
rect 12437 5253 12449 5256
rect 12483 5253 12495 5287
rect 14918 5284 14924 5296
rect 14879 5256 14924 5284
rect 12437 5247 12495 5253
rect 14918 5244 14924 5256
rect 14976 5284 14982 5296
rect 16942 5284 16948 5296
rect 14976 5256 16948 5284
rect 14976 5244 14982 5256
rect 10226 5216 10232 5228
rect 8956 5188 9812 5216
rect 10139 5188 10232 5216
rect 5169 5151 5227 5157
rect 5169 5148 5181 5151
rect 4856 5120 5181 5148
rect 4856 5108 4862 5120
rect 5169 5117 5181 5120
rect 5215 5117 5227 5151
rect 5169 5111 5227 5117
rect 5445 5151 5503 5157
rect 5445 5117 5457 5151
rect 5491 5117 5503 5151
rect 5445 5111 5503 5117
rect 3835 5052 4154 5080
rect 5460 5080 5488 5111
rect 5626 5108 5632 5160
rect 5684 5148 5690 5160
rect 6825 5151 6883 5157
rect 6825 5148 6837 5151
rect 5684 5120 6837 5148
rect 5684 5108 5690 5120
rect 6825 5117 6837 5120
rect 6871 5117 6883 5151
rect 6825 5111 6883 5117
rect 7009 5151 7067 5157
rect 7009 5117 7021 5151
rect 7055 5117 7067 5151
rect 9490 5148 9496 5160
rect 9451 5120 9496 5148
rect 7009 5111 7067 5117
rect 5902 5080 5908 5092
rect 5460 5052 5908 5080
rect 3835 5049 3847 5052
rect 3789 5043 3847 5049
rect 4614 4972 4620 5024
rect 4672 5012 4678 5024
rect 4985 5015 5043 5021
rect 4985 5012 4997 5015
rect 4672 4984 4997 5012
rect 4672 4972 4678 4984
rect 4985 4981 4997 4984
rect 5031 5012 5043 5015
rect 5460 5012 5488 5052
rect 5902 5040 5908 5052
rect 5960 5080 5966 5092
rect 6549 5083 6607 5089
rect 6549 5080 6561 5083
rect 5960 5052 6561 5080
rect 5960 5040 5966 5052
rect 6549 5049 6561 5052
rect 6595 5049 6607 5083
rect 6549 5043 6607 5049
rect 5031 4984 5488 5012
rect 5629 5015 5687 5021
rect 5031 4981 5043 4984
rect 4985 4975 5043 4981
rect 5629 4981 5641 5015
rect 5675 5012 5687 5015
rect 5810 5012 5816 5024
rect 5675 4984 5816 5012
rect 5675 4981 5687 4984
rect 5629 4975 5687 4981
rect 5810 4972 5816 4984
rect 5868 4972 5874 5024
rect 6564 5012 6592 5043
rect 7024 5012 7052 5111
rect 9490 5108 9496 5120
rect 9548 5108 9554 5160
rect 9784 5157 9812 5188
rect 10226 5176 10232 5188
rect 10284 5216 10290 5228
rect 12529 5219 12587 5225
rect 10284 5188 11284 5216
rect 10284 5176 10290 5188
rect 9769 5151 9827 5157
rect 9769 5117 9781 5151
rect 9815 5117 9827 5151
rect 9769 5111 9827 5117
rect 11124 5151 11182 5157
rect 11124 5117 11136 5151
rect 11170 5117 11182 5151
rect 11256 5148 11284 5188
rect 12529 5185 12541 5219
rect 12575 5216 12587 5219
rect 12618 5216 12624 5228
rect 12575 5188 12624 5216
rect 12575 5185 12587 5188
rect 12529 5179 12587 5185
rect 12618 5176 12624 5188
rect 12676 5176 12682 5228
rect 13262 5176 13268 5228
rect 13320 5216 13326 5228
rect 14366 5216 14372 5228
rect 13320 5188 14372 5216
rect 13320 5176 13326 5188
rect 14366 5176 14372 5188
rect 14424 5176 14430 5228
rect 16316 5225 16344 5256
rect 16942 5244 16948 5256
rect 17000 5244 17006 5296
rect 17497 5287 17555 5293
rect 17497 5253 17509 5287
rect 17543 5284 17555 5287
rect 17678 5284 17684 5296
rect 17543 5256 17684 5284
rect 17543 5253 17555 5256
rect 17497 5247 17555 5253
rect 17678 5244 17684 5256
rect 17736 5284 17742 5296
rect 18969 5287 19027 5293
rect 18969 5284 18981 5287
rect 17736 5256 18981 5284
rect 17736 5244 17742 5256
rect 18969 5253 18981 5256
rect 19015 5253 19027 5287
rect 18969 5247 19027 5253
rect 16301 5219 16359 5225
rect 16301 5185 16313 5219
rect 16347 5185 16359 5219
rect 16301 5179 16359 5185
rect 16666 5176 16672 5228
rect 16724 5216 16730 5228
rect 18046 5216 18052 5228
rect 16724 5188 18052 5216
rect 16724 5176 16730 5188
rect 18046 5176 18052 5188
rect 18104 5176 18110 5228
rect 19628 5216 19656 5315
rect 19889 5219 19947 5225
rect 19889 5216 19901 5219
rect 19628 5188 19901 5216
rect 19889 5185 19901 5188
rect 19935 5185 19947 5219
rect 19889 5179 19947 5185
rect 13446 5148 13452 5160
rect 11256 5120 13452 5148
rect 11124 5111 11182 5117
rect 7558 5040 7564 5092
rect 7616 5080 7622 5092
rect 8205 5083 8263 5089
rect 8205 5080 8217 5083
rect 7616 5052 8217 5080
rect 7616 5040 7622 5052
rect 8205 5049 8217 5052
rect 8251 5049 8263 5083
rect 10505 5083 10563 5089
rect 10505 5080 10517 5083
rect 8205 5043 8263 5049
rect 9876 5052 10517 5080
rect 7190 5012 7196 5024
rect 6564 4984 7196 5012
rect 7190 4972 7196 4984
rect 7248 4972 7254 5024
rect 7929 5015 7987 5021
rect 7929 4981 7941 5015
rect 7975 5012 7987 5015
rect 8110 5012 8116 5024
rect 7975 4984 8116 5012
rect 7975 4981 7987 4984
rect 7929 4975 7987 4981
rect 8110 4972 8116 4984
rect 8168 4972 8174 5024
rect 9766 4972 9772 5024
rect 9824 5012 9830 5024
rect 9876 5012 9904 5052
rect 10505 5049 10517 5052
rect 10551 5049 10563 5083
rect 11139 5080 11167 5111
rect 13446 5108 13452 5120
rect 13504 5108 13510 5160
rect 16945 5151 17003 5157
rect 16945 5117 16957 5151
rect 16991 5148 17003 5151
rect 17862 5148 17868 5160
rect 16991 5120 17868 5148
rect 16991 5117 17003 5120
rect 16945 5111 17003 5117
rect 17862 5108 17868 5120
rect 17920 5148 17926 5160
rect 17920 5120 19334 5148
rect 17920 5108 17926 5120
rect 11698 5080 11704 5092
rect 11139 5052 11704 5080
rect 10505 5043 10563 5049
rect 11698 5040 11704 5052
rect 11756 5040 11762 5092
rect 12437 5083 12495 5089
rect 12437 5049 12449 5083
rect 12483 5080 12495 5083
rect 12850 5083 12908 5089
rect 12850 5080 12862 5083
rect 12483 5052 12862 5080
rect 12483 5049 12495 5052
rect 12437 5043 12495 5049
rect 12850 5049 12862 5052
rect 12896 5080 12908 5083
rect 13538 5080 13544 5092
rect 12896 5052 13544 5080
rect 12896 5049 12908 5052
rect 12850 5043 12908 5049
rect 13538 5040 13544 5052
rect 13596 5040 13602 5092
rect 14458 5040 14464 5092
rect 14516 5080 14522 5092
rect 14516 5052 14561 5080
rect 14516 5040 14522 5052
rect 16390 5040 16396 5092
rect 16448 5080 16454 5092
rect 18370 5083 18428 5089
rect 16448 5052 16493 5080
rect 16448 5040 16454 5052
rect 18370 5049 18382 5083
rect 18416 5049 18428 5083
rect 18370 5043 18428 5049
rect 9824 4984 9904 5012
rect 9824 4972 9830 4984
rect 11054 4972 11060 5024
rect 11112 5012 11118 5024
rect 11195 5015 11253 5021
rect 11195 5012 11207 5015
rect 11112 4984 11207 5012
rect 11112 4972 11118 4984
rect 11195 4981 11207 4984
rect 11241 4981 11253 5015
rect 11195 4975 11253 4981
rect 15838 4972 15844 5024
rect 15896 5012 15902 5024
rect 17773 5015 17831 5021
rect 17773 5012 17785 5015
rect 15896 4984 17785 5012
rect 15896 4972 15902 4984
rect 17773 4981 17785 4984
rect 17819 5012 17831 5015
rect 18385 5012 18413 5043
rect 18966 5012 18972 5024
rect 17819 4984 18972 5012
rect 17819 4981 17831 4984
rect 17773 4975 17831 4981
rect 18966 4972 18972 4984
rect 19024 4972 19030 5024
rect 19306 5012 19334 5120
rect 19978 5080 19984 5092
rect 19939 5052 19984 5080
rect 19978 5040 19984 5052
rect 20036 5040 20042 5092
rect 20533 5083 20591 5089
rect 20533 5049 20545 5083
rect 20579 5049 20591 5083
rect 20533 5043 20591 5049
rect 19426 5012 19432 5024
rect 19306 4984 19432 5012
rect 19426 4972 19432 4984
rect 19484 5012 19490 5024
rect 20548 5012 20576 5043
rect 19484 4984 20576 5012
rect 19484 4972 19490 4984
rect 1104 4922 22816 4944
rect 1104 4870 8982 4922
rect 9034 4870 9046 4922
rect 9098 4870 9110 4922
rect 9162 4870 9174 4922
rect 9226 4870 16982 4922
rect 17034 4870 17046 4922
rect 17098 4870 17110 4922
rect 17162 4870 17174 4922
rect 17226 4870 22816 4922
rect 1104 4848 22816 4870
rect 2406 4808 2412 4820
rect 2367 4780 2412 4808
rect 2406 4768 2412 4780
rect 2464 4768 2470 4820
rect 5258 4808 5264 4820
rect 5219 4780 5264 4808
rect 5258 4768 5264 4780
rect 5316 4768 5322 4820
rect 8110 4808 8116 4820
rect 5787 4780 8116 4808
rect 1578 4740 1584 4752
rect 1539 4712 1584 4740
rect 1578 4700 1584 4712
rect 1636 4700 1642 4752
rect 2133 4743 2191 4749
rect 2133 4709 2145 4743
rect 2179 4740 2191 4743
rect 2222 4740 2228 4752
rect 2179 4712 2228 4740
rect 2179 4709 2191 4712
rect 2133 4703 2191 4709
rect 2222 4700 2228 4712
rect 2280 4700 2286 4752
rect 5787 4740 5815 4780
rect 8110 4768 8116 4780
rect 8168 4768 8174 4820
rect 9490 4808 9496 4820
rect 9451 4780 9496 4808
rect 9490 4768 9496 4780
rect 9548 4808 9554 4820
rect 9548 4780 9720 4808
rect 9548 4768 9554 4780
rect 4356 4712 5815 4740
rect 3970 4632 3976 4684
rect 4028 4672 4034 4684
rect 4356 4681 4384 4712
rect 5994 4700 6000 4752
rect 6052 4740 6058 4752
rect 9692 4749 9720 4780
rect 12802 4768 12808 4820
rect 12860 4808 12866 4820
rect 13173 4811 13231 4817
rect 13173 4808 13185 4811
rect 12860 4780 13185 4808
rect 12860 4768 12866 4780
rect 13173 4777 13185 4780
rect 13219 4777 13231 4811
rect 14366 4808 14372 4820
rect 14327 4780 14372 4808
rect 13173 4771 13231 4777
rect 14366 4768 14372 4780
rect 14424 4768 14430 4820
rect 15838 4808 15844 4820
rect 15799 4780 15844 4808
rect 15838 4768 15844 4780
rect 15896 4768 15902 4820
rect 16390 4808 16396 4820
rect 16351 4780 16396 4808
rect 16390 4768 16396 4780
rect 16448 4808 16454 4820
rect 16669 4811 16727 4817
rect 16669 4808 16681 4811
rect 16448 4780 16681 4808
rect 16448 4768 16454 4780
rect 16669 4777 16681 4780
rect 16715 4777 16727 4811
rect 17586 4808 17592 4820
rect 17547 4780 17592 4808
rect 16669 4771 16727 4777
rect 17586 4768 17592 4780
rect 17644 4768 17650 4820
rect 18046 4808 18052 4820
rect 18007 4780 18052 4808
rect 18046 4768 18052 4780
rect 18104 4768 18110 4820
rect 18966 4808 18972 4820
rect 18927 4780 18972 4808
rect 18966 4768 18972 4780
rect 19024 4768 19030 4820
rect 19521 4811 19579 4817
rect 19521 4777 19533 4811
rect 19567 4808 19579 4811
rect 19889 4811 19947 4817
rect 19889 4808 19901 4811
rect 19567 4780 19901 4808
rect 19567 4777 19579 4780
rect 19521 4771 19579 4777
rect 19889 4777 19901 4780
rect 19935 4808 19947 4811
rect 19978 4808 19984 4820
rect 19935 4780 19984 4808
rect 19935 4777 19947 4780
rect 19889 4771 19947 4777
rect 19978 4768 19984 4780
rect 20036 4768 20042 4820
rect 9677 4743 9735 4749
rect 6052 4712 6684 4740
rect 6052 4700 6058 4712
rect 4157 4675 4215 4681
rect 4157 4672 4169 4675
rect 4028 4644 4169 4672
rect 4028 4632 4034 4644
rect 4157 4641 4169 4644
rect 4203 4641 4215 4675
rect 4157 4635 4215 4641
rect 4341 4675 4399 4681
rect 4341 4641 4353 4675
rect 4387 4641 4399 4675
rect 4341 4635 4399 4641
rect 4709 4675 4767 4681
rect 4709 4641 4721 4675
rect 4755 4672 4767 4675
rect 5350 4672 5356 4684
rect 4755 4644 5356 4672
rect 4755 4641 4767 4644
rect 4709 4635 4767 4641
rect 1489 4607 1547 4613
rect 1489 4573 1501 4607
rect 1535 4604 1547 4607
rect 1946 4604 1952 4616
rect 1535 4576 1952 4604
rect 1535 4573 1547 4576
rect 1489 4567 1547 4573
rect 1946 4564 1952 4576
rect 2004 4604 2010 4616
rect 2961 4607 3019 4613
rect 2961 4604 2973 4607
rect 2004 4576 2973 4604
rect 2004 4564 2010 4576
rect 2961 4573 2973 4576
rect 3007 4573 3019 4607
rect 2961 4567 3019 4573
rect 3878 4564 3884 4616
rect 3936 4604 3942 4616
rect 4356 4604 4384 4635
rect 5350 4632 5356 4644
rect 5408 4632 5414 4684
rect 5534 4672 5540 4684
rect 5495 4644 5540 4672
rect 5534 4632 5540 4644
rect 5592 4632 5598 4684
rect 5626 4632 5632 4684
rect 5684 4672 5690 4684
rect 6656 4681 6684 4712
rect 9677 4709 9689 4743
rect 9723 4709 9735 4743
rect 12618 4740 12624 4752
rect 12579 4712 12624 4740
rect 9677 4703 9735 4709
rect 12618 4700 12624 4712
rect 12676 4700 12682 4752
rect 12710 4700 12716 4752
rect 12768 4740 12774 4752
rect 12768 4712 13676 4740
rect 12768 4700 12774 4712
rect 5813 4675 5871 4681
rect 5813 4672 5825 4675
rect 5684 4644 5825 4672
rect 5684 4632 5690 4644
rect 5813 4641 5825 4644
rect 5859 4641 5871 4675
rect 5813 4635 5871 4641
rect 6641 4675 6699 4681
rect 6641 4641 6653 4675
rect 6687 4672 6699 4675
rect 7098 4672 7104 4684
rect 6687 4644 7104 4672
rect 6687 4641 6699 4644
rect 6641 4635 6699 4641
rect 7098 4632 7104 4644
rect 7156 4632 7162 4684
rect 7190 4632 7196 4684
rect 7248 4672 7254 4684
rect 7377 4675 7435 4681
rect 7377 4672 7389 4675
rect 7248 4644 7389 4672
rect 7248 4632 7254 4644
rect 7377 4641 7389 4644
rect 7423 4641 7435 4675
rect 7377 4635 7435 4641
rect 8018 4632 8024 4684
rect 8076 4672 8082 4684
rect 8113 4675 8171 4681
rect 8113 4672 8125 4675
rect 8076 4644 8125 4672
rect 8076 4632 8082 4644
rect 8113 4641 8125 4644
rect 8159 4641 8171 4675
rect 9766 4672 9772 4684
rect 9727 4644 9772 4672
rect 8113 4635 8171 4641
rect 9766 4632 9772 4644
rect 9824 4632 9830 4684
rect 11882 4672 11888 4684
rect 11843 4644 11888 4672
rect 11882 4632 11888 4644
rect 11940 4632 11946 4684
rect 12437 4675 12495 4681
rect 12437 4641 12449 4675
rect 12483 4641 12495 4675
rect 13446 4672 13452 4684
rect 13407 4644 13452 4672
rect 12437 4635 12495 4641
rect 3936 4576 4384 4604
rect 3936 4564 3942 4576
rect 5718 4564 5724 4616
rect 5776 4604 5782 4616
rect 5997 4607 6055 4613
rect 5997 4604 6009 4607
rect 5776 4576 6009 4604
rect 5776 4564 5782 4576
rect 5997 4573 6009 4576
rect 6043 4573 6055 4607
rect 5997 4567 6055 4573
rect 7745 4607 7803 4613
rect 7745 4573 7757 4607
rect 7791 4604 7803 4607
rect 8662 4604 8668 4616
rect 7791 4576 8668 4604
rect 7791 4573 7803 4576
rect 7745 4567 7803 4573
rect 8662 4564 8668 4576
rect 8720 4564 8726 4616
rect 11701 4607 11759 4613
rect 11701 4573 11713 4607
rect 11747 4604 11759 4607
rect 11974 4604 11980 4616
rect 11747 4576 11980 4604
rect 11747 4573 11759 4576
rect 11701 4567 11759 4573
rect 11974 4564 11980 4576
rect 12032 4604 12038 4616
rect 12452 4604 12480 4635
rect 13446 4632 13452 4644
rect 13504 4632 13510 4684
rect 13648 4681 13676 4712
rect 13633 4675 13691 4681
rect 13633 4641 13645 4675
rect 13679 4672 13691 4675
rect 13814 4672 13820 4684
rect 13679 4644 13820 4672
rect 13679 4641 13691 4644
rect 13633 4635 13691 4641
rect 13814 4632 13820 4644
rect 13872 4632 13878 4684
rect 13906 4604 13912 4616
rect 12032 4576 13912 4604
rect 12032 4564 12038 4576
rect 13906 4564 13912 4576
rect 13964 4564 13970 4616
rect 15470 4604 15476 4616
rect 15431 4576 15476 4604
rect 15470 4564 15476 4576
rect 15528 4564 15534 4616
rect 18598 4604 18604 4616
rect 18559 4576 18604 4604
rect 18598 4564 18604 4576
rect 18656 4564 18662 4616
rect 5258 4496 5264 4548
rect 5316 4536 5322 4548
rect 5442 4536 5448 4548
rect 5316 4508 5448 4536
rect 5316 4496 5322 4508
rect 5442 4496 5448 4508
rect 5500 4536 5506 4548
rect 5629 4539 5687 4545
rect 5629 4536 5641 4539
rect 5500 4508 5641 4536
rect 5500 4496 5506 4508
rect 5629 4505 5641 4508
rect 5675 4505 5687 4539
rect 5629 4499 5687 4505
rect 6638 4496 6644 4548
rect 6696 4536 6702 4548
rect 7193 4539 7251 4545
rect 7193 4536 7205 4539
rect 6696 4508 7205 4536
rect 6696 4496 6702 4508
rect 7193 4505 7205 4508
rect 7239 4505 7251 4539
rect 7193 4499 7251 4505
rect 7834 4428 7840 4480
rect 7892 4468 7898 4480
rect 10226 4468 10232 4480
rect 7892 4440 10232 4468
rect 7892 4428 7898 4440
rect 10226 4428 10232 4440
rect 10284 4428 10290 4480
rect 1104 4378 22816 4400
rect 1104 4326 4982 4378
rect 5034 4326 5046 4378
rect 5098 4326 5110 4378
rect 5162 4326 5174 4378
rect 5226 4326 12982 4378
rect 13034 4326 13046 4378
rect 13098 4326 13110 4378
rect 13162 4326 13174 4378
rect 13226 4326 20982 4378
rect 21034 4326 21046 4378
rect 21098 4326 21110 4378
rect 21162 4326 21174 4378
rect 21226 4326 22816 4378
rect 1104 4304 22816 4326
rect 2406 4224 2412 4276
rect 2464 4264 2470 4276
rect 2593 4267 2651 4273
rect 2593 4264 2605 4267
rect 2464 4236 2605 4264
rect 2464 4224 2470 4236
rect 2593 4233 2605 4236
rect 2639 4233 2651 4267
rect 3878 4264 3884 4276
rect 3839 4236 3884 4264
rect 2593 4227 2651 4233
rect 3878 4224 3884 4236
rect 3936 4224 3942 4276
rect 6638 4264 6644 4276
rect 5184 4236 6644 4264
rect 5184 4208 5212 4236
rect 6638 4224 6644 4236
rect 6696 4224 6702 4276
rect 7190 4264 7196 4276
rect 7151 4236 7196 4264
rect 7190 4224 7196 4236
rect 7248 4224 7254 4276
rect 7834 4264 7840 4276
rect 7795 4236 7840 4264
rect 7834 4224 7840 4236
rect 7892 4224 7898 4276
rect 11974 4264 11980 4276
rect 11935 4236 11980 4264
rect 11974 4224 11980 4236
rect 12032 4224 12038 4276
rect 13446 4264 13452 4276
rect 13407 4236 13452 4264
rect 13446 4224 13452 4236
rect 13504 4224 13510 4276
rect 13814 4224 13820 4276
rect 13872 4264 13878 4276
rect 13872 4236 13917 4264
rect 13872 4224 13878 4236
rect 15838 4224 15844 4276
rect 15896 4264 15902 4276
rect 15933 4267 15991 4273
rect 15933 4264 15945 4267
rect 15896 4236 15945 4264
rect 15896 4224 15902 4236
rect 15933 4233 15945 4236
rect 15979 4233 15991 4267
rect 15933 4227 15991 4233
rect 16482 4224 16488 4276
rect 16540 4264 16546 4276
rect 17773 4267 17831 4273
rect 17773 4264 17785 4267
rect 16540 4236 17785 4264
rect 16540 4224 16546 4236
rect 17773 4233 17785 4236
rect 17819 4264 17831 4267
rect 18506 4264 18512 4276
rect 17819 4236 18512 4264
rect 17819 4233 17831 4236
rect 17773 4227 17831 4233
rect 18506 4224 18512 4236
rect 18564 4224 18570 4276
rect 18966 4224 18972 4276
rect 19024 4264 19030 4276
rect 19061 4267 19119 4273
rect 19061 4264 19073 4267
rect 19024 4236 19073 4264
rect 19024 4224 19030 4236
rect 19061 4233 19073 4236
rect 19107 4233 19119 4267
rect 19061 4227 19119 4233
rect 4801 4199 4859 4205
rect 4801 4165 4813 4199
rect 4847 4196 4859 4199
rect 5166 4196 5172 4208
rect 4847 4168 5172 4196
rect 4847 4165 4859 4168
rect 4801 4159 4859 4165
rect 5166 4156 5172 4168
rect 5224 4156 5230 4208
rect 7852 4196 7880 4224
rect 7760 4168 7880 4196
rect 11609 4199 11667 4205
rect 3050 4088 3056 4140
rect 3108 4128 3114 4140
rect 5261 4131 5319 4137
rect 5261 4128 5273 4131
rect 3108 4100 5273 4128
rect 3108 4088 3114 4100
rect 5261 4097 5273 4100
rect 5307 4097 5319 4131
rect 5261 4091 5319 4097
rect 2225 4063 2283 4069
rect 2225 4029 2237 4063
rect 2271 4060 2283 4063
rect 2406 4060 2412 4072
rect 2271 4032 2412 4060
rect 2271 4029 2283 4032
rect 2225 4023 2283 4029
rect 2406 4020 2412 4032
rect 2464 4020 2470 4072
rect 4246 4020 4252 4072
rect 4304 4060 4310 4072
rect 4525 4063 4583 4069
rect 4525 4060 4537 4063
rect 4304 4032 4537 4060
rect 4304 4020 4310 4032
rect 4525 4029 4537 4032
rect 4571 4060 4583 4063
rect 4706 4060 4712 4072
rect 4571 4032 4712 4060
rect 4571 4029 4583 4032
rect 4525 4023 4583 4029
rect 4706 4020 4712 4032
rect 4764 4020 4770 4072
rect 4985 4063 5043 4069
rect 4985 4029 4997 4063
rect 5031 4029 5043 4063
rect 7760 4060 7788 4168
rect 11609 4165 11621 4199
rect 11655 4196 11667 4199
rect 11882 4196 11888 4208
rect 11655 4168 11888 4196
rect 11655 4165 11667 4168
rect 11609 4159 11667 4165
rect 11882 4156 11888 4168
rect 11940 4156 11946 4208
rect 9766 4128 9772 4140
rect 9727 4100 9772 4128
rect 9766 4088 9772 4100
rect 9824 4088 9830 4140
rect 13998 4088 14004 4140
rect 14056 4128 14062 4140
rect 14829 4131 14887 4137
rect 14829 4128 14841 4131
rect 14056 4100 14841 4128
rect 14056 4088 14062 4100
rect 14829 4097 14841 4100
rect 14875 4128 14887 4131
rect 19150 4128 19156 4140
rect 14875 4100 15424 4128
rect 14875 4097 14887 4100
rect 14829 4091 14887 4097
rect 7926 4060 7932 4072
rect 7760 4032 7932 4060
rect 4985 4023 5043 4029
rect 1578 3992 1584 4004
rect 1539 3964 1584 3992
rect 1578 3952 1584 3964
rect 1636 3952 1642 4004
rect 4614 3992 4620 4004
rect 4172 3964 4620 3992
rect 4172 3936 4200 3964
rect 4614 3952 4620 3964
rect 4672 3992 4678 4004
rect 5000 3992 5028 4023
rect 7926 4020 7932 4032
rect 7984 4020 7990 4072
rect 8018 4020 8024 4072
rect 8076 4060 8082 4072
rect 8386 4060 8392 4072
rect 8076 4032 8392 4060
rect 8076 4020 8082 4032
rect 8386 4020 8392 4032
rect 8444 4020 8450 4072
rect 8754 4060 8760 4072
rect 8715 4032 8760 4060
rect 8754 4020 8760 4032
rect 8812 4020 8818 4072
rect 9401 4063 9459 4069
rect 9401 4029 9413 4063
rect 9447 4060 9459 4063
rect 10137 4063 10195 4069
rect 10137 4060 10149 4063
rect 9447 4032 10149 4060
rect 9447 4029 9459 4032
rect 9401 4023 9459 4029
rect 10137 4029 10149 4032
rect 10183 4060 10195 4063
rect 10686 4060 10692 4072
rect 10183 4032 10692 4060
rect 10183 4029 10195 4032
rect 10137 4023 10195 4029
rect 10686 4020 10692 4032
rect 10744 4020 10750 4072
rect 12710 4060 12716 4072
rect 12671 4032 12716 4060
rect 12710 4020 12716 4032
rect 12768 4020 12774 4072
rect 15010 4060 15016 4072
rect 14971 4032 15016 4060
rect 15010 4020 15016 4032
rect 15068 4020 15074 4072
rect 15396 4069 15424 4100
rect 18340 4100 19156 4128
rect 15381 4063 15439 4069
rect 15381 4029 15393 4063
rect 15427 4060 15439 4063
rect 16574 4060 16580 4072
rect 15427 4032 16580 4060
rect 15427 4029 15439 4032
rect 15381 4023 15439 4029
rect 16574 4020 16580 4032
rect 16632 4020 16638 4072
rect 18138 4020 18144 4072
rect 18196 4060 18202 4072
rect 18340 4069 18368 4100
rect 19150 4088 19156 4100
rect 19208 4088 19214 4140
rect 18325 4063 18383 4069
rect 18325 4060 18337 4063
rect 18196 4032 18337 4060
rect 18196 4020 18202 4032
rect 18325 4029 18337 4032
rect 18371 4029 18383 4063
rect 18506 4060 18512 4072
rect 18467 4032 18512 4060
rect 18325 4023 18383 4029
rect 18506 4020 18512 4032
rect 18564 4020 18570 4072
rect 19426 4020 19432 4072
rect 19484 4060 19490 4072
rect 20936 4063 20994 4069
rect 20936 4060 20948 4063
rect 19484 4032 20948 4060
rect 19484 4020 19490 4032
rect 20936 4029 20948 4032
rect 20982 4060 20994 4063
rect 21361 4063 21419 4069
rect 21361 4060 21373 4063
rect 20982 4032 21373 4060
rect 20982 4029 20994 4032
rect 20936 4023 20994 4029
rect 21361 4029 21373 4032
rect 21407 4029 21419 4063
rect 21361 4023 21419 4029
rect 4672 3964 5028 3992
rect 4672 3952 4678 3964
rect 5442 3952 5448 4004
rect 5500 3992 5506 4004
rect 6089 3995 6147 4001
rect 6089 3992 6101 3995
rect 5500 3964 6101 3992
rect 5500 3952 5506 3964
rect 6089 3961 6101 3964
rect 6135 3961 6147 3995
rect 12434 3992 12440 4004
rect 12395 3964 12440 3992
rect 6089 3955 6147 3961
rect 12434 3952 12440 3964
rect 12492 3952 12498 4004
rect 15470 3952 15476 4004
rect 15528 3992 15534 4004
rect 15657 3995 15715 4001
rect 15657 3992 15669 3995
rect 15528 3964 15669 3992
rect 15528 3952 15534 3964
rect 15657 3961 15669 3964
rect 15703 3992 15715 3995
rect 16301 3995 16359 4001
rect 16301 3992 16313 3995
rect 15703 3964 16313 3992
rect 15703 3961 15715 3964
rect 15657 3955 15715 3961
rect 16301 3961 16313 3964
rect 16347 3961 16359 3995
rect 16301 3955 16359 3961
rect 18598 3952 18604 4004
rect 18656 3992 18662 4004
rect 18785 3995 18843 4001
rect 18785 3992 18797 3995
rect 18656 3964 18797 3992
rect 18656 3952 18662 3964
rect 18785 3961 18797 3964
rect 18831 3992 18843 3995
rect 19521 3995 19579 4001
rect 19521 3992 19533 3995
rect 18831 3964 19533 3992
rect 18831 3961 18843 3964
rect 18785 3955 18843 3961
rect 19521 3961 19533 3964
rect 19567 3961 19579 3995
rect 19521 3955 19579 3961
rect 21039 3995 21097 4001
rect 21039 3961 21051 3995
rect 21085 3992 21097 3995
rect 23106 3992 23112 4004
rect 21085 3964 23112 3992
rect 21085 3961 21097 3964
rect 21039 3955 21097 3961
rect 23106 3952 23112 3964
rect 23164 3952 23170 4004
rect 198 3884 204 3936
rect 256 3924 262 3936
rect 3421 3927 3479 3933
rect 3421 3924 3433 3927
rect 256 3896 3433 3924
rect 256 3884 262 3896
rect 3421 3893 3433 3896
rect 3467 3924 3479 3927
rect 3970 3924 3976 3936
rect 3467 3896 3976 3924
rect 3467 3893 3479 3896
rect 3421 3887 3479 3893
rect 3970 3884 3976 3896
rect 4028 3884 4034 3936
rect 4154 3924 4160 3936
rect 4115 3896 4160 3924
rect 4154 3884 4160 3896
rect 4212 3884 4218 3936
rect 4706 3884 4712 3936
rect 4764 3924 4770 3936
rect 5534 3924 5540 3936
rect 4764 3896 5540 3924
rect 4764 3884 4770 3896
rect 5534 3884 5540 3896
rect 5592 3924 5598 3936
rect 5721 3927 5779 3933
rect 5721 3924 5733 3927
rect 5592 3896 5733 3924
rect 5592 3884 5598 3896
rect 5721 3893 5733 3896
rect 5767 3893 5779 3927
rect 8846 3924 8852 3936
rect 8807 3896 8852 3924
rect 5721 3887 5779 3893
rect 8846 3884 8852 3896
rect 8904 3884 8910 3936
rect 10502 3924 10508 3936
rect 10463 3896 10508 3924
rect 10502 3884 10508 3896
rect 10560 3884 10566 3936
rect 1104 3834 22816 3856
rect 1104 3782 8982 3834
rect 9034 3782 9046 3834
rect 9098 3782 9110 3834
rect 9162 3782 9174 3834
rect 9226 3782 16982 3834
rect 17034 3782 17046 3834
rect 17098 3782 17110 3834
rect 17162 3782 17174 3834
rect 17226 3782 22816 3834
rect 1104 3760 22816 3782
rect 1578 3720 1584 3732
rect 1539 3692 1584 3720
rect 1578 3680 1584 3692
rect 1636 3680 1642 3732
rect 1946 3720 1952 3732
rect 1907 3692 1952 3720
rect 1946 3680 1952 3692
rect 2004 3680 2010 3732
rect 5166 3720 5172 3732
rect 5127 3692 5172 3720
rect 5166 3680 5172 3692
rect 5224 3680 5230 3732
rect 5626 3720 5632 3732
rect 5587 3692 5632 3720
rect 5626 3680 5632 3692
rect 5684 3680 5690 3732
rect 7098 3720 7104 3732
rect 7059 3692 7104 3720
rect 7098 3680 7104 3692
rect 7156 3720 7162 3732
rect 8389 3723 8447 3729
rect 8389 3720 8401 3723
rect 7156 3692 8401 3720
rect 7156 3680 7162 3692
rect 8389 3689 8401 3692
rect 8435 3720 8447 3723
rect 8754 3720 8760 3732
rect 8435 3692 8760 3720
rect 8435 3689 8447 3692
rect 8389 3683 8447 3689
rect 8754 3680 8760 3692
rect 8812 3680 8818 3732
rect 11054 3680 11060 3732
rect 11112 3720 11118 3732
rect 11149 3723 11207 3729
rect 11149 3720 11161 3723
rect 11112 3692 11161 3720
rect 11112 3680 11118 3692
rect 11149 3689 11161 3692
rect 11195 3689 11207 3723
rect 12710 3720 12716 3732
rect 11149 3683 11207 3689
rect 11900 3692 12716 3720
rect 3970 3612 3976 3664
rect 4028 3652 4034 3664
rect 4798 3652 4804 3664
rect 4028 3624 4384 3652
rect 4759 3624 4804 3652
rect 4028 3612 4034 3624
rect 4246 3584 4252 3596
rect 4207 3556 4252 3584
rect 4246 3544 4252 3556
rect 4304 3544 4310 3596
rect 4356 3584 4384 3624
rect 4798 3612 4804 3624
rect 4856 3612 4862 3664
rect 9950 3612 9956 3664
rect 10008 3652 10014 3664
rect 10274 3655 10332 3661
rect 10274 3652 10286 3655
rect 10008 3624 10286 3652
rect 10008 3612 10014 3624
rect 10274 3621 10286 3624
rect 10320 3621 10332 3655
rect 11514 3652 11520 3664
rect 10274 3615 10332 3621
rect 10888 3624 11520 3652
rect 5810 3584 5816 3596
rect 4356 3556 5816 3584
rect 5810 3544 5816 3556
rect 5868 3584 5874 3596
rect 5905 3587 5963 3593
rect 5905 3584 5917 3587
rect 5868 3556 5917 3584
rect 5868 3544 5874 3556
rect 5905 3553 5917 3556
rect 5951 3553 5963 3587
rect 5905 3547 5963 3553
rect 6549 3587 6607 3593
rect 6549 3553 6561 3587
rect 6595 3584 6607 3587
rect 6638 3584 6644 3596
rect 6595 3556 6644 3584
rect 6595 3553 6607 3556
rect 6549 3547 6607 3553
rect 6638 3544 6644 3556
rect 6696 3584 6702 3596
rect 7558 3584 7564 3596
rect 6696 3556 7564 3584
rect 6696 3544 6702 3556
rect 7558 3544 7564 3556
rect 7616 3544 7622 3596
rect 8110 3584 8116 3596
rect 8071 3556 8116 3584
rect 8110 3544 8116 3556
rect 8168 3544 8174 3596
rect 10888 3593 10916 3624
rect 11514 3612 11520 3624
rect 11572 3652 11578 3664
rect 11900 3661 11928 3692
rect 12710 3680 12716 3692
rect 12768 3680 12774 3732
rect 13446 3720 13452 3732
rect 13407 3692 13452 3720
rect 13446 3680 13452 3692
rect 13504 3680 13510 3732
rect 15010 3720 15016 3732
rect 14971 3692 15016 3720
rect 15010 3680 15016 3692
rect 15068 3680 15074 3732
rect 18138 3720 18144 3732
rect 18099 3692 18144 3720
rect 18138 3680 18144 3692
rect 18196 3680 18202 3732
rect 11885 3655 11943 3661
rect 11885 3652 11897 3655
rect 11572 3624 11897 3652
rect 11572 3612 11578 3624
rect 11885 3621 11897 3624
rect 11931 3621 11943 3655
rect 11885 3615 11943 3621
rect 10873 3587 10931 3593
rect 10873 3553 10885 3587
rect 10919 3553 10931 3587
rect 10873 3547 10931 3553
rect 13300 3587 13358 3593
rect 13300 3553 13312 3587
rect 13346 3553 13358 3587
rect 13300 3547 13358 3553
rect 8846 3476 8852 3528
rect 8904 3516 8910 3528
rect 9953 3519 10011 3525
rect 9953 3516 9965 3519
rect 8904 3488 9965 3516
rect 8904 3476 8910 3488
rect 9953 3485 9965 3488
rect 9999 3485 10011 3519
rect 11790 3516 11796 3528
rect 11751 3488 11796 3516
rect 9953 3479 10011 3485
rect 11790 3476 11796 3488
rect 11848 3476 11854 3528
rect 12437 3519 12495 3525
rect 12437 3485 12449 3519
rect 12483 3516 12495 3519
rect 12802 3516 12808 3528
rect 12483 3488 12808 3516
rect 12483 3485 12495 3488
rect 12437 3479 12495 3485
rect 12802 3476 12808 3488
rect 12860 3516 12866 3528
rect 13315 3516 13343 3547
rect 12860 3488 13343 3516
rect 12860 3476 12866 3488
rect 7466 3448 7472 3460
rect 7427 3420 7472 3448
rect 7466 3408 7472 3420
rect 7524 3408 7530 3460
rect 1104 3290 22816 3312
rect 1104 3238 4982 3290
rect 5034 3238 5046 3290
rect 5098 3238 5110 3290
rect 5162 3238 5174 3290
rect 5226 3238 12982 3290
rect 13034 3238 13046 3290
rect 13098 3238 13110 3290
rect 13162 3238 13174 3290
rect 13226 3238 20982 3290
rect 21034 3238 21046 3290
rect 21098 3238 21110 3290
rect 21162 3238 21174 3290
rect 21226 3238 22816 3290
rect 1104 3216 22816 3238
rect 5169 3179 5227 3185
rect 5169 3145 5181 3179
rect 5215 3176 5227 3179
rect 5350 3176 5356 3188
rect 5215 3148 5356 3176
rect 5215 3145 5227 3148
rect 5169 3139 5227 3145
rect 5350 3136 5356 3148
rect 5408 3136 5414 3188
rect 5810 3176 5816 3188
rect 5771 3148 5816 3176
rect 5810 3136 5816 3148
rect 5868 3136 5874 3188
rect 6638 3176 6644 3188
rect 6599 3148 6644 3176
rect 6638 3136 6644 3148
rect 6696 3136 6702 3188
rect 8846 3136 8852 3188
rect 8904 3176 8910 3188
rect 9217 3179 9275 3185
rect 9217 3176 9229 3179
rect 8904 3148 9229 3176
rect 8904 3136 8910 3148
rect 9217 3145 9229 3148
rect 9263 3145 9275 3179
rect 11514 3176 11520 3188
rect 11475 3148 11520 3176
rect 9217 3139 9275 3145
rect 11514 3136 11520 3148
rect 11572 3136 11578 3188
rect 12253 3179 12311 3185
rect 12253 3145 12265 3179
rect 12299 3176 12311 3179
rect 12434 3176 12440 3188
rect 12299 3148 12440 3176
rect 12299 3145 12311 3148
rect 12253 3139 12311 3145
rect 12434 3136 12440 3148
rect 12492 3136 12498 3188
rect 13354 3176 13360 3188
rect 12544 3148 13360 3176
rect 5534 3068 5540 3120
rect 5592 3108 5598 3120
rect 7469 3111 7527 3117
rect 7469 3108 7481 3111
rect 5592 3080 7481 3108
rect 5592 3068 5598 3080
rect 7469 3077 7481 3080
rect 7515 3077 7527 3111
rect 11054 3108 11060 3120
rect 7469 3071 7527 3077
rect 10520 3080 11060 3108
rect 7484 3040 7512 3071
rect 8386 3040 8392 3052
rect 7484 3012 8064 3040
rect 8347 3012 8392 3040
rect 4617 2975 4675 2981
rect 4617 2941 4629 2975
rect 4663 2972 4675 2975
rect 5350 2972 5356 2984
rect 4663 2944 5356 2972
rect 4663 2941 4675 2944
rect 4617 2935 4675 2941
rect 5350 2932 5356 2944
rect 5408 2932 5414 2984
rect 7926 2972 7932 2984
rect 7887 2944 7932 2972
rect 7926 2932 7932 2944
rect 7984 2932 7990 2984
rect 8036 2972 8064 3012
rect 8386 3000 8392 3012
rect 8444 3000 8450 3052
rect 10520 3049 10548 3080
rect 11054 3068 11060 3080
rect 11112 3068 11118 3120
rect 12544 3108 12572 3148
rect 13354 3136 13360 3148
rect 13412 3176 13418 3188
rect 13449 3179 13507 3185
rect 13449 3176 13461 3179
rect 13412 3148 13461 3176
rect 13412 3136 13418 3148
rect 13449 3145 13461 3148
rect 13495 3145 13507 3179
rect 13449 3139 13507 3145
rect 11808 3080 12572 3108
rect 11808 3052 11836 3080
rect 12802 3068 12808 3120
rect 12860 3108 12866 3120
rect 13081 3111 13139 3117
rect 13081 3108 13093 3111
rect 12860 3080 13093 3108
rect 12860 3068 12866 3080
rect 13081 3077 13093 3080
rect 13127 3108 13139 3111
rect 13817 3111 13875 3117
rect 13817 3108 13829 3111
rect 13127 3080 13829 3108
rect 13127 3077 13139 3080
rect 13081 3071 13139 3077
rect 13817 3077 13829 3080
rect 13863 3077 13875 3111
rect 13817 3071 13875 3077
rect 10505 3043 10563 3049
rect 10505 3009 10517 3043
rect 10551 3009 10563 3043
rect 10505 3003 10563 3009
rect 11149 3043 11207 3049
rect 11149 3009 11161 3043
rect 11195 3040 11207 3043
rect 11790 3040 11796 3052
rect 11195 3012 11796 3040
rect 11195 3009 11207 3012
rect 11149 3003 11207 3009
rect 11790 3000 11796 3012
rect 11848 3000 11854 3052
rect 11885 3043 11943 3049
rect 11885 3009 11897 3043
rect 11931 3040 11943 3043
rect 12529 3043 12587 3049
rect 12529 3040 12541 3043
rect 11931 3012 12541 3040
rect 11931 3009 11943 3012
rect 11885 3003 11943 3009
rect 12529 3009 12541 3012
rect 12575 3040 12587 3043
rect 14001 3043 14059 3049
rect 14001 3040 14013 3043
rect 12575 3012 14013 3040
rect 12575 3009 12587 3012
rect 12529 3003 12587 3009
rect 14001 3009 14013 3012
rect 14047 3009 14059 3043
rect 14001 3003 14059 3009
rect 8481 2975 8539 2981
rect 8481 2972 8493 2975
rect 8036 2944 8493 2972
rect 8481 2941 8493 2944
rect 8527 2941 8539 2975
rect 8481 2935 8539 2941
rect 7193 2907 7251 2913
rect 7193 2873 7205 2907
rect 7239 2904 7251 2907
rect 8110 2904 8116 2916
rect 7239 2876 8116 2904
rect 7239 2873 7251 2876
rect 7193 2867 7251 2873
rect 8110 2864 8116 2876
rect 8168 2864 8174 2916
rect 9677 2907 9735 2913
rect 9677 2873 9689 2907
rect 9723 2904 9735 2907
rect 10502 2904 10508 2916
rect 9723 2876 10508 2904
rect 9723 2873 9735 2876
rect 9677 2867 9735 2873
rect 10502 2864 10508 2876
rect 10560 2904 10566 2916
rect 10597 2907 10655 2913
rect 10597 2904 10609 2907
rect 10560 2876 10609 2904
rect 10560 2864 10566 2876
rect 10597 2873 10609 2876
rect 10643 2873 10655 2907
rect 10597 2867 10655 2873
rect 12621 2907 12679 2913
rect 12621 2873 12633 2907
rect 12667 2873 12679 2907
rect 12621 2867 12679 2873
rect 4157 2839 4215 2845
rect 4157 2805 4169 2839
rect 4203 2836 4215 2839
rect 4246 2836 4252 2848
rect 4203 2808 4252 2836
rect 4203 2805 4215 2808
rect 4157 2799 4215 2805
rect 4246 2796 4252 2808
rect 4304 2796 4310 2848
rect 8757 2839 8815 2845
rect 8757 2805 8769 2839
rect 8803 2836 8815 2839
rect 9766 2836 9772 2848
rect 8803 2808 9772 2836
rect 8803 2805 8815 2808
rect 8757 2799 8815 2805
rect 9766 2796 9772 2808
rect 9824 2796 9830 2848
rect 9950 2836 9956 2848
rect 9911 2808 9956 2836
rect 9950 2796 9956 2808
rect 10008 2796 10014 2848
rect 12434 2796 12440 2848
rect 12492 2836 12498 2848
rect 12636 2836 12664 2867
rect 12492 2808 12664 2836
rect 12492 2796 12498 2808
rect 1104 2746 22816 2768
rect 1104 2694 8982 2746
rect 9034 2694 9046 2746
rect 9098 2694 9110 2746
rect 9162 2694 9174 2746
rect 9226 2694 16982 2746
rect 17034 2694 17046 2746
rect 17098 2694 17110 2746
rect 17162 2694 17174 2746
rect 17226 2694 22816 2746
rect 1104 2672 22816 2694
rect 6365 2635 6423 2641
rect 6365 2601 6377 2635
rect 6411 2632 6423 2635
rect 6546 2632 6552 2644
rect 6411 2604 6552 2632
rect 6411 2601 6423 2604
rect 6365 2595 6423 2601
rect 5721 2499 5779 2505
rect 5721 2465 5733 2499
rect 5767 2496 5779 2499
rect 6380 2496 6408 2595
rect 6546 2592 6552 2604
rect 6604 2592 6610 2644
rect 7926 2632 7932 2644
rect 7887 2604 7932 2632
rect 7926 2592 7932 2604
rect 7984 2592 7990 2644
rect 8386 2632 8392 2644
rect 8347 2604 8392 2632
rect 8386 2592 8392 2604
rect 8444 2592 8450 2644
rect 9585 2635 9643 2641
rect 9585 2601 9597 2635
rect 9631 2632 9643 2635
rect 9950 2632 9956 2644
rect 9631 2604 9956 2632
rect 9631 2601 9643 2604
rect 9585 2595 9643 2601
rect 9950 2592 9956 2604
rect 10008 2592 10014 2644
rect 10686 2632 10692 2644
rect 10647 2604 10692 2632
rect 10686 2592 10692 2604
rect 10744 2632 10750 2644
rect 12345 2635 12403 2641
rect 12345 2632 12357 2635
rect 10744 2604 12357 2632
rect 10744 2592 10750 2604
rect 12345 2601 12357 2604
rect 12391 2632 12403 2635
rect 12391 2604 12848 2632
rect 12391 2601 12403 2604
rect 12345 2595 12403 2601
rect 6914 2564 6920 2576
rect 6875 2536 6920 2564
rect 6914 2524 6920 2536
rect 6972 2524 6978 2576
rect 9968 2564 9996 2592
rect 12820 2573 12848 2604
rect 10090 2567 10148 2573
rect 10090 2564 10102 2567
rect 9968 2536 10102 2564
rect 10090 2533 10102 2536
rect 10136 2533 10148 2567
rect 10090 2527 10148 2533
rect 12805 2567 12863 2573
rect 12805 2533 12817 2567
rect 12851 2533 12863 2567
rect 13354 2564 13360 2576
rect 13315 2536 13360 2564
rect 12805 2527 12863 2533
rect 13354 2524 13360 2536
rect 13412 2524 13418 2576
rect 7009 2499 7067 2505
rect 7009 2496 7021 2499
rect 5767 2468 6408 2496
rect 6656 2468 7021 2496
rect 5767 2465 5779 2468
rect 5721 2459 5779 2465
rect 1210 2320 1216 2372
rect 1268 2360 1274 2372
rect 6656 2369 6684 2468
rect 7009 2465 7021 2468
rect 7055 2465 7067 2499
rect 7009 2459 7067 2465
rect 8202 2456 8208 2508
rect 8260 2496 8266 2508
rect 8573 2499 8631 2505
rect 8573 2496 8585 2499
rect 8260 2468 8585 2496
rect 8260 2456 8266 2468
rect 8573 2465 8585 2468
rect 8619 2496 8631 2499
rect 9125 2499 9183 2505
rect 9125 2496 9137 2499
rect 8619 2468 9137 2496
rect 8619 2465 8631 2468
rect 8573 2459 8631 2465
rect 9125 2465 9137 2468
rect 9171 2465 9183 2499
rect 9766 2496 9772 2508
rect 9727 2468 9772 2496
rect 9125 2459 9183 2465
rect 9766 2456 9772 2468
rect 9824 2496 9830 2508
rect 10965 2499 11023 2505
rect 10965 2496 10977 2499
rect 9824 2468 10977 2496
rect 9824 2456 9830 2468
rect 10965 2465 10977 2468
rect 11011 2465 11023 2499
rect 11552 2499 11610 2505
rect 11552 2496 11564 2499
rect 10965 2459 11023 2465
rect 11072 2468 11564 2496
rect 6730 2388 6736 2440
rect 6788 2428 6794 2440
rect 9398 2428 9404 2440
rect 6788 2400 9404 2428
rect 6788 2388 6794 2400
rect 9398 2388 9404 2400
rect 9456 2428 9462 2440
rect 11072 2428 11100 2468
rect 11552 2465 11564 2468
rect 11598 2496 11610 2499
rect 11977 2499 12035 2505
rect 11977 2496 11989 2499
rect 11598 2468 11989 2496
rect 11598 2465 11610 2468
rect 11552 2459 11610 2465
rect 11977 2465 11989 2468
rect 12023 2465 12035 2499
rect 11977 2459 12035 2465
rect 14185 2499 14243 2505
rect 14185 2465 14197 2499
rect 14231 2496 14243 2499
rect 17126 2496 17132 2508
rect 14231 2468 14872 2496
rect 17087 2468 17132 2496
rect 14231 2465 14243 2468
rect 14185 2459 14243 2465
rect 9456 2400 11100 2428
rect 11655 2431 11713 2437
rect 9456 2388 9462 2400
rect 11655 2397 11667 2431
rect 11701 2428 11713 2431
rect 12713 2431 12771 2437
rect 12713 2428 12725 2431
rect 11701 2400 12725 2428
rect 11701 2397 11713 2400
rect 11655 2391 11713 2397
rect 12713 2397 12725 2400
rect 12759 2428 12771 2431
rect 13633 2431 13691 2437
rect 13633 2428 13645 2431
rect 12759 2400 13645 2428
rect 12759 2397 12771 2400
rect 12713 2391 12771 2397
rect 13633 2397 13645 2400
rect 13679 2397 13691 2431
rect 13633 2391 13691 2397
rect 6641 2363 6699 2369
rect 6641 2360 6653 2363
rect 1268 2332 6653 2360
rect 1268 2320 1274 2332
rect 6641 2329 6653 2332
rect 6687 2329 6699 2363
rect 6641 2323 6699 2329
rect 8757 2363 8815 2369
rect 8757 2329 8769 2363
rect 8803 2360 8815 2363
rect 12066 2360 12072 2372
rect 8803 2332 12072 2360
rect 8803 2329 8815 2332
rect 8757 2323 8815 2329
rect 12066 2320 12072 2332
rect 12124 2320 12130 2372
rect 5902 2292 5908 2304
rect 5863 2264 5908 2292
rect 5902 2252 5908 2264
rect 5960 2252 5966 2304
rect 14090 2252 14096 2304
rect 14148 2292 14154 2304
rect 14844 2301 14872 2468
rect 17126 2456 17132 2468
rect 17184 2496 17190 2508
rect 17681 2499 17739 2505
rect 17681 2496 17693 2499
rect 17184 2468 17693 2496
rect 17184 2456 17190 2468
rect 17681 2465 17693 2468
rect 17727 2496 17739 2499
rect 17954 2496 17960 2508
rect 17727 2468 17960 2496
rect 17727 2465 17739 2468
rect 17681 2459 17739 2465
rect 17954 2456 17960 2468
rect 18012 2456 18018 2508
rect 17313 2363 17371 2369
rect 17313 2329 17325 2363
rect 17359 2360 17371 2363
rect 19426 2360 19432 2372
rect 17359 2332 19432 2360
rect 17359 2329 17371 2332
rect 17313 2323 17371 2329
rect 19426 2320 19432 2332
rect 19484 2320 19490 2372
rect 14369 2295 14427 2301
rect 14369 2292 14381 2295
rect 14148 2264 14381 2292
rect 14148 2252 14154 2264
rect 14369 2261 14381 2264
rect 14415 2261 14427 2295
rect 14369 2255 14427 2261
rect 14829 2295 14887 2301
rect 14829 2261 14841 2295
rect 14875 2292 14887 2295
rect 15286 2292 15292 2304
rect 14875 2264 15292 2292
rect 14875 2261 14887 2264
rect 14829 2255 14887 2261
rect 15286 2252 15292 2264
rect 15344 2252 15350 2304
rect 1104 2202 22816 2224
rect 1104 2150 4982 2202
rect 5034 2150 5046 2202
rect 5098 2150 5110 2202
rect 5162 2150 5174 2202
rect 5226 2150 12982 2202
rect 13034 2150 13046 2202
rect 13098 2150 13110 2202
rect 13162 2150 13174 2202
rect 13226 2150 20982 2202
rect 21034 2150 21046 2202
rect 21098 2150 21110 2202
rect 21162 2150 21174 2202
rect 21226 2150 22816 2202
rect 1104 2128 22816 2150
<< via1 >>
rect 4982 21734 5034 21786
rect 5046 21734 5098 21786
rect 5110 21734 5162 21786
rect 5174 21734 5226 21786
rect 12982 21734 13034 21786
rect 13046 21734 13098 21786
rect 13110 21734 13162 21786
rect 13174 21734 13226 21786
rect 20982 21734 21034 21786
rect 21046 21734 21098 21786
rect 21110 21734 21162 21786
rect 21174 21734 21226 21786
rect 8982 21190 9034 21242
rect 9046 21190 9098 21242
rect 9110 21190 9162 21242
rect 9174 21190 9226 21242
rect 16982 21190 17034 21242
rect 17046 21190 17098 21242
rect 17110 21190 17162 21242
rect 17174 21190 17226 21242
rect 4982 20646 5034 20698
rect 5046 20646 5098 20698
rect 5110 20646 5162 20698
rect 5174 20646 5226 20698
rect 12982 20646 13034 20698
rect 13046 20646 13098 20698
rect 13110 20646 13162 20698
rect 13174 20646 13226 20698
rect 20982 20646 21034 20698
rect 21046 20646 21098 20698
rect 21110 20646 21162 20698
rect 21174 20646 21226 20698
rect 7012 20544 7064 20596
rect 8668 20544 8720 20596
rect 10784 20544 10836 20596
rect 16580 20544 16632 20596
rect 20628 20544 20680 20596
rect 1308 20408 1360 20460
rect 5632 20383 5684 20392
rect 5632 20349 5641 20383
rect 5641 20349 5675 20383
rect 5675 20349 5684 20383
rect 5632 20340 5684 20349
rect 15108 20383 15160 20392
rect 1768 20204 1820 20256
rect 8392 20204 8444 20256
rect 15108 20349 15117 20383
rect 15117 20349 15151 20383
rect 15151 20349 15160 20383
rect 15108 20340 15160 20349
rect 18236 20340 18288 20392
rect 11980 20204 12032 20256
rect 8982 20102 9034 20154
rect 9046 20102 9098 20154
rect 9110 20102 9162 20154
rect 9174 20102 9226 20154
rect 16982 20102 17034 20154
rect 17046 20102 17098 20154
rect 17110 20102 17162 20154
rect 17174 20102 17226 20154
rect 18972 20000 19024 20052
rect 10232 19864 10284 19916
rect 17684 19864 17736 19916
rect 1216 19660 1268 19712
rect 10232 19703 10284 19712
rect 10232 19669 10241 19703
rect 10241 19669 10275 19703
rect 10275 19669 10284 19703
rect 10232 19660 10284 19669
rect 4982 19558 5034 19610
rect 5046 19558 5098 19610
rect 5110 19558 5162 19610
rect 5174 19558 5226 19610
rect 12982 19558 13034 19610
rect 13046 19558 13098 19610
rect 13110 19558 13162 19610
rect 13174 19558 13226 19610
rect 20982 19558 21034 19610
rect 21046 19558 21098 19610
rect 21110 19558 21162 19610
rect 21174 19558 21226 19610
rect 22652 19456 22704 19508
rect 20812 19252 20864 19304
rect 10232 19184 10284 19236
rect 12808 19184 12860 19236
rect 10508 19116 10560 19168
rect 17684 19116 17736 19168
rect 8982 19014 9034 19066
rect 9046 19014 9098 19066
rect 9110 19014 9162 19066
rect 9174 19014 9226 19066
rect 16982 19014 17034 19066
rect 17046 19014 17098 19066
rect 17110 19014 17162 19066
rect 17174 19014 17226 19066
rect 10508 18912 10560 18964
rect 11520 18912 11572 18964
rect 21272 18912 21324 18964
rect 1308 18844 1360 18896
rect 1676 18776 1728 18828
rect 7472 18844 7524 18896
rect 9772 18844 9824 18896
rect 7104 18819 7156 18828
rect 7104 18785 7113 18819
rect 7113 18785 7147 18819
rect 7147 18785 7156 18819
rect 7104 18776 7156 18785
rect 15200 18776 15252 18828
rect 7196 18751 7248 18760
rect 7196 18717 7205 18751
rect 7205 18717 7239 18751
rect 7239 18717 7248 18751
rect 7196 18708 7248 18717
rect 9680 18751 9732 18760
rect 9680 18717 9689 18751
rect 9689 18717 9723 18751
rect 9723 18717 9732 18751
rect 9680 18708 9732 18717
rect 11796 18708 11848 18760
rect 16672 18776 16724 18828
rect 21548 18776 21600 18828
rect 16856 18708 16908 18760
rect 17316 18751 17368 18760
rect 17316 18717 17325 18751
rect 17325 18717 17359 18751
rect 17359 18717 17368 18751
rect 17316 18708 17368 18717
rect 20352 18708 20404 18760
rect 4804 18572 4856 18624
rect 8300 18615 8352 18624
rect 8300 18581 8309 18615
rect 8309 18581 8343 18615
rect 8343 18581 8352 18615
rect 8300 18572 8352 18581
rect 12348 18615 12400 18624
rect 12348 18581 12357 18615
rect 12357 18581 12391 18615
rect 12391 18581 12400 18615
rect 12348 18572 12400 18581
rect 12624 18615 12676 18624
rect 12624 18581 12633 18615
rect 12633 18581 12667 18615
rect 12667 18581 12676 18615
rect 12624 18572 12676 18581
rect 15568 18572 15620 18624
rect 15752 18615 15804 18624
rect 15752 18581 15761 18615
rect 15761 18581 15795 18615
rect 15795 18581 15804 18615
rect 15752 18572 15804 18581
rect 16120 18615 16172 18624
rect 16120 18581 16129 18615
rect 16129 18581 16163 18615
rect 16163 18581 16172 18615
rect 16120 18572 16172 18581
rect 18788 18615 18840 18624
rect 18788 18581 18797 18615
rect 18797 18581 18831 18615
rect 18831 18581 18840 18615
rect 18788 18572 18840 18581
rect 4982 18470 5034 18522
rect 5046 18470 5098 18522
rect 5110 18470 5162 18522
rect 5174 18470 5226 18522
rect 12982 18470 13034 18522
rect 13046 18470 13098 18522
rect 13110 18470 13162 18522
rect 13174 18470 13226 18522
rect 20982 18470 21034 18522
rect 21046 18470 21098 18522
rect 21110 18470 21162 18522
rect 21174 18470 21226 18522
rect 2412 18368 2464 18420
rect 7472 18368 7524 18420
rect 9772 18368 9824 18420
rect 11520 18411 11572 18420
rect 11520 18377 11529 18411
rect 11529 18377 11563 18411
rect 11563 18377 11572 18411
rect 11520 18368 11572 18377
rect 12348 18368 12400 18420
rect 3424 18207 3476 18216
rect 3424 18173 3433 18207
rect 3433 18173 3467 18207
rect 3467 18173 3476 18207
rect 3424 18164 3476 18173
rect 5540 18300 5592 18352
rect 7104 18300 7156 18352
rect 10876 18300 10928 18352
rect 16856 18368 16908 18420
rect 20352 18411 20404 18420
rect 20352 18377 20361 18411
rect 20361 18377 20395 18411
rect 20395 18377 20404 18411
rect 20352 18368 20404 18377
rect 4804 18232 4856 18284
rect 5356 18275 5408 18284
rect 5356 18241 5365 18275
rect 5365 18241 5399 18275
rect 5399 18241 5408 18275
rect 5356 18232 5408 18241
rect 8576 18275 8628 18284
rect 8576 18241 8585 18275
rect 8585 18241 8619 18275
rect 8619 18241 8628 18275
rect 8576 18232 8628 18241
rect 9680 18232 9732 18284
rect 12624 18232 12676 18284
rect 12808 18275 12860 18284
rect 12808 18241 12817 18275
rect 12817 18241 12851 18275
rect 12851 18241 12860 18275
rect 12808 18232 12860 18241
rect 16120 18232 16172 18284
rect 18788 18275 18840 18284
rect 18788 18241 18797 18275
rect 18797 18241 18831 18275
rect 18831 18241 18840 18275
rect 18788 18232 18840 18241
rect 20812 18232 20864 18284
rect 9864 18207 9916 18216
rect 3148 18096 3200 18148
rect 9864 18173 9873 18207
rect 9873 18173 9907 18207
rect 9907 18173 9916 18207
rect 9864 18164 9916 18173
rect 4068 18139 4120 18148
rect 4068 18105 4077 18139
rect 4077 18105 4111 18139
rect 4111 18105 4120 18139
rect 4068 18096 4120 18105
rect 8300 18139 8352 18148
rect 1676 18071 1728 18080
rect 1676 18037 1685 18071
rect 1685 18037 1719 18071
rect 1719 18037 1728 18071
rect 1676 18028 1728 18037
rect 1952 18071 2004 18080
rect 1952 18037 1961 18071
rect 1961 18037 1995 18071
rect 1995 18037 2004 18071
rect 1952 18028 2004 18037
rect 4436 18071 4488 18080
rect 4436 18037 4445 18071
rect 4445 18037 4479 18071
rect 4479 18037 4488 18071
rect 4436 18028 4488 18037
rect 8300 18105 8309 18139
rect 8309 18105 8343 18139
rect 8343 18105 8352 18139
rect 8300 18096 8352 18105
rect 5172 18028 5224 18080
rect 7472 18071 7524 18080
rect 7472 18037 7481 18071
rect 7481 18037 7515 18071
rect 7515 18037 7524 18071
rect 7472 18028 7524 18037
rect 7932 18028 7984 18080
rect 13176 18164 13228 18216
rect 11060 18028 11112 18080
rect 11796 18071 11848 18080
rect 11796 18037 11805 18071
rect 11805 18037 11839 18071
rect 11839 18037 11848 18071
rect 11796 18028 11848 18037
rect 12348 18028 12400 18080
rect 15752 18096 15804 18148
rect 18420 18096 18472 18148
rect 15200 18071 15252 18080
rect 15200 18037 15209 18071
rect 15209 18037 15243 18071
rect 15243 18037 15252 18071
rect 15200 18028 15252 18037
rect 16672 18071 16724 18080
rect 16672 18037 16681 18071
rect 16681 18037 16715 18071
rect 16715 18037 16724 18071
rect 16672 18028 16724 18037
rect 16856 18028 16908 18080
rect 17408 18028 17460 18080
rect 17500 18028 17552 18080
rect 20536 18028 20588 18080
rect 21548 18071 21600 18080
rect 21548 18037 21557 18071
rect 21557 18037 21591 18071
rect 21591 18037 21600 18071
rect 21548 18028 21600 18037
rect 8982 17926 9034 17978
rect 9046 17926 9098 17978
rect 9110 17926 9162 17978
rect 9174 17926 9226 17978
rect 16982 17926 17034 17978
rect 17046 17926 17098 17978
rect 17110 17926 17162 17978
rect 17174 17926 17226 17978
rect 2228 17867 2280 17876
rect 2228 17833 2237 17867
rect 2237 17833 2271 17867
rect 2271 17833 2280 17867
rect 2228 17824 2280 17833
rect 3424 17867 3476 17876
rect 3424 17833 3433 17867
rect 3433 17833 3467 17867
rect 3467 17833 3476 17867
rect 3424 17824 3476 17833
rect 5172 17867 5224 17876
rect 5172 17833 5181 17867
rect 5181 17833 5215 17867
rect 5215 17833 5224 17867
rect 5172 17824 5224 17833
rect 8392 17824 8444 17876
rect 13176 17824 13228 17876
rect 15660 17867 15712 17876
rect 15660 17833 15669 17867
rect 15669 17833 15703 17867
rect 15703 17833 15712 17867
rect 15660 17824 15712 17833
rect 15752 17824 15804 17876
rect 17500 17867 17552 17876
rect 17500 17833 17509 17867
rect 17509 17833 17543 17867
rect 17543 17833 17552 17867
rect 17500 17824 17552 17833
rect 18788 17824 18840 17876
rect 20536 17867 20588 17876
rect 20536 17833 20545 17867
rect 20545 17833 20579 17867
rect 20579 17833 20588 17867
rect 20536 17824 20588 17833
rect 21088 17867 21140 17876
rect 21088 17833 21097 17867
rect 21097 17833 21131 17867
rect 21131 17833 21140 17867
rect 21088 17824 21140 17833
rect 4160 17756 4212 17808
rect 7748 17756 7800 17808
rect 11796 17756 11848 17808
rect 12256 17756 12308 17808
rect 15200 17756 15252 17808
rect 20720 17756 20772 17808
rect 4068 17688 4120 17740
rect 4712 17688 4764 17740
rect 6000 17731 6052 17740
rect 6000 17697 6044 17731
rect 6044 17697 6052 17731
rect 7196 17731 7248 17740
rect 6000 17688 6052 17697
rect 7196 17697 7205 17731
rect 7205 17697 7239 17731
rect 7239 17697 7248 17731
rect 7196 17688 7248 17697
rect 10876 17731 10928 17740
rect 10876 17697 10885 17731
rect 10885 17697 10919 17731
rect 10919 17697 10928 17731
rect 10876 17688 10928 17697
rect 11060 17731 11112 17740
rect 11060 17697 11069 17731
rect 11069 17697 11103 17731
rect 11103 17697 11112 17731
rect 11060 17688 11112 17697
rect 13268 17688 13320 17740
rect 17316 17688 17368 17740
rect 18880 17731 18932 17740
rect 18880 17697 18889 17731
rect 18889 17697 18923 17731
rect 18923 17697 18932 17731
rect 18880 17688 18932 17697
rect 19064 17688 19116 17740
rect 7472 17552 7524 17604
rect 1860 17484 1912 17536
rect 2780 17527 2832 17536
rect 2780 17493 2789 17527
rect 2789 17493 2823 17527
rect 2823 17493 2832 17527
rect 2780 17484 2832 17493
rect 5908 17484 5960 17536
rect 7932 17484 7984 17536
rect 8852 17484 8904 17536
rect 9864 17527 9916 17536
rect 9864 17493 9873 17527
rect 9873 17493 9907 17527
rect 9907 17493 9916 17527
rect 9864 17484 9916 17493
rect 10784 17484 10836 17536
rect 12624 17620 12676 17672
rect 13360 17620 13412 17672
rect 15292 17663 15344 17672
rect 15292 17629 15301 17663
rect 15301 17629 15335 17663
rect 15335 17629 15344 17663
rect 15292 17620 15344 17629
rect 13820 17552 13872 17604
rect 12716 17484 12768 17536
rect 13360 17484 13412 17536
rect 13452 17484 13504 17536
rect 15476 17484 15528 17536
rect 18052 17527 18104 17536
rect 18052 17493 18061 17527
rect 18061 17493 18095 17527
rect 18095 17493 18104 17527
rect 18052 17484 18104 17493
rect 18420 17527 18472 17536
rect 18420 17493 18429 17527
rect 18429 17493 18463 17527
rect 18463 17493 18472 17527
rect 18420 17484 18472 17493
rect 19708 17484 19760 17536
rect 4982 17382 5034 17434
rect 5046 17382 5098 17434
rect 5110 17382 5162 17434
rect 5174 17382 5226 17434
rect 12982 17382 13034 17434
rect 13046 17382 13098 17434
rect 13110 17382 13162 17434
rect 13174 17382 13226 17434
rect 20982 17382 21034 17434
rect 21046 17382 21098 17434
rect 21110 17382 21162 17434
rect 21174 17382 21226 17434
rect 2228 17280 2280 17332
rect 4068 17280 4120 17332
rect 6000 17323 6052 17332
rect 6000 17289 6009 17323
rect 6009 17289 6043 17323
rect 6043 17289 6052 17323
rect 6000 17280 6052 17289
rect 8300 17280 8352 17332
rect 11980 17280 12032 17332
rect 13452 17280 13504 17332
rect 15292 17280 15344 17332
rect 18052 17280 18104 17332
rect 18880 17280 18932 17332
rect 20720 17280 20772 17332
rect 1676 17212 1728 17264
rect 1952 17144 2004 17196
rect 4712 17212 4764 17264
rect 5356 17144 5408 17196
rect 9772 17212 9824 17264
rect 9496 17119 9548 17128
rect 9496 17085 9514 17119
rect 9514 17085 9548 17119
rect 9496 17076 9548 17085
rect 2780 17008 2832 17060
rect 4436 17051 4488 17060
rect 4436 17017 4445 17051
rect 4445 17017 4479 17051
rect 4479 17017 4488 17051
rect 4436 17008 4488 17017
rect 2228 16940 2280 16992
rect 2596 16940 2648 16992
rect 4160 16983 4212 16992
rect 4160 16949 4169 16983
rect 4169 16949 4203 16983
rect 4203 16949 4212 16983
rect 4160 16940 4212 16949
rect 7932 17008 7984 17060
rect 8116 17008 8168 17060
rect 4988 16940 5040 16992
rect 7748 16983 7800 16992
rect 7748 16949 7757 16983
rect 7757 16949 7791 16983
rect 7791 16949 7800 16983
rect 7748 16940 7800 16949
rect 8484 16940 8536 16992
rect 10784 17076 10836 17128
rect 10416 17008 10468 17060
rect 11060 17076 11112 17128
rect 11152 17051 11204 17060
rect 11152 17017 11161 17051
rect 11161 17017 11195 17051
rect 11195 17017 11204 17051
rect 11152 17008 11204 17017
rect 13268 17212 13320 17264
rect 12532 17187 12584 17196
rect 12532 17153 12541 17187
rect 12541 17153 12575 17187
rect 12575 17153 12584 17187
rect 12532 17144 12584 17153
rect 12808 17187 12860 17196
rect 12808 17153 12817 17187
rect 12817 17153 12851 17187
rect 12851 17153 12860 17187
rect 12808 17144 12860 17153
rect 12900 17144 12952 17196
rect 15568 17144 15620 17196
rect 16212 17144 16264 17196
rect 18420 17144 18472 17196
rect 20812 17144 20864 17196
rect 14096 17119 14148 17128
rect 14096 17085 14105 17119
rect 14105 17085 14139 17119
rect 14139 17085 14148 17119
rect 14096 17076 14148 17085
rect 12624 17051 12676 17060
rect 12624 17017 12633 17051
rect 12633 17017 12667 17051
rect 12667 17017 12676 17051
rect 12624 17008 12676 17017
rect 13728 17008 13780 17060
rect 15844 17051 15896 17060
rect 15844 17017 15853 17051
rect 15853 17017 15887 17051
rect 15887 17017 15896 17051
rect 16396 17051 16448 17060
rect 15844 17008 15896 17017
rect 16396 17017 16405 17051
rect 16405 17017 16439 17051
rect 16439 17017 16448 17051
rect 16396 17008 16448 17017
rect 19708 17051 19760 17060
rect 11796 16983 11848 16992
rect 11796 16949 11805 16983
rect 11805 16949 11839 16983
rect 11839 16949 11848 16983
rect 11796 16940 11848 16949
rect 12256 16983 12308 16992
rect 12256 16949 12265 16983
rect 12265 16949 12299 16983
rect 12299 16949 12308 16983
rect 12256 16940 12308 16949
rect 13268 16940 13320 16992
rect 13544 16940 13596 16992
rect 15660 16940 15712 16992
rect 17500 16940 17552 16992
rect 18052 16940 18104 16992
rect 19708 17017 19717 17051
rect 19717 17017 19751 17051
rect 19751 17017 19760 17051
rect 19708 17008 19760 17017
rect 19800 17051 19852 17060
rect 19800 17017 19809 17051
rect 19809 17017 19843 17051
rect 19843 17017 19852 17051
rect 19800 17008 19852 17017
rect 19064 16983 19116 16992
rect 19064 16949 19073 16983
rect 19073 16949 19107 16983
rect 19107 16949 19116 16983
rect 19064 16940 19116 16949
rect 8982 16838 9034 16890
rect 9046 16838 9098 16890
rect 9110 16838 9162 16890
rect 9174 16838 9226 16890
rect 16982 16838 17034 16890
rect 17046 16838 17098 16890
rect 17110 16838 17162 16890
rect 17174 16838 17226 16890
rect 1860 16779 1912 16788
rect 1860 16745 1869 16779
rect 1869 16745 1903 16779
rect 1903 16745 1912 16779
rect 1860 16736 1912 16745
rect 2780 16779 2832 16788
rect 2780 16745 2789 16779
rect 2789 16745 2823 16779
rect 2823 16745 2832 16779
rect 2780 16736 2832 16745
rect 4988 16779 5040 16788
rect 4988 16745 4997 16779
rect 4997 16745 5031 16779
rect 5031 16745 5040 16779
rect 4988 16736 5040 16745
rect 7196 16779 7248 16788
rect 7196 16745 7205 16779
rect 7205 16745 7239 16779
rect 7239 16745 7248 16779
rect 7196 16736 7248 16745
rect 7932 16779 7984 16788
rect 7932 16745 7941 16779
rect 7941 16745 7975 16779
rect 7975 16745 7984 16779
rect 7932 16736 7984 16745
rect 10692 16779 10744 16788
rect 10692 16745 10701 16779
rect 10701 16745 10735 16779
rect 10735 16745 10744 16779
rect 10692 16736 10744 16745
rect 10876 16736 10928 16788
rect 12256 16736 12308 16788
rect 12716 16779 12768 16788
rect 4160 16668 4212 16720
rect 5908 16711 5960 16720
rect 5908 16677 5917 16711
rect 5917 16677 5951 16711
rect 5951 16677 5960 16711
rect 5908 16668 5960 16677
rect 6000 16711 6052 16720
rect 6000 16677 6009 16711
rect 6009 16677 6043 16711
rect 6043 16677 6052 16711
rect 8208 16711 8260 16720
rect 6000 16668 6052 16677
rect 8208 16677 8217 16711
rect 8217 16677 8251 16711
rect 8251 16677 8260 16711
rect 8208 16668 8260 16677
rect 11520 16668 11572 16720
rect 12716 16745 12725 16779
rect 12725 16745 12759 16779
rect 12759 16745 12768 16779
rect 12716 16736 12768 16745
rect 14096 16736 14148 16788
rect 15844 16736 15896 16788
rect 16212 16736 16264 16788
rect 17316 16736 17368 16788
rect 19800 16779 19852 16788
rect 19800 16745 19809 16779
rect 19809 16745 19843 16779
rect 19843 16745 19852 16779
rect 19800 16736 19852 16745
rect 13268 16668 13320 16720
rect 17500 16668 17552 16720
rect 18972 16668 19024 16720
rect 1676 16600 1728 16652
rect 3148 16600 3200 16652
rect 9588 16643 9640 16652
rect 9588 16609 9597 16643
rect 9597 16609 9631 16643
rect 9631 16609 9640 16643
rect 9588 16600 9640 16609
rect 12532 16600 12584 16652
rect 4068 16575 4120 16584
rect 4068 16541 4077 16575
rect 4077 16541 4111 16575
rect 4111 16541 4120 16575
rect 4068 16532 4120 16541
rect 4804 16532 4856 16584
rect 7932 16532 7984 16584
rect 8576 16532 8628 16584
rect 11152 16532 11204 16584
rect 12164 16532 12216 16584
rect 11888 16464 11940 16516
rect 12900 16464 12952 16516
rect 15476 16600 15528 16652
rect 13360 16532 13412 16584
rect 17316 16600 17368 16652
rect 19064 16600 19116 16652
rect 20812 16600 20864 16652
rect 17500 16532 17552 16584
rect 19432 16532 19484 16584
rect 21088 16507 21140 16516
rect 21088 16473 21097 16507
rect 21097 16473 21131 16507
rect 21131 16473 21140 16507
rect 21088 16464 21140 16473
rect 6920 16439 6972 16448
rect 6920 16405 6929 16439
rect 6929 16405 6963 16439
rect 6963 16405 6972 16439
rect 6920 16396 6972 16405
rect 9312 16396 9364 16448
rect 15844 16396 15896 16448
rect 18328 16439 18380 16448
rect 18328 16405 18337 16439
rect 18337 16405 18371 16439
rect 18371 16405 18380 16439
rect 18328 16396 18380 16405
rect 4982 16294 5034 16346
rect 5046 16294 5098 16346
rect 5110 16294 5162 16346
rect 5174 16294 5226 16346
rect 12982 16294 13034 16346
rect 13046 16294 13098 16346
rect 13110 16294 13162 16346
rect 13174 16294 13226 16346
rect 20982 16294 21034 16346
rect 21046 16294 21098 16346
rect 21110 16294 21162 16346
rect 21174 16294 21226 16346
rect 1584 16167 1636 16176
rect 1584 16133 1593 16167
rect 1593 16133 1627 16167
rect 1627 16133 1636 16167
rect 1584 16124 1636 16133
rect 1952 16056 2004 16108
rect 4068 16192 4120 16244
rect 4160 16235 4212 16244
rect 4160 16201 4169 16235
rect 4169 16201 4203 16235
rect 4203 16201 4212 16235
rect 4804 16235 4856 16244
rect 4160 16192 4212 16201
rect 4804 16201 4813 16235
rect 4813 16201 4847 16235
rect 4847 16201 4856 16235
rect 4804 16192 4856 16201
rect 6000 16192 6052 16244
rect 7012 16192 7064 16244
rect 10968 16192 11020 16244
rect 11428 16192 11480 16244
rect 11796 16192 11848 16244
rect 12164 16235 12216 16244
rect 12164 16201 12173 16235
rect 12173 16201 12207 16235
rect 12207 16201 12216 16235
rect 12164 16192 12216 16201
rect 13360 16192 13412 16244
rect 15476 16235 15528 16244
rect 15476 16201 15485 16235
rect 15485 16201 15519 16235
rect 15519 16201 15528 16235
rect 15476 16192 15528 16201
rect 18972 16192 19024 16244
rect 19432 16235 19484 16244
rect 19432 16201 19441 16235
rect 19441 16201 19475 16235
rect 19475 16201 19484 16235
rect 19432 16192 19484 16201
rect 13268 16167 13320 16176
rect 13268 16133 13277 16167
rect 13277 16133 13311 16167
rect 13311 16133 13320 16167
rect 13268 16124 13320 16133
rect 4436 16056 4488 16108
rect 8116 16056 8168 16108
rect 9312 16056 9364 16108
rect 9588 16056 9640 16108
rect 15016 16124 15068 16176
rect 16396 16167 16448 16176
rect 16396 16133 16405 16167
rect 16405 16133 16439 16167
rect 16439 16133 16448 16167
rect 16396 16124 16448 16133
rect 19708 16124 19760 16176
rect 15844 16099 15896 16108
rect 15844 16065 15853 16099
rect 15853 16065 15887 16099
rect 15887 16065 15896 16099
rect 15844 16056 15896 16065
rect 18144 16099 18196 16108
rect 18144 16065 18153 16099
rect 18153 16065 18187 16099
rect 18187 16065 18196 16099
rect 18144 16056 18196 16065
rect 18328 16056 18380 16108
rect 18420 16099 18472 16108
rect 18420 16065 18429 16099
rect 18429 16065 18463 16099
rect 18463 16065 18472 16099
rect 18420 16056 18472 16065
rect 2320 15988 2372 16040
rect 3148 16031 3200 16040
rect 3148 15997 3157 16031
rect 3157 15997 3191 16031
rect 3191 15997 3200 16031
rect 3148 15988 3200 15997
rect 5448 15988 5500 16040
rect 10232 15988 10284 16040
rect 10784 15988 10836 16040
rect 11796 15988 11848 16040
rect 3608 15920 3660 15972
rect 4712 15920 4764 15972
rect 4804 15920 4856 15972
rect 6920 15963 6972 15972
rect 6920 15929 6929 15963
rect 6929 15929 6963 15963
rect 6963 15929 6972 15963
rect 6920 15920 6972 15929
rect 7012 15963 7064 15972
rect 7012 15929 7021 15963
rect 7021 15929 7055 15963
rect 7055 15929 7064 15963
rect 7012 15920 7064 15929
rect 8208 15920 8260 15972
rect 8760 15920 8812 15972
rect 9772 15920 9824 15972
rect 8668 15852 8720 15904
rect 9588 15852 9640 15904
rect 10968 15895 11020 15904
rect 10968 15861 10977 15895
rect 10977 15861 11011 15895
rect 11011 15861 11020 15895
rect 10968 15852 11020 15861
rect 16212 15920 16264 15972
rect 18328 15920 18380 15972
rect 18512 15920 18564 15972
rect 13268 15852 13320 15904
rect 13728 15852 13780 15904
rect 16672 15852 16724 15904
rect 17316 15852 17368 15904
rect 17500 15852 17552 15904
rect 17960 15852 18012 15904
rect 20812 15920 20864 15972
rect 8982 15750 9034 15802
rect 9046 15750 9098 15802
rect 9110 15750 9162 15802
rect 9174 15750 9226 15802
rect 16982 15750 17034 15802
rect 17046 15750 17098 15802
rect 17110 15750 17162 15802
rect 17174 15750 17226 15802
rect 1952 15691 2004 15700
rect 1952 15657 1961 15691
rect 1961 15657 1995 15691
rect 1995 15657 2004 15691
rect 1952 15648 2004 15657
rect 6920 15648 6972 15700
rect 8760 15691 8812 15700
rect 8760 15657 8769 15691
rect 8769 15657 8803 15691
rect 8803 15657 8812 15691
rect 8760 15648 8812 15657
rect 9312 15648 9364 15700
rect 10232 15691 10284 15700
rect 10232 15657 10241 15691
rect 10241 15657 10275 15691
rect 10275 15657 10284 15691
rect 10232 15648 10284 15657
rect 15660 15691 15712 15700
rect 15660 15657 15669 15691
rect 15669 15657 15703 15691
rect 15703 15657 15712 15691
rect 15660 15648 15712 15657
rect 16212 15691 16264 15700
rect 16212 15657 16221 15691
rect 16221 15657 16255 15691
rect 16255 15657 16264 15691
rect 16212 15648 16264 15657
rect 18144 15648 18196 15700
rect 22008 15648 22060 15700
rect 1308 15580 1360 15632
rect 5540 15580 5592 15632
rect 8484 15580 8536 15632
rect 18512 15580 18564 15632
rect 19708 15580 19760 15632
rect 2136 15512 2188 15564
rect 3056 15512 3108 15564
rect 4804 15512 4856 15564
rect 6000 15555 6052 15564
rect 6000 15521 6009 15555
rect 6009 15521 6043 15555
rect 6043 15521 6052 15555
rect 6000 15512 6052 15521
rect 6184 15555 6236 15564
rect 6184 15521 6193 15555
rect 6193 15521 6227 15555
rect 6227 15521 6236 15555
rect 6184 15512 6236 15521
rect 10416 15555 10468 15564
rect 6460 15487 6512 15496
rect 6460 15453 6469 15487
rect 6469 15453 6503 15487
rect 6503 15453 6512 15487
rect 6460 15444 6512 15453
rect 7840 15487 7892 15496
rect 7840 15453 7849 15487
rect 7849 15453 7883 15487
rect 7883 15453 7892 15487
rect 7840 15444 7892 15453
rect 10416 15521 10425 15555
rect 10425 15521 10459 15555
rect 10459 15521 10468 15555
rect 10416 15512 10468 15521
rect 12072 15512 12124 15564
rect 13544 15512 13596 15564
rect 17132 15555 17184 15564
rect 17132 15521 17150 15555
rect 17150 15521 17184 15555
rect 17132 15512 17184 15521
rect 17960 15512 18012 15564
rect 20812 15512 20864 15564
rect 10600 15444 10652 15496
rect 12624 15444 12676 15496
rect 14740 15444 14792 15496
rect 18696 15444 18748 15496
rect 1676 15376 1728 15428
rect 7932 15376 7984 15428
rect 16120 15376 16172 15428
rect 2320 15308 2372 15360
rect 7656 15308 7708 15360
rect 12532 15308 12584 15360
rect 14004 15351 14056 15360
rect 14004 15317 14013 15351
rect 14013 15317 14047 15351
rect 14047 15317 14056 15351
rect 14004 15308 14056 15317
rect 16488 15351 16540 15360
rect 16488 15317 16497 15351
rect 16497 15317 16531 15351
rect 16531 15317 16540 15351
rect 16488 15308 16540 15317
rect 19524 15351 19576 15360
rect 19524 15317 19533 15351
rect 19533 15317 19567 15351
rect 19567 15317 19576 15351
rect 19524 15308 19576 15317
rect 4982 15206 5034 15258
rect 5046 15206 5098 15258
rect 5110 15206 5162 15258
rect 5174 15206 5226 15258
rect 12982 15206 13034 15258
rect 13046 15206 13098 15258
rect 13110 15206 13162 15258
rect 13174 15206 13226 15258
rect 20982 15206 21034 15258
rect 21046 15206 21098 15258
rect 21110 15206 21162 15258
rect 21174 15206 21226 15258
rect 3056 15147 3108 15156
rect 3056 15113 3065 15147
rect 3065 15113 3099 15147
rect 3099 15113 3108 15147
rect 3056 15104 3108 15113
rect 5540 15104 5592 15156
rect 5908 15104 5960 15156
rect 6184 15011 6236 15020
rect 2320 14943 2372 14952
rect 2320 14909 2329 14943
rect 2329 14909 2363 14943
rect 2363 14909 2372 14943
rect 2320 14900 2372 14909
rect 1952 14807 2004 14816
rect 1952 14773 1961 14807
rect 1961 14773 1995 14807
rect 1995 14773 2004 14807
rect 3424 14900 3476 14952
rect 6184 14977 6193 15011
rect 6193 14977 6227 15011
rect 6227 14977 6236 15011
rect 6184 14968 6236 14977
rect 9772 15104 9824 15156
rect 13544 15147 13596 15156
rect 13544 15113 13553 15147
rect 13553 15113 13587 15147
rect 13587 15113 13596 15147
rect 13544 15104 13596 15113
rect 18328 15104 18380 15156
rect 20812 15104 20864 15156
rect 8208 15036 8260 15088
rect 9496 15036 9548 15088
rect 2780 14875 2832 14884
rect 2780 14841 2789 14875
rect 2789 14841 2823 14875
rect 2823 14841 2832 14875
rect 2780 14832 2832 14841
rect 5356 14832 5408 14884
rect 5540 14900 5592 14952
rect 7656 14943 7708 14952
rect 7656 14909 7665 14943
rect 7665 14909 7699 14943
rect 7699 14909 7708 14943
rect 7656 14900 7708 14909
rect 7840 14968 7892 15020
rect 12532 15011 12584 15020
rect 12532 14977 12541 15011
rect 12541 14977 12575 15011
rect 12575 14977 12584 15011
rect 12532 14968 12584 14977
rect 9496 14943 9548 14952
rect 6000 14832 6052 14884
rect 9496 14909 9505 14943
rect 9505 14909 9539 14943
rect 9539 14909 9548 14943
rect 9496 14900 9548 14909
rect 9772 14900 9824 14952
rect 10416 14900 10468 14952
rect 11244 14943 11296 14952
rect 11244 14909 11253 14943
rect 11253 14909 11287 14943
rect 11287 14909 11296 14943
rect 11244 14900 11296 14909
rect 14004 14943 14056 14952
rect 14004 14909 14013 14943
rect 14013 14909 14047 14943
rect 14047 14909 14056 14943
rect 14004 14900 14056 14909
rect 14556 14943 14608 14952
rect 14556 14909 14565 14943
rect 14565 14909 14599 14943
rect 14599 14909 14608 14943
rect 14556 14900 14608 14909
rect 15476 14900 15528 14952
rect 16488 14900 16540 14952
rect 18604 14900 18656 14952
rect 19524 14943 19576 14952
rect 19524 14909 19533 14943
rect 19533 14909 19567 14943
rect 19567 14909 19576 14943
rect 19524 14900 19576 14909
rect 10232 14875 10284 14884
rect 10232 14841 10241 14875
rect 10241 14841 10275 14875
rect 10275 14841 10284 14875
rect 10232 14832 10284 14841
rect 12624 14875 12676 14884
rect 12624 14841 12633 14875
rect 12633 14841 12667 14875
rect 12667 14841 12676 14875
rect 12624 14832 12676 14841
rect 13820 14832 13872 14884
rect 14740 14875 14792 14884
rect 1952 14764 2004 14773
rect 3884 14807 3936 14816
rect 3884 14773 3893 14807
rect 3893 14773 3927 14807
rect 3927 14773 3936 14807
rect 3884 14764 3936 14773
rect 4804 14807 4856 14816
rect 4804 14773 4813 14807
rect 4813 14773 4847 14807
rect 4847 14773 4856 14807
rect 4804 14764 4856 14773
rect 5448 14807 5500 14816
rect 5448 14773 5457 14807
rect 5457 14773 5491 14807
rect 5491 14773 5500 14807
rect 5448 14764 5500 14773
rect 8484 14764 8536 14816
rect 10968 14764 11020 14816
rect 11888 14764 11940 14816
rect 12072 14764 12124 14816
rect 13728 14764 13780 14816
rect 14740 14841 14749 14875
rect 14749 14841 14783 14875
rect 14783 14841 14792 14875
rect 14740 14832 14792 14841
rect 14648 14764 14700 14816
rect 15660 14764 15712 14816
rect 16580 14832 16632 14884
rect 17132 14832 17184 14884
rect 18696 14807 18748 14816
rect 18696 14773 18705 14807
rect 18705 14773 18739 14807
rect 18739 14773 18748 14807
rect 18696 14764 18748 14773
rect 19432 14807 19484 14816
rect 19432 14773 19441 14807
rect 19441 14773 19475 14807
rect 19475 14773 19484 14807
rect 19432 14764 19484 14773
rect 20444 14807 20496 14816
rect 20444 14773 20453 14807
rect 20453 14773 20487 14807
rect 20487 14773 20496 14807
rect 20444 14764 20496 14773
rect 20996 14764 21048 14816
rect 8982 14662 9034 14714
rect 9046 14662 9098 14714
rect 9110 14662 9162 14714
rect 9174 14662 9226 14714
rect 16982 14662 17034 14714
rect 17046 14662 17098 14714
rect 17110 14662 17162 14714
rect 17174 14662 17226 14714
rect 2596 14603 2648 14612
rect 2596 14569 2605 14603
rect 2605 14569 2639 14603
rect 2639 14569 2648 14603
rect 2596 14560 2648 14569
rect 3424 14560 3476 14612
rect 3700 14560 3752 14612
rect 4160 14560 4212 14612
rect 5356 14603 5408 14612
rect 5356 14569 5365 14603
rect 5365 14569 5399 14603
rect 5399 14569 5408 14603
rect 5356 14560 5408 14569
rect 7840 14603 7892 14612
rect 2320 14492 2372 14544
rect 7012 14535 7064 14544
rect 7012 14501 7021 14535
rect 7021 14501 7055 14535
rect 7055 14501 7064 14535
rect 7012 14492 7064 14501
rect 7840 14569 7849 14603
rect 7849 14569 7883 14603
rect 7883 14569 7892 14603
rect 7840 14560 7892 14569
rect 7932 14560 7984 14612
rect 3884 14424 3936 14476
rect 8760 14424 8812 14476
rect 2780 14356 2832 14408
rect 3792 14288 3844 14340
rect 1584 14263 1636 14272
rect 1584 14229 1593 14263
rect 1593 14229 1627 14263
rect 1627 14229 1636 14263
rect 1584 14220 1636 14229
rect 4528 14220 4580 14272
rect 6368 14220 6420 14272
rect 7472 14331 7524 14340
rect 7472 14297 7481 14331
rect 7481 14297 7515 14331
rect 7515 14297 7524 14331
rect 7472 14288 7524 14297
rect 10968 14492 11020 14544
rect 11888 14492 11940 14544
rect 12808 14560 12860 14612
rect 14740 14560 14792 14612
rect 17408 14560 17460 14612
rect 18512 14560 18564 14612
rect 18696 14560 18748 14612
rect 20444 14560 20496 14612
rect 12256 14535 12308 14544
rect 12256 14501 12265 14535
rect 12265 14501 12299 14535
rect 12299 14501 12308 14535
rect 12256 14492 12308 14501
rect 12624 14492 12676 14544
rect 13820 14535 13872 14544
rect 13820 14501 13829 14535
rect 13829 14501 13863 14535
rect 13863 14501 13872 14535
rect 15844 14535 15896 14544
rect 13820 14492 13872 14501
rect 15844 14501 15853 14535
rect 15853 14501 15887 14535
rect 15887 14501 15896 14535
rect 15844 14492 15896 14501
rect 16212 14492 16264 14544
rect 18420 14492 18472 14544
rect 18604 14535 18656 14544
rect 18604 14501 18613 14535
rect 18613 14501 18647 14535
rect 18647 14501 18656 14535
rect 18604 14492 18656 14501
rect 20720 14492 20772 14544
rect 20996 14535 21048 14544
rect 20996 14501 21005 14535
rect 21005 14501 21039 14535
rect 21039 14501 21048 14535
rect 20996 14492 21048 14501
rect 22192 14492 22244 14544
rect 10232 14467 10284 14476
rect 10232 14433 10241 14467
rect 10241 14433 10275 14467
rect 10275 14433 10284 14467
rect 10232 14424 10284 14433
rect 17868 14467 17920 14476
rect 17868 14433 17877 14467
rect 17877 14433 17911 14467
rect 17911 14433 17920 14467
rect 17868 14424 17920 14433
rect 12440 14399 12492 14408
rect 12440 14365 12449 14399
rect 12449 14365 12483 14399
rect 12483 14365 12492 14399
rect 12440 14356 12492 14365
rect 13728 14399 13780 14408
rect 13728 14365 13737 14399
rect 13737 14365 13771 14399
rect 13771 14365 13780 14399
rect 13728 14356 13780 14365
rect 13912 14356 13964 14408
rect 15752 14399 15804 14408
rect 15752 14365 15761 14399
rect 15761 14365 15795 14399
rect 15795 14365 15804 14399
rect 15752 14356 15804 14365
rect 17500 14356 17552 14408
rect 20352 14424 20404 14476
rect 20812 14356 20864 14408
rect 21272 14399 21324 14408
rect 21272 14365 21281 14399
rect 21281 14365 21315 14399
rect 21315 14365 21324 14399
rect 21272 14356 21324 14365
rect 12256 14288 12308 14340
rect 10600 14220 10652 14272
rect 19064 14263 19116 14272
rect 19064 14229 19073 14263
rect 19073 14229 19107 14263
rect 19107 14229 19116 14263
rect 19064 14220 19116 14229
rect 4982 14118 5034 14170
rect 5046 14118 5098 14170
rect 5110 14118 5162 14170
rect 5174 14118 5226 14170
rect 12982 14118 13034 14170
rect 13046 14118 13098 14170
rect 13110 14118 13162 14170
rect 13174 14118 13226 14170
rect 20982 14118 21034 14170
rect 21046 14118 21098 14170
rect 21110 14118 21162 14170
rect 21174 14118 21226 14170
rect 2596 14059 2648 14068
rect 2596 14025 2605 14059
rect 2605 14025 2639 14059
rect 2639 14025 2648 14059
rect 2596 14016 2648 14025
rect 2780 14016 2832 14068
rect 3884 14016 3936 14068
rect 4160 14016 4212 14068
rect 10232 14016 10284 14068
rect 10324 14059 10376 14068
rect 10324 14025 10333 14059
rect 10333 14025 10367 14059
rect 10367 14025 10376 14059
rect 10324 14016 10376 14025
rect 10968 14016 11020 14068
rect 12256 14016 12308 14068
rect 15752 14016 15804 14068
rect 17868 14059 17920 14068
rect 17868 14025 17877 14059
rect 17877 14025 17911 14059
rect 17911 14025 17920 14059
rect 17868 14016 17920 14025
rect 19156 14016 19208 14068
rect 20720 14059 20772 14068
rect 20720 14025 20729 14059
rect 20729 14025 20763 14059
rect 20763 14025 20772 14059
rect 20720 14016 20772 14025
rect 22192 14059 22244 14068
rect 22192 14025 22201 14059
rect 22201 14025 22235 14059
rect 22235 14025 22244 14059
rect 22192 14016 22244 14025
rect 2136 13991 2188 14000
rect 2136 13957 2145 13991
rect 2145 13957 2179 13991
rect 2179 13957 2188 13991
rect 2136 13948 2188 13957
rect 4252 13948 4304 14000
rect 1584 13923 1636 13932
rect 1584 13889 1593 13923
rect 1593 13889 1627 13923
rect 1627 13889 1636 13923
rect 1584 13880 1636 13889
rect 4620 13948 4672 14000
rect 4896 13812 4948 13864
rect 11244 13948 11296 14000
rect 12624 13948 12676 14000
rect 13820 13948 13872 14000
rect 15844 13991 15896 14000
rect 15844 13957 15853 13991
rect 15853 13957 15887 13991
rect 15887 13957 15896 13991
rect 15844 13948 15896 13957
rect 6460 13880 6512 13932
rect 9956 13923 10008 13932
rect 9956 13889 9965 13923
rect 9965 13889 9999 13923
rect 9999 13889 10008 13923
rect 9956 13880 10008 13889
rect 10324 13880 10376 13932
rect 12532 13880 12584 13932
rect 15476 13923 15528 13932
rect 15476 13889 15485 13923
rect 15485 13889 15519 13923
rect 15519 13889 15528 13923
rect 15476 13880 15528 13889
rect 18788 13880 18840 13932
rect 19064 13923 19116 13932
rect 19064 13889 19073 13923
rect 19073 13889 19107 13923
rect 19107 13889 19116 13923
rect 19064 13880 19116 13889
rect 20352 13923 20404 13932
rect 20352 13889 20361 13923
rect 20361 13889 20395 13923
rect 20395 13889 20404 13923
rect 20352 13880 20404 13889
rect 21272 13923 21324 13932
rect 21272 13889 21281 13923
rect 21281 13889 21315 13923
rect 21315 13889 21324 13923
rect 21272 13880 21324 13889
rect 10416 13855 10468 13864
rect 10416 13821 10425 13855
rect 10425 13821 10459 13855
rect 10459 13821 10468 13855
rect 10416 13812 10468 13821
rect 14740 13855 14792 13864
rect 14740 13821 14749 13855
rect 14749 13821 14783 13855
rect 14783 13821 14792 13855
rect 14740 13812 14792 13821
rect 18052 13855 18104 13864
rect 2044 13744 2096 13796
rect 3884 13787 3936 13796
rect 3884 13753 3893 13787
rect 3893 13753 3927 13787
rect 3927 13753 3936 13787
rect 3884 13744 3936 13753
rect 4252 13744 4304 13796
rect 11336 13744 11388 13796
rect 6276 13676 6328 13728
rect 7840 13676 7892 13728
rect 8668 13719 8720 13728
rect 8668 13685 8677 13719
rect 8677 13685 8711 13719
rect 8711 13685 8720 13719
rect 8668 13676 8720 13685
rect 10140 13676 10192 13728
rect 12440 13676 12492 13728
rect 12624 13787 12676 13796
rect 12624 13753 12633 13787
rect 12633 13753 12667 13787
rect 12667 13753 12676 13787
rect 12624 13744 12676 13753
rect 13176 13676 13228 13728
rect 13728 13676 13780 13728
rect 14556 13719 14608 13728
rect 14556 13685 14565 13719
rect 14565 13685 14599 13719
rect 14599 13685 14608 13719
rect 18052 13821 18096 13855
rect 18096 13821 18104 13855
rect 18052 13812 18104 13821
rect 17500 13719 17552 13728
rect 14556 13676 14608 13685
rect 17500 13685 17509 13719
rect 17509 13685 17543 13719
rect 17543 13685 17552 13719
rect 17500 13676 17552 13685
rect 17592 13676 17644 13728
rect 18880 13719 18932 13728
rect 18880 13685 18889 13719
rect 18889 13685 18923 13719
rect 18923 13685 18932 13719
rect 19432 13812 19484 13864
rect 20628 13744 20680 13796
rect 20996 13787 21048 13796
rect 20996 13753 21005 13787
rect 21005 13753 21039 13787
rect 21039 13753 21048 13787
rect 20996 13744 21048 13753
rect 18880 13676 18932 13685
rect 20812 13676 20864 13728
rect 21088 13676 21140 13728
rect 8982 13574 9034 13626
rect 9046 13574 9098 13626
rect 9110 13574 9162 13626
rect 9174 13574 9226 13626
rect 16982 13574 17034 13626
rect 17046 13574 17098 13626
rect 17110 13574 17162 13626
rect 17174 13574 17226 13626
rect 2044 13472 2096 13524
rect 3884 13472 3936 13524
rect 6368 13472 6420 13524
rect 6460 13472 6512 13524
rect 9956 13472 10008 13524
rect 11336 13472 11388 13524
rect 12808 13515 12860 13524
rect 12808 13481 12817 13515
rect 12817 13481 12851 13515
rect 12851 13481 12860 13515
rect 12808 13472 12860 13481
rect 14740 13515 14792 13524
rect 14740 13481 14749 13515
rect 14749 13481 14783 13515
rect 14783 13481 14792 13515
rect 14740 13472 14792 13481
rect 1860 13404 1912 13456
rect 2504 13404 2556 13456
rect 4528 13447 4580 13456
rect 4528 13413 4537 13447
rect 4537 13413 4571 13447
rect 4571 13413 4580 13447
rect 4528 13404 4580 13413
rect 7012 13404 7064 13456
rect 7840 13404 7892 13456
rect 10416 13447 10468 13456
rect 10416 13413 10425 13447
rect 10425 13413 10459 13447
rect 10459 13413 10468 13447
rect 10416 13404 10468 13413
rect 13176 13404 13228 13456
rect 6184 13336 6236 13388
rect 7656 13336 7708 13388
rect 9588 13336 9640 13388
rect 9772 13336 9824 13388
rect 11888 13379 11940 13388
rect 11888 13345 11897 13379
rect 11897 13345 11931 13379
rect 11931 13345 11940 13379
rect 11888 13336 11940 13345
rect 13728 13379 13780 13388
rect 13728 13345 13737 13379
rect 13737 13345 13771 13379
rect 13771 13345 13780 13379
rect 13728 13336 13780 13345
rect 14188 13379 14240 13388
rect 14188 13345 14197 13379
rect 14197 13345 14231 13379
rect 14231 13345 14240 13379
rect 14188 13336 14240 13345
rect 2136 13268 2188 13320
rect 4436 13311 4488 13320
rect 4436 13277 4445 13311
rect 4445 13277 4479 13311
rect 4479 13277 4488 13311
rect 4436 13268 4488 13277
rect 4252 13200 4304 13252
rect 6276 13268 6328 13320
rect 7288 13311 7340 13320
rect 7288 13277 7297 13311
rect 7297 13277 7331 13311
rect 7331 13277 7340 13311
rect 7288 13268 7340 13277
rect 14280 13311 14332 13320
rect 14280 13277 14289 13311
rect 14289 13277 14323 13311
rect 14323 13277 14332 13311
rect 14280 13268 14332 13277
rect 11888 13200 11940 13252
rect 17684 13472 17736 13524
rect 18512 13515 18564 13524
rect 18512 13481 18521 13515
rect 18521 13481 18555 13515
rect 18555 13481 18564 13515
rect 18512 13472 18564 13481
rect 19340 13472 19392 13524
rect 20996 13472 21048 13524
rect 16028 13447 16080 13456
rect 16028 13413 16037 13447
rect 16037 13413 16071 13447
rect 16071 13413 16080 13447
rect 16028 13404 16080 13413
rect 21088 13447 21140 13456
rect 21088 13413 21097 13447
rect 21097 13413 21131 13447
rect 21131 13413 21140 13447
rect 21088 13404 21140 13413
rect 17500 13379 17552 13388
rect 17500 13345 17509 13379
rect 17509 13345 17543 13379
rect 17543 13345 17552 13379
rect 17500 13336 17552 13345
rect 15936 13311 15988 13320
rect 15936 13277 15945 13311
rect 15945 13277 15979 13311
rect 15979 13277 15988 13311
rect 15936 13268 15988 13277
rect 17592 13268 17644 13320
rect 17960 13200 18012 13252
rect 6460 13175 6512 13184
rect 6460 13141 6469 13175
rect 6469 13141 6503 13175
rect 6503 13141 6512 13175
rect 6460 13132 6512 13141
rect 8668 13175 8720 13184
rect 8668 13141 8677 13175
rect 8677 13141 8711 13175
rect 8711 13141 8720 13175
rect 8668 13132 8720 13141
rect 12440 13175 12492 13184
rect 12440 13141 12449 13175
rect 12449 13141 12483 13175
rect 12483 13141 12492 13175
rect 12440 13132 12492 13141
rect 16120 13132 16172 13184
rect 17408 13132 17460 13184
rect 19064 13311 19116 13320
rect 19064 13277 19073 13311
rect 19073 13277 19107 13311
rect 19107 13277 19116 13311
rect 19064 13268 19116 13277
rect 21272 13311 21324 13320
rect 21272 13277 21281 13311
rect 21281 13277 21315 13311
rect 21315 13277 21324 13311
rect 21272 13268 21324 13277
rect 21364 13200 21416 13252
rect 20628 13175 20680 13184
rect 20628 13141 20637 13175
rect 20637 13141 20671 13175
rect 20671 13141 20680 13175
rect 20628 13132 20680 13141
rect 4982 13030 5034 13082
rect 5046 13030 5098 13082
rect 5110 13030 5162 13082
rect 5174 13030 5226 13082
rect 12982 13030 13034 13082
rect 13046 13030 13098 13082
rect 13110 13030 13162 13082
rect 13174 13030 13226 13082
rect 20982 13030 21034 13082
rect 21046 13030 21098 13082
rect 21110 13030 21162 13082
rect 21174 13030 21226 13082
rect 3608 12971 3660 12980
rect 3608 12937 3617 12971
rect 3617 12937 3651 12971
rect 3651 12937 3660 12971
rect 3608 12928 3660 12937
rect 4528 12928 4580 12980
rect 5632 12928 5684 12980
rect 9588 12928 9640 12980
rect 4436 12860 4488 12912
rect 7472 12903 7524 12912
rect 7472 12869 7481 12903
rect 7481 12869 7515 12903
rect 7515 12869 7524 12903
rect 7472 12860 7524 12869
rect 10140 12860 10192 12912
rect 11888 12903 11940 12912
rect 11888 12869 11897 12903
rect 11897 12869 11931 12903
rect 11931 12869 11940 12903
rect 11888 12860 11940 12869
rect 12440 12928 12492 12980
rect 13728 12928 13780 12980
rect 14188 12860 14240 12912
rect 16028 12928 16080 12980
rect 17500 12860 17552 12912
rect 2136 12835 2188 12844
rect 2136 12801 2145 12835
rect 2145 12801 2179 12835
rect 2179 12801 2188 12835
rect 2136 12792 2188 12801
rect 6460 12792 6512 12844
rect 7932 12792 7984 12844
rect 14280 12835 14332 12844
rect 1676 12767 1728 12776
rect 1676 12733 1685 12767
rect 1685 12733 1719 12767
rect 1719 12733 1728 12767
rect 1676 12724 1728 12733
rect 1952 12767 2004 12776
rect 1952 12733 1961 12767
rect 1961 12733 1995 12767
rect 1995 12733 2004 12767
rect 1952 12724 2004 12733
rect 3608 12724 3660 12776
rect 4804 12724 4856 12776
rect 5632 12767 5684 12776
rect 5632 12733 5641 12767
rect 5641 12733 5675 12767
rect 5675 12733 5684 12767
rect 5632 12724 5684 12733
rect 8668 12767 8720 12776
rect 8668 12733 8677 12767
rect 8677 12733 8711 12767
rect 8711 12733 8720 12767
rect 8668 12724 8720 12733
rect 14280 12801 14289 12835
rect 14289 12801 14323 12835
rect 14323 12801 14332 12835
rect 14280 12792 14332 12801
rect 16120 12835 16172 12844
rect 16120 12801 16129 12835
rect 16129 12801 16163 12835
rect 16163 12801 16172 12835
rect 16120 12792 16172 12801
rect 10600 12767 10652 12776
rect 4252 12699 4304 12708
rect 4252 12665 4261 12699
rect 4261 12665 4295 12699
rect 4295 12665 4304 12699
rect 4252 12656 4304 12665
rect 7012 12699 7064 12708
rect 7012 12665 7021 12699
rect 7021 12665 7055 12699
rect 7055 12665 7064 12699
rect 7012 12656 7064 12665
rect 10600 12733 10609 12767
rect 10609 12733 10643 12767
rect 10643 12733 10652 12767
rect 10600 12724 10652 12733
rect 10232 12656 10284 12708
rect 12348 12724 12400 12776
rect 15844 12724 15896 12776
rect 17960 12860 18012 12912
rect 18788 12835 18840 12844
rect 18788 12801 18797 12835
rect 18797 12801 18831 12835
rect 18831 12801 18840 12835
rect 18788 12792 18840 12801
rect 18512 12767 18564 12776
rect 18512 12733 18521 12767
rect 18521 12733 18555 12767
rect 18555 12733 18564 12767
rect 18512 12724 18564 12733
rect 11244 12656 11296 12708
rect 11336 12656 11388 12708
rect 2872 12588 2924 12640
rect 3424 12588 3476 12640
rect 6184 12631 6236 12640
rect 6184 12597 6193 12631
rect 6193 12597 6227 12631
rect 6227 12597 6236 12631
rect 6184 12588 6236 12597
rect 7196 12588 7248 12640
rect 8852 12631 8904 12640
rect 8852 12597 8861 12631
rect 8861 12597 8895 12631
rect 8895 12597 8904 12631
rect 8852 12588 8904 12597
rect 9680 12631 9732 12640
rect 9680 12597 9689 12631
rect 9689 12597 9723 12631
rect 9723 12597 9732 12631
rect 13728 12631 13780 12640
rect 9680 12588 9732 12597
rect 13728 12597 13737 12631
rect 13737 12597 13771 12631
rect 13771 12597 13780 12631
rect 13728 12588 13780 12597
rect 16764 12699 16816 12708
rect 14648 12631 14700 12640
rect 14648 12597 14657 12631
rect 14657 12597 14691 12631
rect 14691 12597 14700 12631
rect 14648 12588 14700 12597
rect 16028 12588 16080 12640
rect 16764 12665 16773 12699
rect 16773 12665 16807 12699
rect 16807 12665 16816 12699
rect 16764 12656 16816 12665
rect 19800 12699 19852 12708
rect 19800 12665 19809 12699
rect 19809 12665 19843 12699
rect 19843 12665 19852 12699
rect 19800 12656 19852 12665
rect 20812 12928 20864 12980
rect 21916 12971 21968 12980
rect 21916 12937 21925 12971
rect 21925 12937 21959 12971
rect 21959 12937 21968 12971
rect 21916 12928 21968 12937
rect 23572 12860 23624 12912
rect 21916 12724 21968 12776
rect 17408 12588 17460 12640
rect 18880 12588 18932 12640
rect 19432 12588 19484 12640
rect 21364 12656 21416 12708
rect 8982 12486 9034 12538
rect 9046 12486 9098 12538
rect 9110 12486 9162 12538
rect 9174 12486 9226 12538
rect 16982 12486 17034 12538
rect 17046 12486 17098 12538
rect 17110 12486 17162 12538
rect 17174 12486 17226 12538
rect 1584 12384 1636 12436
rect 1676 12384 1728 12436
rect 4436 12384 4488 12436
rect 6276 12427 6328 12436
rect 6276 12393 6285 12427
rect 6285 12393 6319 12427
rect 6319 12393 6328 12427
rect 6276 12384 6328 12393
rect 7840 12427 7892 12436
rect 7840 12393 7849 12427
rect 7849 12393 7883 12427
rect 7883 12393 7892 12427
rect 7840 12384 7892 12393
rect 7932 12384 7984 12436
rect 8852 12427 8904 12436
rect 8852 12393 8861 12427
rect 8861 12393 8895 12427
rect 8895 12393 8904 12427
rect 8852 12384 8904 12393
rect 10600 12384 10652 12436
rect 14280 12427 14332 12436
rect 1860 12359 1912 12368
rect 1860 12325 1869 12359
rect 1869 12325 1903 12359
rect 1903 12325 1912 12359
rect 1860 12316 1912 12325
rect 4252 12359 4304 12368
rect 4252 12325 4261 12359
rect 4261 12325 4295 12359
rect 4295 12325 4304 12359
rect 4252 12316 4304 12325
rect 7196 12316 7248 12368
rect 9588 12316 9640 12368
rect 11336 12316 11388 12368
rect 13452 12316 13504 12368
rect 14280 12393 14289 12427
rect 14289 12393 14323 12427
rect 14323 12393 14332 12427
rect 14280 12384 14332 12393
rect 15936 12427 15988 12436
rect 15936 12393 15945 12427
rect 15945 12393 15979 12427
rect 15979 12393 15988 12427
rect 15936 12384 15988 12393
rect 17408 12384 17460 12436
rect 19064 12427 19116 12436
rect 19064 12393 19073 12427
rect 19073 12393 19107 12427
rect 19107 12393 19116 12427
rect 19064 12384 19116 12393
rect 19800 12384 19852 12436
rect 21364 12427 21416 12436
rect 21364 12393 21373 12427
rect 21373 12393 21407 12427
rect 21407 12393 21416 12427
rect 21364 12384 21416 12393
rect 16212 12359 16264 12368
rect 16212 12325 16221 12359
rect 16221 12325 16255 12359
rect 16255 12325 16264 12359
rect 17776 12359 17828 12368
rect 16212 12316 16264 12325
rect 17776 12325 17785 12359
rect 17785 12325 17819 12359
rect 17819 12325 17828 12359
rect 17776 12316 17828 12325
rect 19432 12359 19484 12368
rect 19432 12325 19441 12359
rect 19441 12325 19475 12359
rect 19475 12325 19484 12359
rect 19432 12316 19484 12325
rect 2872 12291 2924 12300
rect 2872 12257 2881 12291
rect 2881 12257 2915 12291
rect 2915 12257 2924 12291
rect 2872 12248 2924 12257
rect 6000 12248 6052 12300
rect 8392 12248 8444 12300
rect 10416 12291 10468 12300
rect 10416 12257 10425 12291
rect 10425 12257 10459 12291
rect 10459 12257 10468 12291
rect 10416 12248 10468 12257
rect 16764 12291 16816 12300
rect 16764 12257 16773 12291
rect 16773 12257 16807 12291
rect 16807 12257 16816 12291
rect 16764 12248 16816 12257
rect 20352 12248 20404 12300
rect 20812 12248 20864 12300
rect 2596 12180 2648 12232
rect 3148 12223 3200 12232
rect 3148 12189 3157 12223
rect 3157 12189 3191 12223
rect 3191 12189 3200 12223
rect 3148 12180 3200 12189
rect 3424 12180 3476 12232
rect 4160 12223 4212 12232
rect 4160 12189 4169 12223
rect 4169 12189 4203 12223
rect 4203 12189 4212 12223
rect 4620 12223 4672 12232
rect 4160 12180 4212 12189
rect 4620 12189 4629 12223
rect 4629 12189 4663 12223
rect 4663 12189 4672 12223
rect 4620 12180 4672 12189
rect 6276 12180 6328 12232
rect 7288 12180 7340 12232
rect 9772 12223 9824 12232
rect 9772 12189 9781 12223
rect 9781 12189 9815 12223
rect 9815 12189 9824 12223
rect 9772 12180 9824 12189
rect 11244 12223 11296 12232
rect 11244 12189 11253 12223
rect 11253 12189 11287 12223
rect 11287 12189 11296 12223
rect 11244 12180 11296 12189
rect 13820 12180 13872 12232
rect 16120 12223 16172 12232
rect 16120 12189 16129 12223
rect 16129 12189 16163 12223
rect 16163 12189 16172 12223
rect 16120 12180 16172 12189
rect 13636 12155 13688 12164
rect 13636 12121 13645 12155
rect 13645 12121 13679 12155
rect 13679 12121 13688 12155
rect 13636 12112 13688 12121
rect 17684 12223 17736 12232
rect 17684 12189 17693 12223
rect 17693 12189 17727 12223
rect 17727 12189 17736 12223
rect 17684 12180 17736 12189
rect 17960 12223 18012 12232
rect 17960 12189 17969 12223
rect 17969 12189 18003 12223
rect 18003 12189 18012 12223
rect 17960 12180 18012 12189
rect 20076 12180 20128 12232
rect 20628 12112 20680 12164
rect 5540 12044 5592 12096
rect 6552 12087 6604 12096
rect 6552 12053 6561 12087
rect 6561 12053 6595 12087
rect 6595 12053 6604 12087
rect 6552 12044 6604 12053
rect 12164 12087 12216 12096
rect 12164 12053 12173 12087
rect 12173 12053 12207 12087
rect 12207 12053 12216 12087
rect 12164 12044 12216 12053
rect 12532 12087 12584 12096
rect 12532 12053 12541 12087
rect 12541 12053 12575 12087
rect 12575 12053 12584 12087
rect 12532 12044 12584 12053
rect 13360 12044 13412 12096
rect 14556 12044 14608 12096
rect 18420 12044 18472 12096
rect 4982 11942 5034 11994
rect 5046 11942 5098 11994
rect 5110 11942 5162 11994
rect 5174 11942 5226 11994
rect 12982 11942 13034 11994
rect 13046 11942 13098 11994
rect 13110 11942 13162 11994
rect 13174 11942 13226 11994
rect 20982 11942 21034 11994
rect 21046 11942 21098 11994
rect 21110 11942 21162 11994
rect 21174 11942 21226 11994
rect 1860 11840 1912 11892
rect 3516 11840 3568 11892
rect 4252 11840 4304 11892
rect 7196 11840 7248 11892
rect 9588 11883 9640 11892
rect 9588 11849 9597 11883
rect 9597 11849 9631 11883
rect 9631 11849 9640 11883
rect 9588 11840 9640 11849
rect 9772 11840 9824 11892
rect 10232 11883 10284 11892
rect 10232 11849 10241 11883
rect 10241 11849 10275 11883
rect 10275 11849 10284 11883
rect 10232 11840 10284 11849
rect 11244 11840 11296 11892
rect 12164 11883 12216 11892
rect 12164 11849 12173 11883
rect 12173 11849 12207 11883
rect 12207 11849 12216 11883
rect 12164 11840 12216 11849
rect 14648 11883 14700 11892
rect 14648 11849 14657 11883
rect 14657 11849 14691 11883
rect 14691 11849 14700 11883
rect 14648 11840 14700 11849
rect 16120 11840 16172 11892
rect 17776 11840 17828 11892
rect 19432 11883 19484 11892
rect 19432 11849 19441 11883
rect 19441 11849 19475 11883
rect 19475 11849 19484 11883
rect 19432 11840 19484 11849
rect 20076 11883 20128 11892
rect 20076 11849 20085 11883
rect 20085 11849 20119 11883
rect 20119 11849 20128 11883
rect 20076 11840 20128 11849
rect 20812 11840 20864 11892
rect 3148 11747 3200 11756
rect 3148 11713 3157 11747
rect 3157 11713 3191 11747
rect 3191 11713 3200 11747
rect 3148 11704 3200 11713
rect 6000 11772 6052 11824
rect 8576 11772 8628 11824
rect 6552 11704 6604 11756
rect 8852 11704 8904 11756
rect 10416 11772 10468 11824
rect 13636 11772 13688 11824
rect 5540 11636 5592 11688
rect 5724 11679 5776 11688
rect 5724 11645 5733 11679
rect 5733 11645 5767 11679
rect 5767 11645 5776 11679
rect 5724 11636 5776 11645
rect 10508 11679 10560 11688
rect 10508 11645 10517 11679
rect 10517 11645 10551 11679
rect 10551 11645 10560 11679
rect 10508 11636 10560 11645
rect 16212 11704 16264 11756
rect 14832 11679 14884 11688
rect 14832 11645 14841 11679
rect 14841 11645 14875 11679
rect 14875 11645 14884 11679
rect 14832 11636 14884 11645
rect 15844 11636 15896 11688
rect 16856 11636 16908 11688
rect 18420 11636 18472 11688
rect 20720 11679 20772 11688
rect 20720 11645 20729 11679
rect 20729 11645 20763 11679
rect 20763 11645 20772 11679
rect 20720 11636 20772 11645
rect 21548 11636 21600 11688
rect 2872 11568 2924 11620
rect 3516 11611 3568 11620
rect 112 11500 164 11552
rect 3516 11577 3519 11611
rect 3519 11577 3553 11611
rect 3553 11577 3568 11611
rect 3516 11568 3568 11577
rect 11152 11611 11204 11620
rect 8116 11500 8168 11552
rect 8392 11543 8444 11552
rect 8392 11509 8401 11543
rect 8401 11509 8435 11543
rect 8435 11509 8444 11543
rect 8392 11500 8444 11509
rect 11152 11577 11161 11611
rect 11161 11577 11195 11611
rect 11195 11577 11204 11611
rect 11152 11568 11204 11577
rect 12532 11611 12584 11620
rect 12532 11577 12541 11611
rect 12541 11577 12575 11611
rect 12575 11577 12584 11611
rect 12532 11568 12584 11577
rect 11244 11500 11296 11552
rect 12164 11500 12216 11552
rect 14648 11568 14700 11620
rect 15752 11568 15804 11620
rect 18880 11568 18932 11620
rect 13452 11543 13504 11552
rect 13452 11509 13461 11543
rect 13461 11509 13495 11543
rect 13495 11509 13504 11543
rect 13452 11500 13504 11509
rect 13820 11543 13872 11552
rect 13820 11509 13829 11543
rect 13829 11509 13863 11543
rect 13863 11509 13872 11543
rect 13820 11500 13872 11509
rect 8982 11398 9034 11450
rect 9046 11398 9098 11450
rect 9110 11398 9162 11450
rect 9174 11398 9226 11450
rect 16982 11398 17034 11450
rect 17046 11398 17098 11450
rect 17110 11398 17162 11450
rect 17174 11398 17226 11450
rect 3148 11296 3200 11348
rect 4160 11296 4212 11348
rect 6276 11339 6328 11348
rect 6276 11305 6285 11339
rect 6285 11305 6319 11339
rect 6319 11305 6328 11339
rect 6276 11296 6328 11305
rect 7196 11296 7248 11348
rect 8116 11296 8168 11348
rect 9588 11296 9640 11348
rect 9772 11296 9824 11348
rect 13452 11296 13504 11348
rect 17684 11296 17736 11348
rect 2320 11228 2372 11280
rect 3056 11228 3108 11280
rect 5356 11228 5408 11280
rect 2780 11160 2832 11212
rect 4712 11160 4764 11212
rect 5540 11160 5592 11212
rect 6000 11160 6052 11212
rect 7656 11228 7708 11280
rect 11336 11228 11388 11280
rect 14832 11271 14884 11280
rect 14832 11237 14841 11271
rect 14841 11237 14875 11271
rect 14875 11237 14884 11271
rect 14832 11228 14884 11237
rect 18420 11271 18472 11280
rect 18420 11237 18429 11271
rect 18429 11237 18463 11271
rect 18463 11237 18472 11271
rect 18420 11228 18472 11237
rect 6828 11203 6880 11212
rect 6828 11169 6837 11203
rect 6837 11169 6871 11203
rect 6871 11169 6880 11203
rect 6828 11160 6880 11169
rect 8116 11160 8168 11212
rect 8576 11160 8628 11212
rect 11152 11160 11204 11212
rect 13636 11203 13688 11212
rect 13636 11169 13645 11203
rect 13645 11169 13679 11203
rect 13679 11169 13688 11203
rect 13636 11160 13688 11169
rect 14188 11203 14240 11212
rect 14188 11169 14197 11203
rect 14197 11169 14231 11203
rect 14231 11169 14240 11203
rect 14188 11160 14240 11169
rect 15200 11160 15252 11212
rect 16212 11160 16264 11212
rect 17500 11160 17552 11212
rect 18144 11203 18196 11212
rect 18144 11169 18153 11203
rect 18153 11169 18187 11203
rect 18187 11169 18196 11203
rect 18144 11160 18196 11169
rect 19432 11203 19484 11212
rect 19432 11169 19450 11203
rect 19450 11169 19484 11203
rect 19432 11160 19484 11169
rect 20352 11160 20404 11212
rect 3148 11135 3200 11144
rect 3148 11101 3157 11135
rect 3157 11101 3191 11135
rect 3191 11101 3200 11135
rect 3148 11092 3200 11101
rect 6920 11135 6972 11144
rect 6920 11101 6929 11135
rect 6929 11101 6963 11135
rect 6963 11101 6972 11135
rect 6920 11092 6972 11101
rect 4804 11024 4856 11076
rect 5448 11067 5500 11076
rect 5448 11033 5457 11067
rect 5457 11033 5491 11067
rect 5491 11033 5500 11067
rect 5448 11024 5500 11033
rect 1768 10956 1820 11008
rect 2596 10956 2648 11008
rect 3516 10956 3568 11008
rect 4252 10999 4304 11008
rect 4252 10965 4261 10999
rect 4261 10965 4295 10999
rect 4295 10965 4304 10999
rect 4252 10956 4304 10965
rect 7748 10999 7800 11008
rect 7748 10965 7757 10999
rect 7757 10965 7791 10999
rect 7791 10965 7800 10999
rect 7748 10956 7800 10965
rect 7932 10956 7984 11008
rect 10508 10999 10560 11008
rect 10508 10965 10517 10999
rect 10517 10965 10551 10999
rect 10551 10965 10560 10999
rect 10508 10956 10560 10965
rect 12348 10956 12400 11008
rect 13728 10956 13780 11008
rect 16580 10956 16632 11008
rect 19616 10956 19668 11008
rect 19800 10999 19852 11008
rect 19800 10965 19809 10999
rect 19809 10965 19843 10999
rect 19843 10965 19852 10999
rect 19800 10956 19852 10965
rect 4982 10854 5034 10906
rect 5046 10854 5098 10906
rect 5110 10854 5162 10906
rect 5174 10854 5226 10906
rect 12982 10854 13034 10906
rect 13046 10854 13098 10906
rect 13110 10854 13162 10906
rect 13174 10854 13226 10906
rect 20982 10854 21034 10906
rect 21046 10854 21098 10906
rect 21110 10854 21162 10906
rect 21174 10854 21226 10906
rect 2228 10752 2280 10804
rect 3608 10752 3660 10804
rect 5356 10752 5408 10804
rect 8116 10795 8168 10804
rect 8116 10761 8125 10795
rect 8125 10761 8159 10795
rect 8159 10761 8168 10795
rect 8116 10752 8168 10761
rect 2780 10727 2832 10736
rect 2780 10693 2789 10727
rect 2789 10693 2823 10727
rect 2823 10693 2832 10727
rect 2780 10684 2832 10693
rect 4712 10684 4764 10736
rect 6828 10684 6880 10736
rect 1768 10659 1820 10668
rect 1768 10625 1777 10659
rect 1777 10625 1811 10659
rect 1811 10625 1820 10659
rect 1768 10616 1820 10625
rect 3608 10616 3660 10668
rect 4252 10659 4304 10668
rect 4252 10625 4261 10659
rect 4261 10625 4295 10659
rect 4295 10625 4304 10659
rect 4252 10616 4304 10625
rect 7472 10659 7524 10668
rect 7472 10625 7481 10659
rect 7481 10625 7515 10659
rect 7515 10625 7524 10659
rect 7472 10616 7524 10625
rect 5448 10548 5500 10600
rect 9312 10591 9364 10600
rect 9312 10557 9321 10591
rect 9321 10557 9355 10591
rect 9355 10557 9364 10591
rect 9312 10548 9364 10557
rect 10232 10752 10284 10804
rect 11152 10752 11204 10804
rect 11980 10752 12032 10804
rect 13452 10752 13504 10804
rect 16856 10752 16908 10804
rect 17684 10752 17736 10804
rect 19432 10795 19484 10804
rect 19432 10761 19441 10795
rect 19441 10761 19475 10795
rect 19475 10761 19484 10795
rect 19432 10752 19484 10761
rect 21272 10795 21324 10804
rect 21272 10761 21281 10795
rect 21281 10761 21315 10795
rect 21315 10761 21324 10795
rect 21272 10752 21324 10761
rect 12808 10659 12860 10668
rect 12808 10625 12817 10659
rect 12817 10625 12851 10659
rect 12851 10625 12860 10659
rect 12808 10616 12860 10625
rect 13820 10616 13872 10668
rect 2228 10480 2280 10532
rect 4436 10480 4488 10532
rect 7196 10523 7248 10532
rect 7196 10489 7205 10523
rect 7205 10489 7239 10523
rect 7239 10489 7248 10523
rect 7196 10480 7248 10489
rect 7656 10480 7708 10532
rect 10048 10523 10100 10532
rect 10048 10489 10057 10523
rect 10057 10489 10091 10523
rect 10091 10489 10100 10523
rect 10048 10480 10100 10489
rect 12348 10480 12400 10532
rect 3056 10455 3108 10464
rect 3056 10421 3065 10455
rect 3065 10421 3099 10455
rect 3099 10421 3108 10455
rect 3056 10412 3108 10421
rect 6000 10455 6052 10464
rect 6000 10421 6009 10455
rect 6009 10421 6043 10455
rect 6043 10421 6052 10455
rect 6000 10412 6052 10421
rect 11152 10455 11204 10464
rect 11152 10421 11161 10455
rect 11161 10421 11195 10455
rect 11195 10421 11204 10455
rect 11152 10412 11204 10421
rect 11704 10412 11756 10464
rect 12164 10455 12216 10464
rect 12164 10421 12173 10455
rect 12173 10421 12207 10455
rect 12207 10421 12216 10455
rect 13176 10480 13228 10532
rect 14188 10548 14240 10600
rect 16764 10616 16816 10668
rect 17500 10616 17552 10668
rect 19616 10659 19668 10668
rect 19616 10625 19625 10659
rect 19625 10625 19659 10659
rect 19659 10625 19668 10659
rect 19616 10616 19668 10625
rect 19892 10659 19944 10668
rect 19892 10625 19901 10659
rect 19901 10625 19935 10659
rect 19935 10625 19944 10659
rect 19892 10616 19944 10625
rect 14372 10480 14424 10532
rect 16856 10548 16908 10600
rect 17868 10548 17920 10600
rect 15384 10480 15436 10532
rect 16212 10480 16264 10532
rect 12164 10412 12216 10421
rect 12716 10412 12768 10464
rect 13636 10455 13688 10464
rect 13636 10421 13645 10455
rect 13645 10421 13679 10455
rect 13679 10421 13688 10455
rect 13636 10412 13688 10421
rect 16672 10412 16724 10464
rect 17500 10412 17552 10464
rect 18144 10412 18196 10464
rect 19800 10480 19852 10532
rect 8982 10310 9034 10362
rect 9046 10310 9098 10362
rect 9110 10310 9162 10362
rect 9174 10310 9226 10362
rect 16982 10310 17034 10362
rect 17046 10310 17098 10362
rect 17110 10310 17162 10362
rect 17174 10310 17226 10362
rect 1952 10208 2004 10260
rect 2228 10208 2280 10260
rect 4436 10251 4488 10260
rect 4436 10217 4445 10251
rect 4445 10217 4479 10251
rect 4479 10217 4488 10251
rect 4436 10208 4488 10217
rect 4804 10208 4856 10260
rect 7748 10208 7800 10260
rect 13544 10208 13596 10260
rect 15752 10251 15804 10260
rect 7104 10140 7156 10192
rect 7196 10140 7248 10192
rect 8760 10140 8812 10192
rect 9772 10140 9824 10192
rect 11704 10140 11756 10192
rect 12256 10183 12308 10192
rect 12256 10149 12265 10183
rect 12265 10149 12299 10183
rect 12299 10149 12308 10183
rect 13728 10183 13780 10192
rect 12256 10140 12308 10149
rect 13728 10149 13737 10183
rect 13737 10149 13771 10183
rect 13771 10149 13780 10183
rect 13728 10140 13780 10149
rect 15752 10217 15761 10251
rect 15761 10217 15795 10251
rect 15795 10217 15804 10251
rect 15752 10208 15804 10217
rect 19616 10208 19668 10260
rect 17316 10183 17368 10192
rect 17316 10149 17325 10183
rect 17325 10149 17359 10183
rect 17359 10149 17368 10183
rect 17316 10140 17368 10149
rect 18880 10140 18932 10192
rect 3148 10072 3200 10124
rect 3700 10072 3752 10124
rect 6920 10072 6972 10124
rect 8484 10072 8536 10124
rect 8852 10072 8904 10124
rect 10048 10115 10100 10124
rect 10048 10081 10057 10115
rect 10057 10081 10091 10115
rect 10091 10081 10100 10115
rect 10048 10072 10100 10081
rect 19800 10072 19852 10124
rect 20720 10072 20772 10124
rect 1492 10047 1544 10056
rect 1492 10013 1501 10047
rect 1501 10013 1535 10047
rect 1535 10013 1544 10047
rect 1492 10004 1544 10013
rect 12348 10004 12400 10056
rect 12532 10004 12584 10056
rect 13912 10004 13964 10056
rect 15384 10047 15436 10056
rect 15384 10013 15393 10047
rect 15393 10013 15427 10047
rect 15427 10013 15436 10047
rect 15384 10004 15436 10013
rect 16672 10004 16724 10056
rect 17592 10004 17644 10056
rect 18788 10004 18840 10056
rect 13176 9936 13228 9988
rect 17776 9979 17828 9988
rect 17776 9945 17785 9979
rect 17785 9945 17819 9979
rect 17819 9945 17828 9979
rect 17776 9936 17828 9945
rect 4068 9868 4120 9920
rect 5540 9868 5592 9920
rect 9312 9911 9364 9920
rect 9312 9877 9321 9911
rect 9321 9877 9355 9911
rect 9355 9877 9364 9911
rect 9312 9868 9364 9877
rect 9772 9868 9824 9920
rect 10968 9911 11020 9920
rect 10968 9877 10977 9911
rect 10977 9877 11011 9911
rect 11011 9877 11020 9911
rect 10968 9868 11020 9877
rect 16304 9911 16356 9920
rect 16304 9877 16313 9911
rect 16313 9877 16347 9911
rect 16347 9877 16356 9911
rect 16304 9868 16356 9877
rect 18144 9911 18196 9920
rect 18144 9877 18153 9911
rect 18153 9877 18187 9911
rect 18187 9877 18196 9911
rect 18144 9868 18196 9877
rect 20260 9868 20312 9920
rect 4982 9766 5034 9818
rect 5046 9766 5098 9818
rect 5110 9766 5162 9818
rect 5174 9766 5226 9818
rect 12982 9766 13034 9818
rect 13046 9766 13098 9818
rect 13110 9766 13162 9818
rect 13174 9766 13226 9818
rect 20982 9766 21034 9818
rect 21046 9766 21098 9818
rect 21110 9766 21162 9818
rect 21174 9766 21226 9818
rect 1952 9664 2004 9716
rect 3700 9707 3752 9716
rect 3700 9673 3709 9707
rect 3709 9673 3743 9707
rect 3743 9673 3752 9707
rect 3700 9664 3752 9673
rect 4436 9664 4488 9716
rect 5356 9664 5408 9716
rect 8024 9664 8076 9716
rect 10968 9664 11020 9716
rect 12256 9664 12308 9716
rect 13820 9664 13872 9716
rect 14372 9707 14424 9716
rect 14372 9673 14381 9707
rect 14381 9673 14415 9707
rect 14415 9673 14424 9707
rect 14372 9664 14424 9673
rect 15384 9664 15436 9716
rect 16304 9707 16356 9716
rect 16304 9673 16313 9707
rect 16313 9673 16347 9707
rect 16347 9673 16356 9707
rect 16304 9664 16356 9673
rect 17316 9664 17368 9716
rect 18880 9664 18932 9716
rect 19800 9664 19852 9716
rect 20720 9664 20772 9716
rect 7104 9639 7156 9648
rect 1492 9528 1544 9580
rect 7104 9605 7113 9639
rect 7113 9605 7147 9639
rect 7147 9605 7156 9639
rect 7104 9596 7156 9605
rect 12164 9596 12216 9648
rect 13544 9596 13596 9648
rect 14004 9596 14056 9648
rect 5448 9528 5500 9580
rect 7840 9528 7892 9580
rect 8760 9528 8812 9580
rect 12808 9571 12860 9580
rect 12808 9537 12817 9571
rect 12817 9537 12851 9571
rect 12851 9537 12860 9571
rect 12808 9528 12860 9537
rect 13452 9528 13504 9580
rect 13728 9528 13780 9580
rect 1676 9503 1728 9512
rect 1676 9469 1685 9503
rect 1685 9469 1719 9503
rect 1719 9469 1728 9503
rect 1676 9460 1728 9469
rect 2872 9460 2924 9512
rect 8392 9460 8444 9512
rect 9956 9460 10008 9512
rect 14464 9503 14516 9512
rect 14464 9469 14473 9503
rect 14473 9469 14507 9503
rect 14507 9469 14516 9503
rect 14464 9460 14516 9469
rect 16580 9528 16632 9580
rect 18144 9596 18196 9648
rect 21364 9639 21416 9648
rect 21364 9605 21373 9639
rect 21373 9605 21407 9639
rect 21407 9605 21416 9639
rect 21364 9596 21416 9605
rect 20168 9528 20220 9580
rect 20352 9528 20404 9580
rect 2964 9435 3016 9444
rect 2964 9401 2973 9435
rect 2973 9401 3007 9435
rect 3007 9401 3016 9435
rect 2964 9392 3016 9401
rect 4068 9324 4120 9376
rect 7748 9392 7800 9444
rect 8024 9435 8076 9444
rect 8024 9401 8033 9435
rect 8033 9401 8067 9435
rect 8067 9401 8076 9435
rect 8024 9392 8076 9401
rect 9404 9435 9456 9444
rect 9404 9401 9413 9435
rect 9413 9401 9447 9435
rect 9447 9401 9456 9435
rect 9404 9392 9456 9401
rect 9772 9435 9824 9444
rect 9772 9401 9781 9435
rect 9781 9401 9815 9435
rect 9815 9401 9824 9435
rect 9772 9392 9824 9401
rect 11152 9392 11204 9444
rect 12532 9435 12584 9444
rect 12532 9401 12541 9435
rect 12541 9401 12575 9435
rect 12575 9401 12584 9435
rect 12532 9392 12584 9401
rect 15200 9435 15252 9444
rect 8760 9324 8812 9376
rect 12256 9324 12308 9376
rect 15200 9401 15209 9435
rect 15209 9401 15243 9435
rect 15243 9401 15252 9435
rect 15200 9392 15252 9401
rect 15844 9324 15896 9376
rect 16304 9392 16356 9444
rect 17316 9392 17368 9444
rect 18604 9392 18656 9444
rect 18788 9435 18840 9444
rect 18788 9401 18797 9435
rect 18797 9401 18831 9435
rect 18831 9401 18840 9435
rect 18788 9392 18840 9401
rect 19800 9435 19852 9444
rect 19800 9401 19809 9435
rect 19809 9401 19843 9435
rect 19843 9401 19852 9435
rect 19800 9392 19852 9401
rect 20444 9392 20496 9444
rect 8982 9222 9034 9274
rect 9046 9222 9098 9274
rect 9110 9222 9162 9274
rect 9174 9222 9226 9274
rect 16982 9222 17034 9274
rect 17046 9222 17098 9274
rect 17110 9222 17162 9274
rect 17174 9222 17226 9274
rect 1860 9095 1912 9104
rect 20 8984 72 9036
rect 1860 9061 1869 9095
rect 1869 9061 1903 9095
rect 1903 9061 1912 9095
rect 1860 9052 1912 9061
rect 3792 9120 3844 9172
rect 4068 9120 4120 9172
rect 6920 9120 6972 9172
rect 7932 9120 7984 9172
rect 9956 9163 10008 9172
rect 9956 9129 9965 9163
rect 9965 9129 9999 9163
rect 9999 9129 10008 9163
rect 9956 9120 10008 9129
rect 11704 9120 11756 9172
rect 12532 9120 12584 9172
rect 3608 9052 3660 9104
rect 4712 9095 4764 9104
rect 4712 9061 4721 9095
rect 4721 9061 4755 9095
rect 4755 9061 4764 9095
rect 4712 9052 4764 9061
rect 7380 9052 7432 9104
rect 10048 9052 10100 9104
rect 12256 9095 12308 9104
rect 12256 9061 12265 9095
rect 12265 9061 12299 9095
rect 12299 9061 12308 9095
rect 12256 9052 12308 9061
rect 12808 9095 12860 9104
rect 12808 9061 12817 9095
rect 12817 9061 12851 9095
rect 12851 9061 12860 9095
rect 12808 9052 12860 9061
rect 13636 9120 13688 9172
rect 14464 9163 14516 9172
rect 14464 9129 14473 9163
rect 14473 9129 14507 9163
rect 14507 9129 14516 9163
rect 14464 9120 14516 9129
rect 16580 9120 16632 9172
rect 17592 9163 17644 9172
rect 17592 9129 17601 9163
rect 17601 9129 17635 9163
rect 17635 9129 17644 9163
rect 17592 9120 17644 9129
rect 18788 9120 18840 9172
rect 19984 9120 20036 9172
rect 20260 9163 20312 9172
rect 20260 9129 20269 9163
rect 20269 9129 20303 9163
rect 20303 9129 20312 9163
rect 20260 9120 20312 9129
rect 16764 9095 16816 9104
rect 16764 9061 16773 9095
rect 16773 9061 16807 9095
rect 16807 9061 16816 9095
rect 16764 9052 16816 9061
rect 20352 9052 20404 9104
rect 2688 9027 2740 9036
rect 2688 8993 2697 9027
rect 2697 8993 2731 9027
rect 2731 8993 2740 9027
rect 2688 8984 2740 8993
rect 2872 9027 2924 9036
rect 2872 8993 2881 9027
rect 2881 8993 2915 9027
rect 2915 8993 2924 9027
rect 2872 8984 2924 8993
rect 10232 9027 10284 9036
rect 2504 8916 2556 8968
rect 4804 8916 4856 8968
rect 4896 8959 4948 8968
rect 4896 8925 4905 8959
rect 4905 8925 4939 8959
rect 4939 8925 4948 8959
rect 7104 8959 7156 8968
rect 4896 8916 4948 8925
rect 7104 8925 7113 8959
rect 7113 8925 7147 8959
rect 7147 8925 7156 8959
rect 7104 8916 7156 8925
rect 1492 8848 1544 8900
rect 7472 8916 7524 8968
rect 10232 8993 10241 9027
rect 10241 8993 10275 9027
rect 10275 8993 10284 9027
rect 10232 8984 10284 8993
rect 13544 8984 13596 9036
rect 15476 8984 15528 9036
rect 17408 8984 17460 9036
rect 18144 9027 18196 9036
rect 18144 8993 18153 9027
rect 18153 8993 18187 9027
rect 18187 8993 18196 9027
rect 18144 8984 18196 8993
rect 18604 9027 18656 9036
rect 18604 8993 18613 9027
rect 18613 8993 18647 9027
rect 18647 8993 18656 9027
rect 18604 8984 18656 8993
rect 20168 8984 20220 9036
rect 11336 8916 11388 8968
rect 12348 8916 12400 8968
rect 16948 8916 17000 8968
rect 19064 8916 19116 8968
rect 20444 8916 20496 8968
rect 21272 8959 21324 8968
rect 15200 8848 15252 8900
rect 17776 8848 17828 8900
rect 21272 8925 21281 8959
rect 21281 8925 21315 8959
rect 21315 8925 21324 8959
rect 21272 8916 21324 8925
rect 22192 8848 22244 8900
rect 6000 8780 6052 8832
rect 10324 8780 10376 8832
rect 14464 8780 14516 8832
rect 4982 8678 5034 8730
rect 5046 8678 5098 8730
rect 5110 8678 5162 8730
rect 5174 8678 5226 8730
rect 12982 8678 13034 8730
rect 13046 8678 13098 8730
rect 13110 8678 13162 8730
rect 13174 8678 13226 8730
rect 20982 8678 21034 8730
rect 21046 8678 21098 8730
rect 21110 8678 21162 8730
rect 21174 8678 21226 8730
rect 2504 8619 2556 8628
rect 2504 8585 2513 8619
rect 2513 8585 2547 8619
rect 2547 8585 2556 8619
rect 2504 8576 2556 8585
rect 2688 8576 2740 8628
rect 7104 8576 7156 8628
rect 5356 8508 5408 8560
rect 6184 8508 6236 8560
rect 6552 8508 6604 8560
rect 8024 8483 8076 8492
rect 8024 8449 8033 8483
rect 8033 8449 8067 8483
rect 8067 8449 8076 8483
rect 8024 8440 8076 8449
rect 1952 8372 2004 8424
rect 10232 8576 10284 8628
rect 12256 8619 12308 8628
rect 12256 8585 12265 8619
rect 12265 8585 12299 8619
rect 12299 8585 12308 8619
rect 12256 8576 12308 8585
rect 16764 8576 16816 8628
rect 16948 8619 17000 8628
rect 16948 8585 16957 8619
rect 16957 8585 16991 8619
rect 16991 8585 17000 8619
rect 16948 8576 17000 8585
rect 18604 8576 18656 8628
rect 20352 8619 20404 8628
rect 20352 8585 20361 8619
rect 20361 8585 20395 8619
rect 20395 8585 20404 8619
rect 20352 8576 20404 8585
rect 22192 8619 22244 8628
rect 22192 8585 22201 8619
rect 22201 8585 22235 8619
rect 22235 8585 22244 8619
rect 22192 8576 22244 8585
rect 20904 8508 20956 8560
rect 10324 8415 10376 8424
rect 10324 8381 10333 8415
rect 10333 8381 10367 8415
rect 10367 8381 10376 8415
rect 10324 8372 10376 8381
rect 12624 8440 12676 8492
rect 13912 8440 13964 8492
rect 15200 8440 15252 8492
rect 15844 8440 15896 8492
rect 19064 8483 19116 8492
rect 19064 8449 19073 8483
rect 19073 8449 19107 8483
rect 19107 8449 19116 8483
rect 19064 8440 19116 8449
rect 20168 8440 20220 8492
rect 21272 8440 21324 8492
rect 14464 8415 14516 8424
rect 14464 8381 14473 8415
rect 14473 8381 14507 8415
rect 14507 8381 14516 8415
rect 14464 8372 14516 8381
rect 18052 8415 18104 8424
rect 18052 8381 18096 8415
rect 18096 8381 18104 8415
rect 18052 8372 18104 8381
rect 1676 8279 1728 8288
rect 1676 8245 1685 8279
rect 1685 8245 1719 8279
rect 1719 8245 1728 8279
rect 1676 8236 1728 8245
rect 3148 8279 3200 8288
rect 3148 8245 3157 8279
rect 3157 8245 3191 8279
rect 3191 8245 3200 8279
rect 3148 8236 3200 8245
rect 3976 8279 4028 8288
rect 3976 8245 3985 8279
rect 3985 8245 4019 8279
rect 4019 8245 4028 8279
rect 3976 8236 4028 8245
rect 7380 8304 7432 8356
rect 7564 8347 7616 8356
rect 7564 8313 7573 8347
rect 7573 8313 7607 8347
rect 7607 8313 7616 8347
rect 7564 8304 7616 8313
rect 10968 8347 11020 8356
rect 4712 8236 4764 8288
rect 4988 8236 5040 8288
rect 10968 8313 10977 8347
rect 10977 8313 11011 8347
rect 11011 8313 11020 8347
rect 10968 8304 11020 8313
rect 11336 8279 11388 8288
rect 11336 8245 11345 8279
rect 11345 8245 11379 8279
rect 11379 8245 11388 8279
rect 11336 8236 11388 8245
rect 12256 8236 12308 8288
rect 15844 8304 15896 8356
rect 17316 8304 17368 8356
rect 13544 8236 13596 8288
rect 13728 8236 13780 8288
rect 15476 8236 15528 8288
rect 17408 8236 17460 8288
rect 17868 8236 17920 8288
rect 19248 8236 19300 8288
rect 19892 8304 19944 8356
rect 20904 8347 20956 8356
rect 20904 8313 20913 8347
rect 20913 8313 20947 8347
rect 20947 8313 20956 8347
rect 20904 8304 20956 8313
rect 20628 8279 20680 8288
rect 20628 8245 20637 8279
rect 20637 8245 20671 8279
rect 20671 8245 20680 8279
rect 20628 8236 20680 8245
rect 8982 8134 9034 8186
rect 9046 8134 9098 8186
rect 9110 8134 9162 8186
rect 9174 8134 9226 8186
rect 16982 8134 17034 8186
rect 17046 8134 17098 8186
rect 17110 8134 17162 8186
rect 17174 8134 17226 8186
rect 3148 8032 3200 8084
rect 4436 8075 4488 8084
rect 4436 8041 4445 8075
rect 4445 8041 4479 8075
rect 4479 8041 4488 8075
rect 4436 8032 4488 8041
rect 4988 8075 5040 8084
rect 4988 8041 4997 8075
rect 4997 8041 5031 8075
rect 5031 8041 5040 8075
rect 4988 8032 5040 8041
rect 7380 8075 7432 8084
rect 7380 8041 7389 8075
rect 7389 8041 7423 8075
rect 7423 8041 7432 8075
rect 7380 8032 7432 8041
rect 7564 8032 7616 8084
rect 10968 8075 11020 8084
rect 10968 8041 10977 8075
rect 10977 8041 11011 8075
rect 11011 8041 11020 8075
rect 10968 8032 11020 8041
rect 1676 7964 1728 8016
rect 7012 7964 7064 8016
rect 10232 8007 10284 8016
rect 10232 7973 10241 8007
rect 10241 7973 10275 8007
rect 10275 7973 10284 8007
rect 10232 7964 10284 7973
rect 3148 7896 3200 7948
rect 5908 7896 5960 7948
rect 8024 7896 8076 7948
rect 8300 7896 8352 7948
rect 9864 7939 9916 7948
rect 1492 7871 1544 7880
rect 1492 7837 1501 7871
rect 1501 7837 1535 7871
rect 1535 7837 1544 7871
rect 1492 7828 1544 7837
rect 2136 7871 2188 7880
rect 2136 7837 2145 7871
rect 2145 7837 2179 7871
rect 2179 7837 2188 7871
rect 2136 7828 2188 7837
rect 4068 7871 4120 7880
rect 4068 7837 4077 7871
rect 4077 7837 4111 7871
rect 4111 7837 4120 7871
rect 4068 7828 4120 7837
rect 2780 7735 2832 7744
rect 2780 7701 2789 7735
rect 2789 7701 2823 7735
rect 2823 7701 2832 7735
rect 2780 7692 2832 7701
rect 3516 7735 3568 7744
rect 3516 7701 3525 7735
rect 3525 7701 3559 7735
rect 3559 7701 3568 7735
rect 3516 7692 3568 7701
rect 4804 7692 4856 7744
rect 5908 7692 5960 7744
rect 8852 7828 8904 7880
rect 9864 7905 9873 7939
rect 9873 7905 9907 7939
rect 9907 7905 9916 7939
rect 9864 7896 9916 7905
rect 12256 8032 12308 8084
rect 12348 8075 12400 8084
rect 12348 8041 12357 8075
rect 12357 8041 12391 8075
rect 12391 8041 12400 8075
rect 12348 8032 12400 8041
rect 13728 8032 13780 8084
rect 15016 8032 15068 8084
rect 18144 8075 18196 8084
rect 18144 8041 18153 8075
rect 18153 8041 18187 8075
rect 18187 8041 18196 8075
rect 18144 8032 18196 8041
rect 20628 8032 20680 8084
rect 11152 7964 11204 8016
rect 12532 7964 12584 8016
rect 13360 8007 13412 8016
rect 12808 7939 12860 7948
rect 12808 7905 12817 7939
rect 12817 7905 12851 7939
rect 12851 7905 12860 7939
rect 12808 7896 12860 7905
rect 13360 7973 13369 8007
rect 13369 7973 13403 8007
rect 13403 7973 13412 8007
rect 13360 7964 13412 7973
rect 16764 8007 16816 8016
rect 16764 7973 16773 8007
rect 16773 7973 16807 8007
rect 16807 7973 16816 8007
rect 16764 7964 16816 7973
rect 17316 8007 17368 8016
rect 17316 7973 17325 8007
rect 17325 7973 17359 8007
rect 17359 7973 17368 8007
rect 17316 7964 17368 7973
rect 19248 8007 19300 8016
rect 19248 7973 19257 8007
rect 19257 7973 19291 8007
rect 19291 7973 19300 8007
rect 19248 7964 19300 7973
rect 20168 8007 20220 8016
rect 20168 7973 20177 8007
rect 20177 7973 20211 8007
rect 20211 7973 20220 8007
rect 20168 7964 20220 7973
rect 20260 7964 20312 8016
rect 21456 7964 21508 8016
rect 14740 7896 14792 7948
rect 15292 7896 15344 7948
rect 10416 7828 10468 7880
rect 17040 7828 17092 7880
rect 17868 7828 17920 7880
rect 18972 7871 19024 7880
rect 18972 7837 18981 7871
rect 18981 7837 19015 7871
rect 19015 7837 19024 7871
rect 18972 7828 19024 7837
rect 20812 7828 20864 7880
rect 21272 7871 21324 7880
rect 21272 7837 21281 7871
rect 21281 7837 21315 7871
rect 21315 7837 21324 7871
rect 21272 7828 21324 7837
rect 15660 7760 15712 7812
rect 9496 7735 9548 7744
rect 9496 7701 9505 7735
rect 9505 7701 9539 7735
rect 9539 7701 9548 7735
rect 9496 7692 9548 7701
rect 10140 7692 10192 7744
rect 12624 7735 12676 7744
rect 12624 7701 12633 7735
rect 12633 7701 12667 7735
rect 12667 7701 12676 7735
rect 12624 7692 12676 7701
rect 13820 7735 13872 7744
rect 13820 7701 13829 7735
rect 13829 7701 13863 7735
rect 13863 7701 13872 7735
rect 13820 7692 13872 7701
rect 14188 7692 14240 7744
rect 15844 7735 15896 7744
rect 15844 7701 15853 7735
rect 15853 7701 15887 7735
rect 15887 7701 15896 7735
rect 15844 7692 15896 7701
rect 4982 7590 5034 7642
rect 5046 7590 5098 7642
rect 5110 7590 5162 7642
rect 5174 7590 5226 7642
rect 12982 7590 13034 7642
rect 13046 7590 13098 7642
rect 13110 7590 13162 7642
rect 13174 7590 13226 7642
rect 20982 7590 21034 7642
rect 21046 7590 21098 7642
rect 21110 7590 21162 7642
rect 21174 7590 21226 7642
rect 1676 7531 1728 7540
rect 1676 7497 1685 7531
rect 1685 7497 1719 7531
rect 1719 7497 1728 7531
rect 1676 7488 1728 7497
rect 3148 7488 3200 7540
rect 4436 7531 4488 7540
rect 4436 7497 4445 7531
rect 4445 7497 4479 7531
rect 4479 7497 4488 7531
rect 4436 7488 4488 7497
rect 7012 7488 7064 7540
rect 8852 7531 8904 7540
rect 8852 7497 8861 7531
rect 8861 7497 8895 7531
rect 8895 7497 8904 7531
rect 8852 7488 8904 7497
rect 9496 7488 9548 7540
rect 12624 7488 12676 7540
rect 12808 7488 12860 7540
rect 14740 7531 14792 7540
rect 14740 7497 14749 7531
rect 14749 7497 14783 7531
rect 14783 7497 14792 7531
rect 14740 7488 14792 7497
rect 16764 7488 16816 7540
rect 17040 7531 17092 7540
rect 17040 7497 17049 7531
rect 17049 7497 17083 7531
rect 17083 7497 17092 7531
rect 17040 7488 17092 7497
rect 20260 7531 20312 7540
rect 20260 7497 20269 7531
rect 20269 7497 20303 7531
rect 20303 7497 20312 7531
rect 20260 7488 20312 7497
rect 20812 7488 20864 7540
rect 2136 7420 2188 7472
rect 10140 7420 10192 7472
rect 13452 7420 13504 7472
rect 14924 7420 14976 7472
rect 2780 7352 2832 7404
rect 2872 7352 2924 7404
rect 3424 7352 3476 7404
rect 5908 7395 5960 7404
rect 3516 7327 3568 7336
rect 3516 7293 3525 7327
rect 3525 7293 3559 7327
rect 3559 7293 3568 7327
rect 3516 7284 3568 7293
rect 4068 7327 4120 7336
rect 4068 7293 4077 7327
rect 4077 7293 4111 7327
rect 4111 7293 4120 7327
rect 4068 7284 4120 7293
rect 1952 7259 2004 7268
rect 1952 7225 1961 7259
rect 1961 7225 1995 7259
rect 1995 7225 2004 7259
rect 1952 7216 2004 7225
rect 5908 7361 5917 7395
rect 5917 7361 5951 7395
rect 5951 7361 5960 7395
rect 5908 7352 5960 7361
rect 10232 7352 10284 7404
rect 5448 7327 5500 7336
rect 5448 7293 5457 7327
rect 5457 7293 5491 7327
rect 5491 7293 5500 7327
rect 5448 7284 5500 7293
rect 7472 7284 7524 7336
rect 8300 7327 8352 7336
rect 8300 7293 8309 7327
rect 8309 7293 8343 7327
rect 8343 7293 8352 7327
rect 8300 7284 8352 7293
rect 13360 7284 13412 7336
rect 3148 7148 3200 7200
rect 4436 7148 4488 7200
rect 7196 7259 7248 7268
rect 7196 7225 7205 7259
rect 7205 7225 7239 7259
rect 7239 7225 7248 7259
rect 7196 7216 7248 7225
rect 9864 7216 9916 7268
rect 13452 7216 13504 7268
rect 10232 7148 10284 7200
rect 11152 7191 11204 7200
rect 11152 7157 11161 7191
rect 11161 7157 11195 7191
rect 11195 7157 11204 7191
rect 11152 7148 11204 7157
rect 11244 7148 11296 7200
rect 12624 7148 12676 7200
rect 14188 7352 14240 7404
rect 15660 7395 15712 7404
rect 15660 7361 15669 7395
rect 15669 7361 15703 7395
rect 15703 7361 15712 7395
rect 15660 7352 15712 7361
rect 18972 7352 19024 7404
rect 21456 7488 21508 7540
rect 17960 7284 18012 7336
rect 20168 7284 20220 7336
rect 13820 7216 13872 7268
rect 15752 7259 15804 7268
rect 15752 7225 15761 7259
rect 15761 7225 15795 7259
rect 15795 7225 15804 7259
rect 15752 7216 15804 7225
rect 15292 7191 15344 7200
rect 15292 7157 15301 7191
rect 15301 7157 15335 7191
rect 15335 7157 15344 7191
rect 15292 7148 15344 7157
rect 16120 7148 16172 7200
rect 19064 7148 19116 7200
rect 8982 7046 9034 7098
rect 9046 7046 9098 7098
rect 9110 7046 9162 7098
rect 9174 7046 9226 7098
rect 16982 7046 17034 7098
rect 17046 7046 17098 7098
rect 17110 7046 17162 7098
rect 17174 7046 17226 7098
rect 1492 6944 1544 6996
rect 3424 6987 3476 6996
rect 3424 6953 3433 6987
rect 3433 6953 3467 6987
rect 3467 6953 3476 6987
rect 3424 6944 3476 6953
rect 4068 6944 4120 6996
rect 5724 6944 5776 6996
rect 11152 6944 11204 6996
rect 2044 6919 2096 6928
rect 2044 6885 2047 6919
rect 2047 6885 2081 6919
rect 2081 6885 2096 6919
rect 2044 6876 2096 6885
rect 3148 6876 3200 6928
rect 4804 6876 4856 6928
rect 5356 6876 5408 6928
rect 4620 6808 4672 6860
rect 5540 6851 5592 6860
rect 5540 6817 5549 6851
rect 5549 6817 5583 6851
rect 5583 6817 5592 6851
rect 5540 6808 5592 6817
rect 5908 6808 5960 6860
rect 7656 6808 7708 6860
rect 12716 6876 12768 6928
rect 13820 6987 13872 6996
rect 13820 6953 13829 6987
rect 13829 6953 13863 6987
rect 13863 6953 13872 6987
rect 14188 6987 14240 6996
rect 13820 6944 13872 6953
rect 14188 6953 14197 6987
rect 14197 6953 14231 6987
rect 14231 6953 14240 6987
rect 14188 6944 14240 6953
rect 19156 6944 19208 6996
rect 19616 6987 19668 6996
rect 19616 6953 19625 6987
rect 19625 6953 19659 6987
rect 19659 6953 19668 6987
rect 19616 6944 19668 6953
rect 15752 6876 15804 6928
rect 16212 6919 16264 6928
rect 16212 6885 16221 6919
rect 16221 6885 16255 6919
rect 16255 6885 16264 6919
rect 16212 6876 16264 6885
rect 18972 6876 19024 6928
rect 11244 6851 11296 6860
rect 11244 6817 11253 6851
rect 11253 6817 11287 6851
rect 11287 6817 11296 6851
rect 11244 6808 11296 6817
rect 17960 6851 18012 6860
rect 17960 6817 17969 6851
rect 17969 6817 18003 6851
rect 18003 6817 18012 6851
rect 17960 6808 18012 6817
rect 18604 6808 18656 6860
rect 2320 6740 2372 6792
rect 6000 6783 6052 6792
rect 6000 6749 6009 6783
rect 6009 6749 6043 6783
rect 6043 6749 6052 6783
rect 6000 6740 6052 6749
rect 7932 6783 7984 6792
rect 1952 6672 2004 6724
rect 6092 6672 6144 6724
rect 7932 6749 7941 6783
rect 7941 6749 7975 6783
rect 7975 6749 7984 6783
rect 7932 6740 7984 6749
rect 9496 6740 9548 6792
rect 10232 6783 10284 6792
rect 10232 6749 10241 6783
rect 10241 6749 10275 6783
rect 10275 6749 10284 6783
rect 10232 6740 10284 6749
rect 11704 6740 11756 6792
rect 12348 6740 12400 6792
rect 16120 6783 16172 6792
rect 16120 6749 16129 6783
rect 16129 6749 16163 6783
rect 16163 6749 16172 6783
rect 16120 6740 16172 6749
rect 16304 6740 16356 6792
rect 17592 6740 17644 6792
rect 7196 6672 7248 6724
rect 7748 6672 7800 6724
rect 10140 6715 10192 6724
rect 10140 6681 10149 6715
rect 10149 6681 10183 6715
rect 10183 6681 10192 6715
rect 10140 6672 10192 6681
rect 5448 6604 5500 6656
rect 5724 6604 5776 6656
rect 7012 6604 7064 6656
rect 7840 6647 7892 6656
rect 7840 6613 7849 6647
rect 7849 6613 7883 6647
rect 7883 6613 7892 6647
rect 7840 6604 7892 6613
rect 9128 6647 9180 6656
rect 9128 6613 9137 6647
rect 9137 6613 9171 6647
rect 9171 6613 9180 6647
rect 9128 6604 9180 6613
rect 10968 6647 11020 6656
rect 10968 6613 10977 6647
rect 10977 6613 11011 6647
rect 11011 6613 11020 6647
rect 10968 6604 11020 6613
rect 12808 6604 12860 6656
rect 18972 6647 19024 6656
rect 18972 6613 18981 6647
rect 18981 6613 19015 6647
rect 19015 6613 19024 6647
rect 18972 6604 19024 6613
rect 20168 6604 20220 6656
rect 4982 6502 5034 6554
rect 5046 6502 5098 6554
rect 5110 6502 5162 6554
rect 5174 6502 5226 6554
rect 12982 6502 13034 6554
rect 13046 6502 13098 6554
rect 13110 6502 13162 6554
rect 13174 6502 13226 6554
rect 20982 6502 21034 6554
rect 21046 6502 21098 6554
rect 21110 6502 21162 6554
rect 21174 6502 21226 6554
rect 2044 6400 2096 6452
rect 4620 6400 4672 6452
rect 8024 6443 8076 6452
rect 8024 6409 8033 6443
rect 8033 6409 8067 6443
rect 8067 6409 8076 6443
rect 8024 6400 8076 6409
rect 9680 6400 9732 6452
rect 11704 6443 11756 6452
rect 11704 6409 11713 6443
rect 11713 6409 11747 6443
rect 11747 6409 11756 6443
rect 11704 6400 11756 6409
rect 16212 6443 16264 6452
rect 16212 6409 16221 6443
rect 16221 6409 16255 6443
rect 16255 6409 16264 6443
rect 16212 6400 16264 6409
rect 18604 6400 18656 6452
rect 7840 6375 7892 6384
rect 7840 6341 7849 6375
rect 7849 6341 7883 6375
rect 7883 6341 7892 6375
rect 7840 6332 7892 6341
rect 8300 6332 8352 6384
rect 9404 6375 9456 6384
rect 9404 6341 9413 6375
rect 9413 6341 9447 6375
rect 9447 6341 9456 6375
rect 9404 6332 9456 6341
rect 7932 6307 7984 6316
rect 2228 6196 2280 6248
rect 3700 6239 3752 6248
rect 3700 6205 3709 6239
rect 3709 6205 3743 6239
rect 3743 6205 3752 6239
rect 3700 6196 3752 6205
rect 7932 6273 7941 6307
rect 7941 6273 7975 6307
rect 7975 6273 7984 6307
rect 7932 6264 7984 6273
rect 9956 6264 10008 6316
rect 10232 6264 10284 6316
rect 112 6060 164 6112
rect 2320 6103 2372 6112
rect 2320 6069 2329 6103
rect 2329 6069 2363 6103
rect 2363 6069 2372 6103
rect 2320 6060 2372 6069
rect 5540 6196 5592 6248
rect 7656 6196 7708 6248
rect 9772 6196 9824 6248
rect 15936 6332 15988 6384
rect 17960 6332 18012 6384
rect 13452 6264 13504 6316
rect 13912 6264 13964 6316
rect 16304 6264 16356 6316
rect 16488 6264 16540 6316
rect 20168 6307 20220 6316
rect 12532 6196 12584 6248
rect 13544 6196 13596 6248
rect 4804 6060 4856 6112
rect 5540 6103 5592 6112
rect 5540 6069 5549 6103
rect 5549 6069 5583 6103
rect 5583 6069 5592 6103
rect 5540 6060 5592 6069
rect 5908 6103 5960 6112
rect 5908 6069 5917 6103
rect 5917 6069 5951 6103
rect 5951 6069 5960 6103
rect 5908 6060 5960 6069
rect 6092 6060 6144 6112
rect 7472 6060 7524 6112
rect 8024 6128 8076 6180
rect 9128 6171 9180 6180
rect 9128 6137 9137 6171
rect 9137 6137 9171 6171
rect 9171 6137 9180 6171
rect 9128 6128 9180 6137
rect 13268 6128 13320 6180
rect 13820 6171 13872 6180
rect 13820 6137 13829 6171
rect 13829 6137 13863 6171
rect 13863 6137 13872 6171
rect 13820 6128 13872 6137
rect 8300 6060 8352 6112
rect 10968 6103 11020 6112
rect 10968 6069 10977 6103
rect 10977 6069 11011 6103
rect 11011 6069 11020 6103
rect 10968 6060 11020 6069
rect 12348 6060 12400 6112
rect 13544 6103 13596 6112
rect 13544 6069 13553 6103
rect 13553 6069 13587 6103
rect 13587 6069 13596 6103
rect 15844 6128 15896 6180
rect 16856 6196 16908 6248
rect 17868 6196 17920 6248
rect 19616 6239 19668 6248
rect 19616 6205 19625 6239
rect 19625 6205 19659 6239
rect 19659 6205 19668 6239
rect 19616 6196 19668 6205
rect 20168 6273 20177 6307
rect 20177 6273 20211 6307
rect 20211 6273 20220 6307
rect 20168 6264 20220 6273
rect 13544 6060 13596 6069
rect 8982 5958 9034 6010
rect 9046 5958 9098 6010
rect 9110 5958 9162 6010
rect 9174 5958 9226 6010
rect 16982 5958 17034 6010
rect 17046 5958 17098 6010
rect 17110 5958 17162 6010
rect 17174 5958 17226 6010
rect 3240 5856 3292 5908
rect 1952 5831 2004 5840
rect 1952 5797 1961 5831
rect 1961 5797 1995 5831
rect 1995 5797 2004 5831
rect 1952 5788 2004 5797
rect 3700 5720 3752 5772
rect 4160 5720 4212 5772
rect 4988 5856 5040 5908
rect 8024 5856 8076 5908
rect 9496 5856 9548 5908
rect 13452 5856 13504 5908
rect 16120 5856 16172 5908
rect 17868 5856 17920 5908
rect 10416 5831 10468 5840
rect 10416 5797 10425 5831
rect 10425 5797 10459 5831
rect 10459 5797 10468 5831
rect 10416 5788 10468 5797
rect 12348 5831 12400 5840
rect 12348 5797 12357 5831
rect 12357 5797 12391 5831
rect 12391 5797 12400 5831
rect 12348 5788 12400 5797
rect 13360 5831 13412 5840
rect 13360 5797 13369 5831
rect 13369 5797 13403 5831
rect 13403 5797 13412 5831
rect 13360 5788 13412 5797
rect 13912 5831 13964 5840
rect 13912 5797 13921 5831
rect 13921 5797 13955 5831
rect 13955 5797 13964 5831
rect 13912 5788 13964 5797
rect 17684 5831 17736 5840
rect 17684 5797 17693 5831
rect 17693 5797 17727 5831
rect 17727 5797 17736 5831
rect 17684 5788 17736 5797
rect 6000 5763 6052 5772
rect 6000 5729 6009 5763
rect 6009 5729 6043 5763
rect 6043 5729 6052 5763
rect 6000 5720 6052 5729
rect 6092 5763 6144 5772
rect 6092 5729 6101 5763
rect 6101 5729 6135 5763
rect 6135 5729 6144 5763
rect 6092 5720 6144 5729
rect 6736 5763 6788 5772
rect 2136 5652 2188 5704
rect 2228 5695 2280 5704
rect 2228 5661 2237 5695
rect 2237 5661 2271 5695
rect 2271 5661 2280 5695
rect 2228 5652 2280 5661
rect 4804 5695 4856 5704
rect 4804 5661 4813 5695
rect 4813 5661 4847 5695
rect 4847 5661 4856 5695
rect 4804 5652 4856 5661
rect 6736 5729 6745 5763
rect 6745 5729 6779 5763
rect 6779 5729 6788 5763
rect 6736 5720 6788 5729
rect 7564 5763 7616 5772
rect 7564 5729 7573 5763
rect 7573 5729 7607 5763
rect 7607 5729 7616 5763
rect 7564 5720 7616 5729
rect 8116 5720 8168 5772
rect 9772 5720 9824 5772
rect 9956 5763 10008 5772
rect 9956 5729 9965 5763
rect 9965 5729 9999 5763
rect 9999 5729 10008 5763
rect 9956 5720 10008 5729
rect 5632 5516 5684 5568
rect 10324 5652 10376 5704
rect 11980 5720 12032 5772
rect 15936 5763 15988 5772
rect 15936 5729 15945 5763
rect 15945 5729 15979 5763
rect 15979 5729 15988 5763
rect 15936 5720 15988 5729
rect 16488 5763 16540 5772
rect 16488 5729 16497 5763
rect 16497 5729 16531 5763
rect 16531 5729 16540 5763
rect 16488 5720 16540 5729
rect 12808 5652 12860 5704
rect 16672 5695 16724 5704
rect 16672 5661 16681 5695
rect 16681 5661 16715 5695
rect 16715 5661 16724 5695
rect 16672 5652 16724 5661
rect 17592 5695 17644 5704
rect 17592 5661 17601 5695
rect 17601 5661 17635 5695
rect 17635 5661 17644 5695
rect 17592 5652 17644 5661
rect 17868 5695 17920 5704
rect 17868 5661 17877 5695
rect 17877 5661 17911 5695
rect 17911 5661 17920 5695
rect 17868 5652 17920 5661
rect 19340 5695 19392 5704
rect 19340 5661 19349 5695
rect 19349 5661 19383 5695
rect 19383 5661 19392 5695
rect 19340 5652 19392 5661
rect 10968 5584 11020 5636
rect 7012 5559 7064 5568
rect 7012 5525 7021 5559
rect 7021 5525 7055 5559
rect 7055 5525 7064 5559
rect 7012 5516 7064 5525
rect 7472 5559 7524 5568
rect 7472 5525 7481 5559
rect 7481 5525 7515 5559
rect 7515 5525 7524 5559
rect 7472 5516 7524 5525
rect 8300 5516 8352 5568
rect 9312 5516 9364 5568
rect 12624 5559 12676 5568
rect 12624 5525 12633 5559
rect 12633 5525 12667 5559
rect 12667 5525 12676 5559
rect 12624 5516 12676 5525
rect 16948 5559 17000 5568
rect 16948 5525 16957 5559
rect 16957 5525 16991 5559
rect 16991 5525 17000 5559
rect 16948 5516 17000 5525
rect 4982 5414 5034 5466
rect 5046 5414 5098 5466
rect 5110 5414 5162 5466
rect 5174 5414 5226 5466
rect 12982 5414 13034 5466
rect 13046 5414 13098 5466
rect 13110 5414 13162 5466
rect 13174 5414 13226 5466
rect 20982 5414 21034 5466
rect 21046 5414 21098 5466
rect 21110 5414 21162 5466
rect 21174 5414 21226 5466
rect 1952 5312 2004 5364
rect 2412 5312 2464 5364
rect 3240 5355 3292 5364
rect 3240 5321 3249 5355
rect 3249 5321 3283 5355
rect 3283 5321 3292 5355
rect 3240 5312 3292 5321
rect 4160 5355 4212 5364
rect 4160 5321 4169 5355
rect 4169 5321 4203 5355
rect 4203 5321 4212 5355
rect 4160 5312 4212 5321
rect 4804 5312 4856 5364
rect 2044 5244 2096 5296
rect 6092 5312 6144 5364
rect 7012 5312 7064 5364
rect 9312 5355 9364 5364
rect 5264 5287 5316 5296
rect 5264 5253 5273 5287
rect 5273 5253 5307 5287
rect 5307 5253 5316 5287
rect 5264 5244 5316 5253
rect 2044 5040 2096 5092
rect 2872 5040 2924 5092
rect 4804 5108 4856 5160
rect 6000 5176 6052 5228
rect 9312 5321 9321 5355
rect 9321 5321 9355 5355
rect 9355 5321 9364 5355
rect 10968 5355 11020 5364
rect 9312 5312 9364 5321
rect 10968 5321 10977 5355
rect 10977 5321 11011 5355
rect 11011 5321 11020 5355
rect 10968 5312 11020 5321
rect 11704 5312 11756 5364
rect 13360 5312 13412 5364
rect 14464 5312 14516 5364
rect 15936 5312 15988 5364
rect 16488 5312 16540 5364
rect 19340 5312 19392 5364
rect 9956 5244 10008 5296
rect 14924 5287 14976 5296
rect 14924 5253 14933 5287
rect 14933 5253 14967 5287
rect 14967 5253 14976 5287
rect 14924 5244 14976 5253
rect 10232 5219 10284 5228
rect 5632 5108 5684 5160
rect 9496 5151 9548 5160
rect 4620 4972 4672 5024
rect 5908 5040 5960 5092
rect 5816 4972 5868 5024
rect 9496 5117 9505 5151
rect 9505 5117 9539 5151
rect 9539 5117 9548 5151
rect 9496 5108 9548 5117
rect 10232 5185 10241 5219
rect 10241 5185 10275 5219
rect 10275 5185 10284 5219
rect 10232 5176 10284 5185
rect 12624 5176 12676 5228
rect 13268 5176 13320 5228
rect 14372 5219 14424 5228
rect 14372 5185 14381 5219
rect 14381 5185 14415 5219
rect 14415 5185 14424 5219
rect 14372 5176 14424 5185
rect 16948 5244 17000 5296
rect 17684 5244 17736 5296
rect 16672 5176 16724 5228
rect 18052 5219 18104 5228
rect 18052 5185 18061 5219
rect 18061 5185 18095 5219
rect 18095 5185 18104 5219
rect 18052 5176 18104 5185
rect 7564 5040 7616 5092
rect 7196 4972 7248 5024
rect 8116 4972 8168 5024
rect 9772 4972 9824 5024
rect 13452 5108 13504 5160
rect 17868 5108 17920 5160
rect 11704 5040 11756 5092
rect 13544 5040 13596 5092
rect 14464 5083 14516 5092
rect 14464 5049 14473 5083
rect 14473 5049 14507 5083
rect 14507 5049 14516 5083
rect 14464 5040 14516 5049
rect 16396 5083 16448 5092
rect 16396 5049 16405 5083
rect 16405 5049 16439 5083
rect 16439 5049 16448 5083
rect 16396 5040 16448 5049
rect 11060 4972 11112 5024
rect 15844 4972 15896 5024
rect 18972 4972 19024 5024
rect 19984 5083 20036 5092
rect 19984 5049 19993 5083
rect 19993 5049 20027 5083
rect 20027 5049 20036 5083
rect 19984 5040 20036 5049
rect 19432 4972 19484 5024
rect 8982 4870 9034 4922
rect 9046 4870 9098 4922
rect 9110 4870 9162 4922
rect 9174 4870 9226 4922
rect 16982 4870 17034 4922
rect 17046 4870 17098 4922
rect 17110 4870 17162 4922
rect 17174 4870 17226 4922
rect 2412 4811 2464 4820
rect 2412 4777 2421 4811
rect 2421 4777 2455 4811
rect 2455 4777 2464 4811
rect 2412 4768 2464 4777
rect 5264 4811 5316 4820
rect 5264 4777 5273 4811
rect 5273 4777 5307 4811
rect 5307 4777 5316 4811
rect 5264 4768 5316 4777
rect 1584 4743 1636 4752
rect 1584 4709 1593 4743
rect 1593 4709 1627 4743
rect 1627 4709 1636 4743
rect 1584 4700 1636 4709
rect 2228 4700 2280 4752
rect 8116 4768 8168 4820
rect 9496 4811 9548 4820
rect 9496 4777 9505 4811
rect 9505 4777 9539 4811
rect 9539 4777 9548 4811
rect 9496 4768 9548 4777
rect 3976 4632 4028 4684
rect 6000 4700 6052 4752
rect 12808 4768 12860 4820
rect 14372 4811 14424 4820
rect 14372 4777 14381 4811
rect 14381 4777 14415 4811
rect 14415 4777 14424 4811
rect 14372 4768 14424 4777
rect 15844 4811 15896 4820
rect 15844 4777 15853 4811
rect 15853 4777 15887 4811
rect 15887 4777 15896 4811
rect 15844 4768 15896 4777
rect 16396 4811 16448 4820
rect 16396 4777 16405 4811
rect 16405 4777 16439 4811
rect 16439 4777 16448 4811
rect 16396 4768 16448 4777
rect 17592 4811 17644 4820
rect 17592 4777 17601 4811
rect 17601 4777 17635 4811
rect 17635 4777 17644 4811
rect 17592 4768 17644 4777
rect 18052 4811 18104 4820
rect 18052 4777 18061 4811
rect 18061 4777 18095 4811
rect 18095 4777 18104 4811
rect 18052 4768 18104 4777
rect 18972 4811 19024 4820
rect 18972 4777 18981 4811
rect 18981 4777 19015 4811
rect 19015 4777 19024 4811
rect 18972 4768 19024 4777
rect 19984 4768 20036 4820
rect 1952 4564 2004 4616
rect 3884 4564 3936 4616
rect 5356 4632 5408 4684
rect 5540 4675 5592 4684
rect 5540 4641 5549 4675
rect 5549 4641 5583 4675
rect 5583 4641 5592 4675
rect 5540 4632 5592 4641
rect 5632 4632 5684 4684
rect 12624 4743 12676 4752
rect 12624 4709 12633 4743
rect 12633 4709 12667 4743
rect 12667 4709 12676 4743
rect 12624 4700 12676 4709
rect 12716 4700 12768 4752
rect 7104 4675 7156 4684
rect 7104 4641 7113 4675
rect 7113 4641 7147 4675
rect 7147 4641 7156 4675
rect 7104 4632 7156 4641
rect 7196 4632 7248 4684
rect 8024 4632 8076 4684
rect 9772 4675 9824 4684
rect 9772 4641 9781 4675
rect 9781 4641 9815 4675
rect 9815 4641 9824 4675
rect 9772 4632 9824 4641
rect 11888 4675 11940 4684
rect 11888 4641 11897 4675
rect 11897 4641 11931 4675
rect 11931 4641 11940 4675
rect 11888 4632 11940 4641
rect 13452 4675 13504 4684
rect 5724 4564 5776 4616
rect 8668 4564 8720 4616
rect 11980 4564 12032 4616
rect 13452 4641 13461 4675
rect 13461 4641 13495 4675
rect 13495 4641 13504 4675
rect 13452 4632 13504 4641
rect 13820 4632 13872 4684
rect 13912 4607 13964 4616
rect 13912 4573 13921 4607
rect 13921 4573 13955 4607
rect 13955 4573 13964 4607
rect 13912 4564 13964 4573
rect 15476 4607 15528 4616
rect 15476 4573 15485 4607
rect 15485 4573 15519 4607
rect 15519 4573 15528 4607
rect 15476 4564 15528 4573
rect 18604 4607 18656 4616
rect 18604 4573 18613 4607
rect 18613 4573 18647 4607
rect 18647 4573 18656 4607
rect 18604 4564 18656 4573
rect 5264 4496 5316 4548
rect 5448 4496 5500 4548
rect 6644 4496 6696 4548
rect 7840 4428 7892 4480
rect 10232 4428 10284 4480
rect 4982 4326 5034 4378
rect 5046 4326 5098 4378
rect 5110 4326 5162 4378
rect 5174 4326 5226 4378
rect 12982 4326 13034 4378
rect 13046 4326 13098 4378
rect 13110 4326 13162 4378
rect 13174 4326 13226 4378
rect 20982 4326 21034 4378
rect 21046 4326 21098 4378
rect 21110 4326 21162 4378
rect 21174 4326 21226 4378
rect 2412 4224 2464 4276
rect 3884 4267 3936 4276
rect 3884 4233 3893 4267
rect 3893 4233 3927 4267
rect 3927 4233 3936 4267
rect 3884 4224 3936 4233
rect 6644 4267 6696 4276
rect 6644 4233 6653 4267
rect 6653 4233 6687 4267
rect 6687 4233 6696 4267
rect 6644 4224 6696 4233
rect 7196 4267 7248 4276
rect 7196 4233 7205 4267
rect 7205 4233 7239 4267
rect 7239 4233 7248 4267
rect 7196 4224 7248 4233
rect 7840 4267 7892 4276
rect 7840 4233 7849 4267
rect 7849 4233 7883 4267
rect 7883 4233 7892 4267
rect 7840 4224 7892 4233
rect 11980 4267 12032 4276
rect 11980 4233 11989 4267
rect 11989 4233 12023 4267
rect 12023 4233 12032 4267
rect 11980 4224 12032 4233
rect 13452 4267 13504 4276
rect 13452 4233 13461 4267
rect 13461 4233 13495 4267
rect 13495 4233 13504 4267
rect 13452 4224 13504 4233
rect 13820 4267 13872 4276
rect 13820 4233 13829 4267
rect 13829 4233 13863 4267
rect 13863 4233 13872 4267
rect 13820 4224 13872 4233
rect 15844 4224 15896 4276
rect 16488 4224 16540 4276
rect 18512 4224 18564 4276
rect 18972 4224 19024 4276
rect 5172 4156 5224 4208
rect 3056 4088 3108 4140
rect 2412 4020 2464 4072
rect 4252 4020 4304 4072
rect 4712 4063 4764 4072
rect 4712 4029 4721 4063
rect 4721 4029 4755 4063
rect 4755 4029 4764 4063
rect 4712 4020 4764 4029
rect 11888 4156 11940 4208
rect 9772 4131 9824 4140
rect 9772 4097 9781 4131
rect 9781 4097 9815 4131
rect 9815 4097 9824 4131
rect 9772 4088 9824 4097
rect 14004 4088 14056 4140
rect 7932 4063 7984 4072
rect 1584 3995 1636 4004
rect 1584 3961 1593 3995
rect 1593 3961 1627 3995
rect 1627 3961 1636 3995
rect 1584 3952 1636 3961
rect 4620 3952 4672 4004
rect 7932 4029 7941 4063
rect 7941 4029 7975 4063
rect 7975 4029 7984 4063
rect 7932 4020 7984 4029
rect 8024 4020 8076 4072
rect 8392 4063 8444 4072
rect 8392 4029 8401 4063
rect 8401 4029 8435 4063
rect 8435 4029 8444 4063
rect 8392 4020 8444 4029
rect 8760 4063 8812 4072
rect 8760 4029 8769 4063
rect 8769 4029 8803 4063
rect 8803 4029 8812 4063
rect 8760 4020 8812 4029
rect 10692 4020 10744 4072
rect 12716 4063 12768 4072
rect 12716 4029 12725 4063
rect 12725 4029 12759 4063
rect 12759 4029 12768 4063
rect 12716 4020 12768 4029
rect 15016 4063 15068 4072
rect 15016 4029 15025 4063
rect 15025 4029 15059 4063
rect 15059 4029 15068 4063
rect 15016 4020 15068 4029
rect 16580 4020 16632 4072
rect 18144 4020 18196 4072
rect 19156 4088 19208 4140
rect 18512 4063 18564 4072
rect 18512 4029 18521 4063
rect 18521 4029 18555 4063
rect 18555 4029 18564 4063
rect 18512 4020 18564 4029
rect 19432 4020 19484 4072
rect 5448 3952 5500 4004
rect 12440 3995 12492 4004
rect 12440 3961 12449 3995
rect 12449 3961 12483 3995
rect 12483 3961 12492 3995
rect 12440 3952 12492 3961
rect 15476 3952 15528 4004
rect 18604 3952 18656 4004
rect 23112 3952 23164 4004
rect 204 3884 256 3936
rect 3976 3884 4028 3936
rect 4160 3927 4212 3936
rect 4160 3893 4169 3927
rect 4169 3893 4203 3927
rect 4203 3893 4212 3927
rect 4160 3884 4212 3893
rect 4712 3884 4764 3936
rect 5540 3884 5592 3936
rect 8852 3927 8904 3936
rect 8852 3893 8861 3927
rect 8861 3893 8895 3927
rect 8895 3893 8904 3927
rect 8852 3884 8904 3893
rect 10508 3927 10560 3936
rect 10508 3893 10517 3927
rect 10517 3893 10551 3927
rect 10551 3893 10560 3927
rect 10508 3884 10560 3893
rect 8982 3782 9034 3834
rect 9046 3782 9098 3834
rect 9110 3782 9162 3834
rect 9174 3782 9226 3834
rect 16982 3782 17034 3834
rect 17046 3782 17098 3834
rect 17110 3782 17162 3834
rect 17174 3782 17226 3834
rect 1584 3723 1636 3732
rect 1584 3689 1593 3723
rect 1593 3689 1627 3723
rect 1627 3689 1636 3723
rect 1584 3680 1636 3689
rect 1952 3723 2004 3732
rect 1952 3689 1961 3723
rect 1961 3689 1995 3723
rect 1995 3689 2004 3723
rect 1952 3680 2004 3689
rect 5172 3723 5224 3732
rect 5172 3689 5181 3723
rect 5181 3689 5215 3723
rect 5215 3689 5224 3723
rect 5172 3680 5224 3689
rect 5632 3723 5684 3732
rect 5632 3689 5641 3723
rect 5641 3689 5675 3723
rect 5675 3689 5684 3723
rect 5632 3680 5684 3689
rect 7104 3723 7156 3732
rect 7104 3689 7113 3723
rect 7113 3689 7147 3723
rect 7147 3689 7156 3723
rect 7104 3680 7156 3689
rect 8760 3680 8812 3732
rect 11060 3680 11112 3732
rect 12716 3723 12768 3732
rect 3976 3612 4028 3664
rect 4804 3655 4856 3664
rect 4252 3587 4304 3596
rect 4252 3553 4261 3587
rect 4261 3553 4295 3587
rect 4295 3553 4304 3587
rect 4252 3544 4304 3553
rect 4804 3621 4813 3655
rect 4813 3621 4847 3655
rect 4847 3621 4856 3655
rect 4804 3612 4856 3621
rect 9956 3612 10008 3664
rect 5816 3544 5868 3596
rect 6644 3544 6696 3596
rect 7564 3587 7616 3596
rect 7564 3553 7573 3587
rect 7573 3553 7607 3587
rect 7607 3553 7616 3587
rect 7564 3544 7616 3553
rect 8116 3587 8168 3596
rect 8116 3553 8125 3587
rect 8125 3553 8159 3587
rect 8159 3553 8168 3587
rect 8116 3544 8168 3553
rect 11520 3612 11572 3664
rect 12716 3689 12725 3723
rect 12725 3689 12759 3723
rect 12759 3689 12768 3723
rect 12716 3680 12768 3689
rect 13452 3723 13504 3732
rect 13452 3689 13461 3723
rect 13461 3689 13495 3723
rect 13495 3689 13504 3723
rect 13452 3680 13504 3689
rect 15016 3723 15068 3732
rect 15016 3689 15025 3723
rect 15025 3689 15059 3723
rect 15059 3689 15068 3723
rect 15016 3680 15068 3689
rect 18144 3723 18196 3732
rect 18144 3689 18153 3723
rect 18153 3689 18187 3723
rect 18187 3689 18196 3723
rect 18144 3680 18196 3689
rect 8852 3476 8904 3528
rect 11796 3519 11848 3528
rect 11796 3485 11805 3519
rect 11805 3485 11839 3519
rect 11839 3485 11848 3519
rect 11796 3476 11848 3485
rect 12808 3476 12860 3528
rect 7472 3451 7524 3460
rect 7472 3417 7481 3451
rect 7481 3417 7515 3451
rect 7515 3417 7524 3451
rect 7472 3408 7524 3417
rect 4982 3238 5034 3290
rect 5046 3238 5098 3290
rect 5110 3238 5162 3290
rect 5174 3238 5226 3290
rect 12982 3238 13034 3290
rect 13046 3238 13098 3290
rect 13110 3238 13162 3290
rect 13174 3238 13226 3290
rect 20982 3238 21034 3290
rect 21046 3238 21098 3290
rect 21110 3238 21162 3290
rect 21174 3238 21226 3290
rect 5356 3136 5408 3188
rect 5816 3179 5868 3188
rect 5816 3145 5825 3179
rect 5825 3145 5859 3179
rect 5859 3145 5868 3179
rect 5816 3136 5868 3145
rect 6644 3179 6696 3188
rect 6644 3145 6653 3179
rect 6653 3145 6687 3179
rect 6687 3145 6696 3179
rect 6644 3136 6696 3145
rect 8852 3136 8904 3188
rect 11520 3179 11572 3188
rect 11520 3145 11529 3179
rect 11529 3145 11563 3179
rect 11563 3145 11572 3179
rect 11520 3136 11572 3145
rect 12440 3136 12492 3188
rect 5540 3068 5592 3120
rect 8392 3043 8444 3052
rect 5356 2975 5408 2984
rect 5356 2941 5365 2975
rect 5365 2941 5399 2975
rect 5399 2941 5408 2975
rect 5356 2932 5408 2941
rect 7932 2975 7984 2984
rect 7932 2941 7941 2975
rect 7941 2941 7975 2975
rect 7975 2941 7984 2975
rect 7932 2932 7984 2941
rect 8392 3009 8401 3043
rect 8401 3009 8435 3043
rect 8435 3009 8444 3043
rect 8392 3000 8444 3009
rect 11060 3068 11112 3120
rect 13360 3136 13412 3188
rect 12808 3068 12860 3120
rect 11796 3000 11848 3052
rect 8116 2864 8168 2916
rect 10508 2864 10560 2916
rect 4252 2796 4304 2848
rect 9772 2796 9824 2848
rect 9956 2839 10008 2848
rect 9956 2805 9965 2839
rect 9965 2805 9999 2839
rect 9999 2805 10008 2839
rect 9956 2796 10008 2805
rect 12440 2796 12492 2848
rect 8982 2694 9034 2746
rect 9046 2694 9098 2746
rect 9110 2694 9162 2746
rect 9174 2694 9226 2746
rect 16982 2694 17034 2746
rect 17046 2694 17098 2746
rect 17110 2694 17162 2746
rect 17174 2694 17226 2746
rect 6552 2592 6604 2644
rect 7932 2635 7984 2644
rect 7932 2601 7941 2635
rect 7941 2601 7975 2635
rect 7975 2601 7984 2635
rect 7932 2592 7984 2601
rect 8392 2635 8444 2644
rect 8392 2601 8401 2635
rect 8401 2601 8435 2635
rect 8435 2601 8444 2635
rect 8392 2592 8444 2601
rect 9956 2592 10008 2644
rect 10692 2635 10744 2644
rect 10692 2601 10701 2635
rect 10701 2601 10735 2635
rect 10735 2601 10744 2635
rect 10692 2592 10744 2601
rect 6920 2567 6972 2576
rect 6920 2533 6929 2567
rect 6929 2533 6963 2567
rect 6963 2533 6972 2567
rect 6920 2524 6972 2533
rect 13360 2567 13412 2576
rect 13360 2533 13369 2567
rect 13369 2533 13403 2567
rect 13403 2533 13412 2567
rect 13360 2524 13412 2533
rect 1216 2320 1268 2372
rect 8208 2456 8260 2508
rect 9772 2499 9824 2508
rect 9772 2465 9781 2499
rect 9781 2465 9815 2499
rect 9815 2465 9824 2499
rect 9772 2456 9824 2465
rect 6736 2388 6788 2440
rect 9404 2388 9456 2440
rect 17132 2499 17184 2508
rect 12072 2320 12124 2372
rect 5908 2295 5960 2304
rect 5908 2261 5917 2295
rect 5917 2261 5951 2295
rect 5951 2261 5960 2295
rect 5908 2252 5960 2261
rect 14096 2252 14148 2304
rect 17132 2465 17141 2499
rect 17141 2465 17175 2499
rect 17175 2465 17184 2499
rect 17132 2456 17184 2465
rect 17960 2456 18012 2508
rect 19432 2320 19484 2372
rect 15292 2252 15344 2304
rect 4982 2150 5034 2202
rect 5046 2150 5098 2202
rect 5110 2150 5162 2202
rect 5174 2150 5226 2202
rect 12982 2150 13034 2202
rect 13046 2150 13098 2202
rect 13110 2150 13162 2202
rect 13174 2150 13226 2202
rect 20982 2150 21034 2202
rect 21046 2150 21098 2202
rect 21110 2150 21162 2202
rect 21174 2150 21226 2202
<< metal2 >>
rect 938 23610 994 24000
rect 2870 23610 2926 24000
rect 4894 23610 4950 24000
rect 938 23582 1256 23610
rect 938 23520 994 23582
rect 1228 19718 1256 23582
rect 2870 23582 3280 23610
rect 2870 23520 2926 23582
rect 1306 22536 1362 22545
rect 1306 22471 1362 22480
rect 1320 20466 1348 22471
rect 2134 20904 2190 20913
rect 2134 20839 2190 20848
rect 1308 20460 1360 20466
rect 1308 20402 1360 20408
rect 1768 20256 1820 20262
rect 1768 20198 1820 20204
rect 1216 19712 1268 19718
rect 1216 19654 1268 19660
rect 1306 19272 1362 19281
rect 1306 19207 1362 19216
rect 1320 18902 1348 19207
rect 1308 18896 1360 18902
rect 1308 18838 1360 18844
rect 1676 18828 1728 18834
rect 1676 18770 1728 18776
rect 1688 18086 1716 18770
rect 1676 18080 1728 18086
rect 1676 18022 1728 18028
rect 1306 17776 1362 17785
rect 1306 17711 1362 17720
rect 1320 15638 1348 17711
rect 1688 17270 1716 18022
rect 1676 17264 1728 17270
rect 1676 17206 1728 17212
rect 1676 16652 1728 16658
rect 1676 16594 1728 16600
rect 1582 16280 1638 16289
rect 1582 16215 1638 16224
rect 1596 16182 1624 16215
rect 1584 16176 1636 16182
rect 1584 16118 1636 16124
rect 1308 15632 1360 15638
rect 1308 15574 1360 15580
rect 1688 15434 1716 16594
rect 1676 15428 1728 15434
rect 1676 15370 1728 15376
rect 1584 14272 1636 14278
rect 1584 14214 1636 14220
rect 1596 13938 1624 14214
rect 1584 13932 1636 13938
rect 1584 13874 1636 13880
rect 18 13424 74 13433
rect 18 13359 74 13368
rect 32 9042 60 13359
rect 1596 12442 1624 13874
rect 1688 12782 1716 15370
rect 1676 12776 1728 12782
rect 1676 12718 1728 12724
rect 1688 12442 1716 12718
rect 1584 12436 1636 12442
rect 1584 12378 1636 12384
rect 1676 12436 1728 12442
rect 1676 12378 1728 12384
rect 112 11552 164 11558
rect 112 11494 164 11500
rect 124 10305 152 11494
rect 110 10296 166 10305
rect 110 10231 166 10240
rect 1492 10056 1544 10062
rect 1492 9998 1544 10004
rect 110 9616 166 9625
rect 1504 9586 1532 9998
rect 110 9551 166 9560
rect 1492 9580 1544 9586
rect 20 9036 72 9042
rect 20 8978 72 8984
rect 124 8673 152 9551
rect 1492 9522 1544 9528
rect 1688 9518 1716 12378
rect 1780 12209 1808 20198
rect 1952 18080 2004 18086
rect 1952 18022 2004 18028
rect 1860 17536 1912 17542
rect 1860 17478 1912 17484
rect 1872 16794 1900 17478
rect 1964 17202 1992 18022
rect 1952 17196 2004 17202
rect 1952 17138 2004 17144
rect 2148 16810 2176 20839
rect 2412 18420 2464 18426
rect 2412 18362 2464 18368
rect 2228 17876 2280 17882
rect 2228 17818 2280 17824
rect 2240 17338 2268 17818
rect 2228 17332 2280 17338
rect 2228 17274 2280 17280
rect 2240 16998 2268 17274
rect 2228 16992 2280 16998
rect 2228 16934 2280 16940
rect 1860 16788 1912 16794
rect 2148 16782 2268 16810
rect 1860 16730 1912 16736
rect 1952 16108 2004 16114
rect 1952 16050 2004 16056
rect 1964 15706 1992 16050
rect 1952 15700 2004 15706
rect 1952 15642 2004 15648
rect 2136 15564 2188 15570
rect 2136 15506 2188 15512
rect 1952 14816 2004 14822
rect 1952 14758 2004 14764
rect 1860 13456 1912 13462
rect 1860 13398 1912 13404
rect 1872 12374 1900 13398
rect 1964 12782 1992 14758
rect 2148 14006 2176 15506
rect 2136 14000 2188 14006
rect 2136 13942 2188 13948
rect 2044 13796 2096 13802
rect 2044 13738 2096 13744
rect 2056 13530 2084 13738
rect 2044 13524 2096 13530
rect 2044 13466 2096 13472
rect 2136 13320 2188 13326
rect 2136 13262 2188 13268
rect 2148 12850 2176 13262
rect 2136 12844 2188 12850
rect 2136 12786 2188 12792
rect 1952 12776 2004 12782
rect 1952 12718 2004 12724
rect 1860 12368 1912 12374
rect 1860 12310 1912 12316
rect 1766 12200 1822 12209
rect 1766 12135 1822 12144
rect 1872 11898 1900 12310
rect 1860 11892 1912 11898
rect 1912 11852 1992 11880
rect 1860 11834 1912 11840
rect 1768 11008 1820 11014
rect 1768 10950 1820 10956
rect 1780 10674 1808 10950
rect 1768 10668 1820 10674
rect 1768 10610 1820 10616
rect 1858 10296 1914 10305
rect 1964 10266 1992 11852
rect 2240 10810 2268 16782
rect 2320 16040 2372 16046
rect 2320 15982 2372 15988
rect 2332 15366 2360 15982
rect 2320 15360 2372 15366
rect 2320 15302 2372 15308
rect 2332 14958 2360 15302
rect 2320 14952 2372 14958
rect 2320 14894 2372 14900
rect 2332 14550 2360 14894
rect 2320 14544 2372 14550
rect 2320 14486 2372 14492
rect 2332 11286 2360 14486
rect 2424 12866 2452 18362
rect 3148 18148 3200 18154
rect 3148 18090 3200 18096
rect 2780 17536 2832 17542
rect 2780 17478 2832 17484
rect 2792 17066 2820 17478
rect 2780 17060 2832 17066
rect 2780 17002 2832 17008
rect 2596 16992 2648 16998
rect 2596 16934 2648 16940
rect 2608 14618 2636 16934
rect 2792 16794 2820 17002
rect 2780 16788 2832 16794
rect 2780 16730 2832 16736
rect 3160 16658 3188 18090
rect 3148 16652 3200 16658
rect 3148 16594 3200 16600
rect 3160 16046 3188 16594
rect 3148 16040 3200 16046
rect 3148 15982 3200 15988
rect 3056 15564 3108 15570
rect 3056 15506 3108 15512
rect 3068 15162 3096 15506
rect 3056 15156 3108 15162
rect 3056 15098 3108 15104
rect 2780 14884 2832 14890
rect 2780 14826 2832 14832
rect 2596 14612 2648 14618
rect 2596 14554 2648 14560
rect 2608 14074 2636 14554
rect 2792 14414 2820 14826
rect 2780 14408 2832 14414
rect 2780 14350 2832 14356
rect 2792 14074 2820 14350
rect 2596 14068 2648 14074
rect 2596 14010 2648 14016
rect 2780 14068 2832 14074
rect 2780 14010 2832 14016
rect 2504 13456 2556 13462
rect 2608 13444 2636 14010
rect 2556 13416 2636 13444
rect 2504 13398 2556 13404
rect 2424 12838 2544 12866
rect 2516 12594 2544 12838
rect 2872 12640 2924 12646
rect 2516 12566 2636 12594
rect 2872 12582 2924 12588
rect 2608 12238 2636 12566
rect 2884 12306 2912 12582
rect 2872 12300 2924 12306
rect 2872 12242 2924 12248
rect 2596 12232 2648 12238
rect 2596 12174 2648 12180
rect 2320 11280 2372 11286
rect 2320 11222 2372 11228
rect 2608 11014 2636 12174
rect 2884 11626 2912 12242
rect 3148 12232 3200 12238
rect 3148 12174 3200 12180
rect 3160 11762 3188 12174
rect 3148 11756 3200 11762
rect 3148 11698 3200 11704
rect 2872 11620 2924 11626
rect 2872 11562 2924 11568
rect 3160 11354 3188 11698
rect 3148 11348 3200 11354
rect 3148 11290 3200 11296
rect 3056 11280 3108 11286
rect 3056 11222 3108 11228
rect 2780 11212 2832 11218
rect 2780 11154 2832 11160
rect 2596 11008 2648 11014
rect 2596 10950 2648 10956
rect 2228 10804 2280 10810
rect 2228 10746 2280 10752
rect 2792 10742 2820 11154
rect 2780 10736 2832 10742
rect 2832 10696 2912 10724
rect 2780 10678 2832 10684
rect 2228 10532 2280 10538
rect 2228 10474 2280 10480
rect 2240 10266 2268 10474
rect 1858 10231 1914 10240
rect 1952 10260 2004 10266
rect 1676 9512 1728 9518
rect 1676 9454 1728 9460
rect 1872 9110 1900 10231
rect 1952 10202 2004 10208
rect 2228 10260 2280 10266
rect 2228 10202 2280 10208
rect 1964 9722 1992 10202
rect 1952 9716 2004 9722
rect 1952 9658 2004 9664
rect 2884 9518 2912 10696
rect 3068 10470 3096 11222
rect 3148 11144 3200 11150
rect 3148 11086 3200 11092
rect 3056 10464 3108 10470
rect 3056 10406 3108 10412
rect 2872 9512 2924 9518
rect 2872 9454 2924 9460
rect 1860 9104 1912 9110
rect 1860 9046 1912 9052
rect 2884 9042 2912 9454
rect 2964 9444 3016 9450
rect 2964 9386 3016 9392
rect 2976 9353 3004 9386
rect 2962 9344 3018 9353
rect 2962 9279 3018 9288
rect 2688 9036 2740 9042
rect 2688 8978 2740 8984
rect 2872 9036 2924 9042
rect 2872 8978 2924 8984
rect 2504 8968 2556 8974
rect 2504 8910 2556 8916
rect 1492 8900 1544 8906
rect 1492 8842 1544 8848
rect 110 8664 166 8673
rect 110 8599 166 8608
rect 1504 7886 1532 8842
rect 2516 8634 2544 8910
rect 2700 8634 2728 8978
rect 2504 8628 2556 8634
rect 2504 8570 2556 8576
rect 2688 8628 2740 8634
rect 2688 8570 2740 8576
rect 1952 8424 2004 8430
rect 1952 8366 2004 8372
rect 1676 8288 1728 8294
rect 1676 8230 1728 8236
rect 1688 8022 1716 8230
rect 1676 8016 1728 8022
rect 1676 7958 1728 7964
rect 1492 7880 1544 7886
rect 1492 7822 1544 7828
rect 1504 7002 1532 7822
rect 1688 7546 1716 7958
rect 1676 7540 1728 7546
rect 1676 7482 1728 7488
rect 1964 7274 1992 8366
rect 2136 7880 2188 7886
rect 2136 7822 2188 7828
rect 2148 7478 2176 7822
rect 2780 7744 2832 7750
rect 2780 7686 2832 7692
rect 2136 7472 2188 7478
rect 2136 7414 2188 7420
rect 1952 7268 2004 7274
rect 1952 7210 2004 7216
rect 1492 6996 1544 7002
rect 1492 6938 1544 6944
rect 1964 6730 1992 7210
rect 2044 6928 2096 6934
rect 2044 6870 2096 6876
rect 1952 6724 2004 6730
rect 1952 6666 2004 6672
rect 2056 6458 2084 6870
rect 2044 6452 2096 6458
rect 2044 6394 2096 6400
rect 112 6112 164 6118
rect 112 6054 164 6060
rect 124 5545 152 6054
rect 1952 5840 2004 5846
rect 1952 5782 2004 5788
rect 110 5536 166 5545
rect 110 5471 166 5480
rect 1964 5370 1992 5782
rect 1952 5364 2004 5370
rect 1952 5306 2004 5312
rect 2056 5302 2084 6394
rect 2148 5710 2176 7414
rect 2792 7410 2820 7686
rect 2884 7410 2912 8978
rect 2780 7404 2832 7410
rect 2780 7346 2832 7352
rect 2872 7404 2924 7410
rect 2872 7346 2924 7352
rect 2320 6792 2372 6798
rect 2320 6734 2372 6740
rect 2228 6248 2280 6254
rect 2228 6190 2280 6196
rect 2240 5710 2268 6190
rect 2332 6118 2360 6734
rect 2320 6112 2372 6118
rect 2320 6054 2372 6060
rect 2136 5704 2188 5710
rect 2136 5646 2188 5652
rect 2228 5704 2280 5710
rect 2228 5646 2280 5652
rect 2044 5296 2096 5302
rect 2044 5238 2096 5244
rect 2056 5098 2084 5238
rect 2044 5092 2096 5098
rect 2044 5034 2096 5040
rect 2240 4758 2268 5646
rect 2412 5364 2464 5370
rect 2412 5306 2464 5312
rect 2424 4826 2452 5306
rect 2872 5092 2924 5098
rect 2872 5034 2924 5040
rect 2412 4820 2464 4826
rect 2412 4762 2464 4768
rect 1584 4752 1636 4758
rect 1584 4694 1636 4700
rect 2228 4752 2280 4758
rect 2228 4694 2280 4700
rect 1596 4010 1624 4694
rect 1952 4616 2004 4622
rect 1952 4558 2004 4564
rect 1584 4004 1636 4010
rect 1584 3946 1636 3952
rect 204 3936 256 3942
rect 110 3904 166 3913
rect 166 3884 204 3890
rect 166 3878 256 3884
rect 166 3862 244 3878
rect 110 3839 166 3848
rect 1596 3738 1624 3946
rect 1964 3738 1992 4558
rect 2424 4282 2452 4762
rect 2412 4276 2464 4282
rect 2412 4218 2464 4224
rect 2424 4078 2452 4218
rect 2412 4072 2464 4078
rect 2412 4014 2464 4020
rect 1584 3732 1636 3738
rect 1584 3674 1636 3680
rect 1952 3732 2004 3738
rect 1952 3674 2004 3680
rect 1216 2372 1268 2378
rect 1216 2314 1268 2320
rect 938 82 994 480
rect 1228 82 1256 2314
rect 938 54 1256 82
rect 2778 82 2834 480
rect 2884 82 2912 5034
rect 3068 4146 3096 10406
rect 3160 10130 3188 11086
rect 3148 10124 3200 10130
rect 3148 10066 3200 10072
rect 3148 8288 3200 8294
rect 3148 8230 3200 8236
rect 3160 8090 3188 8230
rect 3148 8084 3200 8090
rect 3148 8026 3200 8032
rect 3148 7948 3200 7954
rect 3252 7936 3280 23582
rect 4724 23582 4950 23610
rect 3424 18216 3476 18222
rect 3424 18158 3476 18164
rect 3436 17882 3464 18158
rect 4068 18148 4120 18154
rect 4068 18090 4120 18096
rect 3424 17876 3476 17882
rect 3424 17818 3476 17824
rect 3436 14958 3464 17818
rect 4080 17746 4108 18090
rect 4436 18080 4488 18086
rect 4436 18022 4488 18028
rect 4160 17808 4212 17814
rect 4160 17750 4212 17756
rect 4068 17740 4120 17746
rect 4068 17682 4120 17688
rect 4080 17338 4108 17682
rect 4068 17332 4120 17338
rect 4068 17274 4120 17280
rect 4172 16998 4200 17750
rect 4448 17066 4476 18022
rect 4724 17746 4752 23582
rect 4894 23520 4950 23582
rect 6918 23610 6974 24000
rect 8942 23610 8998 24000
rect 10874 23610 10930 24000
rect 6918 23582 7052 23610
rect 6918 23520 6974 23582
rect 4956 21788 5252 21808
rect 5012 21786 5036 21788
rect 5092 21786 5116 21788
rect 5172 21786 5196 21788
rect 5034 21734 5036 21786
rect 5098 21734 5110 21786
rect 5172 21734 5174 21786
rect 5012 21732 5036 21734
rect 5092 21732 5116 21734
rect 5172 21732 5196 21734
rect 4956 21712 5252 21732
rect 4956 20700 5252 20720
rect 5012 20698 5036 20700
rect 5092 20698 5116 20700
rect 5172 20698 5196 20700
rect 5034 20646 5036 20698
rect 5098 20646 5110 20698
rect 5172 20646 5174 20698
rect 5012 20644 5036 20646
rect 5092 20644 5116 20646
rect 5172 20644 5196 20646
rect 4956 20624 5252 20644
rect 7024 20602 7052 23582
rect 8680 23582 8998 23610
rect 8680 20602 8708 23582
rect 8942 23520 8998 23582
rect 10796 23582 10930 23610
rect 8956 21244 9252 21264
rect 9012 21242 9036 21244
rect 9092 21242 9116 21244
rect 9172 21242 9196 21244
rect 9034 21190 9036 21242
rect 9098 21190 9110 21242
rect 9172 21190 9174 21242
rect 9012 21188 9036 21190
rect 9092 21188 9116 21190
rect 9172 21188 9196 21190
rect 8956 21168 9252 21188
rect 10796 20602 10824 23582
rect 10874 23520 10930 23582
rect 12898 23610 12954 24000
rect 14922 23610 14978 24000
rect 16946 23610 17002 24000
rect 12898 23582 13308 23610
rect 12898 23520 12954 23582
rect 12956 21788 13252 21808
rect 13012 21786 13036 21788
rect 13092 21786 13116 21788
rect 13172 21786 13196 21788
rect 13034 21734 13036 21786
rect 13098 21734 13110 21786
rect 13172 21734 13174 21786
rect 13012 21732 13036 21734
rect 13092 21732 13116 21734
rect 13172 21732 13196 21734
rect 12956 21712 13252 21732
rect 12956 20700 13252 20720
rect 13012 20698 13036 20700
rect 13092 20698 13116 20700
rect 13172 20698 13196 20700
rect 13034 20646 13036 20698
rect 13098 20646 13110 20698
rect 13172 20646 13174 20698
rect 13012 20644 13036 20646
rect 13092 20644 13116 20646
rect 13172 20644 13196 20646
rect 12956 20624 13252 20644
rect 7012 20596 7064 20602
rect 7012 20538 7064 20544
rect 8668 20596 8720 20602
rect 8668 20538 8720 20544
rect 10784 20596 10836 20602
rect 10784 20538 10836 20544
rect 5632 20392 5684 20398
rect 5632 20334 5684 20340
rect 4956 19612 5252 19632
rect 5012 19610 5036 19612
rect 5092 19610 5116 19612
rect 5172 19610 5196 19612
rect 5034 19558 5036 19610
rect 5098 19558 5110 19610
rect 5172 19558 5174 19610
rect 5012 19556 5036 19558
rect 5092 19556 5116 19558
rect 5172 19556 5196 19558
rect 4956 19536 5252 19556
rect 4804 18624 4856 18630
rect 4804 18566 4856 18572
rect 4816 18290 4844 18566
rect 4956 18524 5252 18544
rect 5012 18522 5036 18524
rect 5092 18522 5116 18524
rect 5172 18522 5196 18524
rect 5034 18470 5036 18522
rect 5098 18470 5110 18522
rect 5172 18470 5174 18522
rect 5012 18468 5036 18470
rect 5092 18468 5116 18470
rect 5172 18468 5196 18470
rect 4956 18448 5252 18468
rect 5540 18352 5592 18358
rect 5540 18294 5592 18300
rect 4804 18284 4856 18290
rect 4804 18226 4856 18232
rect 5356 18284 5408 18290
rect 5356 18226 5408 18232
rect 4712 17740 4764 17746
rect 4712 17682 4764 17688
rect 4712 17264 4764 17270
rect 4712 17206 4764 17212
rect 4436 17060 4488 17066
rect 4436 17002 4488 17008
rect 4160 16992 4212 16998
rect 4160 16934 4212 16940
rect 4172 16726 4200 16934
rect 4160 16720 4212 16726
rect 4160 16662 4212 16668
rect 4068 16584 4120 16590
rect 4068 16526 4120 16532
rect 4080 16250 4108 16526
rect 4172 16250 4200 16662
rect 4068 16244 4120 16250
rect 4068 16186 4120 16192
rect 4160 16244 4212 16250
rect 4160 16186 4212 16192
rect 3608 15972 3660 15978
rect 3608 15914 3660 15920
rect 3424 14952 3476 14958
rect 3424 14894 3476 14900
rect 3436 14618 3464 14894
rect 3424 14612 3476 14618
rect 3424 14554 3476 14560
rect 3620 12986 3648 15914
rect 3884 14816 3936 14822
rect 3884 14758 3936 14764
rect 3700 14612 3752 14618
rect 3700 14554 3752 14560
rect 3712 13814 3740 14554
rect 3896 14482 3924 14758
rect 4172 14618 4200 16186
rect 4448 16114 4476 17002
rect 4436 16108 4488 16114
rect 4436 16050 4488 16056
rect 4724 15978 4752 17206
rect 4816 16590 4844 18226
rect 5172 18080 5224 18086
rect 5172 18022 5224 18028
rect 5184 17882 5212 18022
rect 5172 17876 5224 17882
rect 5172 17818 5224 17824
rect 4956 17436 5252 17456
rect 5012 17434 5036 17436
rect 5092 17434 5116 17436
rect 5172 17434 5196 17436
rect 5034 17382 5036 17434
rect 5098 17382 5110 17434
rect 5172 17382 5174 17434
rect 5012 17380 5036 17382
rect 5092 17380 5116 17382
rect 5172 17380 5196 17382
rect 4956 17360 5252 17380
rect 5368 17202 5396 18226
rect 5356 17196 5408 17202
rect 5356 17138 5408 17144
rect 4988 16992 5040 16998
rect 4988 16934 5040 16940
rect 5000 16794 5028 16934
rect 4988 16788 5040 16794
rect 4988 16730 5040 16736
rect 4804 16584 4856 16590
rect 4804 16526 4856 16532
rect 4956 16348 5252 16368
rect 5012 16346 5036 16348
rect 5092 16346 5116 16348
rect 5172 16346 5196 16348
rect 5034 16294 5036 16346
rect 5098 16294 5110 16346
rect 5172 16294 5174 16346
rect 5012 16292 5036 16294
rect 5092 16292 5116 16294
rect 5172 16292 5196 16294
rect 4956 16272 5252 16292
rect 4804 16244 4856 16250
rect 4804 16186 4856 16192
rect 4816 15978 4844 16186
rect 5448 16040 5500 16046
rect 5448 15982 5500 15988
rect 4712 15972 4764 15978
rect 4712 15914 4764 15920
rect 4804 15972 4856 15978
rect 4804 15914 4856 15920
rect 4804 15564 4856 15570
rect 4804 15506 4856 15512
rect 4816 14822 4844 15506
rect 4956 15260 5252 15280
rect 5012 15258 5036 15260
rect 5092 15258 5116 15260
rect 5172 15258 5196 15260
rect 5034 15206 5036 15258
rect 5098 15206 5110 15258
rect 5172 15206 5174 15258
rect 5012 15204 5036 15206
rect 5092 15204 5116 15206
rect 5172 15204 5196 15206
rect 4956 15184 5252 15204
rect 5356 14884 5408 14890
rect 5356 14826 5408 14832
rect 4804 14816 4856 14822
rect 4804 14758 4856 14764
rect 4160 14612 4212 14618
rect 4160 14554 4212 14560
rect 3884 14476 3936 14482
rect 3884 14418 3936 14424
rect 3792 14340 3844 14346
rect 3792 14282 3844 14288
rect 3804 13954 3832 14282
rect 3896 14074 3924 14418
rect 4172 14074 4200 14554
rect 4710 14512 4766 14521
rect 4710 14447 4766 14456
rect 4528 14272 4580 14278
rect 4528 14214 4580 14220
rect 3884 14068 3936 14074
rect 3884 14010 3936 14016
rect 4160 14068 4212 14074
rect 4160 14010 4212 14016
rect 4252 14000 4304 14006
rect 3804 13926 3924 13954
rect 4252 13942 4304 13948
rect 3712 13786 3832 13814
rect 3896 13802 3924 13926
rect 4264 13802 4292 13942
rect 3608 12980 3660 12986
rect 3608 12922 3660 12928
rect 3620 12782 3648 12922
rect 3608 12776 3660 12782
rect 3608 12718 3660 12724
rect 3424 12640 3476 12646
rect 3424 12582 3476 12588
rect 3436 12238 3464 12582
rect 3424 12232 3476 12238
rect 3424 12174 3476 12180
rect 3516 11892 3568 11898
rect 3516 11834 3568 11840
rect 3528 11626 3556 11834
rect 3516 11620 3568 11626
rect 3568 11580 3648 11608
rect 3516 11562 3568 11568
rect 3516 11008 3568 11014
rect 3516 10950 3568 10956
rect 3200 7908 3280 7936
rect 3148 7890 3200 7896
rect 3160 7857 3188 7890
rect 3146 7848 3202 7857
rect 3146 7783 3202 7792
rect 3160 7546 3188 7783
rect 3528 7750 3556 10950
rect 3620 10810 3648 11580
rect 3608 10804 3660 10810
rect 3608 10746 3660 10752
rect 3608 10668 3660 10674
rect 3608 10610 3660 10616
rect 3620 9110 3648 10610
rect 3700 10124 3752 10130
rect 3700 10066 3752 10072
rect 3712 9722 3740 10066
rect 3700 9716 3752 9722
rect 3700 9658 3752 9664
rect 3804 9178 3832 13786
rect 3884 13796 3936 13802
rect 3884 13738 3936 13744
rect 4252 13796 4304 13802
rect 4252 13738 4304 13744
rect 3896 13530 3924 13738
rect 3884 13524 3936 13530
rect 3884 13466 3936 13472
rect 4264 13258 4292 13738
rect 4540 13462 4568 14214
rect 4620 14000 4672 14006
rect 4620 13942 4672 13948
rect 4528 13456 4580 13462
rect 4528 13398 4580 13404
rect 4436 13320 4488 13326
rect 4436 13262 4488 13268
rect 4252 13252 4304 13258
rect 4252 13194 4304 13200
rect 4448 12918 4476 13262
rect 4540 12986 4568 13398
rect 4528 12980 4580 12986
rect 4528 12922 4580 12928
rect 4436 12912 4488 12918
rect 4436 12854 4488 12860
rect 4252 12708 4304 12714
rect 4252 12650 4304 12656
rect 4264 12374 4292 12650
rect 4448 12442 4476 12854
rect 4436 12436 4488 12442
rect 4436 12378 4488 12384
rect 4252 12368 4304 12374
rect 4252 12310 4304 12316
rect 4160 12232 4212 12238
rect 4160 12174 4212 12180
rect 4172 11354 4200 12174
rect 4264 11898 4292 12310
rect 4632 12238 4660 13942
rect 4724 13297 4752 14447
rect 4816 14056 4844 14758
rect 5368 14618 5396 14826
rect 5460 14822 5488 15982
rect 5552 15638 5580 18294
rect 5540 15632 5592 15638
rect 5540 15574 5592 15580
rect 5552 15162 5580 15574
rect 5540 15156 5592 15162
rect 5540 15098 5592 15104
rect 5552 14958 5580 15098
rect 5540 14952 5592 14958
rect 5540 14894 5592 14900
rect 5448 14816 5500 14822
rect 5448 14758 5500 14764
rect 5356 14612 5408 14618
rect 5356 14554 5408 14560
rect 4956 14172 5252 14192
rect 5012 14170 5036 14172
rect 5092 14170 5116 14172
rect 5172 14170 5196 14172
rect 5034 14118 5036 14170
rect 5098 14118 5110 14170
rect 5172 14118 5174 14170
rect 5012 14116 5036 14118
rect 5092 14116 5116 14118
rect 5172 14116 5196 14118
rect 4956 14096 5252 14116
rect 4816 14028 4936 14056
rect 4908 13870 4936 14028
rect 4896 13864 4948 13870
rect 4896 13806 4948 13812
rect 4710 13288 4766 13297
rect 4710 13223 4766 13232
rect 4956 13084 5252 13104
rect 5012 13082 5036 13084
rect 5092 13082 5116 13084
rect 5172 13082 5196 13084
rect 5034 13030 5036 13082
rect 5098 13030 5110 13082
rect 5172 13030 5174 13082
rect 5012 13028 5036 13030
rect 5092 13028 5116 13030
rect 5172 13028 5196 13030
rect 4956 13008 5252 13028
rect 5644 12986 5672 20334
rect 8392 20256 8444 20262
rect 8392 20198 8444 20204
rect 11980 20256 12032 20262
rect 11980 20198 12032 20204
rect 7472 18896 7524 18902
rect 7472 18838 7524 18844
rect 7104 18828 7156 18834
rect 7104 18770 7156 18776
rect 7116 18358 7144 18770
rect 7196 18760 7248 18766
rect 7196 18702 7248 18708
rect 7104 18352 7156 18358
rect 7104 18294 7156 18300
rect 7208 17746 7236 18702
rect 7484 18426 7512 18838
rect 8300 18624 8352 18630
rect 8300 18566 8352 18572
rect 7472 18420 7524 18426
rect 7472 18362 7524 18368
rect 7484 18086 7512 18362
rect 8312 18154 8340 18566
rect 8300 18148 8352 18154
rect 8300 18090 8352 18096
rect 7472 18080 7524 18086
rect 7472 18022 7524 18028
rect 7932 18080 7984 18086
rect 7932 18022 7984 18028
rect 6000 17740 6052 17746
rect 6000 17682 6052 17688
rect 7196 17740 7248 17746
rect 7196 17682 7248 17688
rect 5908 17536 5960 17542
rect 5908 17478 5960 17484
rect 5920 16726 5948 17478
rect 6012 17338 6040 17682
rect 6000 17332 6052 17338
rect 6052 17292 6132 17320
rect 6000 17274 6052 17280
rect 5908 16720 5960 16726
rect 5908 16662 5960 16668
rect 6000 16720 6052 16726
rect 6000 16662 6052 16668
rect 6012 16250 6040 16662
rect 6000 16244 6052 16250
rect 6000 16186 6052 16192
rect 6000 15564 6052 15570
rect 6000 15506 6052 15512
rect 5908 15156 5960 15162
rect 5908 15098 5960 15104
rect 5632 12980 5684 12986
rect 5632 12922 5684 12928
rect 5644 12782 5672 12922
rect 4804 12776 4856 12782
rect 4804 12718 4856 12724
rect 5632 12776 5684 12782
rect 5632 12718 5684 12724
rect 4620 12232 4672 12238
rect 4620 12174 4672 12180
rect 4252 11892 4304 11898
rect 4252 11834 4304 11840
rect 4816 11665 4844 12718
rect 5540 12096 5592 12102
rect 5540 12038 5592 12044
rect 4956 11996 5252 12016
rect 5012 11994 5036 11996
rect 5092 11994 5116 11996
rect 5172 11994 5196 11996
rect 5034 11942 5036 11994
rect 5098 11942 5110 11994
rect 5172 11942 5174 11994
rect 5012 11940 5036 11942
rect 5092 11940 5116 11942
rect 5172 11940 5196 11942
rect 4956 11920 5252 11940
rect 5552 11694 5580 12038
rect 5540 11688 5592 11694
rect 4802 11656 4858 11665
rect 5540 11630 5592 11636
rect 5724 11688 5776 11694
rect 5724 11630 5776 11636
rect 4802 11591 4858 11600
rect 4160 11348 4212 11354
rect 4816 11336 4844 11591
rect 4160 11290 4212 11296
rect 4632 11308 4844 11336
rect 4252 11008 4304 11014
rect 4252 10950 4304 10956
rect 4264 10674 4292 10950
rect 4252 10668 4304 10674
rect 4252 10610 4304 10616
rect 4436 10532 4488 10538
rect 4436 10474 4488 10480
rect 4448 10266 4476 10474
rect 4436 10260 4488 10266
rect 4436 10202 4488 10208
rect 4068 9920 4120 9926
rect 4068 9862 4120 9868
rect 4080 9382 4108 9862
rect 4448 9722 4476 10202
rect 4436 9716 4488 9722
rect 4436 9658 4488 9664
rect 4068 9376 4120 9382
rect 4068 9318 4120 9324
rect 4080 9178 4108 9318
rect 3792 9172 3844 9178
rect 3792 9114 3844 9120
rect 4068 9172 4120 9178
rect 4068 9114 4120 9120
rect 3608 9104 3660 9110
rect 3608 9046 3660 9052
rect 3804 7993 3832 9114
rect 3976 8288 4028 8294
rect 3976 8230 4028 8236
rect 3790 7984 3846 7993
rect 3790 7919 3846 7928
rect 3516 7744 3568 7750
rect 3516 7686 3568 7692
rect 3148 7540 3200 7546
rect 3148 7482 3200 7488
rect 3424 7404 3476 7410
rect 3424 7346 3476 7352
rect 3148 7200 3200 7206
rect 3148 7142 3200 7148
rect 3160 6934 3188 7142
rect 3436 7002 3464 7346
rect 3528 7342 3556 7686
rect 3516 7336 3568 7342
rect 3516 7278 3568 7284
rect 3424 6996 3476 7002
rect 3424 6938 3476 6944
rect 3148 6928 3200 6934
rect 3148 6870 3200 6876
rect 3240 5908 3292 5914
rect 3240 5850 3292 5856
rect 3252 5370 3280 5850
rect 3240 5364 3292 5370
rect 3240 5306 3292 5312
rect 3528 5137 3556 7278
rect 3988 6905 4016 8230
rect 4436 8084 4488 8090
rect 4436 8026 4488 8032
rect 4068 7880 4120 7886
rect 4068 7822 4120 7828
rect 4080 7342 4108 7822
rect 4448 7546 4476 8026
rect 4436 7540 4488 7546
rect 4436 7482 4488 7488
rect 4068 7336 4120 7342
rect 4068 7278 4120 7284
rect 4080 7002 4108 7278
rect 4448 7206 4476 7482
rect 4436 7200 4488 7206
rect 4436 7142 4488 7148
rect 4068 6996 4120 7002
rect 4068 6938 4120 6944
rect 3974 6896 4030 6905
rect 4632 6866 4660 11308
rect 5356 11280 5408 11286
rect 5356 11222 5408 11228
rect 4712 11212 4764 11218
rect 4712 11154 4764 11160
rect 4724 10742 4752 11154
rect 4804 11076 4856 11082
rect 4804 11018 4856 11024
rect 4712 10736 4764 10742
rect 4712 10678 4764 10684
rect 4816 10266 4844 11018
rect 4956 10908 5252 10928
rect 5012 10906 5036 10908
rect 5092 10906 5116 10908
rect 5172 10906 5196 10908
rect 5034 10854 5036 10906
rect 5098 10854 5110 10906
rect 5172 10854 5174 10906
rect 5012 10852 5036 10854
rect 5092 10852 5116 10854
rect 5172 10852 5196 10854
rect 4956 10832 5252 10852
rect 5368 10810 5396 11222
rect 5552 11218 5580 11630
rect 5540 11212 5592 11218
rect 5540 11154 5592 11160
rect 5448 11076 5500 11082
rect 5448 11018 5500 11024
rect 5356 10804 5408 10810
rect 5356 10746 5408 10752
rect 5460 10606 5488 11018
rect 5448 10600 5500 10606
rect 5448 10542 5500 10548
rect 4804 10260 4856 10266
rect 4804 10202 4856 10208
rect 4712 9104 4764 9110
rect 4712 9046 4764 9052
rect 4816 9058 4844 10202
rect 4956 9820 5252 9840
rect 5012 9818 5036 9820
rect 5092 9818 5116 9820
rect 5172 9818 5196 9820
rect 5034 9766 5036 9818
rect 5098 9766 5110 9818
rect 5172 9766 5174 9818
rect 5012 9764 5036 9766
rect 5092 9764 5116 9766
rect 5172 9764 5196 9766
rect 4956 9744 5252 9764
rect 5356 9716 5408 9722
rect 5356 9658 5408 9664
rect 4724 8294 4752 9046
rect 4816 9030 4936 9058
rect 4908 8974 4936 9030
rect 4804 8968 4856 8974
rect 4804 8910 4856 8916
rect 4896 8968 4948 8974
rect 4896 8910 4948 8916
rect 4712 8288 4764 8294
rect 4712 8230 4764 8236
rect 4816 7750 4844 8910
rect 4956 8732 5252 8752
rect 5012 8730 5036 8732
rect 5092 8730 5116 8732
rect 5172 8730 5196 8732
rect 5034 8678 5036 8730
rect 5098 8678 5110 8730
rect 5172 8678 5174 8730
rect 5012 8676 5036 8678
rect 5092 8676 5116 8678
rect 5172 8676 5196 8678
rect 4956 8656 5252 8676
rect 5368 8566 5396 9658
rect 5460 9586 5488 10542
rect 5540 9920 5592 9926
rect 5540 9862 5592 9868
rect 5448 9580 5500 9586
rect 5448 9522 5500 9528
rect 5356 8560 5408 8566
rect 5356 8502 5408 8508
rect 4988 8288 5040 8294
rect 4988 8230 5040 8236
rect 5000 8090 5028 8230
rect 4988 8084 5040 8090
rect 4988 8026 5040 8032
rect 4804 7744 4856 7750
rect 4804 7686 4856 7692
rect 4816 6934 4844 7686
rect 4956 7644 5252 7664
rect 5012 7642 5036 7644
rect 5092 7642 5116 7644
rect 5172 7642 5196 7644
rect 5034 7590 5036 7642
rect 5098 7590 5110 7642
rect 5172 7590 5174 7642
rect 5012 7588 5036 7590
rect 5092 7588 5116 7590
rect 5172 7588 5196 7590
rect 4956 7568 5252 7588
rect 5448 7336 5500 7342
rect 5552 7324 5580 9862
rect 5500 7296 5580 7324
rect 5448 7278 5500 7284
rect 4804 6928 4856 6934
rect 4804 6870 4856 6876
rect 5356 6928 5408 6934
rect 5356 6870 5408 6876
rect 3974 6831 4030 6840
rect 4620 6860 4672 6866
rect 4620 6802 4672 6808
rect 4632 6458 4660 6802
rect 4956 6556 5252 6576
rect 5012 6554 5036 6556
rect 5092 6554 5116 6556
rect 5172 6554 5196 6556
rect 5034 6502 5036 6554
rect 5098 6502 5110 6554
rect 5172 6502 5174 6554
rect 5012 6500 5036 6502
rect 5092 6500 5116 6502
rect 5172 6500 5196 6502
rect 4956 6480 5252 6500
rect 4620 6452 4672 6458
rect 4620 6394 4672 6400
rect 4632 6361 4660 6394
rect 4618 6352 4674 6361
rect 4618 6287 4674 6296
rect 3700 6248 3752 6254
rect 3700 6190 3752 6196
rect 3712 5778 3740 6190
rect 4804 6112 4856 6118
rect 4804 6054 4856 6060
rect 4816 5896 4844 6054
rect 4988 5908 5040 5914
rect 4816 5868 4988 5896
rect 3700 5772 3752 5778
rect 3700 5714 3752 5720
rect 4160 5772 4212 5778
rect 4160 5714 4212 5720
rect 4172 5370 4200 5714
rect 4816 5710 4844 5868
rect 4988 5850 5040 5856
rect 4804 5704 4856 5710
rect 4804 5646 4856 5652
rect 4816 5370 4844 5646
rect 4956 5468 5252 5488
rect 5012 5466 5036 5468
rect 5092 5466 5116 5468
rect 5172 5466 5196 5468
rect 5034 5414 5036 5466
rect 5098 5414 5110 5466
rect 5172 5414 5174 5466
rect 5012 5412 5036 5414
rect 5092 5412 5116 5414
rect 5172 5412 5196 5414
rect 4956 5392 5252 5412
rect 4160 5364 4212 5370
rect 4160 5306 4212 5312
rect 4804 5364 4856 5370
rect 4804 5306 4856 5312
rect 5264 5296 5316 5302
rect 5264 5238 5316 5244
rect 4804 5160 4856 5166
rect 3514 5128 3570 5137
rect 4804 5102 4856 5108
rect 3514 5063 3570 5072
rect 4620 5024 4672 5030
rect 4620 4966 4672 4972
rect 3976 4684 4028 4690
rect 3976 4626 4028 4632
rect 3884 4616 3936 4622
rect 3884 4558 3936 4564
rect 3896 4282 3924 4558
rect 3884 4276 3936 4282
rect 3884 4218 3936 4224
rect 3056 4140 3108 4146
rect 3056 4082 3108 4088
rect 3988 3942 4016 4626
rect 4252 4072 4304 4078
rect 4252 4014 4304 4020
rect 3976 3936 4028 3942
rect 3976 3878 4028 3884
rect 4160 3936 4212 3942
rect 4160 3878 4212 3884
rect 3988 3670 4016 3878
rect 3976 3664 4028 3670
rect 3976 3606 4028 3612
rect 4172 1329 4200 3878
rect 4264 3602 4292 4014
rect 4632 4010 4660 4966
rect 4712 4072 4764 4078
rect 4712 4014 4764 4020
rect 4620 4004 4672 4010
rect 4620 3946 4672 3952
rect 4724 3942 4752 4014
rect 4712 3936 4764 3942
rect 4712 3878 4764 3884
rect 4816 3670 4844 5102
rect 5276 4826 5304 5238
rect 5264 4820 5316 4826
rect 5264 4762 5316 4768
rect 5276 4554 5304 4762
rect 5368 4690 5396 6870
rect 5460 6662 5488 7278
rect 5736 7002 5764 11630
rect 5920 7954 5948 15098
rect 6012 14890 6040 15506
rect 6000 14884 6052 14890
rect 6000 14826 6052 14832
rect 6104 13814 6132 17292
rect 7208 16794 7236 17682
rect 7484 17610 7512 18022
rect 7748 17808 7800 17814
rect 7748 17750 7800 17756
rect 7472 17604 7524 17610
rect 7472 17546 7524 17552
rect 7760 16998 7788 17750
rect 7944 17542 7972 18022
rect 7932 17536 7984 17542
rect 7932 17478 7984 17484
rect 7944 17066 7972 17478
rect 8312 17338 8340 18090
rect 8404 17882 8432 20198
rect 8956 20156 9252 20176
rect 9012 20154 9036 20156
rect 9092 20154 9116 20156
rect 9172 20154 9196 20156
rect 9034 20102 9036 20154
rect 9098 20102 9110 20154
rect 9172 20102 9174 20154
rect 9012 20100 9036 20102
rect 9092 20100 9116 20102
rect 9172 20100 9196 20102
rect 8956 20080 9252 20100
rect 10232 19916 10284 19922
rect 10232 19858 10284 19864
rect 10244 19718 10272 19858
rect 10232 19712 10284 19718
rect 10232 19654 10284 19660
rect 10244 19242 10272 19654
rect 10232 19236 10284 19242
rect 10232 19178 10284 19184
rect 10508 19168 10560 19174
rect 10508 19110 10560 19116
rect 8956 19068 9252 19088
rect 9012 19066 9036 19068
rect 9092 19066 9116 19068
rect 9172 19066 9196 19068
rect 9034 19014 9036 19066
rect 9098 19014 9110 19066
rect 9172 19014 9174 19066
rect 9012 19012 9036 19014
rect 9092 19012 9116 19014
rect 9172 19012 9196 19014
rect 8956 18992 9252 19012
rect 10520 18970 10548 19110
rect 10508 18964 10560 18970
rect 10508 18906 10560 18912
rect 11520 18964 11572 18970
rect 11520 18906 11572 18912
rect 9772 18896 9824 18902
rect 9772 18838 9824 18844
rect 9680 18760 9732 18766
rect 9680 18702 9732 18708
rect 9692 18290 9720 18702
rect 9784 18426 9812 18838
rect 11532 18426 11560 18906
rect 11796 18760 11848 18766
rect 11796 18702 11848 18708
rect 9772 18420 9824 18426
rect 9772 18362 9824 18368
rect 11520 18420 11572 18426
rect 11520 18362 11572 18368
rect 10876 18352 10928 18358
rect 10876 18294 10928 18300
rect 8576 18284 8628 18290
rect 8576 18226 8628 18232
rect 9680 18284 9732 18290
rect 9680 18226 9732 18232
rect 8392 17876 8444 17882
rect 8392 17818 8444 17824
rect 8300 17332 8352 17338
rect 8300 17274 8352 17280
rect 7932 17060 7984 17066
rect 7932 17002 7984 17008
rect 8116 17060 8168 17066
rect 8116 17002 8168 17008
rect 7748 16992 7800 16998
rect 7748 16934 7800 16940
rect 7944 16794 7972 17002
rect 7196 16788 7248 16794
rect 7196 16730 7248 16736
rect 7932 16788 7984 16794
rect 7932 16730 7984 16736
rect 7932 16584 7984 16590
rect 7932 16526 7984 16532
rect 6920 16448 6972 16454
rect 6920 16390 6972 16396
rect 6932 15978 6960 16390
rect 7012 16244 7064 16250
rect 7012 16186 7064 16192
rect 7024 15978 7052 16186
rect 6920 15972 6972 15978
rect 6920 15914 6972 15920
rect 7012 15972 7064 15978
rect 7012 15914 7064 15920
rect 6932 15706 6960 15914
rect 6920 15700 6972 15706
rect 6920 15642 6972 15648
rect 6184 15564 6236 15570
rect 6184 15506 6236 15512
rect 6196 15026 6224 15506
rect 6460 15496 6512 15502
rect 6460 15438 6512 15444
rect 7840 15496 7892 15502
rect 7840 15438 7892 15444
rect 6184 15020 6236 15026
rect 6184 14962 6236 14968
rect 6368 14272 6420 14278
rect 6368 14214 6420 14220
rect 6104 13786 6224 13814
rect 6196 13394 6224 13786
rect 6276 13728 6328 13734
rect 6276 13670 6328 13676
rect 6184 13388 6236 13394
rect 6184 13330 6236 13336
rect 6196 12646 6224 13330
rect 6288 13326 6316 13670
rect 6380 13530 6408 14214
rect 6472 13938 6500 15438
rect 7656 15360 7708 15366
rect 7656 15302 7708 15308
rect 7668 14958 7696 15302
rect 7852 15026 7880 15438
rect 7944 15434 7972 16526
rect 8128 16114 8156 17002
rect 8208 16720 8260 16726
rect 8208 16662 8260 16668
rect 8116 16108 8168 16114
rect 8116 16050 8168 16056
rect 8220 15978 8248 16662
rect 8208 15972 8260 15978
rect 8208 15914 8260 15920
rect 7932 15428 7984 15434
rect 7932 15370 7984 15376
rect 7840 15020 7892 15026
rect 7840 14962 7892 14968
rect 7656 14952 7708 14958
rect 7656 14894 7708 14900
rect 7012 14544 7064 14550
rect 7012 14486 7064 14492
rect 6460 13932 6512 13938
rect 6460 13874 6512 13880
rect 6472 13530 6500 13874
rect 6368 13524 6420 13530
rect 6368 13466 6420 13472
rect 6460 13524 6512 13530
rect 6460 13466 6512 13472
rect 7024 13462 7052 14486
rect 7472 14340 7524 14346
rect 7472 14282 7524 14288
rect 7012 13456 7064 13462
rect 7012 13398 7064 13404
rect 6276 13320 6328 13326
rect 6276 13262 6328 13268
rect 7288 13320 7340 13326
rect 7288 13262 7340 13268
rect 6184 12640 6236 12646
rect 6184 12582 6236 12588
rect 6000 12300 6052 12306
rect 6000 12242 6052 12248
rect 6012 11830 6040 12242
rect 6000 11824 6052 11830
rect 6000 11766 6052 11772
rect 6000 11212 6052 11218
rect 6000 11154 6052 11160
rect 6012 10470 6040 11154
rect 6000 10464 6052 10470
rect 6000 10406 6052 10412
rect 6012 8838 6040 10406
rect 6000 8832 6052 8838
rect 6000 8774 6052 8780
rect 5908 7948 5960 7954
rect 5908 7890 5960 7896
rect 5908 7744 5960 7750
rect 5908 7686 5960 7692
rect 5920 7410 5948 7686
rect 5908 7404 5960 7410
rect 5908 7346 5960 7352
rect 5724 6996 5776 7002
rect 5724 6938 5776 6944
rect 5540 6860 5592 6866
rect 5540 6802 5592 6808
rect 5908 6860 5960 6866
rect 5908 6802 5960 6808
rect 5448 6656 5500 6662
rect 5448 6598 5500 6604
rect 5552 6254 5580 6802
rect 5724 6656 5776 6662
rect 5724 6598 5776 6604
rect 5540 6248 5592 6254
rect 5540 6190 5592 6196
rect 5552 6118 5580 6190
rect 5540 6112 5592 6118
rect 5540 6054 5592 6060
rect 5552 4690 5580 6054
rect 5632 5568 5684 5574
rect 5632 5510 5684 5516
rect 5644 5166 5672 5510
rect 5632 5160 5684 5166
rect 5632 5102 5684 5108
rect 5644 4690 5672 5102
rect 5356 4684 5408 4690
rect 5356 4626 5408 4632
rect 5540 4684 5592 4690
rect 5540 4626 5592 4632
rect 5632 4684 5684 4690
rect 5632 4626 5684 4632
rect 5264 4548 5316 4554
rect 5264 4490 5316 4496
rect 5448 4548 5500 4554
rect 5448 4490 5500 4496
rect 4956 4380 5252 4400
rect 5012 4378 5036 4380
rect 5092 4378 5116 4380
rect 5172 4378 5196 4380
rect 5034 4326 5036 4378
rect 5098 4326 5110 4378
rect 5172 4326 5174 4378
rect 5012 4324 5036 4326
rect 5092 4324 5116 4326
rect 5172 4324 5196 4326
rect 4956 4304 5252 4324
rect 5172 4208 5224 4214
rect 5172 4150 5224 4156
rect 5184 3738 5212 4150
rect 5460 4010 5488 4490
rect 5448 4004 5500 4010
rect 5448 3946 5500 3952
rect 5172 3732 5224 3738
rect 5224 3692 5396 3720
rect 5172 3674 5224 3680
rect 4804 3664 4856 3670
rect 4804 3606 4856 3612
rect 4252 3596 4304 3602
rect 4252 3538 4304 3544
rect 4264 2854 4292 3538
rect 4956 3292 5252 3312
rect 5012 3290 5036 3292
rect 5092 3290 5116 3292
rect 5172 3290 5196 3292
rect 5034 3238 5036 3290
rect 5098 3238 5110 3290
rect 5172 3238 5174 3290
rect 5012 3236 5036 3238
rect 5092 3236 5116 3238
rect 5172 3236 5196 3238
rect 4956 3216 5252 3236
rect 5368 3194 5396 3692
rect 5356 3188 5408 3194
rect 5356 3130 5408 3136
rect 5356 2984 5408 2990
rect 5460 2972 5488 3946
rect 5552 3942 5580 4626
rect 5540 3936 5592 3942
rect 5540 3878 5592 3884
rect 5552 3126 5580 3878
rect 5644 3738 5672 4626
rect 5736 4622 5764 6598
rect 5920 6118 5948 6802
rect 6012 6798 6040 8774
rect 6196 8566 6224 12582
rect 6288 12442 6316 13262
rect 6460 13184 6512 13190
rect 6460 13126 6512 13132
rect 6472 12850 6500 13126
rect 6460 12844 6512 12850
rect 6460 12786 6512 12792
rect 7012 12708 7064 12714
rect 7012 12650 7064 12656
rect 7024 12594 7052 12650
rect 7196 12640 7248 12646
rect 7024 12588 7196 12594
rect 7024 12582 7248 12588
rect 7024 12566 7236 12582
rect 6276 12436 6328 12442
rect 6276 12378 6328 12384
rect 7208 12374 7236 12566
rect 7196 12368 7248 12374
rect 7196 12310 7248 12316
rect 6276 12232 6328 12238
rect 6276 12174 6328 12180
rect 6288 11354 6316 12174
rect 6552 12096 6604 12102
rect 6552 12038 6604 12044
rect 6564 11762 6592 12038
rect 7208 11898 7236 12310
rect 7300 12238 7328 13262
rect 7484 12918 7512 14282
rect 7668 13394 7696 14894
rect 7852 14618 7880 14962
rect 7944 14618 7972 15370
rect 8208 15088 8260 15094
rect 8208 15030 8260 15036
rect 7840 14612 7892 14618
rect 7840 14554 7892 14560
rect 7932 14612 7984 14618
rect 7932 14554 7984 14560
rect 7840 13728 7892 13734
rect 7840 13670 7892 13676
rect 7852 13462 7880 13670
rect 7840 13456 7892 13462
rect 7840 13398 7892 13404
rect 7656 13388 7708 13394
rect 7656 13330 7708 13336
rect 7472 12912 7524 12918
rect 7472 12854 7524 12860
rect 7288 12232 7340 12238
rect 7288 12174 7340 12180
rect 7196 11892 7248 11898
rect 7196 11834 7248 11840
rect 6552 11756 6604 11762
rect 6552 11698 6604 11704
rect 7208 11354 7236 11834
rect 6276 11348 6328 11354
rect 6276 11290 6328 11296
rect 7196 11348 7248 11354
rect 7196 11290 7248 11296
rect 7668 11286 7696 13330
rect 7852 12442 7880 13398
rect 7932 12844 7984 12850
rect 7932 12786 7984 12792
rect 7944 12442 7972 12786
rect 7840 12436 7892 12442
rect 7840 12378 7892 12384
rect 7932 12436 7984 12442
rect 7932 12378 7984 12384
rect 8116 11552 8168 11558
rect 8116 11494 8168 11500
rect 8128 11354 8156 11494
rect 8116 11348 8168 11354
rect 8116 11290 8168 11296
rect 7656 11280 7708 11286
rect 7656 11222 7708 11228
rect 6828 11212 6880 11218
rect 6828 11154 6880 11160
rect 8116 11212 8168 11218
rect 8116 11154 8168 11160
rect 6840 10742 6868 11154
rect 6920 11144 6972 11150
rect 6920 11086 6972 11092
rect 6828 10736 6880 10742
rect 6828 10678 6880 10684
rect 6932 10130 6960 11086
rect 7748 11008 7800 11014
rect 7748 10950 7800 10956
rect 7932 11008 7984 11014
rect 7932 10950 7984 10956
rect 7472 10668 7524 10674
rect 7472 10610 7524 10616
rect 7196 10532 7248 10538
rect 7196 10474 7248 10480
rect 7208 10198 7236 10474
rect 7104 10192 7156 10198
rect 7104 10134 7156 10140
rect 7196 10192 7248 10198
rect 7196 10134 7248 10140
rect 6920 10124 6972 10130
rect 6920 10066 6972 10072
rect 6932 9178 6960 10066
rect 7116 9654 7144 10134
rect 7104 9648 7156 9654
rect 7024 9608 7104 9636
rect 6920 9172 6972 9178
rect 6920 9114 6972 9120
rect 6184 8560 6236 8566
rect 6184 8502 6236 8508
rect 6552 8560 6604 8566
rect 6552 8502 6604 8508
rect 6000 6792 6052 6798
rect 6000 6734 6052 6740
rect 6092 6724 6144 6730
rect 6092 6666 6144 6672
rect 6104 6118 6132 6666
rect 5908 6112 5960 6118
rect 5908 6054 5960 6060
rect 6092 6112 6144 6118
rect 6092 6054 6144 6060
rect 5814 5128 5870 5137
rect 5920 5098 5948 6054
rect 6104 5778 6132 6054
rect 6000 5772 6052 5778
rect 6000 5714 6052 5720
rect 6092 5772 6144 5778
rect 6092 5714 6144 5720
rect 6012 5234 6040 5714
rect 6104 5370 6132 5714
rect 6092 5364 6144 5370
rect 6092 5306 6144 5312
rect 6000 5228 6052 5234
rect 6000 5170 6052 5176
rect 5814 5063 5870 5072
rect 5908 5092 5960 5098
rect 5828 5030 5856 5063
rect 5908 5034 5960 5040
rect 5816 5024 5868 5030
rect 5816 4966 5868 4972
rect 6012 4758 6040 5170
rect 6000 4752 6052 4758
rect 6000 4694 6052 4700
rect 5724 4616 5776 4622
rect 5724 4558 5776 4564
rect 5632 3732 5684 3738
rect 5632 3674 5684 3680
rect 5816 3596 5868 3602
rect 5816 3538 5868 3544
rect 5828 3194 5856 3538
rect 5816 3188 5868 3194
rect 5816 3130 5868 3136
rect 5540 3120 5592 3126
rect 5540 3062 5592 3068
rect 5408 2944 5488 2972
rect 5356 2926 5408 2932
rect 4252 2848 4304 2854
rect 4252 2790 4304 2796
rect 4158 1320 4214 1329
rect 4158 1255 4214 1264
rect 2778 54 2912 82
rect 4264 82 4292 2790
rect 4956 2204 5252 2224
rect 5012 2202 5036 2204
rect 5092 2202 5116 2204
rect 5172 2202 5196 2204
rect 5034 2150 5036 2202
rect 5098 2150 5110 2202
rect 5172 2150 5174 2202
rect 5012 2148 5036 2150
rect 5092 2148 5116 2150
rect 5172 2148 5196 2150
rect 4956 2128 5252 2148
rect 4618 82 4674 480
rect 5368 241 5396 2926
rect 6564 2650 6592 8502
rect 7024 8022 7052 9608
rect 7104 9590 7156 9596
rect 7380 9104 7432 9110
rect 7380 9046 7432 9052
rect 7104 8968 7156 8974
rect 7104 8910 7156 8916
rect 7116 8634 7144 8910
rect 7104 8628 7156 8634
rect 7104 8570 7156 8576
rect 7392 8362 7420 9046
rect 7484 8974 7512 10610
rect 7656 10532 7708 10538
rect 7760 10520 7788 10950
rect 7708 10492 7788 10520
rect 7656 10474 7708 10480
rect 7760 10266 7788 10492
rect 7748 10260 7800 10266
rect 7748 10202 7800 10208
rect 7760 9450 7788 10202
rect 7840 9580 7892 9586
rect 7944 9568 7972 10950
rect 8128 10810 8156 11154
rect 8116 10804 8168 10810
rect 8116 10746 8168 10752
rect 8024 9716 8076 9722
rect 8024 9658 8076 9664
rect 7892 9540 7972 9568
rect 7840 9522 7892 9528
rect 7748 9444 7800 9450
rect 7748 9386 7800 9392
rect 7944 9178 7972 9540
rect 8036 9450 8064 9658
rect 8024 9444 8076 9450
rect 8024 9386 8076 9392
rect 7932 9172 7984 9178
rect 7932 9114 7984 9120
rect 7472 8968 7524 8974
rect 7472 8910 7524 8916
rect 8036 8498 8064 9386
rect 8024 8492 8076 8498
rect 8024 8434 8076 8440
rect 7380 8356 7432 8362
rect 7380 8298 7432 8304
rect 7564 8356 7616 8362
rect 7564 8298 7616 8304
rect 7392 8090 7420 8298
rect 7576 8090 7604 8298
rect 7380 8084 7432 8090
rect 7380 8026 7432 8032
rect 7564 8084 7616 8090
rect 7564 8026 7616 8032
rect 7012 8016 7064 8022
rect 6734 7984 6790 7993
rect 7012 7958 7064 7964
rect 6734 7919 6790 7928
rect 6748 5778 6776 7919
rect 7024 7546 7052 7958
rect 8024 7948 8076 7954
rect 8024 7890 8076 7896
rect 7012 7540 7064 7546
rect 7012 7482 7064 7488
rect 7472 7336 7524 7342
rect 7472 7278 7524 7284
rect 7196 7268 7248 7274
rect 7196 7210 7248 7216
rect 7208 6730 7236 7210
rect 7196 6724 7248 6730
rect 7196 6666 7248 6672
rect 7012 6656 7064 6662
rect 7012 6598 7064 6604
rect 6736 5772 6788 5778
rect 6736 5714 6788 5720
rect 7024 5574 7052 6598
rect 7484 6118 7512 7278
rect 7656 6860 7708 6866
rect 7656 6802 7708 6808
rect 7668 6254 7696 6802
rect 7932 6792 7984 6798
rect 7932 6734 7984 6740
rect 7748 6724 7800 6730
rect 7748 6666 7800 6672
rect 7656 6248 7708 6254
rect 7656 6190 7708 6196
rect 7472 6112 7524 6118
rect 7472 6054 7524 6060
rect 7484 5574 7512 6054
rect 7564 5772 7616 5778
rect 7564 5714 7616 5720
rect 7012 5568 7064 5574
rect 7012 5510 7064 5516
rect 7472 5568 7524 5574
rect 7472 5510 7524 5516
rect 7024 5370 7052 5510
rect 7012 5364 7064 5370
rect 7012 5306 7064 5312
rect 6644 4548 6696 4554
rect 6644 4490 6696 4496
rect 6656 4282 6684 4490
rect 6644 4276 6696 4282
rect 6644 4218 6696 4224
rect 7024 4154 7052 5306
rect 7196 5024 7248 5030
rect 7196 4966 7248 4972
rect 7208 4690 7236 4966
rect 7104 4684 7156 4690
rect 7104 4626 7156 4632
rect 7196 4684 7248 4690
rect 7196 4626 7248 4632
rect 6932 4126 7052 4154
rect 6644 3596 6696 3602
rect 6644 3538 6696 3544
rect 6656 3194 6684 3538
rect 6644 3188 6696 3194
rect 6644 3130 6696 3136
rect 6552 2644 6604 2650
rect 6552 2586 6604 2592
rect 6932 2582 6960 4126
rect 7116 3738 7144 4626
rect 7208 4282 7236 4626
rect 7196 4276 7248 4282
rect 7196 4218 7248 4224
rect 7104 3732 7156 3738
rect 7104 3674 7156 3680
rect 7484 3466 7512 5510
rect 7576 5098 7604 5714
rect 7564 5092 7616 5098
rect 7564 5034 7616 5040
rect 7576 3602 7604 5034
rect 7760 4468 7788 6666
rect 7840 6656 7892 6662
rect 7840 6598 7892 6604
rect 7852 6390 7880 6598
rect 7840 6384 7892 6390
rect 7840 6326 7892 6332
rect 7944 6322 7972 6734
rect 8036 6458 8064 7890
rect 8024 6452 8076 6458
rect 8024 6394 8076 6400
rect 7932 6316 7984 6322
rect 7932 6258 7984 6264
rect 8024 6180 8076 6186
rect 8024 6122 8076 6128
rect 8036 5914 8064 6122
rect 8024 5908 8076 5914
rect 8024 5850 8076 5856
rect 8036 4690 8064 5850
rect 8116 5772 8168 5778
rect 8116 5714 8168 5720
rect 8128 5030 8156 5714
rect 8116 5024 8168 5030
rect 8116 4966 8168 4972
rect 8128 4826 8156 4966
rect 8116 4820 8168 4826
rect 8116 4762 8168 4768
rect 8024 4684 8076 4690
rect 8024 4626 8076 4632
rect 7840 4480 7892 4486
rect 7760 4440 7840 4468
rect 7840 4422 7892 4428
rect 7852 4282 7880 4422
rect 7840 4276 7892 4282
rect 7840 4218 7892 4224
rect 8036 4078 8064 4626
rect 7932 4072 7984 4078
rect 7932 4014 7984 4020
rect 8024 4072 8076 4078
rect 8024 4014 8076 4020
rect 7564 3596 7616 3602
rect 7564 3538 7616 3544
rect 7472 3460 7524 3466
rect 7472 3402 7524 3408
rect 7944 2990 7972 4014
rect 8128 3602 8156 4762
rect 8116 3596 8168 3602
rect 8116 3538 8168 3544
rect 7932 2984 7984 2990
rect 8128 2961 8156 3538
rect 7932 2926 7984 2932
rect 8114 2952 8170 2961
rect 7944 2650 7972 2926
rect 8114 2887 8116 2896
rect 8168 2887 8170 2896
rect 8116 2858 8168 2864
rect 8128 2827 8156 2858
rect 7932 2644 7984 2650
rect 7932 2586 7984 2592
rect 6920 2576 6972 2582
rect 6920 2518 6972 2524
rect 8220 2514 8248 15030
rect 8404 12424 8432 17818
rect 8484 16992 8536 16998
rect 8484 16934 8536 16940
rect 8496 15638 8524 16934
rect 8588 16590 8616 18226
rect 9864 18216 9916 18222
rect 9864 18158 9916 18164
rect 8956 17980 9252 18000
rect 9012 17978 9036 17980
rect 9092 17978 9116 17980
rect 9172 17978 9196 17980
rect 9034 17926 9036 17978
rect 9098 17926 9110 17978
rect 9172 17926 9174 17978
rect 9012 17924 9036 17926
rect 9092 17924 9116 17926
rect 9172 17924 9196 17926
rect 8956 17904 9252 17924
rect 9876 17649 9904 18158
rect 10888 17746 10916 18294
rect 11060 18080 11112 18086
rect 11060 18022 11112 18028
rect 11072 17746 11100 18022
rect 10876 17740 10928 17746
rect 10876 17682 10928 17688
rect 11060 17740 11112 17746
rect 11060 17682 11112 17688
rect 9862 17640 9918 17649
rect 9862 17575 9918 17584
rect 9876 17542 9904 17575
rect 8852 17536 8904 17542
rect 8852 17478 8904 17484
rect 9864 17536 9916 17542
rect 9864 17478 9916 17484
rect 10784 17536 10836 17542
rect 10784 17478 10836 17484
rect 8576 16584 8628 16590
rect 8576 16526 8628 16532
rect 8760 15972 8812 15978
rect 8760 15914 8812 15920
rect 8668 15904 8720 15910
rect 8588 15864 8668 15892
rect 8484 15632 8536 15638
rect 8484 15574 8536 15580
rect 8496 14822 8524 15574
rect 8484 14816 8536 14822
rect 8484 14758 8536 14764
rect 8404 12396 8524 12424
rect 8392 12300 8444 12306
rect 8392 12242 8444 12248
rect 8404 11558 8432 12242
rect 8392 11552 8444 11558
rect 8392 11494 8444 11500
rect 8404 9518 8432 11494
rect 8496 10305 8524 12396
rect 8588 11830 8616 15864
rect 8668 15846 8720 15852
rect 8772 15706 8800 15914
rect 8760 15700 8812 15706
rect 8760 15642 8812 15648
rect 8760 14476 8812 14482
rect 8680 14436 8760 14464
rect 8680 13734 8708 14436
rect 8760 14418 8812 14424
rect 8864 13814 8892 17478
rect 9772 17264 9824 17270
rect 9772 17206 9824 17212
rect 9496 17128 9548 17134
rect 9496 17070 9548 17076
rect 8956 16892 9252 16912
rect 9012 16890 9036 16892
rect 9092 16890 9116 16892
rect 9172 16890 9196 16892
rect 9034 16838 9036 16890
rect 9098 16838 9110 16890
rect 9172 16838 9174 16890
rect 9012 16836 9036 16838
rect 9092 16836 9116 16838
rect 9172 16836 9196 16838
rect 8956 16816 9252 16836
rect 9312 16448 9364 16454
rect 9312 16390 9364 16396
rect 9324 16114 9352 16390
rect 9312 16108 9364 16114
rect 9312 16050 9364 16056
rect 8956 15804 9252 15824
rect 9012 15802 9036 15804
rect 9092 15802 9116 15804
rect 9172 15802 9196 15804
rect 9034 15750 9036 15802
rect 9098 15750 9110 15802
rect 9172 15750 9174 15802
rect 9012 15748 9036 15750
rect 9092 15748 9116 15750
rect 9172 15748 9196 15750
rect 8956 15728 9252 15748
rect 9324 15706 9352 16050
rect 9312 15700 9364 15706
rect 9312 15642 9364 15648
rect 9508 15094 9536 17070
rect 9588 16652 9640 16658
rect 9588 16594 9640 16600
rect 9600 16114 9628 16594
rect 9588 16108 9640 16114
rect 9588 16050 9640 16056
rect 9600 15910 9628 16050
rect 9784 15978 9812 17206
rect 10796 17134 10824 17478
rect 10784 17128 10836 17134
rect 10784 17070 10836 17076
rect 10416 17060 10468 17066
rect 10416 17002 10468 17008
rect 10232 16040 10284 16046
rect 10232 15982 10284 15988
rect 9772 15972 9824 15978
rect 9772 15914 9824 15920
rect 9588 15904 9640 15910
rect 9588 15846 9640 15852
rect 10244 15706 10272 15982
rect 10232 15700 10284 15706
rect 10232 15642 10284 15648
rect 10428 15570 10456 17002
rect 10692 16788 10744 16794
rect 10692 16730 10744 16736
rect 10416 15564 10468 15570
rect 10416 15506 10468 15512
rect 9772 15156 9824 15162
rect 9772 15098 9824 15104
rect 9496 15088 9548 15094
rect 9496 15030 9548 15036
rect 9784 14958 9812 15098
rect 10428 14958 10456 15506
rect 10600 15496 10652 15502
rect 10600 15438 10652 15444
rect 9496 14952 9548 14958
rect 9496 14894 9548 14900
rect 9772 14952 9824 14958
rect 9772 14894 9824 14900
rect 10416 14952 10468 14958
rect 10416 14894 10468 14900
rect 8956 14716 9252 14736
rect 9012 14714 9036 14716
rect 9092 14714 9116 14716
rect 9172 14714 9196 14716
rect 9034 14662 9036 14714
rect 9098 14662 9110 14714
rect 9172 14662 9174 14714
rect 9012 14660 9036 14662
rect 9092 14660 9116 14662
rect 9172 14660 9196 14662
rect 8956 14640 9252 14660
rect 8772 13786 8892 13814
rect 8668 13728 8720 13734
rect 8668 13670 8720 13676
rect 8668 13184 8720 13190
rect 8772 13172 8800 13786
rect 8956 13628 9252 13648
rect 9012 13626 9036 13628
rect 9092 13626 9116 13628
rect 9172 13626 9196 13628
rect 9034 13574 9036 13626
rect 9098 13574 9110 13626
rect 9172 13574 9174 13626
rect 9012 13572 9036 13574
rect 9092 13572 9116 13574
rect 9172 13572 9196 13574
rect 8956 13552 9252 13572
rect 8720 13144 8800 13172
rect 8668 13126 8720 13132
rect 8680 12782 8708 13126
rect 8668 12776 8720 12782
rect 8668 12718 8720 12724
rect 8576 11824 8628 11830
rect 8576 11766 8628 11772
rect 8588 11218 8616 11766
rect 8576 11212 8628 11218
rect 8576 11154 8628 11160
rect 8482 10296 8538 10305
rect 8482 10231 8538 10240
rect 8496 10130 8524 10231
rect 8484 10124 8536 10130
rect 8484 10066 8536 10072
rect 8392 9512 8444 9518
rect 8392 9454 8444 9460
rect 8680 9353 8708 12718
rect 8852 12640 8904 12646
rect 8852 12582 8904 12588
rect 8864 12442 8892 12582
rect 8956 12540 9252 12560
rect 9012 12538 9036 12540
rect 9092 12538 9116 12540
rect 9172 12538 9196 12540
rect 9034 12486 9036 12538
rect 9098 12486 9110 12538
rect 9172 12486 9174 12538
rect 9012 12484 9036 12486
rect 9092 12484 9116 12486
rect 9172 12484 9196 12486
rect 8956 12464 9252 12484
rect 8852 12436 8904 12442
rect 8852 12378 8904 12384
rect 8864 11762 8892 12378
rect 8852 11756 8904 11762
rect 8852 11698 8904 11704
rect 8956 11452 9252 11472
rect 9012 11450 9036 11452
rect 9092 11450 9116 11452
rect 9172 11450 9196 11452
rect 9034 11398 9036 11450
rect 9098 11398 9110 11450
rect 9172 11398 9174 11450
rect 9012 11396 9036 11398
rect 9092 11396 9116 11398
rect 9172 11396 9196 11398
rect 8956 11376 9252 11396
rect 9312 10600 9364 10606
rect 9508 10588 9536 14894
rect 9784 13394 9812 14894
rect 10232 14884 10284 14890
rect 10232 14826 10284 14832
rect 10244 14482 10272 14826
rect 10232 14476 10284 14482
rect 10232 14418 10284 14424
rect 10244 14074 10272 14418
rect 10612 14278 10640 15438
rect 10600 14272 10652 14278
rect 10600 14214 10652 14220
rect 10232 14068 10284 14074
rect 10232 14010 10284 14016
rect 10324 14068 10376 14074
rect 10324 14010 10376 14016
rect 10336 13938 10364 14010
rect 9956 13932 10008 13938
rect 9956 13874 10008 13880
rect 10324 13932 10376 13938
rect 10324 13874 10376 13880
rect 9968 13530 9996 13874
rect 10416 13864 10468 13870
rect 10416 13806 10468 13812
rect 10140 13728 10192 13734
rect 10140 13670 10192 13676
rect 9956 13524 10008 13530
rect 9956 13466 10008 13472
rect 9588 13388 9640 13394
rect 9772 13388 9824 13394
rect 9588 13330 9640 13336
rect 9692 13348 9772 13376
rect 9600 12986 9628 13330
rect 9588 12980 9640 12986
rect 9588 12922 9640 12928
rect 9692 12646 9720 13348
rect 9772 13330 9824 13336
rect 10152 12918 10180 13670
rect 10428 13462 10456 13806
rect 10416 13456 10468 13462
rect 10416 13398 10468 13404
rect 10140 12912 10192 12918
rect 10140 12854 10192 12860
rect 9680 12640 9732 12646
rect 9680 12582 9732 12588
rect 9588 12368 9640 12374
rect 9588 12310 9640 12316
rect 9600 11898 9628 12310
rect 9588 11892 9640 11898
rect 9588 11834 9640 11840
rect 9600 11354 9628 11834
rect 9588 11348 9640 11354
rect 9588 11290 9640 11296
rect 9364 10560 9536 10588
rect 9312 10542 9364 10548
rect 8956 10364 9252 10384
rect 9012 10362 9036 10364
rect 9092 10362 9116 10364
rect 9172 10362 9196 10364
rect 9034 10310 9036 10362
rect 9098 10310 9110 10362
rect 9172 10310 9174 10362
rect 9012 10308 9036 10310
rect 9092 10308 9116 10310
rect 9172 10308 9196 10310
rect 8956 10288 9252 10308
rect 8760 10192 8812 10198
rect 8760 10134 8812 10140
rect 8772 9586 8800 10134
rect 8852 10124 8904 10130
rect 8852 10066 8904 10072
rect 8760 9580 8812 9586
rect 8760 9522 8812 9528
rect 8760 9376 8812 9382
rect 8666 9344 8722 9353
rect 8864 9364 8892 10066
rect 9324 9926 9352 10542
rect 9312 9920 9364 9926
rect 9312 9862 9364 9868
rect 9404 9444 9456 9450
rect 9404 9386 9456 9392
rect 8812 9336 8892 9364
rect 9416 9353 9444 9386
rect 9402 9344 9458 9353
rect 8760 9318 8812 9324
rect 8666 9279 8722 9288
rect 8300 7948 8352 7954
rect 8300 7890 8352 7896
rect 8312 7342 8340 7890
rect 8300 7336 8352 7342
rect 8300 7278 8352 7284
rect 8300 6384 8352 6390
rect 8300 6326 8352 6332
rect 8312 6118 8340 6326
rect 8300 6112 8352 6118
rect 8300 6054 8352 6060
rect 8312 5574 8340 6054
rect 8300 5568 8352 5574
rect 8300 5510 8352 5516
rect 8312 2825 8340 5510
rect 8680 4622 8708 9279
rect 8772 8945 8800 9318
rect 8956 9276 9252 9296
rect 9402 9279 9458 9288
rect 9586 9344 9642 9353
rect 9586 9279 9642 9288
rect 9012 9274 9036 9276
rect 9092 9274 9116 9276
rect 9172 9274 9196 9276
rect 9034 9222 9036 9274
rect 9098 9222 9110 9274
rect 9172 9222 9174 9274
rect 9012 9220 9036 9222
rect 9092 9220 9116 9222
rect 9172 9220 9196 9222
rect 8956 9200 9252 9220
rect 8758 8936 8814 8945
rect 8758 8871 8814 8880
rect 8956 8188 9252 8208
rect 9012 8186 9036 8188
rect 9092 8186 9116 8188
rect 9172 8186 9196 8188
rect 9034 8134 9036 8186
rect 9098 8134 9110 8186
rect 9172 8134 9174 8186
rect 9012 8132 9036 8134
rect 9092 8132 9116 8134
rect 9172 8132 9196 8134
rect 8956 8112 9252 8132
rect 8852 7880 8904 7886
rect 8852 7822 8904 7828
rect 8864 7546 8892 7822
rect 9496 7744 9548 7750
rect 9496 7686 9548 7692
rect 9508 7546 9536 7686
rect 8852 7540 8904 7546
rect 8852 7482 8904 7488
rect 9496 7540 9548 7546
rect 9496 7482 9548 7488
rect 8956 7100 9252 7120
rect 9012 7098 9036 7100
rect 9092 7098 9116 7100
rect 9172 7098 9196 7100
rect 9034 7046 9036 7098
rect 9098 7046 9110 7098
rect 9172 7046 9174 7098
rect 9012 7044 9036 7046
rect 9092 7044 9116 7046
rect 9172 7044 9196 7046
rect 8956 7024 9252 7044
rect 9508 6798 9536 7482
rect 9496 6792 9548 6798
rect 9496 6734 9548 6740
rect 9128 6656 9180 6662
rect 9128 6598 9180 6604
rect 9140 6186 9168 6598
rect 9404 6384 9456 6390
rect 9324 6344 9404 6372
rect 9128 6180 9180 6186
rect 9128 6122 9180 6128
rect 8956 6012 9252 6032
rect 9012 6010 9036 6012
rect 9092 6010 9116 6012
rect 9172 6010 9196 6012
rect 9034 5958 9036 6010
rect 9098 5958 9110 6010
rect 9172 5958 9174 6010
rect 9012 5956 9036 5958
rect 9092 5956 9116 5958
rect 9172 5956 9196 5958
rect 8956 5936 9252 5956
rect 9324 5574 9352 6344
rect 9404 6326 9456 6332
rect 9508 5914 9536 6734
rect 9496 5908 9548 5914
rect 9496 5850 9548 5856
rect 9312 5568 9364 5574
rect 9312 5510 9364 5516
rect 9324 5370 9352 5510
rect 9312 5364 9364 5370
rect 9312 5306 9364 5312
rect 9508 5166 9536 5850
rect 9496 5160 9548 5166
rect 9496 5102 9548 5108
rect 8956 4924 9252 4944
rect 9012 4922 9036 4924
rect 9092 4922 9116 4924
rect 9172 4922 9196 4924
rect 9034 4870 9036 4922
rect 9098 4870 9110 4922
rect 9172 4870 9174 4922
rect 9012 4868 9036 4870
rect 9092 4868 9116 4870
rect 9172 4868 9196 4870
rect 8956 4848 9252 4868
rect 9508 4826 9536 5102
rect 9496 4820 9548 4826
rect 9496 4762 9548 4768
rect 8668 4616 8720 4622
rect 8668 4558 8720 4564
rect 9600 4154 9628 9279
rect 9692 6458 9720 12582
rect 9772 12232 9824 12238
rect 9772 12174 9824 12180
rect 9784 11898 9812 12174
rect 9772 11892 9824 11898
rect 9772 11834 9824 11840
rect 9784 11354 9812 11834
rect 9954 11792 10010 11801
rect 9954 11727 10010 11736
rect 9772 11348 9824 11354
rect 9772 11290 9824 11296
rect 9772 10192 9824 10198
rect 9772 10134 9824 10140
rect 9784 9926 9812 10134
rect 9772 9920 9824 9926
rect 9772 9862 9824 9868
rect 9784 9450 9812 9862
rect 9968 9625 9996 11727
rect 10048 10532 10100 10538
rect 10048 10474 10100 10480
rect 10060 10130 10088 10474
rect 10048 10124 10100 10130
rect 10048 10066 10100 10072
rect 9954 9616 10010 9625
rect 9954 9551 10010 9560
rect 9956 9512 10008 9518
rect 9956 9454 10008 9460
rect 9772 9444 9824 9450
rect 9772 9386 9824 9392
rect 9968 9178 9996 9454
rect 9956 9172 10008 9178
rect 9956 9114 10008 9120
rect 10060 9110 10088 10066
rect 10048 9104 10100 9110
rect 10048 9046 10100 9052
rect 10152 8956 10180 12854
rect 10612 12782 10640 14214
rect 10600 12776 10652 12782
rect 10600 12718 10652 12724
rect 10232 12708 10284 12714
rect 10232 12650 10284 12656
rect 10244 11898 10272 12650
rect 10612 12442 10640 12718
rect 10600 12436 10652 12442
rect 10600 12378 10652 12384
rect 10416 12300 10468 12306
rect 10416 12242 10468 12248
rect 10428 12209 10456 12242
rect 10414 12200 10470 12209
rect 10414 12135 10470 12144
rect 10232 11892 10284 11898
rect 10232 11834 10284 11840
rect 10244 10810 10272 11834
rect 10428 11830 10456 12135
rect 10416 11824 10468 11830
rect 10416 11766 10468 11772
rect 10508 11688 10560 11694
rect 10704 11676 10732 16730
rect 10796 16046 10824 17070
rect 10888 16794 10916 17682
rect 11072 17134 11100 17682
rect 11060 17128 11112 17134
rect 11060 17070 11112 17076
rect 11152 17060 11204 17066
rect 11152 17002 11204 17008
rect 10876 16788 10928 16794
rect 10876 16730 10928 16736
rect 11164 16590 11192 17002
rect 11532 16726 11560 18362
rect 11808 18086 11836 18702
rect 11796 18080 11848 18086
rect 11796 18022 11848 18028
rect 11808 17814 11836 18022
rect 11796 17808 11848 17814
rect 11796 17750 11848 17756
rect 11992 17338 12020 20198
rect 12956 19612 13252 19632
rect 13012 19610 13036 19612
rect 13092 19610 13116 19612
rect 13172 19610 13196 19612
rect 13034 19558 13036 19610
rect 13098 19558 13110 19610
rect 13172 19558 13174 19610
rect 13012 19556 13036 19558
rect 13092 19556 13116 19558
rect 13172 19556 13196 19558
rect 12956 19536 13252 19556
rect 12808 19236 12860 19242
rect 12808 19178 12860 19184
rect 12348 18624 12400 18630
rect 12348 18566 12400 18572
rect 12624 18624 12676 18630
rect 12624 18566 12676 18572
rect 12360 18426 12388 18566
rect 12348 18420 12400 18426
rect 12348 18362 12400 18368
rect 12360 18086 12388 18362
rect 12636 18290 12664 18566
rect 12820 18290 12848 19178
rect 12956 18524 13252 18544
rect 13012 18522 13036 18524
rect 13092 18522 13116 18524
rect 13172 18522 13196 18524
rect 13034 18470 13036 18522
rect 13098 18470 13110 18522
rect 13172 18470 13174 18522
rect 13012 18468 13036 18470
rect 13092 18468 13116 18470
rect 13172 18468 13196 18470
rect 12956 18448 13252 18468
rect 12624 18284 12676 18290
rect 12624 18226 12676 18232
rect 12808 18284 12860 18290
rect 12808 18226 12860 18232
rect 12348 18080 12400 18086
rect 12348 18022 12400 18028
rect 12256 17808 12308 17814
rect 12256 17750 12308 17756
rect 11980 17332 12032 17338
rect 11980 17274 12032 17280
rect 11796 16992 11848 16998
rect 11794 16960 11796 16969
rect 11848 16960 11850 16969
rect 11794 16895 11850 16904
rect 11520 16720 11572 16726
rect 11520 16662 11572 16668
rect 11152 16584 11204 16590
rect 11152 16526 11204 16532
rect 10968 16244 11020 16250
rect 10968 16186 11020 16192
rect 11428 16244 11480 16250
rect 11532 16232 11560 16662
rect 11808 16250 11836 16895
rect 11888 16516 11940 16522
rect 11888 16458 11940 16464
rect 11480 16204 11560 16232
rect 11796 16244 11848 16250
rect 11428 16186 11480 16192
rect 11796 16186 11848 16192
rect 10784 16040 10836 16046
rect 10784 15982 10836 15988
rect 10980 15910 11008 16186
rect 11796 16040 11848 16046
rect 11900 16028 11928 16458
rect 11848 16000 11928 16028
rect 11796 15982 11848 15988
rect 10968 15904 11020 15910
rect 10968 15846 11020 15852
rect 10980 14822 11008 15846
rect 11244 14952 11296 14958
rect 11244 14894 11296 14900
rect 10968 14816 11020 14822
rect 10968 14758 11020 14764
rect 10980 14550 11008 14758
rect 10968 14544 11020 14550
rect 10968 14486 11020 14492
rect 10980 14074 11008 14486
rect 10968 14068 11020 14074
rect 10968 14010 11020 14016
rect 11256 14006 11284 14894
rect 11888 14816 11940 14822
rect 11888 14758 11940 14764
rect 11900 14550 11928 14758
rect 11888 14544 11940 14550
rect 11888 14486 11940 14492
rect 11244 14000 11296 14006
rect 11244 13942 11296 13948
rect 11256 13841 11284 13942
rect 11242 13832 11298 13841
rect 11242 13767 11298 13776
rect 11336 13796 11388 13802
rect 11336 13738 11388 13744
rect 11348 13530 11376 13738
rect 11336 13524 11388 13530
rect 11336 13466 11388 13472
rect 11348 12714 11376 13466
rect 11888 13388 11940 13394
rect 11888 13330 11940 13336
rect 11900 13258 11928 13330
rect 11888 13252 11940 13258
rect 11888 13194 11940 13200
rect 11900 12918 11928 13194
rect 11888 12912 11940 12918
rect 11888 12854 11940 12860
rect 11244 12708 11296 12714
rect 11244 12650 11296 12656
rect 11336 12708 11388 12714
rect 11336 12650 11388 12656
rect 11256 12238 11284 12650
rect 11348 12374 11376 12650
rect 11336 12368 11388 12374
rect 11336 12310 11388 12316
rect 11244 12232 11296 12238
rect 11244 12174 11296 12180
rect 11256 11898 11284 12174
rect 11244 11892 11296 11898
rect 11244 11834 11296 11840
rect 10560 11648 10732 11676
rect 10508 11630 10560 11636
rect 10520 11014 10548 11630
rect 11152 11620 11204 11626
rect 11152 11562 11204 11568
rect 11164 11218 11192 11562
rect 11244 11552 11296 11558
rect 11244 11494 11296 11500
rect 11256 11268 11284 11494
rect 11348 11286 11376 12310
rect 11336 11280 11388 11286
rect 11256 11240 11336 11268
rect 11152 11212 11204 11218
rect 11152 11154 11204 11160
rect 10508 11008 10560 11014
rect 10508 10950 10560 10956
rect 10232 10804 10284 10810
rect 10232 10746 10284 10752
rect 10244 9042 10272 10746
rect 10232 9036 10284 9042
rect 10232 8978 10284 8984
rect 10060 8928 10180 8956
rect 9864 7948 9916 7954
rect 9864 7890 9916 7896
rect 9876 7274 9904 7890
rect 9864 7268 9916 7274
rect 9864 7210 9916 7216
rect 9680 6452 9732 6458
rect 9680 6394 9732 6400
rect 9956 6316 10008 6322
rect 9956 6258 10008 6264
rect 9772 6248 9824 6254
rect 9772 6190 9824 6196
rect 9784 5778 9812 6190
rect 9968 5778 9996 6258
rect 9772 5772 9824 5778
rect 9772 5714 9824 5720
rect 9956 5772 10008 5778
rect 9956 5714 10008 5720
rect 9784 5030 9812 5714
rect 9956 5296 10008 5302
rect 9956 5238 10008 5244
rect 9772 5024 9824 5030
rect 9772 4966 9824 4972
rect 9784 4690 9812 4966
rect 9772 4684 9824 4690
rect 9772 4626 9824 4632
rect 9416 4126 9628 4154
rect 9784 4154 9812 4626
rect 9784 4146 9904 4154
rect 9772 4140 9904 4146
rect 8392 4072 8444 4078
rect 8392 4014 8444 4020
rect 8760 4072 8812 4078
rect 8760 4014 8812 4020
rect 8404 3058 8432 4014
rect 8772 3738 8800 4014
rect 8852 3936 8904 3942
rect 8852 3878 8904 3884
rect 8760 3732 8812 3738
rect 8760 3674 8812 3680
rect 8864 3534 8892 3878
rect 8956 3836 9252 3856
rect 9012 3834 9036 3836
rect 9092 3834 9116 3836
rect 9172 3834 9196 3836
rect 9034 3782 9036 3834
rect 9098 3782 9110 3834
rect 9172 3782 9174 3834
rect 9012 3780 9036 3782
rect 9092 3780 9116 3782
rect 9172 3780 9196 3782
rect 8956 3760 9252 3780
rect 8852 3528 8904 3534
rect 8852 3470 8904 3476
rect 8864 3194 8892 3470
rect 8852 3188 8904 3194
rect 8852 3130 8904 3136
rect 8392 3052 8444 3058
rect 8392 2994 8444 3000
rect 8298 2816 8354 2825
rect 8298 2751 8354 2760
rect 8404 2650 8432 2994
rect 8956 2748 9252 2768
rect 9012 2746 9036 2748
rect 9092 2746 9116 2748
rect 9172 2746 9196 2748
rect 9034 2694 9036 2746
rect 9098 2694 9110 2746
rect 9172 2694 9174 2746
rect 9012 2692 9036 2694
rect 9092 2692 9116 2694
rect 9172 2692 9196 2694
rect 8956 2672 9252 2692
rect 8392 2644 8444 2650
rect 8392 2586 8444 2592
rect 8208 2508 8260 2514
rect 8208 2450 8260 2456
rect 9416 2446 9444 4126
rect 9824 4126 9904 4140
rect 9772 4082 9824 4088
rect 9772 2848 9824 2854
rect 9772 2790 9824 2796
rect 9784 2514 9812 2790
rect 9772 2508 9824 2514
rect 9772 2450 9824 2456
rect 6736 2440 6788 2446
rect 6736 2382 6788 2388
rect 9404 2440 9456 2446
rect 9404 2382 9456 2388
rect 5908 2304 5960 2310
rect 5908 2246 5960 2252
rect 5920 1329 5948 2246
rect 5906 1320 5962 1329
rect 5906 1255 5962 1264
rect 5354 232 5410 241
rect 5354 167 5410 176
rect 4264 54 4674 82
rect 938 0 994 54
rect 2778 0 2834 54
rect 4618 0 4674 54
rect 6458 82 6514 480
rect 6748 82 6776 2382
rect 9876 1737 9904 4126
rect 9968 3670 9996 5238
rect 9956 3664 10008 3670
rect 9956 3606 10008 3612
rect 9968 2854 9996 3606
rect 9956 2848 10008 2854
rect 9956 2790 10008 2796
rect 9968 2650 9996 2790
rect 9956 2644 10008 2650
rect 9956 2586 10008 2592
rect 9862 1728 9918 1737
rect 9862 1663 9918 1672
rect 8574 1592 8630 1601
rect 8574 1527 8630 1536
rect 6458 54 6776 82
rect 8298 82 8354 480
rect 8588 82 8616 1527
rect 8298 54 8616 82
rect 10060 82 10088 8928
rect 10244 8634 10272 8978
rect 10324 8832 10376 8838
rect 10324 8774 10376 8780
rect 10232 8628 10284 8634
rect 10232 8570 10284 8576
rect 10244 8022 10272 8570
rect 10336 8430 10364 8774
rect 10324 8424 10376 8430
rect 10324 8366 10376 8372
rect 10232 8016 10284 8022
rect 10232 7958 10284 7964
rect 10140 7744 10192 7750
rect 10140 7686 10192 7692
rect 10152 7478 10180 7686
rect 10140 7472 10192 7478
rect 10140 7414 10192 7420
rect 10152 6730 10180 7414
rect 10232 7404 10284 7410
rect 10232 7346 10284 7352
rect 10244 7206 10272 7346
rect 10232 7200 10284 7206
rect 10232 7142 10284 7148
rect 10244 6798 10272 7142
rect 10232 6792 10284 6798
rect 10232 6734 10284 6740
rect 10140 6724 10192 6730
rect 10140 6666 10192 6672
rect 10244 6322 10272 6734
rect 10232 6316 10284 6322
rect 10232 6258 10284 6264
rect 10336 5710 10364 8366
rect 10520 7993 10548 10950
rect 11164 10810 11192 11154
rect 11152 10804 11204 10810
rect 11152 10746 11204 10752
rect 11152 10464 11204 10470
rect 11256 10452 11284 11240
rect 11336 11222 11388 11228
rect 11992 10810 12020 17274
rect 12268 16998 12296 17750
rect 12636 17678 12664 18226
rect 12624 17672 12676 17678
rect 12624 17614 12676 17620
rect 12716 17536 12768 17542
rect 12716 17478 12768 17484
rect 12532 17196 12584 17202
rect 12532 17138 12584 17144
rect 12256 16992 12308 16998
rect 12256 16934 12308 16940
rect 12268 16794 12296 16934
rect 12256 16788 12308 16794
rect 12256 16730 12308 16736
rect 12544 16658 12572 17138
rect 12624 17060 12676 17066
rect 12624 17002 12676 17008
rect 12636 16969 12664 17002
rect 12622 16960 12678 16969
rect 12622 16895 12678 16904
rect 12728 16794 12756 17478
rect 12820 17202 12848 18226
rect 13176 18216 13228 18222
rect 13176 18158 13228 18164
rect 13188 17882 13216 18158
rect 13176 17876 13228 17882
rect 13176 17818 13228 17824
rect 13280 17746 13308 23582
rect 14922 23582 15056 23610
rect 14922 23520 14978 23582
rect 13268 17740 13320 17746
rect 13268 17682 13320 17688
rect 12956 17436 13252 17456
rect 13012 17434 13036 17436
rect 13092 17434 13116 17436
rect 13172 17434 13196 17436
rect 13034 17382 13036 17434
rect 13098 17382 13110 17434
rect 13172 17382 13174 17434
rect 13012 17380 13036 17382
rect 13092 17380 13116 17382
rect 13172 17380 13196 17382
rect 12956 17360 13252 17380
rect 13280 17270 13308 17682
rect 13360 17672 13412 17678
rect 13360 17614 13412 17620
rect 13372 17542 13400 17614
rect 13820 17604 13872 17610
rect 13820 17546 13872 17552
rect 13360 17536 13412 17542
rect 13360 17478 13412 17484
rect 13452 17536 13504 17542
rect 13452 17478 13504 17484
rect 13464 17338 13492 17478
rect 13452 17332 13504 17338
rect 13452 17274 13504 17280
rect 13268 17264 13320 17270
rect 13268 17206 13320 17212
rect 12808 17196 12860 17202
rect 12808 17138 12860 17144
rect 12900 17196 12952 17202
rect 12900 17138 12952 17144
rect 12716 16788 12768 16794
rect 12716 16730 12768 16736
rect 12532 16652 12584 16658
rect 12452 16612 12532 16640
rect 12164 16584 12216 16590
rect 12164 16526 12216 16532
rect 12176 16250 12204 16526
rect 12164 16244 12216 16250
rect 12164 16186 12216 16192
rect 12072 15564 12124 15570
rect 12072 15506 12124 15512
rect 12084 14822 12112 15506
rect 12072 14816 12124 14822
rect 12072 14758 12124 14764
rect 12084 11801 12112 14758
rect 12256 14544 12308 14550
rect 12256 14486 12308 14492
rect 12268 14346 12296 14486
rect 12452 14414 12480 16612
rect 12532 16594 12584 16600
rect 12912 16522 12940 17138
rect 13280 16998 13308 17206
rect 13728 17060 13780 17066
rect 13728 17002 13780 17008
rect 13268 16992 13320 16998
rect 13268 16934 13320 16940
rect 13544 16992 13596 16998
rect 13544 16934 13596 16940
rect 13268 16720 13320 16726
rect 13268 16662 13320 16668
rect 12900 16516 12952 16522
rect 12900 16458 12952 16464
rect 12956 16348 13252 16368
rect 13012 16346 13036 16348
rect 13092 16346 13116 16348
rect 13172 16346 13196 16348
rect 13034 16294 13036 16346
rect 13098 16294 13110 16346
rect 13172 16294 13174 16346
rect 13012 16292 13036 16294
rect 13092 16292 13116 16294
rect 13172 16292 13196 16294
rect 12956 16272 13252 16292
rect 13280 16182 13308 16662
rect 13360 16584 13412 16590
rect 13360 16526 13412 16532
rect 13372 16250 13400 16526
rect 13360 16244 13412 16250
rect 13360 16186 13412 16192
rect 13268 16176 13320 16182
rect 13268 16118 13320 16124
rect 13268 15904 13320 15910
rect 13268 15846 13320 15852
rect 12624 15496 12676 15502
rect 12624 15438 12676 15444
rect 12532 15360 12584 15366
rect 12532 15302 12584 15308
rect 12544 15026 12572 15302
rect 12532 15020 12584 15026
rect 12532 14962 12584 14968
rect 12636 14890 12664 15438
rect 12956 15260 13252 15280
rect 13012 15258 13036 15260
rect 13092 15258 13116 15260
rect 13172 15258 13196 15260
rect 13034 15206 13036 15258
rect 13098 15206 13110 15258
rect 13172 15206 13174 15258
rect 13012 15204 13036 15206
rect 13092 15204 13116 15206
rect 13172 15204 13196 15206
rect 12956 15184 13252 15204
rect 12624 14884 12676 14890
rect 12624 14826 12676 14832
rect 12636 14550 12664 14826
rect 12808 14612 12860 14618
rect 12808 14554 12860 14560
rect 12624 14544 12676 14550
rect 12624 14486 12676 14492
rect 12440 14408 12492 14414
rect 12440 14350 12492 14356
rect 12256 14340 12308 14346
rect 12256 14282 12308 14288
rect 12268 14074 12296 14282
rect 12256 14068 12308 14074
rect 12256 14010 12308 14016
rect 12452 13920 12480 14350
rect 12624 14000 12676 14006
rect 12624 13942 12676 13948
rect 12532 13932 12584 13938
rect 12452 13892 12532 13920
rect 12532 13874 12584 13880
rect 12636 13802 12664 13942
rect 12624 13796 12676 13802
rect 12624 13738 12676 13744
rect 12440 13728 12492 13734
rect 12440 13670 12492 13676
rect 12346 13288 12402 13297
rect 12346 13223 12402 13232
rect 12360 12782 12388 13223
rect 12452 13190 12480 13670
rect 12820 13530 12848 14554
rect 12956 14172 13252 14192
rect 13012 14170 13036 14172
rect 13092 14170 13116 14172
rect 13172 14170 13196 14172
rect 13034 14118 13036 14170
rect 13098 14118 13110 14170
rect 13172 14118 13174 14170
rect 13012 14116 13036 14118
rect 13092 14116 13116 14118
rect 13172 14116 13196 14118
rect 12956 14096 13252 14116
rect 13176 13728 13228 13734
rect 13176 13670 13228 13676
rect 12808 13524 12860 13530
rect 12808 13466 12860 13472
rect 13188 13462 13216 13670
rect 13176 13456 13228 13462
rect 13176 13398 13228 13404
rect 12440 13184 12492 13190
rect 12440 13126 12492 13132
rect 12452 12986 12480 13126
rect 12956 13084 13252 13104
rect 13012 13082 13036 13084
rect 13092 13082 13116 13084
rect 13172 13082 13196 13084
rect 13034 13030 13036 13082
rect 13098 13030 13110 13082
rect 13172 13030 13174 13082
rect 13012 13028 13036 13030
rect 13092 13028 13116 13030
rect 13172 13028 13196 13030
rect 12956 13008 13252 13028
rect 12440 12980 12492 12986
rect 12440 12922 12492 12928
rect 12348 12776 12400 12782
rect 12348 12718 12400 12724
rect 12164 12096 12216 12102
rect 12164 12038 12216 12044
rect 12532 12096 12584 12102
rect 12532 12038 12584 12044
rect 12176 11898 12204 12038
rect 12164 11892 12216 11898
rect 12164 11834 12216 11840
rect 12070 11792 12126 11801
rect 12070 11727 12126 11736
rect 12176 11558 12204 11834
rect 12544 11626 12572 12038
rect 12956 11996 13252 12016
rect 13012 11994 13036 11996
rect 13092 11994 13116 11996
rect 13172 11994 13196 11996
rect 13034 11942 13036 11994
rect 13098 11942 13110 11994
rect 13172 11942 13174 11994
rect 13012 11940 13036 11942
rect 13092 11940 13116 11942
rect 13172 11940 13196 11942
rect 12956 11920 13252 11940
rect 12532 11620 12584 11626
rect 12532 11562 12584 11568
rect 12164 11552 12216 11558
rect 12164 11494 12216 11500
rect 12348 11008 12400 11014
rect 12348 10950 12400 10956
rect 11980 10804 12032 10810
rect 11980 10746 12032 10752
rect 12360 10538 12388 10950
rect 12348 10532 12400 10538
rect 12348 10474 12400 10480
rect 11204 10424 11284 10452
rect 11704 10464 11756 10470
rect 11152 10406 11204 10412
rect 11704 10406 11756 10412
rect 12164 10464 12216 10470
rect 12164 10406 12216 10412
rect 10968 9920 11020 9926
rect 10968 9862 11020 9868
rect 10980 9722 11008 9862
rect 10968 9716 11020 9722
rect 10968 9658 11020 9664
rect 11164 9450 11192 10406
rect 11716 10198 11744 10406
rect 11704 10192 11756 10198
rect 11704 10134 11756 10140
rect 11152 9444 11204 9450
rect 11152 9386 11204 9392
rect 10968 8356 11020 8362
rect 10968 8298 11020 8304
rect 10980 8090 11008 8298
rect 10968 8084 11020 8090
rect 10968 8026 11020 8032
rect 11164 8022 11192 9386
rect 11334 9208 11390 9217
rect 11716 9178 11744 10134
rect 12176 9654 12204 10406
rect 12256 10192 12308 10198
rect 12256 10134 12308 10140
rect 12268 9722 12296 10134
rect 12360 10062 12388 10474
rect 12544 10062 12572 11562
rect 12956 10908 13252 10928
rect 13012 10906 13036 10908
rect 13092 10906 13116 10908
rect 13172 10906 13196 10908
rect 13034 10854 13036 10906
rect 13098 10854 13110 10906
rect 13172 10854 13174 10906
rect 13012 10852 13036 10854
rect 13092 10852 13116 10854
rect 13172 10852 13196 10854
rect 12956 10832 13252 10852
rect 12808 10668 12860 10674
rect 12808 10610 12860 10616
rect 12716 10464 12768 10470
rect 12716 10406 12768 10412
rect 12348 10056 12400 10062
rect 12348 9998 12400 10004
rect 12532 10056 12584 10062
rect 12532 9998 12584 10004
rect 12256 9716 12308 9722
rect 12256 9658 12308 9664
rect 12164 9648 12216 9654
rect 12164 9590 12216 9596
rect 12268 9382 12296 9658
rect 12532 9444 12584 9450
rect 12532 9386 12584 9392
rect 12256 9376 12308 9382
rect 12256 9318 12308 9324
rect 12544 9178 12572 9386
rect 11334 9143 11390 9152
rect 11704 9172 11756 9178
rect 11348 8974 11376 9143
rect 11704 9114 11756 9120
rect 12532 9172 12584 9178
rect 12532 9114 12584 9120
rect 12256 9104 12308 9110
rect 12256 9046 12308 9052
rect 11336 8968 11388 8974
rect 11336 8910 11388 8916
rect 11348 8294 11376 8910
rect 12268 8634 12296 9046
rect 12348 8968 12400 8974
rect 12348 8910 12400 8916
rect 12256 8628 12308 8634
rect 12256 8570 12308 8576
rect 12268 8294 12296 8570
rect 11336 8288 11388 8294
rect 11336 8230 11388 8236
rect 12256 8288 12308 8294
rect 12256 8230 12308 8236
rect 11152 8016 11204 8022
rect 10506 7984 10562 7993
rect 11152 7958 11204 7964
rect 10506 7919 10562 7928
rect 10416 7880 10468 7886
rect 10416 7822 10468 7828
rect 10428 5846 10456 7822
rect 11164 7206 11192 7958
rect 11152 7200 11204 7206
rect 11152 7142 11204 7148
rect 11244 7200 11296 7206
rect 11244 7142 11296 7148
rect 11164 7002 11192 7142
rect 11152 6996 11204 7002
rect 11152 6938 11204 6944
rect 11256 6866 11284 7142
rect 11244 6860 11296 6866
rect 11244 6802 11296 6808
rect 10968 6656 11020 6662
rect 10968 6598 11020 6604
rect 10980 6118 11008 6598
rect 10968 6112 11020 6118
rect 10968 6054 11020 6060
rect 10416 5840 10468 5846
rect 10416 5782 10468 5788
rect 10324 5704 10376 5710
rect 10324 5646 10376 5652
rect 10980 5642 11008 6054
rect 10968 5636 11020 5642
rect 10968 5578 11020 5584
rect 10980 5370 11008 5578
rect 10968 5364 11020 5370
rect 10968 5306 11020 5312
rect 10232 5228 10284 5234
rect 10232 5170 10284 5176
rect 10244 4486 10272 5170
rect 11348 5137 11376 8230
rect 12268 8090 12296 8230
rect 12360 8090 12388 8910
rect 12624 8492 12676 8498
rect 12624 8434 12676 8440
rect 12256 8084 12308 8090
rect 12256 8026 12308 8032
rect 12348 8084 12400 8090
rect 12348 8026 12400 8032
rect 12532 8016 12584 8022
rect 12532 7958 12584 7964
rect 12544 7188 12572 7958
rect 12636 7750 12664 8434
rect 12624 7744 12676 7750
rect 12624 7686 12676 7692
rect 12636 7546 12664 7686
rect 12624 7540 12676 7546
rect 12624 7482 12676 7488
rect 12624 7200 12676 7206
rect 12544 7160 12624 7188
rect 12624 7142 12676 7148
rect 12530 6896 12586 6905
rect 12530 6831 12586 6840
rect 11704 6792 11756 6798
rect 11704 6734 11756 6740
rect 12348 6792 12400 6798
rect 12348 6734 12400 6740
rect 11716 6458 11744 6734
rect 11704 6452 11756 6458
rect 11704 6394 11756 6400
rect 11716 6361 11744 6394
rect 11702 6352 11758 6361
rect 11702 6287 11758 6296
rect 11716 5370 11744 6287
rect 12360 6118 12388 6734
rect 12544 6254 12572 6831
rect 12532 6248 12584 6254
rect 12532 6190 12584 6196
rect 12348 6112 12400 6118
rect 12348 6054 12400 6060
rect 12360 5846 12388 6054
rect 12348 5840 12400 5846
rect 12348 5782 12400 5788
rect 11980 5772 12032 5778
rect 11980 5714 12032 5720
rect 11704 5364 11756 5370
rect 11704 5306 11756 5312
rect 11334 5128 11390 5137
rect 11716 5098 11744 5306
rect 11886 5128 11942 5137
rect 11334 5063 11390 5072
rect 11704 5092 11756 5098
rect 11886 5063 11942 5072
rect 11704 5034 11756 5040
rect 11060 5024 11112 5030
rect 11060 4966 11112 4972
rect 10232 4480 10284 4486
rect 10232 4422 10284 4428
rect 10692 4072 10744 4078
rect 10692 4014 10744 4020
rect 10508 3936 10560 3942
rect 10508 3878 10560 3884
rect 10520 2922 10548 3878
rect 10508 2916 10560 2922
rect 10508 2858 10560 2864
rect 10704 2650 10732 4014
rect 11072 3738 11100 4966
rect 11900 4690 11928 5063
rect 11888 4684 11940 4690
rect 11888 4626 11940 4632
rect 11900 4214 11928 4626
rect 11992 4622 12020 5714
rect 12636 5692 12664 7142
rect 12728 6934 12756 10406
rect 12820 9586 12848 10610
rect 13176 10532 13228 10538
rect 13176 10474 13228 10480
rect 13188 9994 13216 10474
rect 13176 9988 13228 9994
rect 13176 9930 13228 9936
rect 12956 9820 13252 9840
rect 13012 9818 13036 9820
rect 13092 9818 13116 9820
rect 13172 9818 13196 9820
rect 13034 9766 13036 9818
rect 13098 9766 13110 9818
rect 13172 9766 13174 9818
rect 13012 9764 13036 9766
rect 13092 9764 13116 9766
rect 13172 9764 13196 9766
rect 12956 9744 13252 9764
rect 12808 9580 12860 9586
rect 12808 9522 12860 9528
rect 12820 9110 12848 9522
rect 12808 9104 12860 9110
rect 12808 9046 12860 9052
rect 12956 8732 13252 8752
rect 13012 8730 13036 8732
rect 13092 8730 13116 8732
rect 13172 8730 13196 8732
rect 13034 8678 13036 8730
rect 13098 8678 13110 8730
rect 13172 8678 13174 8730
rect 13012 8676 13036 8678
rect 13092 8676 13116 8678
rect 13172 8676 13196 8678
rect 12956 8656 13252 8676
rect 12808 7948 12860 7954
rect 12808 7890 12860 7896
rect 12820 7546 12848 7890
rect 12956 7644 13252 7664
rect 13012 7642 13036 7644
rect 13092 7642 13116 7644
rect 13172 7642 13196 7644
rect 13034 7590 13036 7642
rect 13098 7590 13110 7642
rect 13172 7590 13174 7642
rect 13012 7588 13036 7590
rect 13092 7588 13116 7590
rect 13172 7588 13196 7590
rect 12956 7568 13252 7588
rect 12808 7540 12860 7546
rect 12808 7482 12860 7488
rect 13280 7313 13308 15846
rect 13556 15570 13584 16934
rect 13740 15910 13768 17002
rect 13728 15904 13780 15910
rect 13728 15846 13780 15852
rect 13544 15564 13596 15570
rect 13544 15506 13596 15512
rect 13556 15162 13584 15506
rect 13544 15156 13596 15162
rect 13544 15098 13596 15104
rect 13740 14822 13768 15846
rect 13832 14890 13860 17546
rect 14096 17128 14148 17134
rect 14096 17070 14148 17076
rect 14108 16794 14136 17070
rect 14096 16788 14148 16794
rect 14096 16730 14148 16736
rect 15028 16182 15056 23582
rect 16592 23582 17002 23610
rect 16592 20602 16620 23582
rect 16946 23520 17002 23582
rect 18878 23610 18934 24000
rect 20902 23610 20958 24000
rect 22926 23610 22982 24000
rect 18878 23582 19012 23610
rect 18878 23520 18934 23582
rect 16956 21244 17252 21264
rect 17012 21242 17036 21244
rect 17092 21242 17116 21244
rect 17172 21242 17196 21244
rect 17034 21190 17036 21242
rect 17098 21190 17110 21242
rect 17172 21190 17174 21242
rect 17012 21188 17036 21190
rect 17092 21188 17116 21190
rect 17172 21188 17196 21190
rect 16956 21168 17252 21188
rect 16580 20596 16632 20602
rect 16580 20538 16632 20544
rect 15108 20392 15160 20398
rect 15108 20334 15160 20340
rect 18236 20392 18288 20398
rect 18236 20334 18288 20340
rect 15016 16176 15068 16182
rect 15016 16118 15068 16124
rect 14740 15496 14792 15502
rect 14740 15438 14792 15444
rect 14004 15360 14056 15366
rect 14004 15302 14056 15308
rect 14016 14958 14044 15302
rect 14004 14952 14056 14958
rect 14004 14894 14056 14900
rect 14556 14952 14608 14958
rect 14556 14894 14608 14900
rect 13820 14884 13872 14890
rect 13872 14844 13952 14872
rect 13820 14826 13872 14832
rect 13728 14816 13780 14822
rect 13728 14758 13780 14764
rect 13820 14544 13872 14550
rect 13820 14486 13872 14492
rect 13728 14408 13780 14414
rect 13728 14350 13780 14356
rect 13740 13734 13768 14350
rect 13832 14006 13860 14486
rect 13924 14414 13952 14844
rect 13912 14408 13964 14414
rect 13912 14350 13964 14356
rect 13820 14000 13872 14006
rect 13820 13942 13872 13948
rect 13728 13728 13780 13734
rect 13728 13670 13780 13676
rect 13728 13388 13780 13394
rect 13728 13330 13780 13336
rect 13740 12986 13768 13330
rect 13728 12980 13780 12986
rect 13728 12922 13780 12928
rect 13740 12646 13768 12922
rect 13728 12640 13780 12646
rect 13728 12582 13780 12588
rect 13452 12368 13504 12374
rect 13452 12310 13504 12316
rect 13360 12096 13412 12102
rect 13360 12038 13412 12044
rect 13372 8022 13400 12038
rect 13464 11558 13492 12310
rect 13636 12164 13688 12170
rect 13636 12106 13688 12112
rect 13648 11830 13676 12106
rect 13636 11824 13688 11830
rect 13636 11766 13688 11772
rect 13452 11552 13504 11558
rect 13452 11494 13504 11500
rect 13464 11354 13492 11494
rect 13452 11348 13504 11354
rect 13452 11290 13504 11296
rect 13636 11212 13688 11218
rect 13740 11200 13768 12582
rect 13820 12232 13872 12238
rect 13820 12174 13872 12180
rect 13832 11558 13860 12174
rect 13820 11552 13872 11558
rect 13820 11494 13872 11500
rect 13688 11172 13768 11200
rect 13636 11154 13688 11160
rect 13452 10804 13504 10810
rect 13452 10746 13504 10752
rect 13464 9761 13492 10746
rect 13648 10470 13676 11154
rect 13728 11008 13780 11014
rect 13728 10950 13780 10956
rect 13636 10464 13688 10470
rect 13636 10406 13688 10412
rect 13544 10260 13596 10266
rect 13544 10202 13596 10208
rect 13450 9752 13506 9761
rect 13450 9687 13506 9696
rect 13556 9654 13584 10202
rect 13740 10198 13768 10950
rect 13832 10674 13860 11494
rect 14016 11200 14044 14894
rect 14568 13734 14596 14894
rect 14752 14890 14780 15438
rect 14740 14884 14792 14890
rect 14740 14826 14792 14832
rect 14648 14816 14700 14822
rect 14648 14758 14700 14764
rect 14556 13728 14608 13734
rect 14556 13670 14608 13676
rect 14188 13388 14240 13394
rect 14188 13330 14240 13336
rect 14200 12918 14228 13330
rect 14280 13320 14332 13326
rect 14280 13262 14332 13268
rect 14188 12912 14240 12918
rect 14188 12854 14240 12860
rect 14292 12850 14320 13262
rect 14280 12844 14332 12850
rect 14280 12786 14332 12792
rect 14292 12442 14320 12786
rect 14280 12436 14332 12442
rect 14280 12378 14332 12384
rect 14568 12102 14596 13670
rect 14660 12646 14688 14758
rect 14752 14618 14780 14826
rect 14740 14612 14792 14618
rect 14740 14554 14792 14560
rect 14740 13864 14792 13870
rect 14740 13806 14792 13812
rect 14752 13530 14780 13806
rect 14740 13524 14792 13530
rect 14740 13466 14792 13472
rect 14648 12640 14700 12646
rect 14648 12582 14700 12588
rect 14556 12096 14608 12102
rect 14556 12038 14608 12044
rect 14660 11898 14688 12582
rect 15120 12345 15148 20334
rect 16956 20156 17252 20176
rect 17012 20154 17036 20156
rect 17092 20154 17116 20156
rect 17172 20154 17196 20156
rect 17034 20102 17036 20154
rect 17098 20102 17110 20154
rect 17172 20102 17174 20154
rect 17012 20100 17036 20102
rect 17092 20100 17116 20102
rect 17172 20100 17196 20102
rect 16956 20080 17252 20100
rect 17684 19916 17736 19922
rect 17684 19858 17736 19864
rect 17696 19174 17724 19858
rect 17684 19168 17736 19174
rect 17684 19110 17736 19116
rect 16956 19068 17252 19088
rect 17012 19066 17036 19068
rect 17092 19066 17116 19068
rect 17172 19066 17196 19068
rect 17034 19014 17036 19066
rect 17098 19014 17110 19066
rect 17172 19014 17174 19066
rect 17012 19012 17036 19014
rect 17092 19012 17116 19014
rect 17172 19012 17196 19014
rect 16956 18992 17252 19012
rect 15200 18828 15252 18834
rect 15200 18770 15252 18776
rect 16672 18828 16724 18834
rect 16672 18770 16724 18776
rect 15212 18086 15240 18770
rect 15568 18624 15620 18630
rect 15568 18566 15620 18572
rect 15752 18624 15804 18630
rect 15752 18566 15804 18572
rect 16120 18624 16172 18630
rect 16120 18566 16172 18572
rect 15200 18080 15252 18086
rect 15200 18022 15252 18028
rect 15212 17814 15240 18022
rect 15200 17808 15252 17814
rect 15200 17750 15252 17756
rect 15106 12336 15162 12345
rect 15106 12271 15162 12280
rect 14648 11892 14700 11898
rect 14648 11834 14700 11840
rect 14660 11626 14688 11834
rect 14832 11688 14884 11694
rect 14832 11630 14884 11636
rect 14648 11620 14700 11626
rect 14648 11562 14700 11568
rect 14844 11286 14872 11630
rect 14832 11280 14884 11286
rect 14832 11222 14884 11228
rect 15212 11218 15240 17750
rect 15292 17672 15344 17678
rect 15292 17614 15344 17620
rect 15304 17338 15332 17614
rect 15476 17536 15528 17542
rect 15476 17478 15528 17484
rect 15292 17332 15344 17338
rect 15292 17274 15344 17280
rect 15488 16658 15516 17478
rect 15580 17202 15608 18566
rect 15764 18154 15792 18566
rect 16132 18290 16160 18566
rect 16120 18284 16172 18290
rect 16120 18226 16172 18232
rect 15752 18148 15804 18154
rect 15752 18090 15804 18096
rect 15764 17882 15792 18090
rect 16684 18086 16712 18770
rect 16856 18760 16908 18766
rect 16856 18702 16908 18708
rect 17316 18760 17368 18766
rect 17316 18702 17368 18708
rect 16868 18426 16896 18702
rect 16856 18420 16908 18426
rect 16856 18362 16908 18368
rect 16868 18086 16896 18362
rect 16672 18080 16724 18086
rect 16672 18022 16724 18028
rect 16856 18080 16908 18086
rect 16856 18022 16908 18028
rect 15660 17876 15712 17882
rect 15660 17818 15712 17824
rect 15752 17876 15804 17882
rect 15752 17818 15804 17824
rect 15568 17196 15620 17202
rect 15568 17138 15620 17144
rect 15672 16998 15700 17818
rect 15764 17048 15792 17818
rect 16212 17196 16264 17202
rect 16212 17138 16264 17144
rect 15844 17060 15896 17066
rect 15764 17020 15844 17048
rect 15844 17002 15896 17008
rect 15660 16992 15712 16998
rect 15660 16934 15712 16940
rect 15476 16652 15528 16658
rect 15476 16594 15528 16600
rect 15488 16250 15516 16594
rect 15476 16244 15528 16250
rect 15476 16186 15528 16192
rect 15672 15706 15700 16934
rect 15856 16794 15884 17002
rect 16224 16794 16252 17138
rect 16396 17060 16448 17066
rect 16396 17002 16448 17008
rect 15844 16788 15896 16794
rect 15844 16730 15896 16736
rect 16212 16788 16264 16794
rect 16212 16730 16264 16736
rect 15844 16448 15896 16454
rect 15844 16390 15896 16396
rect 15856 16114 15884 16390
rect 16408 16182 16436 17002
rect 16396 16176 16448 16182
rect 16396 16118 16448 16124
rect 15844 16108 15896 16114
rect 15844 16050 15896 16056
rect 16212 15972 16264 15978
rect 16212 15914 16264 15920
rect 16224 15706 16252 15914
rect 16684 15910 16712 18022
rect 16956 17980 17252 18000
rect 17012 17978 17036 17980
rect 17092 17978 17116 17980
rect 17172 17978 17196 17980
rect 17034 17926 17036 17978
rect 17098 17926 17110 17978
rect 17172 17926 17174 17978
rect 17012 17924 17036 17926
rect 17092 17924 17116 17926
rect 17172 17924 17196 17926
rect 16956 17904 17252 17924
rect 17328 17746 17356 18702
rect 17408 18080 17460 18086
rect 17408 18022 17460 18028
rect 17500 18080 17552 18086
rect 17500 18022 17552 18028
rect 17316 17740 17368 17746
rect 17316 17682 17368 17688
rect 16956 16892 17252 16912
rect 17012 16890 17036 16892
rect 17092 16890 17116 16892
rect 17172 16890 17196 16892
rect 17034 16838 17036 16890
rect 17098 16838 17110 16890
rect 17172 16838 17174 16890
rect 17012 16836 17036 16838
rect 17092 16836 17116 16838
rect 17172 16836 17196 16838
rect 16956 16816 17252 16836
rect 17328 16794 17356 17682
rect 17316 16788 17368 16794
rect 17316 16730 17368 16736
rect 17316 16652 17368 16658
rect 17316 16594 17368 16600
rect 17328 15910 17356 16594
rect 16672 15904 16724 15910
rect 16672 15846 16724 15852
rect 17316 15904 17368 15910
rect 17316 15846 17368 15852
rect 16956 15804 17252 15824
rect 17012 15802 17036 15804
rect 17092 15802 17116 15804
rect 17172 15802 17196 15804
rect 17034 15750 17036 15802
rect 17098 15750 17110 15802
rect 17172 15750 17174 15802
rect 17012 15748 17036 15750
rect 17092 15748 17116 15750
rect 17172 15748 17196 15750
rect 16956 15728 17252 15748
rect 15660 15700 15712 15706
rect 15660 15642 15712 15648
rect 16212 15700 16264 15706
rect 16212 15642 16264 15648
rect 15476 14952 15528 14958
rect 15476 14894 15528 14900
rect 15488 13938 15516 14894
rect 15672 14822 15700 15642
rect 16120 15428 16172 15434
rect 16120 15370 16172 15376
rect 15660 14816 15712 14822
rect 15660 14758 15712 14764
rect 15844 14544 15896 14550
rect 15844 14486 15896 14492
rect 15752 14408 15804 14414
rect 15752 14350 15804 14356
rect 15764 14074 15792 14350
rect 15752 14068 15804 14074
rect 15752 14010 15804 14016
rect 15856 14006 15884 14486
rect 15844 14000 15896 14006
rect 15844 13942 15896 13948
rect 15476 13932 15528 13938
rect 15476 13874 15528 13880
rect 16028 13456 16080 13462
rect 16028 13398 16080 13404
rect 15936 13320 15988 13326
rect 15936 13262 15988 13268
rect 15844 12776 15896 12782
rect 15844 12718 15896 12724
rect 15856 11694 15884 12718
rect 15948 12442 15976 13262
rect 16040 12986 16068 13398
rect 16132 13190 16160 15370
rect 16224 14550 16252 15642
rect 17132 15564 17184 15570
rect 17132 15506 17184 15512
rect 16488 15360 16540 15366
rect 16488 15302 16540 15308
rect 16500 14958 16528 15302
rect 16488 14952 16540 14958
rect 16488 14894 16540 14900
rect 17144 14890 17172 15506
rect 16580 14884 16632 14890
rect 16580 14826 16632 14832
rect 17132 14884 17184 14890
rect 17132 14826 17184 14832
rect 16592 14770 16620 14826
rect 16500 14742 16620 14770
rect 16212 14544 16264 14550
rect 16212 14486 16264 14492
rect 16120 13184 16172 13190
rect 16120 13126 16172 13132
rect 16028 12980 16080 12986
rect 16028 12922 16080 12928
rect 16040 12646 16068 12922
rect 16132 12850 16160 13126
rect 16120 12844 16172 12850
rect 16120 12786 16172 12792
rect 16028 12640 16080 12646
rect 16028 12582 16080 12588
rect 15936 12436 15988 12442
rect 15936 12378 15988 12384
rect 16212 12368 16264 12374
rect 16212 12310 16264 12316
rect 16120 12232 16172 12238
rect 16120 12174 16172 12180
rect 16132 11898 16160 12174
rect 16120 11892 16172 11898
rect 16120 11834 16172 11840
rect 16224 11762 16252 12310
rect 16212 11756 16264 11762
rect 16212 11698 16264 11704
rect 15844 11688 15896 11694
rect 15844 11630 15896 11636
rect 15752 11620 15804 11626
rect 15752 11562 15804 11568
rect 14188 11212 14240 11218
rect 14016 11172 14188 11200
rect 14188 11154 14240 11160
rect 15200 11212 15252 11218
rect 15200 11154 15252 11160
rect 13820 10668 13872 10674
rect 13820 10610 13872 10616
rect 14200 10606 14228 11154
rect 14188 10600 14240 10606
rect 14188 10542 14240 10548
rect 14372 10532 14424 10538
rect 14372 10474 14424 10480
rect 15384 10532 15436 10538
rect 15384 10474 15436 10480
rect 13728 10192 13780 10198
rect 13648 10152 13728 10180
rect 13544 9648 13596 9654
rect 13544 9590 13596 9596
rect 13452 9580 13504 9586
rect 13452 9522 13504 9528
rect 13360 8016 13412 8022
rect 13360 7958 13412 7964
rect 13464 7478 13492 9522
rect 13542 9480 13598 9489
rect 13542 9415 13598 9424
rect 13556 9042 13584 9415
rect 13648 9178 13676 10152
rect 13728 10134 13780 10140
rect 13912 10056 13964 10062
rect 13912 9998 13964 10004
rect 13740 9722 13860 9738
rect 13740 9716 13872 9722
rect 13740 9710 13820 9716
rect 13740 9586 13768 9710
rect 13820 9658 13872 9664
rect 13728 9580 13780 9586
rect 13728 9522 13780 9528
rect 13636 9172 13688 9178
rect 13636 9114 13688 9120
rect 13544 9036 13596 9042
rect 13544 8978 13596 8984
rect 13556 8294 13584 8978
rect 13924 8498 13952 9998
rect 14384 9722 14412 10474
rect 15396 10062 15424 10474
rect 15764 10266 15792 11562
rect 16212 11212 16264 11218
rect 16212 11154 16264 11160
rect 16224 10538 16252 11154
rect 16212 10532 16264 10538
rect 16212 10474 16264 10480
rect 15752 10260 15804 10266
rect 15752 10202 15804 10208
rect 15384 10056 15436 10062
rect 15384 9998 15436 10004
rect 15396 9722 15424 9998
rect 15474 9752 15530 9761
rect 14372 9716 14424 9722
rect 14372 9658 14424 9664
rect 15384 9716 15436 9722
rect 15474 9687 15530 9696
rect 15384 9658 15436 9664
rect 14004 9648 14056 9654
rect 14004 9590 14056 9596
rect 14016 9217 14044 9590
rect 14464 9512 14516 9518
rect 14464 9454 14516 9460
rect 14002 9208 14058 9217
rect 14476 9178 14504 9454
rect 15200 9444 15252 9450
rect 15200 9386 15252 9392
rect 14002 9143 14058 9152
rect 14464 9172 14516 9178
rect 14464 9114 14516 9120
rect 14476 8838 14504 9114
rect 14738 8936 14794 8945
rect 15212 8906 15240 9386
rect 15488 9042 15516 9687
rect 15764 9674 15792 10202
rect 16304 9920 16356 9926
rect 16304 9862 16356 9868
rect 16316 9722 16344 9862
rect 16304 9716 16356 9722
rect 15764 9646 15884 9674
rect 16304 9658 16356 9664
rect 15856 9382 15884 9646
rect 16316 9450 16344 9658
rect 16304 9444 16356 9450
rect 16304 9386 16356 9392
rect 15844 9376 15896 9382
rect 15844 9318 15896 9324
rect 15476 9036 15528 9042
rect 15476 8978 15528 8984
rect 14738 8871 14794 8880
rect 15200 8900 15252 8906
rect 14464 8832 14516 8838
rect 14464 8774 14516 8780
rect 13912 8492 13964 8498
rect 13912 8434 13964 8440
rect 14464 8424 14516 8430
rect 14464 8366 14516 8372
rect 13544 8288 13596 8294
rect 13544 8230 13596 8236
rect 13728 8288 13780 8294
rect 13728 8230 13780 8236
rect 13452 7472 13504 7478
rect 13358 7440 13414 7449
rect 13452 7414 13504 7420
rect 13358 7375 13414 7384
rect 13372 7342 13400 7375
rect 13360 7336 13412 7342
rect 13266 7304 13322 7313
rect 13360 7278 13412 7284
rect 13266 7239 13322 7248
rect 13452 7268 13504 7274
rect 13452 7210 13504 7216
rect 12716 6928 12768 6934
rect 12716 6870 12768 6876
rect 12808 6656 12860 6662
rect 12808 6598 12860 6604
rect 12820 5710 12848 6598
rect 12956 6556 13252 6576
rect 13012 6554 13036 6556
rect 13092 6554 13116 6556
rect 13172 6554 13196 6556
rect 13034 6502 13036 6554
rect 13098 6502 13110 6554
rect 13172 6502 13174 6554
rect 13012 6500 13036 6502
rect 13092 6500 13116 6502
rect 13172 6500 13196 6502
rect 12956 6480 13252 6500
rect 13464 6322 13492 7210
rect 13452 6316 13504 6322
rect 13452 6258 13504 6264
rect 13268 6180 13320 6186
rect 13268 6122 13320 6128
rect 12808 5704 12860 5710
rect 12636 5664 12756 5692
rect 12624 5568 12676 5574
rect 12624 5510 12676 5516
rect 12636 5234 12664 5510
rect 12624 5228 12676 5234
rect 12624 5170 12676 5176
rect 12636 4758 12664 5170
rect 12728 4758 12756 5664
rect 12808 5646 12860 5652
rect 12820 4826 12848 5646
rect 12956 5468 13252 5488
rect 13012 5466 13036 5468
rect 13092 5466 13116 5468
rect 13172 5466 13196 5468
rect 13034 5414 13036 5466
rect 13098 5414 13110 5466
rect 13172 5414 13174 5466
rect 13012 5412 13036 5414
rect 13092 5412 13116 5414
rect 13172 5412 13196 5414
rect 12956 5392 13252 5412
rect 13280 5234 13308 6122
rect 13464 5914 13492 6258
rect 13556 6254 13584 8230
rect 13740 8090 13768 8230
rect 13728 8084 13780 8090
rect 13728 8026 13780 8032
rect 14476 7857 14504 8366
rect 14752 7954 14780 8871
rect 15200 8842 15252 8848
rect 15212 8498 15240 8842
rect 15200 8492 15252 8498
rect 15200 8434 15252 8440
rect 15488 8294 15516 8978
rect 15856 8498 15884 9318
rect 15844 8492 15896 8498
rect 15844 8434 15896 8440
rect 15856 8362 15884 8434
rect 15844 8356 15896 8362
rect 15844 8298 15896 8304
rect 15476 8288 15528 8294
rect 15476 8230 15528 8236
rect 15016 8084 15068 8090
rect 15016 8026 15068 8032
rect 14740 7948 14792 7954
rect 14740 7890 14792 7896
rect 14462 7848 14518 7857
rect 14462 7783 14518 7792
rect 13820 7744 13872 7750
rect 13820 7686 13872 7692
rect 14188 7744 14240 7750
rect 14188 7686 14240 7692
rect 13832 7274 13860 7686
rect 14200 7410 14228 7686
rect 14752 7546 14780 7890
rect 14740 7540 14792 7546
rect 14740 7482 14792 7488
rect 14924 7472 14976 7478
rect 14924 7414 14976 7420
rect 14188 7404 14240 7410
rect 14188 7346 14240 7352
rect 13820 7268 13872 7274
rect 13820 7210 13872 7216
rect 13832 7002 13860 7210
rect 14200 7002 14228 7346
rect 13820 6996 13872 7002
rect 13820 6938 13872 6944
rect 14188 6996 14240 7002
rect 14188 6938 14240 6944
rect 13544 6248 13596 6254
rect 13544 6190 13596 6196
rect 13832 6186 13860 6938
rect 13912 6316 13964 6322
rect 13912 6258 13964 6264
rect 13820 6180 13872 6186
rect 13820 6122 13872 6128
rect 13544 6112 13596 6118
rect 13544 6054 13596 6060
rect 13452 5908 13504 5914
rect 13452 5850 13504 5856
rect 13360 5840 13412 5846
rect 13360 5782 13412 5788
rect 13372 5370 13400 5782
rect 13360 5364 13412 5370
rect 13360 5306 13412 5312
rect 13268 5228 13320 5234
rect 13268 5170 13320 5176
rect 13452 5160 13504 5166
rect 13452 5102 13504 5108
rect 12808 4820 12860 4826
rect 12808 4762 12860 4768
rect 12624 4752 12676 4758
rect 12624 4694 12676 4700
rect 12716 4752 12768 4758
rect 12716 4694 12768 4700
rect 13464 4690 13492 5102
rect 13556 5098 13584 6054
rect 13924 5846 13952 6258
rect 13912 5840 13964 5846
rect 13912 5782 13964 5788
rect 14464 5364 14516 5370
rect 14464 5306 14516 5312
rect 14372 5228 14424 5234
rect 14372 5170 14424 5176
rect 13544 5092 13596 5098
rect 13544 5034 13596 5040
rect 14384 4826 14412 5170
rect 14476 5098 14504 5306
rect 14936 5302 14964 7414
rect 14924 5296 14976 5302
rect 14924 5238 14976 5244
rect 14464 5092 14516 5098
rect 14464 5034 14516 5040
rect 14372 4820 14424 4826
rect 14372 4762 14424 4768
rect 13452 4684 13504 4690
rect 13452 4626 13504 4632
rect 13820 4684 13872 4690
rect 13820 4626 13872 4632
rect 11980 4616 12032 4622
rect 11980 4558 12032 4564
rect 11992 4282 12020 4558
rect 12956 4380 13252 4400
rect 13012 4378 13036 4380
rect 13092 4378 13116 4380
rect 13172 4378 13196 4380
rect 13034 4326 13036 4378
rect 13098 4326 13110 4378
rect 13172 4326 13174 4378
rect 13012 4324 13036 4326
rect 13092 4324 13116 4326
rect 13172 4324 13196 4326
rect 12956 4304 13252 4324
rect 13464 4282 13492 4626
rect 13832 4282 13860 4626
rect 13912 4616 13964 4622
rect 13912 4558 13964 4564
rect 11980 4276 12032 4282
rect 11980 4218 12032 4224
rect 13452 4276 13504 4282
rect 13452 4218 13504 4224
rect 13820 4276 13872 4282
rect 13820 4218 13872 4224
rect 11888 4208 11940 4214
rect 11888 4150 11940 4156
rect 13924 4154 13952 4558
rect 13924 4146 14044 4154
rect 13924 4140 14056 4146
rect 13924 4126 14004 4140
rect 14004 4082 14056 4088
rect 15028 4078 15056 8026
rect 15292 7948 15344 7954
rect 15292 7890 15344 7896
rect 15304 7206 15332 7890
rect 15660 7812 15712 7818
rect 15660 7754 15712 7760
rect 15672 7410 15700 7754
rect 15856 7750 15884 8298
rect 15934 7984 15990 7993
rect 15934 7919 15990 7928
rect 15844 7744 15896 7750
rect 15844 7686 15896 7692
rect 15660 7404 15712 7410
rect 15660 7346 15712 7352
rect 15752 7268 15804 7274
rect 15752 7210 15804 7216
rect 15292 7200 15344 7206
rect 15292 7142 15344 7148
rect 12716 4072 12768 4078
rect 15016 4072 15068 4078
rect 12716 4014 12768 4020
rect 13450 4040 13506 4049
rect 12440 4004 12492 4010
rect 12440 3946 12492 3952
rect 11060 3732 11112 3738
rect 11060 3674 11112 3680
rect 11072 3126 11100 3674
rect 11520 3664 11572 3670
rect 11520 3606 11572 3612
rect 11532 3194 11560 3606
rect 11796 3528 11848 3534
rect 11796 3470 11848 3476
rect 11520 3188 11572 3194
rect 11520 3130 11572 3136
rect 11060 3120 11112 3126
rect 11060 3062 11112 3068
rect 11808 3058 11836 3470
rect 12452 3194 12480 3946
rect 12728 3738 12756 4014
rect 15016 4014 15068 4020
rect 13450 3975 13506 3984
rect 13464 3738 13492 3975
rect 15028 3738 15056 4014
rect 12716 3732 12768 3738
rect 12716 3674 12768 3680
rect 13452 3732 13504 3738
rect 13452 3674 13504 3680
rect 15016 3732 15068 3738
rect 15016 3674 15068 3680
rect 12808 3528 12860 3534
rect 12808 3470 12860 3476
rect 12440 3188 12492 3194
rect 12440 3130 12492 3136
rect 11796 3052 11848 3058
rect 11796 2994 11848 3000
rect 12452 2854 12480 3130
rect 12820 3126 12848 3470
rect 12956 3292 13252 3312
rect 13012 3290 13036 3292
rect 13092 3290 13116 3292
rect 13172 3290 13196 3292
rect 13034 3238 13036 3290
rect 13098 3238 13110 3290
rect 13172 3238 13174 3290
rect 13012 3236 13036 3238
rect 13092 3236 13116 3238
rect 13172 3236 13196 3238
rect 12956 3216 13252 3236
rect 13360 3188 13412 3194
rect 13360 3130 13412 3136
rect 12808 3120 12860 3126
rect 12808 3062 12860 3068
rect 12440 2848 12492 2854
rect 12440 2790 12492 2796
rect 10692 2644 10744 2650
rect 10692 2586 10744 2592
rect 13372 2582 13400 3130
rect 13360 2576 13412 2582
rect 13360 2518 13412 2524
rect 12072 2372 12124 2378
rect 12072 2314 12124 2320
rect 10138 82 10194 480
rect 10060 54 10194 82
rect 6458 0 6514 54
rect 8298 0 8354 54
rect 10138 0 10194 54
rect 11978 82 12034 480
rect 12084 82 12112 2314
rect 15304 2310 15332 7142
rect 15764 6934 15792 7210
rect 15752 6928 15804 6934
rect 15752 6870 15804 6876
rect 15856 6186 15884 7686
rect 15948 6390 15976 7919
rect 16500 7857 16528 14742
rect 16956 14716 17252 14736
rect 17012 14714 17036 14716
rect 17092 14714 17116 14716
rect 17172 14714 17196 14716
rect 17034 14662 17036 14714
rect 17098 14662 17110 14714
rect 17172 14662 17174 14714
rect 17012 14660 17036 14662
rect 17092 14660 17116 14662
rect 17172 14660 17196 14662
rect 16956 14640 17252 14660
rect 17420 14618 17448 18022
rect 17512 17882 17540 18022
rect 17500 17876 17552 17882
rect 17500 17818 17552 17824
rect 17512 16998 17540 17818
rect 17500 16992 17552 16998
rect 17500 16934 17552 16940
rect 17512 16726 17540 16934
rect 17500 16720 17552 16726
rect 17500 16662 17552 16668
rect 17500 16584 17552 16590
rect 17500 16526 17552 16532
rect 17512 15910 17540 16526
rect 17500 15904 17552 15910
rect 17500 15846 17552 15852
rect 17408 14612 17460 14618
rect 17408 14554 17460 14560
rect 17512 14498 17540 15846
rect 17420 14470 17540 14498
rect 16956 13628 17252 13648
rect 17012 13626 17036 13628
rect 17092 13626 17116 13628
rect 17172 13626 17196 13628
rect 17034 13574 17036 13626
rect 17098 13574 17110 13626
rect 17172 13574 17174 13626
rect 17012 13572 17036 13574
rect 17092 13572 17116 13574
rect 17172 13572 17196 13574
rect 16956 13552 17252 13572
rect 17420 13190 17448 14470
rect 17500 14408 17552 14414
rect 17500 14350 17552 14356
rect 17512 13734 17540 14350
rect 17500 13728 17552 13734
rect 17500 13670 17552 13676
rect 17592 13728 17644 13734
rect 17592 13670 17644 13676
rect 17512 13394 17540 13670
rect 17500 13388 17552 13394
rect 17500 13330 17552 13336
rect 17408 13184 17460 13190
rect 17408 13126 17460 13132
rect 16764 12708 16816 12714
rect 16764 12650 16816 12656
rect 16776 12306 16804 12650
rect 17420 12646 17448 13126
rect 17512 12918 17540 13330
rect 17604 13326 17632 13670
rect 17696 13530 17724 19110
rect 17866 17640 17922 17649
rect 17866 17575 17922 17584
rect 17880 14482 17908 17575
rect 18052 17536 18104 17542
rect 18052 17478 18104 17484
rect 18064 17338 18092 17478
rect 18052 17332 18104 17338
rect 18052 17274 18104 17280
rect 18064 16998 18092 17274
rect 18052 16992 18104 16998
rect 18052 16934 18104 16940
rect 18144 16108 18196 16114
rect 18144 16050 18196 16056
rect 17960 15904 18012 15910
rect 17960 15846 18012 15852
rect 17972 15570 18000 15846
rect 18156 15706 18184 16050
rect 18144 15700 18196 15706
rect 18144 15642 18196 15648
rect 17960 15564 18012 15570
rect 17960 15506 18012 15512
rect 17868 14476 17920 14482
rect 17868 14418 17920 14424
rect 17880 14074 17908 14418
rect 17868 14068 17920 14074
rect 17868 14010 17920 14016
rect 18052 13864 18104 13870
rect 18052 13806 18104 13812
rect 17684 13524 17736 13530
rect 17736 13484 17908 13512
rect 17684 13466 17736 13472
rect 17592 13320 17644 13326
rect 17592 13262 17644 13268
rect 17500 12912 17552 12918
rect 17500 12854 17552 12860
rect 17408 12640 17460 12646
rect 17408 12582 17460 12588
rect 16956 12540 17252 12560
rect 17012 12538 17036 12540
rect 17092 12538 17116 12540
rect 17172 12538 17196 12540
rect 17034 12486 17036 12538
rect 17098 12486 17110 12538
rect 17172 12486 17174 12538
rect 17012 12484 17036 12486
rect 17092 12484 17116 12486
rect 17172 12484 17196 12486
rect 16956 12464 17252 12484
rect 17420 12442 17448 12582
rect 17408 12436 17460 12442
rect 17408 12378 17460 12384
rect 16764 12300 16816 12306
rect 16764 12242 16816 12248
rect 16856 11688 16908 11694
rect 16856 11630 16908 11636
rect 16580 11008 16632 11014
rect 16580 10950 16632 10956
rect 16592 9586 16620 10950
rect 16868 10810 16896 11630
rect 16956 11452 17252 11472
rect 17012 11450 17036 11452
rect 17092 11450 17116 11452
rect 17172 11450 17196 11452
rect 17034 11398 17036 11450
rect 17098 11398 17110 11450
rect 17172 11398 17174 11450
rect 17012 11396 17036 11398
rect 17092 11396 17116 11398
rect 17172 11396 17196 11398
rect 16956 11376 17252 11396
rect 16856 10804 16908 10810
rect 16856 10746 16908 10752
rect 16764 10668 16816 10674
rect 16764 10610 16816 10616
rect 16672 10464 16724 10470
rect 16776 10452 16804 10610
rect 16868 10606 16896 10746
rect 16856 10600 16908 10606
rect 16856 10542 16908 10548
rect 16776 10424 16896 10452
rect 16672 10406 16724 10412
rect 16684 10062 16712 10406
rect 16672 10056 16724 10062
rect 16672 9998 16724 10004
rect 16580 9580 16632 9586
rect 16580 9522 16632 9528
rect 16592 9178 16620 9522
rect 16580 9172 16632 9178
rect 16580 9114 16632 9120
rect 16764 9104 16816 9110
rect 16764 9046 16816 9052
rect 16776 8634 16804 9046
rect 16764 8628 16816 8634
rect 16764 8570 16816 8576
rect 16776 8022 16804 8570
rect 16764 8016 16816 8022
rect 16764 7958 16816 7964
rect 16486 7848 16542 7857
rect 16486 7783 16542 7792
rect 16776 7546 16804 7958
rect 16764 7540 16816 7546
rect 16764 7482 16816 7488
rect 16120 7200 16172 7206
rect 16120 7142 16172 7148
rect 16132 6798 16160 7142
rect 16212 6928 16264 6934
rect 16212 6870 16264 6876
rect 16120 6792 16172 6798
rect 16120 6734 16172 6740
rect 15936 6384 15988 6390
rect 15936 6326 15988 6332
rect 15844 6180 15896 6186
rect 15844 6122 15896 6128
rect 15856 5030 15884 6122
rect 15948 5778 15976 6326
rect 16132 5914 16160 6734
rect 16224 6458 16252 6870
rect 16304 6792 16356 6798
rect 16304 6734 16356 6740
rect 16212 6452 16264 6458
rect 16212 6394 16264 6400
rect 16316 6322 16344 6734
rect 16304 6316 16356 6322
rect 16304 6258 16356 6264
rect 16488 6316 16540 6322
rect 16488 6258 16540 6264
rect 16120 5908 16172 5914
rect 16120 5850 16172 5856
rect 16500 5778 16528 6258
rect 16868 6254 16896 10424
rect 16956 10364 17252 10384
rect 17012 10362 17036 10364
rect 17092 10362 17116 10364
rect 17172 10362 17196 10364
rect 17034 10310 17036 10362
rect 17098 10310 17110 10362
rect 17172 10310 17174 10362
rect 17012 10308 17036 10310
rect 17092 10308 17116 10310
rect 17172 10308 17196 10310
rect 16956 10288 17252 10308
rect 17316 10192 17368 10198
rect 17316 10134 17368 10140
rect 17328 9722 17356 10134
rect 17316 9716 17368 9722
rect 17316 9658 17368 9664
rect 17316 9444 17368 9450
rect 17316 9386 17368 9392
rect 16956 9276 17252 9296
rect 17012 9274 17036 9276
rect 17092 9274 17116 9276
rect 17172 9274 17196 9276
rect 17034 9222 17036 9274
rect 17098 9222 17110 9274
rect 17172 9222 17174 9274
rect 17012 9220 17036 9222
rect 17092 9220 17116 9222
rect 17172 9220 17196 9222
rect 16956 9200 17252 9220
rect 16948 8968 17000 8974
rect 16948 8910 17000 8916
rect 16960 8634 16988 8910
rect 16948 8628 17000 8634
rect 16948 8570 17000 8576
rect 17328 8362 17356 9386
rect 17420 9042 17448 12378
rect 17512 11218 17540 12854
rect 17776 12368 17828 12374
rect 17776 12310 17828 12316
rect 17684 12232 17736 12238
rect 17684 12174 17736 12180
rect 17696 11354 17724 12174
rect 17788 11898 17816 12310
rect 17776 11892 17828 11898
rect 17776 11834 17828 11840
rect 17684 11348 17736 11354
rect 17684 11290 17736 11296
rect 17500 11212 17552 11218
rect 17500 11154 17552 11160
rect 17512 10674 17540 11154
rect 17696 10810 17724 11290
rect 17684 10804 17736 10810
rect 17684 10746 17736 10752
rect 17500 10668 17552 10674
rect 17500 10610 17552 10616
rect 17880 10606 17908 13484
rect 17960 13252 18012 13258
rect 17960 13194 18012 13200
rect 17972 12918 18000 13194
rect 17960 12912 18012 12918
rect 17960 12854 18012 12860
rect 17972 12238 18000 12854
rect 17960 12232 18012 12238
rect 17960 12174 18012 12180
rect 17868 10600 17920 10606
rect 17868 10542 17920 10548
rect 17500 10464 17552 10470
rect 17500 10406 17552 10412
rect 17408 9036 17460 9042
rect 17408 8978 17460 8984
rect 17316 8356 17368 8362
rect 17316 8298 17368 8304
rect 16956 8188 17252 8208
rect 17012 8186 17036 8188
rect 17092 8186 17116 8188
rect 17172 8186 17196 8188
rect 17034 8134 17036 8186
rect 17098 8134 17110 8186
rect 17172 8134 17174 8186
rect 17012 8132 17036 8134
rect 17092 8132 17116 8134
rect 17172 8132 17196 8134
rect 16956 8112 17252 8132
rect 17328 8022 17356 8298
rect 17408 8288 17460 8294
rect 17408 8230 17460 8236
rect 17316 8016 17368 8022
rect 17316 7958 17368 7964
rect 17040 7880 17092 7886
rect 17040 7822 17092 7828
rect 17052 7546 17080 7822
rect 17040 7540 17092 7546
rect 17040 7482 17092 7488
rect 16956 7100 17252 7120
rect 17012 7098 17036 7100
rect 17092 7098 17116 7100
rect 17172 7098 17196 7100
rect 17034 7046 17036 7098
rect 17098 7046 17110 7098
rect 17172 7046 17174 7098
rect 17012 7044 17036 7046
rect 17092 7044 17116 7046
rect 17172 7044 17196 7046
rect 16956 7024 17252 7044
rect 16856 6248 16908 6254
rect 16856 6190 16908 6196
rect 16956 6012 17252 6032
rect 17012 6010 17036 6012
rect 17092 6010 17116 6012
rect 17172 6010 17196 6012
rect 17034 5958 17036 6010
rect 17098 5958 17110 6010
rect 17172 5958 17174 6010
rect 17012 5956 17036 5958
rect 17092 5956 17116 5958
rect 17172 5956 17196 5958
rect 16956 5936 17252 5956
rect 15936 5772 15988 5778
rect 15936 5714 15988 5720
rect 16488 5772 16540 5778
rect 16488 5714 16540 5720
rect 15948 5370 15976 5714
rect 16500 5370 16528 5714
rect 16672 5704 16724 5710
rect 16672 5646 16724 5652
rect 15936 5364 15988 5370
rect 15936 5306 15988 5312
rect 16488 5364 16540 5370
rect 16488 5306 16540 5312
rect 16396 5092 16448 5098
rect 16396 5034 16448 5040
rect 15844 5024 15896 5030
rect 15844 4966 15896 4972
rect 15856 4826 15884 4966
rect 16408 4826 16436 5034
rect 15844 4820 15896 4826
rect 15844 4762 15896 4768
rect 16396 4820 16448 4826
rect 16396 4762 16448 4768
rect 15476 4616 15528 4622
rect 15476 4558 15528 4564
rect 15488 4010 15516 4558
rect 15856 4282 15884 4762
rect 16500 4282 16528 5306
rect 16684 5234 16712 5646
rect 16948 5568 17000 5574
rect 16948 5510 17000 5516
rect 16960 5302 16988 5510
rect 16948 5296 17000 5302
rect 16948 5238 17000 5244
rect 16672 5228 16724 5234
rect 16672 5170 16724 5176
rect 16956 4924 17252 4944
rect 17012 4922 17036 4924
rect 17092 4922 17116 4924
rect 17172 4922 17196 4924
rect 17034 4870 17036 4922
rect 17098 4870 17110 4922
rect 17172 4870 17174 4922
rect 17012 4868 17036 4870
rect 17092 4868 17116 4870
rect 17172 4868 17196 4870
rect 16956 4848 17252 4868
rect 15844 4276 15896 4282
rect 15844 4218 15896 4224
rect 16488 4276 16540 4282
rect 16488 4218 16540 4224
rect 16500 4154 16528 4218
rect 16500 4126 16620 4154
rect 16592 4078 16620 4126
rect 16580 4072 16632 4078
rect 16580 4014 16632 4020
rect 15476 4004 15528 4010
rect 15476 3946 15528 3952
rect 16956 3836 17252 3856
rect 17012 3834 17036 3836
rect 17092 3834 17116 3836
rect 17172 3834 17196 3836
rect 17034 3782 17036 3834
rect 17098 3782 17110 3834
rect 17172 3782 17174 3834
rect 17012 3780 17036 3782
rect 17092 3780 17116 3782
rect 17172 3780 17196 3782
rect 16956 3760 17252 3780
rect 16956 2748 17252 2768
rect 17012 2746 17036 2748
rect 17092 2746 17116 2748
rect 17172 2746 17196 2748
rect 17034 2694 17036 2746
rect 17098 2694 17110 2746
rect 17172 2694 17174 2746
rect 17012 2692 17036 2694
rect 17092 2692 17116 2694
rect 17172 2692 17196 2694
rect 16956 2672 17252 2692
rect 17132 2508 17184 2514
rect 17132 2450 17184 2456
rect 14096 2304 14148 2310
rect 14096 2246 14148 2252
rect 15292 2304 15344 2310
rect 15292 2246 15344 2252
rect 12956 2204 13252 2224
rect 13012 2202 13036 2204
rect 13092 2202 13116 2204
rect 13172 2202 13196 2204
rect 13034 2150 13036 2202
rect 13098 2150 13110 2202
rect 13172 2150 13174 2202
rect 13012 2148 13036 2150
rect 13092 2148 13116 2150
rect 13172 2148 13196 2150
rect 12956 2128 13252 2148
rect 11978 54 12112 82
rect 13818 82 13874 480
rect 14108 82 14136 2246
rect 13818 54 14136 82
rect 15304 82 15332 2246
rect 17144 1601 17172 2450
rect 17130 1592 17186 1601
rect 17130 1527 17186 1536
rect 15658 82 15714 480
rect 15304 54 15714 82
rect 17420 82 17448 8230
rect 17512 7177 17540 10406
rect 17592 10056 17644 10062
rect 17592 9998 17644 10004
rect 17604 9178 17632 9998
rect 17776 9988 17828 9994
rect 17776 9930 17828 9936
rect 17592 9172 17644 9178
rect 17592 9114 17644 9120
rect 17788 8906 17816 9930
rect 17776 8900 17828 8906
rect 17776 8842 17828 8848
rect 18064 8430 18092 13806
rect 18144 11212 18196 11218
rect 18144 11154 18196 11160
rect 18156 10470 18184 11154
rect 18144 10464 18196 10470
rect 18144 10406 18196 10412
rect 18156 9926 18184 10406
rect 18144 9920 18196 9926
rect 18144 9862 18196 9868
rect 18156 9654 18184 9862
rect 18144 9648 18196 9654
rect 18144 9590 18196 9596
rect 18248 9489 18276 20334
rect 18984 20058 19012 23582
rect 20640 23582 20958 23610
rect 19982 22672 20038 22681
rect 19982 22607 20038 22616
rect 18972 20052 19024 20058
rect 18972 19994 19024 20000
rect 18788 18624 18840 18630
rect 18788 18566 18840 18572
rect 18800 18290 18828 18566
rect 18788 18284 18840 18290
rect 18788 18226 18840 18232
rect 18420 18148 18472 18154
rect 18420 18090 18472 18096
rect 18432 17542 18460 18090
rect 18800 17882 18828 18226
rect 18788 17876 18840 17882
rect 18788 17818 18840 17824
rect 18880 17740 18932 17746
rect 18880 17682 18932 17688
rect 19064 17740 19116 17746
rect 19064 17682 19116 17688
rect 18892 17649 18920 17682
rect 18878 17640 18934 17649
rect 18878 17575 18934 17584
rect 18420 17536 18472 17542
rect 18420 17478 18472 17484
rect 18432 17202 18460 17478
rect 18892 17338 18920 17575
rect 18880 17332 18932 17338
rect 18880 17274 18932 17280
rect 18420 17196 18472 17202
rect 18420 17138 18472 17144
rect 18328 16448 18380 16454
rect 18328 16390 18380 16396
rect 18340 16114 18368 16390
rect 18432 16114 18460 17138
rect 19076 16998 19104 17682
rect 19708 17536 19760 17542
rect 19708 17478 19760 17484
rect 19720 17066 19748 17478
rect 19708 17060 19760 17066
rect 19708 17002 19760 17008
rect 19800 17060 19852 17066
rect 19800 17002 19852 17008
rect 19064 16992 19116 16998
rect 19064 16934 19116 16940
rect 18972 16720 19024 16726
rect 18972 16662 19024 16668
rect 18984 16250 19012 16662
rect 19076 16658 19104 16934
rect 19064 16652 19116 16658
rect 19064 16594 19116 16600
rect 19432 16584 19484 16590
rect 19432 16526 19484 16532
rect 19444 16250 19472 16526
rect 18972 16244 19024 16250
rect 18972 16186 19024 16192
rect 19432 16244 19484 16250
rect 19432 16186 19484 16192
rect 19720 16182 19748 17002
rect 19812 16794 19840 17002
rect 19800 16788 19852 16794
rect 19800 16730 19852 16736
rect 19708 16176 19760 16182
rect 19708 16118 19760 16124
rect 18328 16108 18380 16114
rect 18328 16050 18380 16056
rect 18420 16108 18472 16114
rect 18420 16050 18472 16056
rect 18328 15972 18380 15978
rect 18328 15914 18380 15920
rect 18340 15162 18368 15914
rect 18328 15156 18380 15162
rect 18328 15098 18380 15104
rect 18432 14550 18460 16050
rect 18512 15972 18564 15978
rect 18512 15914 18564 15920
rect 18524 15638 18552 15914
rect 19720 15638 19748 16118
rect 18512 15632 18564 15638
rect 18512 15574 18564 15580
rect 19708 15632 19760 15638
rect 19708 15574 19760 15580
rect 18696 15496 18748 15502
rect 18696 15438 18748 15444
rect 18604 14952 18656 14958
rect 18604 14894 18656 14900
rect 18512 14612 18564 14618
rect 18512 14554 18564 14560
rect 18420 14544 18472 14550
rect 18420 14486 18472 14492
rect 18524 13530 18552 14554
rect 18616 14550 18644 14894
rect 18708 14822 18736 15438
rect 19524 15360 19576 15366
rect 19524 15302 19576 15308
rect 19536 14958 19564 15302
rect 19524 14952 19576 14958
rect 19524 14894 19576 14900
rect 18696 14816 18748 14822
rect 18696 14758 18748 14764
rect 19432 14816 19484 14822
rect 19432 14758 19484 14764
rect 18708 14618 18736 14758
rect 18696 14612 18748 14618
rect 18696 14554 18748 14560
rect 18604 14544 18656 14550
rect 18604 14486 18656 14492
rect 19064 14272 19116 14278
rect 19064 14214 19116 14220
rect 19076 13938 19104 14214
rect 19156 14068 19208 14074
rect 19156 14010 19208 14016
rect 18788 13932 18840 13938
rect 18788 13874 18840 13880
rect 19064 13932 19116 13938
rect 19064 13874 19116 13880
rect 18512 13524 18564 13530
rect 18512 13466 18564 13472
rect 18524 12782 18552 13466
rect 18800 12850 18828 13874
rect 18880 13728 18932 13734
rect 18880 13670 18932 13676
rect 18788 12844 18840 12850
rect 18788 12786 18840 12792
rect 18512 12776 18564 12782
rect 18512 12718 18564 12724
rect 18892 12646 18920 13670
rect 19064 13320 19116 13326
rect 19064 13262 19116 13268
rect 18880 12640 18932 12646
rect 18880 12582 18932 12588
rect 18420 12096 18472 12102
rect 18420 12038 18472 12044
rect 18432 11694 18460 12038
rect 18420 11688 18472 11694
rect 18420 11630 18472 11636
rect 18432 11286 18460 11630
rect 18892 11626 18920 12582
rect 19076 12442 19104 13262
rect 19064 12436 19116 12442
rect 19064 12378 19116 12384
rect 18880 11620 18932 11626
rect 18880 11562 18932 11568
rect 18420 11280 18472 11286
rect 18420 11222 18472 11228
rect 18892 10198 18920 11562
rect 18880 10192 18932 10198
rect 18880 10134 18932 10140
rect 18788 10056 18840 10062
rect 18788 9998 18840 10004
rect 18234 9480 18290 9489
rect 18800 9450 18828 9998
rect 18892 9722 18920 10134
rect 18880 9716 18932 9722
rect 18880 9658 18932 9664
rect 18234 9415 18290 9424
rect 18604 9444 18656 9450
rect 18604 9386 18656 9392
rect 18788 9444 18840 9450
rect 18788 9386 18840 9392
rect 18616 9042 18644 9386
rect 18800 9178 18828 9386
rect 18788 9172 18840 9178
rect 18788 9114 18840 9120
rect 18144 9036 18196 9042
rect 18144 8978 18196 8984
rect 18604 9036 18656 9042
rect 18604 8978 18656 8984
rect 18052 8424 18104 8430
rect 18052 8366 18104 8372
rect 17868 8288 17920 8294
rect 17868 8230 17920 8236
rect 17880 7886 17908 8230
rect 17868 7880 17920 7886
rect 17868 7822 17920 7828
rect 17958 7848 18014 7857
rect 17958 7783 18014 7792
rect 17972 7342 18000 7783
rect 17960 7336 18012 7342
rect 17960 7278 18012 7284
rect 17498 7168 17554 7177
rect 17498 7103 17554 7112
rect 17960 6860 18012 6866
rect 17960 6802 18012 6808
rect 17592 6792 17644 6798
rect 17592 6734 17644 6740
rect 17604 5710 17632 6734
rect 17972 6390 18000 6802
rect 17960 6384 18012 6390
rect 17960 6326 18012 6332
rect 17868 6248 17920 6254
rect 18064 6236 18092 8366
rect 18156 8090 18184 8978
rect 18616 8634 18644 8978
rect 19064 8968 19116 8974
rect 19064 8910 19116 8916
rect 18604 8628 18656 8634
rect 18604 8570 18656 8576
rect 18144 8084 18196 8090
rect 18144 8026 18196 8032
rect 18616 6866 18644 8570
rect 19076 8498 19104 8910
rect 19064 8492 19116 8498
rect 19064 8434 19116 8440
rect 18972 7880 19024 7886
rect 18972 7822 19024 7828
rect 18984 7410 19012 7822
rect 18972 7404 19024 7410
rect 18972 7346 19024 7352
rect 18984 6934 19012 7346
rect 19064 7200 19116 7206
rect 19064 7142 19116 7148
rect 18972 6928 19024 6934
rect 18972 6870 19024 6876
rect 18604 6860 18656 6866
rect 18604 6802 18656 6808
rect 18616 6458 18644 6802
rect 18972 6656 19024 6662
rect 19076 6644 19104 7142
rect 19168 7002 19196 14010
rect 19444 13870 19472 14758
rect 19432 13864 19484 13870
rect 19352 13824 19432 13852
rect 19352 13530 19380 13824
rect 19432 13806 19484 13812
rect 19340 13524 19392 13530
rect 19340 13466 19392 13472
rect 19800 12708 19852 12714
rect 19800 12650 19852 12656
rect 19432 12640 19484 12646
rect 19432 12582 19484 12588
rect 19444 12374 19472 12582
rect 19812 12442 19840 12650
rect 19800 12436 19852 12442
rect 19800 12378 19852 12384
rect 19432 12368 19484 12374
rect 19432 12310 19484 12316
rect 19444 11898 19472 12310
rect 19432 11892 19484 11898
rect 19432 11834 19484 11840
rect 19432 11212 19484 11218
rect 19432 11154 19484 11160
rect 19444 10810 19472 11154
rect 19616 11008 19668 11014
rect 19616 10950 19668 10956
rect 19800 11008 19852 11014
rect 19800 10950 19852 10956
rect 19432 10804 19484 10810
rect 19432 10746 19484 10752
rect 19628 10674 19656 10950
rect 19616 10668 19668 10674
rect 19616 10610 19668 10616
rect 19628 10266 19656 10610
rect 19812 10538 19840 10950
rect 19892 10668 19944 10674
rect 19892 10610 19944 10616
rect 19800 10532 19852 10538
rect 19800 10474 19852 10480
rect 19616 10260 19668 10266
rect 19616 10202 19668 10208
rect 19812 10130 19840 10474
rect 19800 10124 19852 10130
rect 19800 10066 19852 10072
rect 19812 9722 19840 10066
rect 19800 9716 19852 9722
rect 19800 9658 19852 9664
rect 19812 9450 19840 9658
rect 19800 9444 19852 9450
rect 19800 9386 19852 9392
rect 19904 8362 19932 10610
rect 19996 9178 20024 22607
rect 20640 20602 20668 23582
rect 20902 23520 20958 23582
rect 22664 23582 22982 23610
rect 20956 21788 21252 21808
rect 21012 21786 21036 21788
rect 21092 21786 21116 21788
rect 21172 21786 21196 21788
rect 21034 21734 21036 21786
rect 21098 21734 21110 21786
rect 21172 21734 21174 21786
rect 21012 21732 21036 21734
rect 21092 21732 21116 21734
rect 21172 21732 21196 21734
rect 20956 21712 21252 21732
rect 22006 21176 22062 21185
rect 22006 21111 22062 21120
rect 20956 20700 21252 20720
rect 21012 20698 21036 20700
rect 21092 20698 21116 20700
rect 21172 20698 21196 20700
rect 21034 20646 21036 20698
rect 21098 20646 21110 20698
rect 21172 20646 21174 20698
rect 21012 20644 21036 20646
rect 21092 20644 21116 20646
rect 21172 20644 21196 20646
rect 20956 20624 21252 20644
rect 20628 20596 20680 20602
rect 20628 20538 20680 20544
rect 21270 19816 21326 19825
rect 21270 19751 21326 19760
rect 20956 19612 21252 19632
rect 21012 19610 21036 19612
rect 21092 19610 21116 19612
rect 21172 19610 21196 19612
rect 21034 19558 21036 19610
rect 21098 19558 21110 19610
rect 21172 19558 21174 19610
rect 21012 19556 21036 19558
rect 21092 19556 21116 19558
rect 21172 19556 21196 19558
rect 20956 19536 21252 19556
rect 20812 19304 20864 19310
rect 20812 19246 20864 19252
rect 20352 18760 20404 18766
rect 20352 18702 20404 18708
rect 20364 18426 20392 18702
rect 20352 18420 20404 18426
rect 20352 18362 20404 18368
rect 20824 18290 20852 19246
rect 21284 18970 21312 19751
rect 21272 18964 21324 18970
rect 21272 18906 21324 18912
rect 21548 18828 21600 18834
rect 21548 18770 21600 18776
rect 20956 18524 21252 18544
rect 21012 18522 21036 18524
rect 21092 18522 21116 18524
rect 21172 18522 21196 18524
rect 21034 18470 21036 18522
rect 21098 18470 21110 18522
rect 21172 18470 21174 18522
rect 21012 18468 21036 18470
rect 21092 18468 21116 18470
rect 21172 18468 21196 18470
rect 20956 18448 21252 18468
rect 20812 18284 20864 18290
rect 20812 18226 20864 18232
rect 20536 18080 20588 18086
rect 20536 18022 20588 18028
rect 20548 17882 20576 18022
rect 20536 17876 20588 17882
rect 20536 17818 20588 17824
rect 20720 17808 20772 17814
rect 20720 17750 20772 17756
rect 20732 17338 20760 17750
rect 20720 17332 20772 17338
rect 20720 17274 20772 17280
rect 20824 17202 20852 18226
rect 21086 18184 21142 18193
rect 21086 18119 21142 18128
rect 21100 17882 21128 18119
rect 21560 18086 21588 18770
rect 21548 18080 21600 18086
rect 21548 18022 21600 18028
rect 21088 17876 21140 17882
rect 21088 17818 21140 17824
rect 20956 17436 21252 17456
rect 21012 17434 21036 17436
rect 21092 17434 21116 17436
rect 21172 17434 21196 17436
rect 21034 17382 21036 17434
rect 21098 17382 21110 17434
rect 21172 17382 21174 17434
rect 21012 17380 21036 17382
rect 21092 17380 21116 17382
rect 21172 17380 21196 17382
rect 20956 17360 21252 17380
rect 20812 17196 20864 17202
rect 20812 17138 20864 17144
rect 21086 16688 21142 16697
rect 20812 16652 20864 16658
rect 21086 16623 21142 16632
rect 20812 16594 20864 16600
rect 20824 15978 20852 16594
rect 21100 16522 21128 16623
rect 21088 16516 21140 16522
rect 21088 16458 21140 16464
rect 20956 16348 21252 16368
rect 21012 16346 21036 16348
rect 21092 16346 21116 16348
rect 21172 16346 21196 16348
rect 21034 16294 21036 16346
rect 21098 16294 21110 16346
rect 21172 16294 21174 16346
rect 21012 16292 21036 16294
rect 21092 16292 21116 16294
rect 21172 16292 21196 16294
rect 20956 16272 21252 16292
rect 20812 15972 20864 15978
rect 20812 15914 20864 15920
rect 20812 15564 20864 15570
rect 20812 15506 20864 15512
rect 20824 15162 20852 15506
rect 20956 15260 21252 15280
rect 21012 15258 21036 15260
rect 21092 15258 21116 15260
rect 21172 15258 21196 15260
rect 21034 15206 21036 15258
rect 21098 15206 21110 15258
rect 21172 15206 21174 15258
rect 21012 15204 21036 15206
rect 21092 15204 21116 15206
rect 21172 15204 21196 15206
rect 20956 15184 21252 15204
rect 20812 15156 20864 15162
rect 20812 15098 20864 15104
rect 20444 14816 20496 14822
rect 20444 14758 20496 14764
rect 20456 14618 20484 14758
rect 20444 14612 20496 14618
rect 20444 14554 20496 14560
rect 20720 14544 20772 14550
rect 20720 14486 20772 14492
rect 20352 14476 20404 14482
rect 20352 14418 20404 14424
rect 20364 13977 20392 14418
rect 20732 14074 20760 14486
rect 20824 14414 20852 15098
rect 20996 14816 21048 14822
rect 20996 14758 21048 14764
rect 21008 14550 21036 14758
rect 20996 14544 21048 14550
rect 20996 14486 21048 14492
rect 20812 14408 20864 14414
rect 20812 14350 20864 14356
rect 21272 14408 21324 14414
rect 21272 14350 21324 14356
rect 20956 14172 21252 14192
rect 21012 14170 21036 14172
rect 21092 14170 21116 14172
rect 21172 14170 21196 14172
rect 21034 14118 21036 14170
rect 21098 14118 21110 14170
rect 21172 14118 21174 14170
rect 21012 14116 21036 14118
rect 21092 14116 21116 14118
rect 21172 14116 21196 14118
rect 20956 14096 21252 14116
rect 20720 14068 20772 14074
rect 20720 14010 20772 14016
rect 20350 13968 20406 13977
rect 21284 13938 21312 14350
rect 20350 13903 20352 13912
rect 20404 13903 20406 13912
rect 21272 13932 21324 13938
rect 20352 13874 20404 13880
rect 21272 13874 21324 13880
rect 20364 12306 20392 13874
rect 20628 13796 20680 13802
rect 20628 13738 20680 13744
rect 20996 13796 21048 13802
rect 20996 13738 21048 13744
rect 20640 13190 20668 13738
rect 20812 13728 20864 13734
rect 20812 13670 20864 13676
rect 20628 13184 20680 13190
rect 20628 13126 20680 13132
rect 20352 12300 20404 12306
rect 20352 12242 20404 12248
rect 20076 12232 20128 12238
rect 20076 12174 20128 12180
rect 20088 11898 20116 12174
rect 20076 11892 20128 11898
rect 20076 11834 20128 11840
rect 20364 11218 20392 12242
rect 20640 12170 20668 13126
rect 20824 12986 20852 13670
rect 21008 13530 21036 13738
rect 21088 13728 21140 13734
rect 21088 13670 21140 13676
rect 20996 13524 21048 13530
rect 20996 13466 21048 13472
rect 21100 13462 21128 13670
rect 21088 13456 21140 13462
rect 21088 13398 21140 13404
rect 21284 13326 21312 13874
rect 21272 13320 21324 13326
rect 21272 13262 21324 13268
rect 21364 13252 21416 13258
rect 21364 13194 21416 13200
rect 20956 13084 21252 13104
rect 21012 13082 21036 13084
rect 21092 13082 21116 13084
rect 21172 13082 21196 13084
rect 21034 13030 21036 13082
rect 21098 13030 21110 13082
rect 21172 13030 21174 13082
rect 21012 13028 21036 13030
rect 21092 13028 21116 13030
rect 21172 13028 21196 13030
rect 20956 13008 21252 13028
rect 20812 12980 20864 12986
rect 20812 12922 20864 12928
rect 21376 12714 21404 13194
rect 21364 12708 21416 12714
rect 21364 12650 21416 12656
rect 21376 12442 21404 12650
rect 21364 12436 21416 12442
rect 21364 12378 21416 12384
rect 20812 12300 20864 12306
rect 20812 12242 20864 12248
rect 20628 12164 20680 12170
rect 20628 12106 20680 12112
rect 20824 11898 20852 12242
rect 20956 11996 21252 12016
rect 21012 11994 21036 11996
rect 21092 11994 21116 11996
rect 21172 11994 21196 11996
rect 21034 11942 21036 11994
rect 21098 11942 21110 11994
rect 21172 11942 21174 11994
rect 21012 11940 21036 11942
rect 21092 11940 21116 11942
rect 21172 11940 21196 11942
rect 20956 11920 21252 11940
rect 20812 11892 20864 11898
rect 20812 11834 20864 11840
rect 20718 11792 20774 11801
rect 20718 11727 20774 11736
rect 20732 11694 20760 11727
rect 21560 11694 21588 18022
rect 22020 15706 22048 21111
rect 22664 19514 22692 23582
rect 22926 23520 22982 23582
rect 22652 19508 22704 19514
rect 22652 19450 22704 19456
rect 22008 15700 22060 15706
rect 22008 15642 22060 15648
rect 21914 15192 21970 15201
rect 21914 15127 21970 15136
rect 21928 13705 21956 15127
rect 22192 14544 22244 14550
rect 22192 14486 22244 14492
rect 22204 14074 22232 14486
rect 22192 14068 22244 14074
rect 22192 14010 22244 14016
rect 21914 13696 21970 13705
rect 21914 13631 21970 13640
rect 21928 12986 21956 13631
rect 21916 12980 21968 12986
rect 21916 12922 21968 12928
rect 21928 12782 21956 12922
rect 23572 12912 23624 12918
rect 23572 12854 23624 12860
rect 21916 12776 21968 12782
rect 23584 12753 23612 12854
rect 21916 12718 21968 12724
rect 23570 12744 23626 12753
rect 23570 12679 23626 12688
rect 20720 11688 20772 11694
rect 20720 11630 20772 11636
rect 21548 11688 21600 11694
rect 21548 11630 21600 11636
rect 20352 11212 20404 11218
rect 20352 11154 20404 11160
rect 20260 9920 20312 9926
rect 20260 9862 20312 9868
rect 20168 9580 20220 9586
rect 20272 9568 20300 9862
rect 20364 9586 20392 11154
rect 20732 10130 20760 11630
rect 21270 11248 21326 11257
rect 21270 11183 21326 11192
rect 20956 10908 21252 10928
rect 21012 10906 21036 10908
rect 21092 10906 21116 10908
rect 21172 10906 21196 10908
rect 21034 10854 21036 10906
rect 21098 10854 21110 10906
rect 21172 10854 21174 10906
rect 21012 10852 21036 10854
rect 21092 10852 21116 10854
rect 21172 10852 21196 10854
rect 20956 10832 21252 10852
rect 21284 10810 21312 11183
rect 21272 10804 21324 10810
rect 21272 10746 21324 10752
rect 20720 10124 20772 10130
rect 20720 10066 20772 10072
rect 20732 9722 20760 10066
rect 20956 9820 21252 9840
rect 21012 9818 21036 9820
rect 21092 9818 21116 9820
rect 21172 9818 21196 9820
rect 21034 9766 21036 9818
rect 21098 9766 21110 9818
rect 21172 9766 21174 9818
rect 21012 9764 21036 9766
rect 21092 9764 21116 9766
rect 21172 9764 21196 9766
rect 20956 9744 21252 9764
rect 21362 9752 21418 9761
rect 20720 9716 20772 9722
rect 21362 9687 21418 9696
rect 20720 9658 20772 9664
rect 21376 9654 21404 9687
rect 21364 9648 21416 9654
rect 21364 9590 21416 9596
rect 20220 9540 20300 9568
rect 20168 9522 20220 9528
rect 20272 9178 20300 9540
rect 20352 9580 20404 9586
rect 20352 9522 20404 9528
rect 20444 9444 20496 9450
rect 20444 9386 20496 9392
rect 19984 9172 20036 9178
rect 19984 9114 20036 9120
rect 20260 9172 20312 9178
rect 20260 9114 20312 9120
rect 20352 9104 20404 9110
rect 20352 9046 20404 9052
rect 20168 9036 20220 9042
rect 20168 8978 20220 8984
rect 20180 8498 20208 8978
rect 20364 8634 20392 9046
rect 20456 8974 20484 9386
rect 20444 8968 20496 8974
rect 20444 8910 20496 8916
rect 21272 8968 21324 8974
rect 21272 8910 21324 8916
rect 20956 8732 21252 8752
rect 21012 8730 21036 8732
rect 21092 8730 21116 8732
rect 21172 8730 21196 8732
rect 21034 8678 21036 8730
rect 21098 8678 21110 8730
rect 21172 8678 21174 8730
rect 21012 8676 21036 8678
rect 21092 8676 21116 8678
rect 21172 8676 21196 8678
rect 20956 8656 21252 8676
rect 20352 8628 20404 8634
rect 20352 8570 20404 8576
rect 20904 8560 20956 8566
rect 20904 8502 20956 8508
rect 20168 8492 20220 8498
rect 20168 8434 20220 8440
rect 19892 8356 19944 8362
rect 19892 8298 19944 8304
rect 19248 8288 19300 8294
rect 19248 8230 19300 8236
rect 19260 8022 19288 8230
rect 20180 8022 20208 8434
rect 20916 8362 20944 8502
rect 21284 8498 21312 8910
rect 22192 8900 22244 8906
rect 22192 8842 22244 8848
rect 22204 8634 22232 8842
rect 22192 8628 22244 8634
rect 22192 8570 22244 8576
rect 21272 8492 21324 8498
rect 21272 8434 21324 8440
rect 20904 8356 20956 8362
rect 20904 8298 20956 8304
rect 20628 8288 20680 8294
rect 20628 8230 20680 8236
rect 20640 8090 20668 8230
rect 20628 8084 20680 8090
rect 20628 8026 20680 8032
rect 19248 8016 19300 8022
rect 19248 7958 19300 7964
rect 20168 8016 20220 8022
rect 20168 7958 20220 7964
rect 20260 8016 20312 8022
rect 20260 7958 20312 7964
rect 20272 7546 20300 7958
rect 21284 7886 21312 8434
rect 23570 8256 23626 8265
rect 23570 8191 23626 8200
rect 21456 8016 21508 8022
rect 21456 7958 21508 7964
rect 20812 7880 20864 7886
rect 20812 7822 20864 7828
rect 21272 7880 21324 7886
rect 21272 7822 21324 7828
rect 20824 7546 20852 7822
rect 20956 7644 21252 7664
rect 21012 7642 21036 7644
rect 21092 7642 21116 7644
rect 21172 7642 21196 7644
rect 21034 7590 21036 7642
rect 21098 7590 21110 7642
rect 21172 7590 21174 7642
rect 21012 7588 21036 7590
rect 21092 7588 21116 7590
rect 21172 7588 21196 7590
rect 20956 7568 21252 7588
rect 21468 7546 21496 7958
rect 20260 7540 20312 7546
rect 20260 7482 20312 7488
rect 20812 7540 20864 7546
rect 20812 7482 20864 7488
rect 21456 7540 21508 7546
rect 21456 7482 21508 7488
rect 20168 7336 20220 7342
rect 23584 7313 23612 8191
rect 20168 7278 20220 7284
rect 23570 7304 23626 7313
rect 19156 6996 19208 7002
rect 19156 6938 19208 6944
rect 19616 6996 19668 7002
rect 19616 6938 19668 6944
rect 19024 6616 19104 6644
rect 18972 6598 19024 6604
rect 18604 6452 18656 6458
rect 18604 6394 18656 6400
rect 17868 6190 17920 6196
rect 17972 6208 18092 6236
rect 17880 5914 17908 6190
rect 17868 5908 17920 5914
rect 17868 5850 17920 5856
rect 17684 5840 17736 5846
rect 17684 5782 17736 5788
rect 17592 5704 17644 5710
rect 17592 5646 17644 5652
rect 17604 4826 17632 5646
rect 17696 5302 17724 5782
rect 17868 5704 17920 5710
rect 17868 5646 17920 5652
rect 17684 5296 17736 5302
rect 17684 5238 17736 5244
rect 17880 5166 17908 5646
rect 17868 5160 17920 5166
rect 17868 5102 17920 5108
rect 17592 4820 17644 4826
rect 17592 4762 17644 4768
rect 17972 2514 18000 6208
rect 18052 5228 18104 5234
rect 18052 5170 18104 5176
rect 18064 4826 18092 5170
rect 18984 5030 19012 6598
rect 18972 5024 19024 5030
rect 18972 4966 19024 4972
rect 18984 4826 19012 4966
rect 18052 4820 18104 4826
rect 18052 4762 18104 4768
rect 18972 4820 19024 4826
rect 18972 4762 19024 4768
rect 18604 4616 18656 4622
rect 18604 4558 18656 4564
rect 18512 4276 18564 4282
rect 18512 4218 18564 4224
rect 18524 4078 18552 4218
rect 18144 4072 18196 4078
rect 18144 4014 18196 4020
rect 18512 4072 18564 4078
rect 18512 4014 18564 4020
rect 18156 3738 18184 4014
rect 18616 4010 18644 4558
rect 18984 4282 19012 4762
rect 18972 4276 19024 4282
rect 18972 4218 19024 4224
rect 19168 4146 19196 6938
rect 19628 6254 19656 6938
rect 20180 6662 20208 7278
rect 23570 7239 23626 7248
rect 20168 6656 20220 6662
rect 20168 6598 20220 6604
rect 20180 6322 20208 6598
rect 20956 6556 21252 6576
rect 21012 6554 21036 6556
rect 21092 6554 21116 6556
rect 21172 6554 21196 6556
rect 21034 6502 21036 6554
rect 21098 6502 21110 6554
rect 21172 6502 21174 6554
rect 21012 6500 21036 6502
rect 21092 6500 21116 6502
rect 21172 6500 21196 6502
rect 20956 6480 21252 6500
rect 20168 6316 20220 6322
rect 20168 6258 20220 6264
rect 19616 6248 19668 6254
rect 19616 6190 19668 6196
rect 19340 5704 19392 5710
rect 19340 5646 19392 5652
rect 19352 5370 19380 5646
rect 20956 5468 21252 5488
rect 21012 5466 21036 5468
rect 21092 5466 21116 5468
rect 21172 5466 21196 5468
rect 21034 5414 21036 5466
rect 21098 5414 21110 5466
rect 21172 5414 21174 5466
rect 21012 5412 21036 5414
rect 21092 5412 21116 5414
rect 21172 5412 21196 5414
rect 20956 5392 21252 5412
rect 19340 5364 19392 5370
rect 19340 5306 19392 5312
rect 23570 5264 23626 5273
rect 23570 5199 23626 5208
rect 19984 5092 20036 5098
rect 19984 5034 20036 5040
rect 19432 5024 19484 5030
rect 19432 4966 19484 4972
rect 19156 4140 19208 4146
rect 19156 4082 19208 4088
rect 19444 4078 19472 4966
rect 19996 4826 20024 5034
rect 19984 4820 20036 4826
rect 19984 4762 20036 4768
rect 20956 4380 21252 4400
rect 21012 4378 21036 4380
rect 21092 4378 21116 4380
rect 21172 4378 21196 4380
rect 21034 4326 21036 4378
rect 21098 4326 21110 4378
rect 21172 4326 21174 4378
rect 21012 4324 21036 4326
rect 21092 4324 21116 4326
rect 21172 4324 21196 4326
rect 20956 4304 21252 4324
rect 19432 4072 19484 4078
rect 23584 4049 23612 5199
rect 19432 4014 19484 4020
rect 23570 4040 23626 4049
rect 18604 4004 18656 4010
rect 18604 3946 18656 3952
rect 23112 4004 23164 4010
rect 23570 3975 23626 3984
rect 23112 3946 23164 3952
rect 18144 3732 18196 3738
rect 18144 3674 18196 3680
rect 20956 3292 21252 3312
rect 21012 3290 21036 3292
rect 21092 3290 21116 3292
rect 21172 3290 21196 3292
rect 21034 3238 21036 3290
rect 21098 3238 21110 3290
rect 21172 3238 21174 3290
rect 21012 3236 21036 3238
rect 21092 3236 21116 3238
rect 21172 3236 21196 3238
rect 20956 3216 21252 3236
rect 17960 2508 18012 2514
rect 17960 2450 18012 2456
rect 19432 2372 19484 2378
rect 19432 2314 19484 2320
rect 17498 82 17554 480
rect 17420 54 17554 82
rect 11978 0 12034 54
rect 13818 0 13874 54
rect 15658 0 15714 54
rect 17498 0 17554 54
rect 19338 82 19394 480
rect 19444 82 19472 2314
rect 20956 2204 21252 2224
rect 21012 2202 21036 2204
rect 21092 2202 21116 2204
rect 21172 2202 21196 2204
rect 21034 2150 21036 2202
rect 21098 2150 21110 2202
rect 21172 2150 21174 2202
rect 21012 2148 21036 2150
rect 21092 2148 21116 2150
rect 21172 2148 21196 2150
rect 20956 2128 21252 2148
rect 21270 1320 21326 1329
rect 21270 1255 21326 1264
rect 19338 54 19472 82
rect 21178 82 21234 480
rect 21284 82 21312 1255
rect 21178 54 21312 82
rect 23018 82 23074 480
rect 23124 82 23152 3946
rect 23018 54 23152 82
rect 19338 0 19394 54
rect 21178 0 21234 54
rect 23018 0 23074 54
<< via2 >>
rect 1306 22480 1362 22536
rect 2134 20848 2190 20904
rect 1306 19216 1362 19272
rect 1306 17720 1362 17776
rect 1582 16224 1638 16280
rect 18 13368 74 13424
rect 110 10240 166 10296
rect 110 9560 166 9616
rect 1766 12144 1822 12200
rect 1858 10240 1914 10296
rect 2962 9288 3018 9344
rect 110 8608 166 8664
rect 110 5480 166 5536
rect 110 3848 166 3904
rect 4956 21786 5012 21788
rect 5036 21786 5092 21788
rect 5116 21786 5172 21788
rect 5196 21786 5252 21788
rect 4956 21734 4982 21786
rect 4982 21734 5012 21786
rect 5036 21734 5046 21786
rect 5046 21734 5092 21786
rect 5116 21734 5162 21786
rect 5162 21734 5172 21786
rect 5196 21734 5226 21786
rect 5226 21734 5252 21786
rect 4956 21732 5012 21734
rect 5036 21732 5092 21734
rect 5116 21732 5172 21734
rect 5196 21732 5252 21734
rect 4956 20698 5012 20700
rect 5036 20698 5092 20700
rect 5116 20698 5172 20700
rect 5196 20698 5252 20700
rect 4956 20646 4982 20698
rect 4982 20646 5012 20698
rect 5036 20646 5046 20698
rect 5046 20646 5092 20698
rect 5116 20646 5162 20698
rect 5162 20646 5172 20698
rect 5196 20646 5226 20698
rect 5226 20646 5252 20698
rect 4956 20644 5012 20646
rect 5036 20644 5092 20646
rect 5116 20644 5172 20646
rect 5196 20644 5252 20646
rect 8956 21242 9012 21244
rect 9036 21242 9092 21244
rect 9116 21242 9172 21244
rect 9196 21242 9252 21244
rect 8956 21190 8982 21242
rect 8982 21190 9012 21242
rect 9036 21190 9046 21242
rect 9046 21190 9092 21242
rect 9116 21190 9162 21242
rect 9162 21190 9172 21242
rect 9196 21190 9226 21242
rect 9226 21190 9252 21242
rect 8956 21188 9012 21190
rect 9036 21188 9092 21190
rect 9116 21188 9172 21190
rect 9196 21188 9252 21190
rect 12956 21786 13012 21788
rect 13036 21786 13092 21788
rect 13116 21786 13172 21788
rect 13196 21786 13252 21788
rect 12956 21734 12982 21786
rect 12982 21734 13012 21786
rect 13036 21734 13046 21786
rect 13046 21734 13092 21786
rect 13116 21734 13162 21786
rect 13162 21734 13172 21786
rect 13196 21734 13226 21786
rect 13226 21734 13252 21786
rect 12956 21732 13012 21734
rect 13036 21732 13092 21734
rect 13116 21732 13172 21734
rect 13196 21732 13252 21734
rect 12956 20698 13012 20700
rect 13036 20698 13092 20700
rect 13116 20698 13172 20700
rect 13196 20698 13252 20700
rect 12956 20646 12982 20698
rect 12982 20646 13012 20698
rect 13036 20646 13046 20698
rect 13046 20646 13092 20698
rect 13116 20646 13162 20698
rect 13162 20646 13172 20698
rect 13196 20646 13226 20698
rect 13226 20646 13252 20698
rect 12956 20644 13012 20646
rect 13036 20644 13092 20646
rect 13116 20644 13172 20646
rect 13196 20644 13252 20646
rect 4956 19610 5012 19612
rect 5036 19610 5092 19612
rect 5116 19610 5172 19612
rect 5196 19610 5252 19612
rect 4956 19558 4982 19610
rect 4982 19558 5012 19610
rect 5036 19558 5046 19610
rect 5046 19558 5092 19610
rect 5116 19558 5162 19610
rect 5162 19558 5172 19610
rect 5196 19558 5226 19610
rect 5226 19558 5252 19610
rect 4956 19556 5012 19558
rect 5036 19556 5092 19558
rect 5116 19556 5172 19558
rect 5196 19556 5252 19558
rect 4956 18522 5012 18524
rect 5036 18522 5092 18524
rect 5116 18522 5172 18524
rect 5196 18522 5252 18524
rect 4956 18470 4982 18522
rect 4982 18470 5012 18522
rect 5036 18470 5046 18522
rect 5046 18470 5092 18522
rect 5116 18470 5162 18522
rect 5162 18470 5172 18522
rect 5196 18470 5226 18522
rect 5226 18470 5252 18522
rect 4956 18468 5012 18470
rect 5036 18468 5092 18470
rect 5116 18468 5172 18470
rect 5196 18468 5252 18470
rect 4956 17434 5012 17436
rect 5036 17434 5092 17436
rect 5116 17434 5172 17436
rect 5196 17434 5252 17436
rect 4956 17382 4982 17434
rect 4982 17382 5012 17434
rect 5036 17382 5046 17434
rect 5046 17382 5092 17434
rect 5116 17382 5162 17434
rect 5162 17382 5172 17434
rect 5196 17382 5226 17434
rect 5226 17382 5252 17434
rect 4956 17380 5012 17382
rect 5036 17380 5092 17382
rect 5116 17380 5172 17382
rect 5196 17380 5252 17382
rect 4956 16346 5012 16348
rect 5036 16346 5092 16348
rect 5116 16346 5172 16348
rect 5196 16346 5252 16348
rect 4956 16294 4982 16346
rect 4982 16294 5012 16346
rect 5036 16294 5046 16346
rect 5046 16294 5092 16346
rect 5116 16294 5162 16346
rect 5162 16294 5172 16346
rect 5196 16294 5226 16346
rect 5226 16294 5252 16346
rect 4956 16292 5012 16294
rect 5036 16292 5092 16294
rect 5116 16292 5172 16294
rect 5196 16292 5252 16294
rect 4956 15258 5012 15260
rect 5036 15258 5092 15260
rect 5116 15258 5172 15260
rect 5196 15258 5252 15260
rect 4956 15206 4982 15258
rect 4982 15206 5012 15258
rect 5036 15206 5046 15258
rect 5046 15206 5092 15258
rect 5116 15206 5162 15258
rect 5162 15206 5172 15258
rect 5196 15206 5226 15258
rect 5226 15206 5252 15258
rect 4956 15204 5012 15206
rect 5036 15204 5092 15206
rect 5116 15204 5172 15206
rect 5196 15204 5252 15206
rect 4710 14456 4766 14512
rect 3146 7792 3202 7848
rect 4956 14170 5012 14172
rect 5036 14170 5092 14172
rect 5116 14170 5172 14172
rect 5196 14170 5252 14172
rect 4956 14118 4982 14170
rect 4982 14118 5012 14170
rect 5036 14118 5046 14170
rect 5046 14118 5092 14170
rect 5116 14118 5162 14170
rect 5162 14118 5172 14170
rect 5196 14118 5226 14170
rect 5226 14118 5252 14170
rect 4956 14116 5012 14118
rect 5036 14116 5092 14118
rect 5116 14116 5172 14118
rect 5196 14116 5252 14118
rect 4710 13232 4766 13288
rect 4956 13082 5012 13084
rect 5036 13082 5092 13084
rect 5116 13082 5172 13084
rect 5196 13082 5252 13084
rect 4956 13030 4982 13082
rect 4982 13030 5012 13082
rect 5036 13030 5046 13082
rect 5046 13030 5092 13082
rect 5116 13030 5162 13082
rect 5162 13030 5172 13082
rect 5196 13030 5226 13082
rect 5226 13030 5252 13082
rect 4956 13028 5012 13030
rect 5036 13028 5092 13030
rect 5116 13028 5172 13030
rect 5196 13028 5252 13030
rect 4956 11994 5012 11996
rect 5036 11994 5092 11996
rect 5116 11994 5172 11996
rect 5196 11994 5252 11996
rect 4956 11942 4982 11994
rect 4982 11942 5012 11994
rect 5036 11942 5046 11994
rect 5046 11942 5092 11994
rect 5116 11942 5162 11994
rect 5162 11942 5172 11994
rect 5196 11942 5226 11994
rect 5226 11942 5252 11994
rect 4956 11940 5012 11942
rect 5036 11940 5092 11942
rect 5116 11940 5172 11942
rect 5196 11940 5252 11942
rect 4802 11600 4858 11656
rect 3790 7928 3846 7984
rect 3974 6840 4030 6896
rect 4956 10906 5012 10908
rect 5036 10906 5092 10908
rect 5116 10906 5172 10908
rect 5196 10906 5252 10908
rect 4956 10854 4982 10906
rect 4982 10854 5012 10906
rect 5036 10854 5046 10906
rect 5046 10854 5092 10906
rect 5116 10854 5162 10906
rect 5162 10854 5172 10906
rect 5196 10854 5226 10906
rect 5226 10854 5252 10906
rect 4956 10852 5012 10854
rect 5036 10852 5092 10854
rect 5116 10852 5172 10854
rect 5196 10852 5252 10854
rect 4956 9818 5012 9820
rect 5036 9818 5092 9820
rect 5116 9818 5172 9820
rect 5196 9818 5252 9820
rect 4956 9766 4982 9818
rect 4982 9766 5012 9818
rect 5036 9766 5046 9818
rect 5046 9766 5092 9818
rect 5116 9766 5162 9818
rect 5162 9766 5172 9818
rect 5196 9766 5226 9818
rect 5226 9766 5252 9818
rect 4956 9764 5012 9766
rect 5036 9764 5092 9766
rect 5116 9764 5172 9766
rect 5196 9764 5252 9766
rect 4956 8730 5012 8732
rect 5036 8730 5092 8732
rect 5116 8730 5172 8732
rect 5196 8730 5252 8732
rect 4956 8678 4982 8730
rect 4982 8678 5012 8730
rect 5036 8678 5046 8730
rect 5046 8678 5092 8730
rect 5116 8678 5162 8730
rect 5162 8678 5172 8730
rect 5196 8678 5226 8730
rect 5226 8678 5252 8730
rect 4956 8676 5012 8678
rect 5036 8676 5092 8678
rect 5116 8676 5172 8678
rect 5196 8676 5252 8678
rect 4956 7642 5012 7644
rect 5036 7642 5092 7644
rect 5116 7642 5172 7644
rect 5196 7642 5252 7644
rect 4956 7590 4982 7642
rect 4982 7590 5012 7642
rect 5036 7590 5046 7642
rect 5046 7590 5092 7642
rect 5116 7590 5162 7642
rect 5162 7590 5172 7642
rect 5196 7590 5226 7642
rect 5226 7590 5252 7642
rect 4956 7588 5012 7590
rect 5036 7588 5092 7590
rect 5116 7588 5172 7590
rect 5196 7588 5252 7590
rect 4956 6554 5012 6556
rect 5036 6554 5092 6556
rect 5116 6554 5172 6556
rect 5196 6554 5252 6556
rect 4956 6502 4982 6554
rect 4982 6502 5012 6554
rect 5036 6502 5046 6554
rect 5046 6502 5092 6554
rect 5116 6502 5162 6554
rect 5162 6502 5172 6554
rect 5196 6502 5226 6554
rect 5226 6502 5252 6554
rect 4956 6500 5012 6502
rect 5036 6500 5092 6502
rect 5116 6500 5172 6502
rect 5196 6500 5252 6502
rect 4618 6296 4674 6352
rect 4956 5466 5012 5468
rect 5036 5466 5092 5468
rect 5116 5466 5172 5468
rect 5196 5466 5252 5468
rect 4956 5414 4982 5466
rect 4982 5414 5012 5466
rect 5036 5414 5046 5466
rect 5046 5414 5092 5466
rect 5116 5414 5162 5466
rect 5162 5414 5172 5466
rect 5196 5414 5226 5466
rect 5226 5414 5252 5466
rect 4956 5412 5012 5414
rect 5036 5412 5092 5414
rect 5116 5412 5172 5414
rect 5196 5412 5252 5414
rect 3514 5072 3570 5128
rect 8956 20154 9012 20156
rect 9036 20154 9092 20156
rect 9116 20154 9172 20156
rect 9196 20154 9252 20156
rect 8956 20102 8982 20154
rect 8982 20102 9012 20154
rect 9036 20102 9046 20154
rect 9046 20102 9092 20154
rect 9116 20102 9162 20154
rect 9162 20102 9172 20154
rect 9196 20102 9226 20154
rect 9226 20102 9252 20154
rect 8956 20100 9012 20102
rect 9036 20100 9092 20102
rect 9116 20100 9172 20102
rect 9196 20100 9252 20102
rect 8956 19066 9012 19068
rect 9036 19066 9092 19068
rect 9116 19066 9172 19068
rect 9196 19066 9252 19068
rect 8956 19014 8982 19066
rect 8982 19014 9012 19066
rect 9036 19014 9046 19066
rect 9046 19014 9092 19066
rect 9116 19014 9162 19066
rect 9162 19014 9172 19066
rect 9196 19014 9226 19066
rect 9226 19014 9252 19066
rect 8956 19012 9012 19014
rect 9036 19012 9092 19014
rect 9116 19012 9172 19014
rect 9196 19012 9252 19014
rect 4956 4378 5012 4380
rect 5036 4378 5092 4380
rect 5116 4378 5172 4380
rect 5196 4378 5252 4380
rect 4956 4326 4982 4378
rect 4982 4326 5012 4378
rect 5036 4326 5046 4378
rect 5046 4326 5092 4378
rect 5116 4326 5162 4378
rect 5162 4326 5172 4378
rect 5196 4326 5226 4378
rect 5226 4326 5252 4378
rect 4956 4324 5012 4326
rect 5036 4324 5092 4326
rect 5116 4324 5172 4326
rect 5196 4324 5252 4326
rect 4956 3290 5012 3292
rect 5036 3290 5092 3292
rect 5116 3290 5172 3292
rect 5196 3290 5252 3292
rect 4956 3238 4982 3290
rect 4982 3238 5012 3290
rect 5036 3238 5046 3290
rect 5046 3238 5092 3290
rect 5116 3238 5162 3290
rect 5162 3238 5172 3290
rect 5196 3238 5226 3290
rect 5226 3238 5252 3290
rect 4956 3236 5012 3238
rect 5036 3236 5092 3238
rect 5116 3236 5172 3238
rect 5196 3236 5252 3238
rect 5814 5072 5870 5128
rect 4158 1264 4214 1320
rect 4956 2202 5012 2204
rect 5036 2202 5092 2204
rect 5116 2202 5172 2204
rect 5196 2202 5252 2204
rect 4956 2150 4982 2202
rect 4982 2150 5012 2202
rect 5036 2150 5046 2202
rect 5046 2150 5092 2202
rect 5116 2150 5162 2202
rect 5162 2150 5172 2202
rect 5196 2150 5226 2202
rect 5226 2150 5252 2202
rect 4956 2148 5012 2150
rect 5036 2148 5092 2150
rect 5116 2148 5172 2150
rect 5196 2148 5252 2150
rect 6734 7928 6790 7984
rect 8114 2916 8170 2952
rect 8114 2896 8116 2916
rect 8116 2896 8168 2916
rect 8168 2896 8170 2916
rect 8956 17978 9012 17980
rect 9036 17978 9092 17980
rect 9116 17978 9172 17980
rect 9196 17978 9252 17980
rect 8956 17926 8982 17978
rect 8982 17926 9012 17978
rect 9036 17926 9046 17978
rect 9046 17926 9092 17978
rect 9116 17926 9162 17978
rect 9162 17926 9172 17978
rect 9196 17926 9226 17978
rect 9226 17926 9252 17978
rect 8956 17924 9012 17926
rect 9036 17924 9092 17926
rect 9116 17924 9172 17926
rect 9196 17924 9252 17926
rect 9862 17584 9918 17640
rect 8956 16890 9012 16892
rect 9036 16890 9092 16892
rect 9116 16890 9172 16892
rect 9196 16890 9252 16892
rect 8956 16838 8982 16890
rect 8982 16838 9012 16890
rect 9036 16838 9046 16890
rect 9046 16838 9092 16890
rect 9116 16838 9162 16890
rect 9162 16838 9172 16890
rect 9196 16838 9226 16890
rect 9226 16838 9252 16890
rect 8956 16836 9012 16838
rect 9036 16836 9092 16838
rect 9116 16836 9172 16838
rect 9196 16836 9252 16838
rect 8956 15802 9012 15804
rect 9036 15802 9092 15804
rect 9116 15802 9172 15804
rect 9196 15802 9252 15804
rect 8956 15750 8982 15802
rect 8982 15750 9012 15802
rect 9036 15750 9046 15802
rect 9046 15750 9092 15802
rect 9116 15750 9162 15802
rect 9162 15750 9172 15802
rect 9196 15750 9226 15802
rect 9226 15750 9252 15802
rect 8956 15748 9012 15750
rect 9036 15748 9092 15750
rect 9116 15748 9172 15750
rect 9196 15748 9252 15750
rect 8956 14714 9012 14716
rect 9036 14714 9092 14716
rect 9116 14714 9172 14716
rect 9196 14714 9252 14716
rect 8956 14662 8982 14714
rect 8982 14662 9012 14714
rect 9036 14662 9046 14714
rect 9046 14662 9092 14714
rect 9116 14662 9162 14714
rect 9162 14662 9172 14714
rect 9196 14662 9226 14714
rect 9226 14662 9252 14714
rect 8956 14660 9012 14662
rect 9036 14660 9092 14662
rect 9116 14660 9172 14662
rect 9196 14660 9252 14662
rect 8956 13626 9012 13628
rect 9036 13626 9092 13628
rect 9116 13626 9172 13628
rect 9196 13626 9252 13628
rect 8956 13574 8982 13626
rect 8982 13574 9012 13626
rect 9036 13574 9046 13626
rect 9046 13574 9092 13626
rect 9116 13574 9162 13626
rect 9162 13574 9172 13626
rect 9196 13574 9226 13626
rect 9226 13574 9252 13626
rect 8956 13572 9012 13574
rect 9036 13572 9092 13574
rect 9116 13572 9172 13574
rect 9196 13572 9252 13574
rect 8482 10240 8538 10296
rect 8956 12538 9012 12540
rect 9036 12538 9092 12540
rect 9116 12538 9172 12540
rect 9196 12538 9252 12540
rect 8956 12486 8982 12538
rect 8982 12486 9012 12538
rect 9036 12486 9046 12538
rect 9046 12486 9092 12538
rect 9116 12486 9162 12538
rect 9162 12486 9172 12538
rect 9196 12486 9226 12538
rect 9226 12486 9252 12538
rect 8956 12484 9012 12486
rect 9036 12484 9092 12486
rect 9116 12484 9172 12486
rect 9196 12484 9252 12486
rect 8956 11450 9012 11452
rect 9036 11450 9092 11452
rect 9116 11450 9172 11452
rect 9196 11450 9252 11452
rect 8956 11398 8982 11450
rect 8982 11398 9012 11450
rect 9036 11398 9046 11450
rect 9046 11398 9092 11450
rect 9116 11398 9162 11450
rect 9162 11398 9172 11450
rect 9196 11398 9226 11450
rect 9226 11398 9252 11450
rect 8956 11396 9012 11398
rect 9036 11396 9092 11398
rect 9116 11396 9172 11398
rect 9196 11396 9252 11398
rect 8956 10362 9012 10364
rect 9036 10362 9092 10364
rect 9116 10362 9172 10364
rect 9196 10362 9252 10364
rect 8956 10310 8982 10362
rect 8982 10310 9012 10362
rect 9036 10310 9046 10362
rect 9046 10310 9092 10362
rect 9116 10310 9162 10362
rect 9162 10310 9172 10362
rect 9196 10310 9226 10362
rect 9226 10310 9252 10362
rect 8956 10308 9012 10310
rect 9036 10308 9092 10310
rect 9116 10308 9172 10310
rect 9196 10308 9252 10310
rect 8666 9288 8722 9344
rect 9402 9288 9458 9344
rect 9586 9288 9642 9344
rect 8956 9274 9012 9276
rect 9036 9274 9092 9276
rect 9116 9274 9172 9276
rect 9196 9274 9252 9276
rect 8956 9222 8982 9274
rect 8982 9222 9012 9274
rect 9036 9222 9046 9274
rect 9046 9222 9092 9274
rect 9116 9222 9162 9274
rect 9162 9222 9172 9274
rect 9196 9222 9226 9274
rect 9226 9222 9252 9274
rect 8956 9220 9012 9222
rect 9036 9220 9092 9222
rect 9116 9220 9172 9222
rect 9196 9220 9252 9222
rect 8758 8880 8814 8936
rect 8956 8186 9012 8188
rect 9036 8186 9092 8188
rect 9116 8186 9172 8188
rect 9196 8186 9252 8188
rect 8956 8134 8982 8186
rect 8982 8134 9012 8186
rect 9036 8134 9046 8186
rect 9046 8134 9092 8186
rect 9116 8134 9162 8186
rect 9162 8134 9172 8186
rect 9196 8134 9226 8186
rect 9226 8134 9252 8186
rect 8956 8132 9012 8134
rect 9036 8132 9092 8134
rect 9116 8132 9172 8134
rect 9196 8132 9252 8134
rect 8956 7098 9012 7100
rect 9036 7098 9092 7100
rect 9116 7098 9172 7100
rect 9196 7098 9252 7100
rect 8956 7046 8982 7098
rect 8982 7046 9012 7098
rect 9036 7046 9046 7098
rect 9046 7046 9092 7098
rect 9116 7046 9162 7098
rect 9162 7046 9172 7098
rect 9196 7046 9226 7098
rect 9226 7046 9252 7098
rect 8956 7044 9012 7046
rect 9036 7044 9092 7046
rect 9116 7044 9172 7046
rect 9196 7044 9252 7046
rect 8956 6010 9012 6012
rect 9036 6010 9092 6012
rect 9116 6010 9172 6012
rect 9196 6010 9252 6012
rect 8956 5958 8982 6010
rect 8982 5958 9012 6010
rect 9036 5958 9046 6010
rect 9046 5958 9092 6010
rect 9116 5958 9162 6010
rect 9162 5958 9172 6010
rect 9196 5958 9226 6010
rect 9226 5958 9252 6010
rect 8956 5956 9012 5958
rect 9036 5956 9092 5958
rect 9116 5956 9172 5958
rect 9196 5956 9252 5958
rect 8956 4922 9012 4924
rect 9036 4922 9092 4924
rect 9116 4922 9172 4924
rect 9196 4922 9252 4924
rect 8956 4870 8982 4922
rect 8982 4870 9012 4922
rect 9036 4870 9046 4922
rect 9046 4870 9092 4922
rect 9116 4870 9162 4922
rect 9162 4870 9172 4922
rect 9196 4870 9226 4922
rect 9226 4870 9252 4922
rect 8956 4868 9012 4870
rect 9036 4868 9092 4870
rect 9116 4868 9172 4870
rect 9196 4868 9252 4870
rect 9954 11736 10010 11792
rect 9954 9560 10010 9616
rect 10414 12144 10470 12200
rect 12956 19610 13012 19612
rect 13036 19610 13092 19612
rect 13116 19610 13172 19612
rect 13196 19610 13252 19612
rect 12956 19558 12982 19610
rect 12982 19558 13012 19610
rect 13036 19558 13046 19610
rect 13046 19558 13092 19610
rect 13116 19558 13162 19610
rect 13162 19558 13172 19610
rect 13196 19558 13226 19610
rect 13226 19558 13252 19610
rect 12956 19556 13012 19558
rect 13036 19556 13092 19558
rect 13116 19556 13172 19558
rect 13196 19556 13252 19558
rect 12956 18522 13012 18524
rect 13036 18522 13092 18524
rect 13116 18522 13172 18524
rect 13196 18522 13252 18524
rect 12956 18470 12982 18522
rect 12982 18470 13012 18522
rect 13036 18470 13046 18522
rect 13046 18470 13092 18522
rect 13116 18470 13162 18522
rect 13162 18470 13172 18522
rect 13196 18470 13226 18522
rect 13226 18470 13252 18522
rect 12956 18468 13012 18470
rect 13036 18468 13092 18470
rect 13116 18468 13172 18470
rect 13196 18468 13252 18470
rect 11794 16940 11796 16960
rect 11796 16940 11848 16960
rect 11848 16940 11850 16960
rect 11794 16904 11850 16940
rect 11242 13776 11298 13832
rect 8956 3834 9012 3836
rect 9036 3834 9092 3836
rect 9116 3834 9172 3836
rect 9196 3834 9252 3836
rect 8956 3782 8982 3834
rect 8982 3782 9012 3834
rect 9036 3782 9046 3834
rect 9046 3782 9092 3834
rect 9116 3782 9162 3834
rect 9162 3782 9172 3834
rect 9196 3782 9226 3834
rect 9226 3782 9252 3834
rect 8956 3780 9012 3782
rect 9036 3780 9092 3782
rect 9116 3780 9172 3782
rect 9196 3780 9252 3782
rect 8298 2760 8354 2816
rect 8956 2746 9012 2748
rect 9036 2746 9092 2748
rect 9116 2746 9172 2748
rect 9196 2746 9252 2748
rect 8956 2694 8982 2746
rect 8982 2694 9012 2746
rect 9036 2694 9046 2746
rect 9046 2694 9092 2746
rect 9116 2694 9162 2746
rect 9162 2694 9172 2746
rect 9196 2694 9226 2746
rect 9226 2694 9252 2746
rect 8956 2692 9012 2694
rect 9036 2692 9092 2694
rect 9116 2692 9172 2694
rect 9196 2692 9252 2694
rect 5906 1264 5962 1320
rect 5354 176 5410 232
rect 9862 1672 9918 1728
rect 8574 1536 8630 1592
rect 12622 16904 12678 16960
rect 12956 17434 13012 17436
rect 13036 17434 13092 17436
rect 13116 17434 13172 17436
rect 13196 17434 13252 17436
rect 12956 17382 12982 17434
rect 12982 17382 13012 17434
rect 13036 17382 13046 17434
rect 13046 17382 13092 17434
rect 13116 17382 13162 17434
rect 13162 17382 13172 17434
rect 13196 17382 13226 17434
rect 13226 17382 13252 17434
rect 12956 17380 13012 17382
rect 13036 17380 13092 17382
rect 13116 17380 13172 17382
rect 13196 17380 13252 17382
rect 12956 16346 13012 16348
rect 13036 16346 13092 16348
rect 13116 16346 13172 16348
rect 13196 16346 13252 16348
rect 12956 16294 12982 16346
rect 12982 16294 13012 16346
rect 13036 16294 13046 16346
rect 13046 16294 13092 16346
rect 13116 16294 13162 16346
rect 13162 16294 13172 16346
rect 13196 16294 13226 16346
rect 13226 16294 13252 16346
rect 12956 16292 13012 16294
rect 13036 16292 13092 16294
rect 13116 16292 13172 16294
rect 13196 16292 13252 16294
rect 12956 15258 13012 15260
rect 13036 15258 13092 15260
rect 13116 15258 13172 15260
rect 13196 15258 13252 15260
rect 12956 15206 12982 15258
rect 12982 15206 13012 15258
rect 13036 15206 13046 15258
rect 13046 15206 13092 15258
rect 13116 15206 13162 15258
rect 13162 15206 13172 15258
rect 13196 15206 13226 15258
rect 13226 15206 13252 15258
rect 12956 15204 13012 15206
rect 13036 15204 13092 15206
rect 13116 15204 13172 15206
rect 13196 15204 13252 15206
rect 12346 13232 12402 13288
rect 12956 14170 13012 14172
rect 13036 14170 13092 14172
rect 13116 14170 13172 14172
rect 13196 14170 13252 14172
rect 12956 14118 12982 14170
rect 12982 14118 13012 14170
rect 13036 14118 13046 14170
rect 13046 14118 13092 14170
rect 13116 14118 13162 14170
rect 13162 14118 13172 14170
rect 13196 14118 13226 14170
rect 13226 14118 13252 14170
rect 12956 14116 13012 14118
rect 13036 14116 13092 14118
rect 13116 14116 13172 14118
rect 13196 14116 13252 14118
rect 12956 13082 13012 13084
rect 13036 13082 13092 13084
rect 13116 13082 13172 13084
rect 13196 13082 13252 13084
rect 12956 13030 12982 13082
rect 12982 13030 13012 13082
rect 13036 13030 13046 13082
rect 13046 13030 13092 13082
rect 13116 13030 13162 13082
rect 13162 13030 13172 13082
rect 13196 13030 13226 13082
rect 13226 13030 13252 13082
rect 12956 13028 13012 13030
rect 13036 13028 13092 13030
rect 13116 13028 13172 13030
rect 13196 13028 13252 13030
rect 12070 11736 12126 11792
rect 12956 11994 13012 11996
rect 13036 11994 13092 11996
rect 13116 11994 13172 11996
rect 13196 11994 13252 11996
rect 12956 11942 12982 11994
rect 12982 11942 13012 11994
rect 13036 11942 13046 11994
rect 13046 11942 13092 11994
rect 13116 11942 13162 11994
rect 13162 11942 13172 11994
rect 13196 11942 13226 11994
rect 13226 11942 13252 11994
rect 12956 11940 13012 11942
rect 13036 11940 13092 11942
rect 13116 11940 13172 11942
rect 13196 11940 13252 11942
rect 11334 9152 11390 9208
rect 12956 10906 13012 10908
rect 13036 10906 13092 10908
rect 13116 10906 13172 10908
rect 13196 10906 13252 10908
rect 12956 10854 12982 10906
rect 12982 10854 13012 10906
rect 13036 10854 13046 10906
rect 13046 10854 13092 10906
rect 13116 10854 13162 10906
rect 13162 10854 13172 10906
rect 13196 10854 13226 10906
rect 13226 10854 13252 10906
rect 12956 10852 13012 10854
rect 13036 10852 13092 10854
rect 13116 10852 13172 10854
rect 13196 10852 13252 10854
rect 10506 7928 10562 7984
rect 12530 6840 12586 6896
rect 11702 6296 11758 6352
rect 11334 5072 11390 5128
rect 11886 5072 11942 5128
rect 12956 9818 13012 9820
rect 13036 9818 13092 9820
rect 13116 9818 13172 9820
rect 13196 9818 13252 9820
rect 12956 9766 12982 9818
rect 12982 9766 13012 9818
rect 13036 9766 13046 9818
rect 13046 9766 13092 9818
rect 13116 9766 13162 9818
rect 13162 9766 13172 9818
rect 13196 9766 13226 9818
rect 13226 9766 13252 9818
rect 12956 9764 13012 9766
rect 13036 9764 13092 9766
rect 13116 9764 13172 9766
rect 13196 9764 13252 9766
rect 12956 8730 13012 8732
rect 13036 8730 13092 8732
rect 13116 8730 13172 8732
rect 13196 8730 13252 8732
rect 12956 8678 12982 8730
rect 12982 8678 13012 8730
rect 13036 8678 13046 8730
rect 13046 8678 13092 8730
rect 13116 8678 13162 8730
rect 13162 8678 13172 8730
rect 13196 8678 13226 8730
rect 13226 8678 13252 8730
rect 12956 8676 13012 8678
rect 13036 8676 13092 8678
rect 13116 8676 13172 8678
rect 13196 8676 13252 8678
rect 12956 7642 13012 7644
rect 13036 7642 13092 7644
rect 13116 7642 13172 7644
rect 13196 7642 13252 7644
rect 12956 7590 12982 7642
rect 12982 7590 13012 7642
rect 13036 7590 13046 7642
rect 13046 7590 13092 7642
rect 13116 7590 13162 7642
rect 13162 7590 13172 7642
rect 13196 7590 13226 7642
rect 13226 7590 13252 7642
rect 12956 7588 13012 7590
rect 13036 7588 13092 7590
rect 13116 7588 13172 7590
rect 13196 7588 13252 7590
rect 16956 21242 17012 21244
rect 17036 21242 17092 21244
rect 17116 21242 17172 21244
rect 17196 21242 17252 21244
rect 16956 21190 16982 21242
rect 16982 21190 17012 21242
rect 17036 21190 17046 21242
rect 17046 21190 17092 21242
rect 17116 21190 17162 21242
rect 17162 21190 17172 21242
rect 17196 21190 17226 21242
rect 17226 21190 17252 21242
rect 16956 21188 17012 21190
rect 17036 21188 17092 21190
rect 17116 21188 17172 21190
rect 17196 21188 17252 21190
rect 13450 9696 13506 9752
rect 16956 20154 17012 20156
rect 17036 20154 17092 20156
rect 17116 20154 17172 20156
rect 17196 20154 17252 20156
rect 16956 20102 16982 20154
rect 16982 20102 17012 20154
rect 17036 20102 17046 20154
rect 17046 20102 17092 20154
rect 17116 20102 17162 20154
rect 17162 20102 17172 20154
rect 17196 20102 17226 20154
rect 17226 20102 17252 20154
rect 16956 20100 17012 20102
rect 17036 20100 17092 20102
rect 17116 20100 17172 20102
rect 17196 20100 17252 20102
rect 16956 19066 17012 19068
rect 17036 19066 17092 19068
rect 17116 19066 17172 19068
rect 17196 19066 17252 19068
rect 16956 19014 16982 19066
rect 16982 19014 17012 19066
rect 17036 19014 17046 19066
rect 17046 19014 17092 19066
rect 17116 19014 17162 19066
rect 17162 19014 17172 19066
rect 17196 19014 17226 19066
rect 17226 19014 17252 19066
rect 16956 19012 17012 19014
rect 17036 19012 17092 19014
rect 17116 19012 17172 19014
rect 17196 19012 17252 19014
rect 15106 12280 15162 12336
rect 16956 17978 17012 17980
rect 17036 17978 17092 17980
rect 17116 17978 17172 17980
rect 17196 17978 17252 17980
rect 16956 17926 16982 17978
rect 16982 17926 17012 17978
rect 17036 17926 17046 17978
rect 17046 17926 17092 17978
rect 17116 17926 17162 17978
rect 17162 17926 17172 17978
rect 17196 17926 17226 17978
rect 17226 17926 17252 17978
rect 16956 17924 17012 17926
rect 17036 17924 17092 17926
rect 17116 17924 17172 17926
rect 17196 17924 17252 17926
rect 16956 16890 17012 16892
rect 17036 16890 17092 16892
rect 17116 16890 17172 16892
rect 17196 16890 17252 16892
rect 16956 16838 16982 16890
rect 16982 16838 17012 16890
rect 17036 16838 17046 16890
rect 17046 16838 17092 16890
rect 17116 16838 17162 16890
rect 17162 16838 17172 16890
rect 17196 16838 17226 16890
rect 17226 16838 17252 16890
rect 16956 16836 17012 16838
rect 17036 16836 17092 16838
rect 17116 16836 17172 16838
rect 17196 16836 17252 16838
rect 16956 15802 17012 15804
rect 17036 15802 17092 15804
rect 17116 15802 17172 15804
rect 17196 15802 17252 15804
rect 16956 15750 16982 15802
rect 16982 15750 17012 15802
rect 17036 15750 17046 15802
rect 17046 15750 17092 15802
rect 17116 15750 17162 15802
rect 17162 15750 17172 15802
rect 17196 15750 17226 15802
rect 17226 15750 17252 15802
rect 16956 15748 17012 15750
rect 17036 15748 17092 15750
rect 17116 15748 17172 15750
rect 17196 15748 17252 15750
rect 13542 9424 13598 9480
rect 15474 9696 15530 9752
rect 14002 9152 14058 9208
rect 14738 8880 14794 8936
rect 13358 7384 13414 7440
rect 13266 7248 13322 7304
rect 12956 6554 13012 6556
rect 13036 6554 13092 6556
rect 13116 6554 13172 6556
rect 13196 6554 13252 6556
rect 12956 6502 12982 6554
rect 12982 6502 13012 6554
rect 13036 6502 13046 6554
rect 13046 6502 13092 6554
rect 13116 6502 13162 6554
rect 13162 6502 13172 6554
rect 13196 6502 13226 6554
rect 13226 6502 13252 6554
rect 12956 6500 13012 6502
rect 13036 6500 13092 6502
rect 13116 6500 13172 6502
rect 13196 6500 13252 6502
rect 12956 5466 13012 5468
rect 13036 5466 13092 5468
rect 13116 5466 13172 5468
rect 13196 5466 13252 5468
rect 12956 5414 12982 5466
rect 12982 5414 13012 5466
rect 13036 5414 13046 5466
rect 13046 5414 13092 5466
rect 13116 5414 13162 5466
rect 13162 5414 13172 5466
rect 13196 5414 13226 5466
rect 13226 5414 13252 5466
rect 12956 5412 13012 5414
rect 13036 5412 13092 5414
rect 13116 5412 13172 5414
rect 13196 5412 13252 5414
rect 14462 7792 14518 7848
rect 12956 4378 13012 4380
rect 13036 4378 13092 4380
rect 13116 4378 13172 4380
rect 13196 4378 13252 4380
rect 12956 4326 12982 4378
rect 12982 4326 13012 4378
rect 13036 4326 13046 4378
rect 13046 4326 13092 4378
rect 13116 4326 13162 4378
rect 13162 4326 13172 4378
rect 13196 4326 13226 4378
rect 13226 4326 13252 4378
rect 12956 4324 13012 4326
rect 13036 4324 13092 4326
rect 13116 4324 13172 4326
rect 13196 4324 13252 4326
rect 15934 7928 15990 7984
rect 13450 3984 13506 4040
rect 12956 3290 13012 3292
rect 13036 3290 13092 3292
rect 13116 3290 13172 3292
rect 13196 3290 13252 3292
rect 12956 3238 12982 3290
rect 12982 3238 13012 3290
rect 13036 3238 13046 3290
rect 13046 3238 13092 3290
rect 13116 3238 13162 3290
rect 13162 3238 13172 3290
rect 13196 3238 13226 3290
rect 13226 3238 13252 3290
rect 12956 3236 13012 3238
rect 13036 3236 13092 3238
rect 13116 3236 13172 3238
rect 13196 3236 13252 3238
rect 16956 14714 17012 14716
rect 17036 14714 17092 14716
rect 17116 14714 17172 14716
rect 17196 14714 17252 14716
rect 16956 14662 16982 14714
rect 16982 14662 17012 14714
rect 17036 14662 17046 14714
rect 17046 14662 17092 14714
rect 17116 14662 17162 14714
rect 17162 14662 17172 14714
rect 17196 14662 17226 14714
rect 17226 14662 17252 14714
rect 16956 14660 17012 14662
rect 17036 14660 17092 14662
rect 17116 14660 17172 14662
rect 17196 14660 17252 14662
rect 16956 13626 17012 13628
rect 17036 13626 17092 13628
rect 17116 13626 17172 13628
rect 17196 13626 17252 13628
rect 16956 13574 16982 13626
rect 16982 13574 17012 13626
rect 17036 13574 17046 13626
rect 17046 13574 17092 13626
rect 17116 13574 17162 13626
rect 17162 13574 17172 13626
rect 17196 13574 17226 13626
rect 17226 13574 17252 13626
rect 16956 13572 17012 13574
rect 17036 13572 17092 13574
rect 17116 13572 17172 13574
rect 17196 13572 17252 13574
rect 17866 17584 17922 17640
rect 16956 12538 17012 12540
rect 17036 12538 17092 12540
rect 17116 12538 17172 12540
rect 17196 12538 17252 12540
rect 16956 12486 16982 12538
rect 16982 12486 17012 12538
rect 17036 12486 17046 12538
rect 17046 12486 17092 12538
rect 17116 12486 17162 12538
rect 17162 12486 17172 12538
rect 17196 12486 17226 12538
rect 17226 12486 17252 12538
rect 16956 12484 17012 12486
rect 17036 12484 17092 12486
rect 17116 12484 17172 12486
rect 17196 12484 17252 12486
rect 16956 11450 17012 11452
rect 17036 11450 17092 11452
rect 17116 11450 17172 11452
rect 17196 11450 17252 11452
rect 16956 11398 16982 11450
rect 16982 11398 17012 11450
rect 17036 11398 17046 11450
rect 17046 11398 17092 11450
rect 17116 11398 17162 11450
rect 17162 11398 17172 11450
rect 17196 11398 17226 11450
rect 17226 11398 17252 11450
rect 16956 11396 17012 11398
rect 17036 11396 17092 11398
rect 17116 11396 17172 11398
rect 17196 11396 17252 11398
rect 16486 7792 16542 7848
rect 16956 10362 17012 10364
rect 17036 10362 17092 10364
rect 17116 10362 17172 10364
rect 17196 10362 17252 10364
rect 16956 10310 16982 10362
rect 16982 10310 17012 10362
rect 17036 10310 17046 10362
rect 17046 10310 17092 10362
rect 17116 10310 17162 10362
rect 17162 10310 17172 10362
rect 17196 10310 17226 10362
rect 17226 10310 17252 10362
rect 16956 10308 17012 10310
rect 17036 10308 17092 10310
rect 17116 10308 17172 10310
rect 17196 10308 17252 10310
rect 16956 9274 17012 9276
rect 17036 9274 17092 9276
rect 17116 9274 17172 9276
rect 17196 9274 17252 9276
rect 16956 9222 16982 9274
rect 16982 9222 17012 9274
rect 17036 9222 17046 9274
rect 17046 9222 17092 9274
rect 17116 9222 17162 9274
rect 17162 9222 17172 9274
rect 17196 9222 17226 9274
rect 17226 9222 17252 9274
rect 16956 9220 17012 9222
rect 17036 9220 17092 9222
rect 17116 9220 17172 9222
rect 17196 9220 17252 9222
rect 16956 8186 17012 8188
rect 17036 8186 17092 8188
rect 17116 8186 17172 8188
rect 17196 8186 17252 8188
rect 16956 8134 16982 8186
rect 16982 8134 17012 8186
rect 17036 8134 17046 8186
rect 17046 8134 17092 8186
rect 17116 8134 17162 8186
rect 17162 8134 17172 8186
rect 17196 8134 17226 8186
rect 17226 8134 17252 8186
rect 16956 8132 17012 8134
rect 17036 8132 17092 8134
rect 17116 8132 17172 8134
rect 17196 8132 17252 8134
rect 16956 7098 17012 7100
rect 17036 7098 17092 7100
rect 17116 7098 17172 7100
rect 17196 7098 17252 7100
rect 16956 7046 16982 7098
rect 16982 7046 17012 7098
rect 17036 7046 17046 7098
rect 17046 7046 17092 7098
rect 17116 7046 17162 7098
rect 17162 7046 17172 7098
rect 17196 7046 17226 7098
rect 17226 7046 17252 7098
rect 16956 7044 17012 7046
rect 17036 7044 17092 7046
rect 17116 7044 17172 7046
rect 17196 7044 17252 7046
rect 16956 6010 17012 6012
rect 17036 6010 17092 6012
rect 17116 6010 17172 6012
rect 17196 6010 17252 6012
rect 16956 5958 16982 6010
rect 16982 5958 17012 6010
rect 17036 5958 17046 6010
rect 17046 5958 17092 6010
rect 17116 5958 17162 6010
rect 17162 5958 17172 6010
rect 17196 5958 17226 6010
rect 17226 5958 17252 6010
rect 16956 5956 17012 5958
rect 17036 5956 17092 5958
rect 17116 5956 17172 5958
rect 17196 5956 17252 5958
rect 16956 4922 17012 4924
rect 17036 4922 17092 4924
rect 17116 4922 17172 4924
rect 17196 4922 17252 4924
rect 16956 4870 16982 4922
rect 16982 4870 17012 4922
rect 17036 4870 17046 4922
rect 17046 4870 17092 4922
rect 17116 4870 17162 4922
rect 17162 4870 17172 4922
rect 17196 4870 17226 4922
rect 17226 4870 17252 4922
rect 16956 4868 17012 4870
rect 17036 4868 17092 4870
rect 17116 4868 17172 4870
rect 17196 4868 17252 4870
rect 16956 3834 17012 3836
rect 17036 3834 17092 3836
rect 17116 3834 17172 3836
rect 17196 3834 17252 3836
rect 16956 3782 16982 3834
rect 16982 3782 17012 3834
rect 17036 3782 17046 3834
rect 17046 3782 17092 3834
rect 17116 3782 17162 3834
rect 17162 3782 17172 3834
rect 17196 3782 17226 3834
rect 17226 3782 17252 3834
rect 16956 3780 17012 3782
rect 17036 3780 17092 3782
rect 17116 3780 17172 3782
rect 17196 3780 17252 3782
rect 16956 2746 17012 2748
rect 17036 2746 17092 2748
rect 17116 2746 17172 2748
rect 17196 2746 17252 2748
rect 16956 2694 16982 2746
rect 16982 2694 17012 2746
rect 17036 2694 17046 2746
rect 17046 2694 17092 2746
rect 17116 2694 17162 2746
rect 17162 2694 17172 2746
rect 17196 2694 17226 2746
rect 17226 2694 17252 2746
rect 16956 2692 17012 2694
rect 17036 2692 17092 2694
rect 17116 2692 17172 2694
rect 17196 2692 17252 2694
rect 12956 2202 13012 2204
rect 13036 2202 13092 2204
rect 13116 2202 13172 2204
rect 13196 2202 13252 2204
rect 12956 2150 12982 2202
rect 12982 2150 13012 2202
rect 13036 2150 13046 2202
rect 13046 2150 13092 2202
rect 13116 2150 13162 2202
rect 13162 2150 13172 2202
rect 13196 2150 13226 2202
rect 13226 2150 13252 2202
rect 12956 2148 13012 2150
rect 13036 2148 13092 2150
rect 13116 2148 13172 2150
rect 13196 2148 13252 2150
rect 17130 1536 17186 1592
rect 19982 22616 20038 22672
rect 18878 17584 18934 17640
rect 18234 9424 18290 9480
rect 17958 7792 18014 7848
rect 17498 7112 17554 7168
rect 20956 21786 21012 21788
rect 21036 21786 21092 21788
rect 21116 21786 21172 21788
rect 21196 21786 21252 21788
rect 20956 21734 20982 21786
rect 20982 21734 21012 21786
rect 21036 21734 21046 21786
rect 21046 21734 21092 21786
rect 21116 21734 21162 21786
rect 21162 21734 21172 21786
rect 21196 21734 21226 21786
rect 21226 21734 21252 21786
rect 20956 21732 21012 21734
rect 21036 21732 21092 21734
rect 21116 21732 21172 21734
rect 21196 21732 21252 21734
rect 22006 21120 22062 21176
rect 20956 20698 21012 20700
rect 21036 20698 21092 20700
rect 21116 20698 21172 20700
rect 21196 20698 21252 20700
rect 20956 20646 20982 20698
rect 20982 20646 21012 20698
rect 21036 20646 21046 20698
rect 21046 20646 21092 20698
rect 21116 20646 21162 20698
rect 21162 20646 21172 20698
rect 21196 20646 21226 20698
rect 21226 20646 21252 20698
rect 20956 20644 21012 20646
rect 21036 20644 21092 20646
rect 21116 20644 21172 20646
rect 21196 20644 21252 20646
rect 21270 19760 21326 19816
rect 20956 19610 21012 19612
rect 21036 19610 21092 19612
rect 21116 19610 21172 19612
rect 21196 19610 21252 19612
rect 20956 19558 20982 19610
rect 20982 19558 21012 19610
rect 21036 19558 21046 19610
rect 21046 19558 21092 19610
rect 21116 19558 21162 19610
rect 21162 19558 21172 19610
rect 21196 19558 21226 19610
rect 21226 19558 21252 19610
rect 20956 19556 21012 19558
rect 21036 19556 21092 19558
rect 21116 19556 21172 19558
rect 21196 19556 21252 19558
rect 20956 18522 21012 18524
rect 21036 18522 21092 18524
rect 21116 18522 21172 18524
rect 21196 18522 21252 18524
rect 20956 18470 20982 18522
rect 20982 18470 21012 18522
rect 21036 18470 21046 18522
rect 21046 18470 21092 18522
rect 21116 18470 21162 18522
rect 21162 18470 21172 18522
rect 21196 18470 21226 18522
rect 21226 18470 21252 18522
rect 20956 18468 21012 18470
rect 21036 18468 21092 18470
rect 21116 18468 21172 18470
rect 21196 18468 21252 18470
rect 21086 18128 21142 18184
rect 20956 17434 21012 17436
rect 21036 17434 21092 17436
rect 21116 17434 21172 17436
rect 21196 17434 21252 17436
rect 20956 17382 20982 17434
rect 20982 17382 21012 17434
rect 21036 17382 21046 17434
rect 21046 17382 21092 17434
rect 21116 17382 21162 17434
rect 21162 17382 21172 17434
rect 21196 17382 21226 17434
rect 21226 17382 21252 17434
rect 20956 17380 21012 17382
rect 21036 17380 21092 17382
rect 21116 17380 21172 17382
rect 21196 17380 21252 17382
rect 21086 16632 21142 16688
rect 20956 16346 21012 16348
rect 21036 16346 21092 16348
rect 21116 16346 21172 16348
rect 21196 16346 21252 16348
rect 20956 16294 20982 16346
rect 20982 16294 21012 16346
rect 21036 16294 21046 16346
rect 21046 16294 21092 16346
rect 21116 16294 21162 16346
rect 21162 16294 21172 16346
rect 21196 16294 21226 16346
rect 21226 16294 21252 16346
rect 20956 16292 21012 16294
rect 21036 16292 21092 16294
rect 21116 16292 21172 16294
rect 21196 16292 21252 16294
rect 20956 15258 21012 15260
rect 21036 15258 21092 15260
rect 21116 15258 21172 15260
rect 21196 15258 21252 15260
rect 20956 15206 20982 15258
rect 20982 15206 21012 15258
rect 21036 15206 21046 15258
rect 21046 15206 21092 15258
rect 21116 15206 21162 15258
rect 21162 15206 21172 15258
rect 21196 15206 21226 15258
rect 21226 15206 21252 15258
rect 20956 15204 21012 15206
rect 21036 15204 21092 15206
rect 21116 15204 21172 15206
rect 21196 15204 21252 15206
rect 20956 14170 21012 14172
rect 21036 14170 21092 14172
rect 21116 14170 21172 14172
rect 21196 14170 21252 14172
rect 20956 14118 20982 14170
rect 20982 14118 21012 14170
rect 21036 14118 21046 14170
rect 21046 14118 21092 14170
rect 21116 14118 21162 14170
rect 21162 14118 21172 14170
rect 21196 14118 21226 14170
rect 21226 14118 21252 14170
rect 20956 14116 21012 14118
rect 21036 14116 21092 14118
rect 21116 14116 21172 14118
rect 21196 14116 21252 14118
rect 20350 13932 20406 13968
rect 20350 13912 20352 13932
rect 20352 13912 20404 13932
rect 20404 13912 20406 13932
rect 20956 13082 21012 13084
rect 21036 13082 21092 13084
rect 21116 13082 21172 13084
rect 21196 13082 21252 13084
rect 20956 13030 20982 13082
rect 20982 13030 21012 13082
rect 21036 13030 21046 13082
rect 21046 13030 21092 13082
rect 21116 13030 21162 13082
rect 21162 13030 21172 13082
rect 21196 13030 21226 13082
rect 21226 13030 21252 13082
rect 20956 13028 21012 13030
rect 21036 13028 21092 13030
rect 21116 13028 21172 13030
rect 21196 13028 21252 13030
rect 20956 11994 21012 11996
rect 21036 11994 21092 11996
rect 21116 11994 21172 11996
rect 21196 11994 21252 11996
rect 20956 11942 20982 11994
rect 20982 11942 21012 11994
rect 21036 11942 21046 11994
rect 21046 11942 21092 11994
rect 21116 11942 21162 11994
rect 21162 11942 21172 11994
rect 21196 11942 21226 11994
rect 21226 11942 21252 11994
rect 20956 11940 21012 11942
rect 21036 11940 21092 11942
rect 21116 11940 21172 11942
rect 21196 11940 21252 11942
rect 20718 11736 20774 11792
rect 21914 15136 21970 15192
rect 21914 13640 21970 13696
rect 23570 12688 23626 12744
rect 21270 11192 21326 11248
rect 20956 10906 21012 10908
rect 21036 10906 21092 10908
rect 21116 10906 21172 10908
rect 21196 10906 21252 10908
rect 20956 10854 20982 10906
rect 20982 10854 21012 10906
rect 21036 10854 21046 10906
rect 21046 10854 21092 10906
rect 21116 10854 21162 10906
rect 21162 10854 21172 10906
rect 21196 10854 21226 10906
rect 21226 10854 21252 10906
rect 20956 10852 21012 10854
rect 21036 10852 21092 10854
rect 21116 10852 21172 10854
rect 21196 10852 21252 10854
rect 20956 9818 21012 9820
rect 21036 9818 21092 9820
rect 21116 9818 21172 9820
rect 21196 9818 21252 9820
rect 20956 9766 20982 9818
rect 20982 9766 21012 9818
rect 21036 9766 21046 9818
rect 21046 9766 21092 9818
rect 21116 9766 21162 9818
rect 21162 9766 21172 9818
rect 21196 9766 21226 9818
rect 21226 9766 21252 9818
rect 20956 9764 21012 9766
rect 21036 9764 21092 9766
rect 21116 9764 21172 9766
rect 21196 9764 21252 9766
rect 21362 9696 21418 9752
rect 20956 8730 21012 8732
rect 21036 8730 21092 8732
rect 21116 8730 21172 8732
rect 21196 8730 21252 8732
rect 20956 8678 20982 8730
rect 20982 8678 21012 8730
rect 21036 8678 21046 8730
rect 21046 8678 21092 8730
rect 21116 8678 21162 8730
rect 21162 8678 21172 8730
rect 21196 8678 21226 8730
rect 21226 8678 21252 8730
rect 20956 8676 21012 8678
rect 21036 8676 21092 8678
rect 21116 8676 21172 8678
rect 21196 8676 21252 8678
rect 23570 8200 23626 8256
rect 20956 7642 21012 7644
rect 21036 7642 21092 7644
rect 21116 7642 21172 7644
rect 21196 7642 21252 7644
rect 20956 7590 20982 7642
rect 20982 7590 21012 7642
rect 21036 7590 21046 7642
rect 21046 7590 21092 7642
rect 21116 7590 21162 7642
rect 21162 7590 21172 7642
rect 21196 7590 21226 7642
rect 21226 7590 21252 7642
rect 20956 7588 21012 7590
rect 21036 7588 21092 7590
rect 21116 7588 21172 7590
rect 21196 7588 21252 7590
rect 23570 7248 23626 7304
rect 20956 6554 21012 6556
rect 21036 6554 21092 6556
rect 21116 6554 21172 6556
rect 21196 6554 21252 6556
rect 20956 6502 20982 6554
rect 20982 6502 21012 6554
rect 21036 6502 21046 6554
rect 21046 6502 21092 6554
rect 21116 6502 21162 6554
rect 21162 6502 21172 6554
rect 21196 6502 21226 6554
rect 21226 6502 21252 6554
rect 20956 6500 21012 6502
rect 21036 6500 21092 6502
rect 21116 6500 21172 6502
rect 21196 6500 21252 6502
rect 20956 5466 21012 5468
rect 21036 5466 21092 5468
rect 21116 5466 21172 5468
rect 21196 5466 21252 5468
rect 20956 5414 20982 5466
rect 20982 5414 21012 5466
rect 21036 5414 21046 5466
rect 21046 5414 21092 5466
rect 21116 5414 21162 5466
rect 21162 5414 21172 5466
rect 21196 5414 21226 5466
rect 21226 5414 21252 5466
rect 20956 5412 21012 5414
rect 21036 5412 21092 5414
rect 21116 5412 21172 5414
rect 21196 5412 21252 5414
rect 23570 5208 23626 5264
rect 20956 4378 21012 4380
rect 21036 4378 21092 4380
rect 21116 4378 21172 4380
rect 21196 4378 21252 4380
rect 20956 4326 20982 4378
rect 20982 4326 21012 4378
rect 21036 4326 21046 4378
rect 21046 4326 21092 4378
rect 21116 4326 21162 4378
rect 21162 4326 21172 4378
rect 21196 4326 21226 4378
rect 21226 4326 21252 4378
rect 20956 4324 21012 4326
rect 21036 4324 21092 4326
rect 21116 4324 21172 4326
rect 21196 4324 21252 4326
rect 23570 3984 23626 4040
rect 20956 3290 21012 3292
rect 21036 3290 21092 3292
rect 21116 3290 21172 3292
rect 21196 3290 21252 3292
rect 20956 3238 20982 3290
rect 20982 3238 21012 3290
rect 21036 3238 21046 3290
rect 21046 3238 21092 3290
rect 21116 3238 21162 3290
rect 21162 3238 21172 3290
rect 21196 3238 21226 3290
rect 21226 3238 21252 3290
rect 20956 3236 21012 3238
rect 21036 3236 21092 3238
rect 21116 3236 21172 3238
rect 21196 3236 21252 3238
rect 20956 2202 21012 2204
rect 21036 2202 21092 2204
rect 21116 2202 21172 2204
rect 21196 2202 21252 2204
rect 20956 2150 20982 2202
rect 20982 2150 21012 2202
rect 21036 2150 21046 2202
rect 21046 2150 21092 2202
rect 21116 2150 21162 2202
rect 21162 2150 21172 2202
rect 21196 2150 21226 2202
rect 21226 2150 21252 2202
rect 20956 2148 21012 2150
rect 21036 2148 21092 2150
rect 21116 2148 21172 2150
rect 21196 2148 21252 2150
rect 21270 1264 21326 1320
<< metal3 >>
rect 23520 23128 24000 23248
rect 0 22992 480 23112
rect 62 22538 122 22992
rect 19977 22674 20043 22677
rect 23614 22674 23674 23128
rect 19977 22672 23674 22674
rect 19977 22616 19982 22672
rect 20038 22616 23674 22672
rect 19977 22614 23674 22616
rect 19977 22611 20043 22614
rect 1301 22538 1367 22541
rect 62 22536 1367 22538
rect 62 22480 1306 22536
rect 1362 22480 1367 22536
rect 62 22478 1367 22480
rect 1301 22475 1367 22478
rect 4944 21792 5264 21793
rect 4944 21728 4952 21792
rect 5016 21728 5032 21792
rect 5096 21728 5112 21792
rect 5176 21728 5192 21792
rect 5256 21728 5264 21792
rect 4944 21727 5264 21728
rect 12944 21792 13264 21793
rect 12944 21728 12952 21792
rect 13016 21728 13032 21792
rect 13096 21728 13112 21792
rect 13176 21728 13192 21792
rect 13256 21728 13264 21792
rect 12944 21727 13264 21728
rect 20944 21792 21264 21793
rect 20944 21728 20952 21792
rect 21016 21728 21032 21792
rect 21096 21728 21112 21792
rect 21176 21728 21192 21792
rect 21256 21728 21264 21792
rect 20944 21727 21264 21728
rect 23520 21632 24000 21752
rect 0 21360 480 21480
rect 62 20906 122 21360
rect 8944 21248 9264 21249
rect 8944 21184 8952 21248
rect 9016 21184 9032 21248
rect 9096 21184 9112 21248
rect 9176 21184 9192 21248
rect 9256 21184 9264 21248
rect 8944 21183 9264 21184
rect 16944 21248 17264 21249
rect 16944 21184 16952 21248
rect 17016 21184 17032 21248
rect 17096 21184 17112 21248
rect 17176 21184 17192 21248
rect 17256 21184 17264 21248
rect 16944 21183 17264 21184
rect 22001 21178 22067 21181
rect 23614 21178 23674 21632
rect 22001 21176 23674 21178
rect 22001 21120 22006 21176
rect 22062 21120 23674 21176
rect 22001 21118 23674 21120
rect 22001 21115 22067 21118
rect 2129 20906 2195 20909
rect 62 20904 2195 20906
rect 62 20848 2134 20904
rect 2190 20848 2195 20904
rect 62 20846 2195 20848
rect 2129 20843 2195 20846
rect 4944 20704 5264 20705
rect 4944 20640 4952 20704
rect 5016 20640 5032 20704
rect 5096 20640 5112 20704
rect 5176 20640 5192 20704
rect 5256 20640 5264 20704
rect 4944 20639 5264 20640
rect 12944 20704 13264 20705
rect 12944 20640 12952 20704
rect 13016 20640 13032 20704
rect 13096 20640 13112 20704
rect 13176 20640 13192 20704
rect 13256 20640 13264 20704
rect 12944 20639 13264 20640
rect 20944 20704 21264 20705
rect 20944 20640 20952 20704
rect 21016 20640 21032 20704
rect 21096 20640 21112 20704
rect 21176 20640 21192 20704
rect 21256 20640 21264 20704
rect 20944 20639 21264 20640
rect 8944 20160 9264 20161
rect 8944 20096 8952 20160
rect 9016 20096 9032 20160
rect 9096 20096 9112 20160
rect 9176 20096 9192 20160
rect 9256 20096 9264 20160
rect 8944 20095 9264 20096
rect 16944 20160 17264 20161
rect 16944 20096 16952 20160
rect 17016 20096 17032 20160
rect 17096 20096 17112 20160
rect 17176 20096 17192 20160
rect 17256 20096 17264 20160
rect 23520 20136 24000 20256
rect 16944 20095 17264 20096
rect 0 19728 480 19848
rect 21265 19818 21331 19821
rect 23614 19818 23674 20136
rect 21265 19816 23674 19818
rect 21265 19760 21270 19816
rect 21326 19760 23674 19816
rect 21265 19758 23674 19760
rect 21265 19755 21331 19758
rect 62 19274 122 19728
rect 4944 19616 5264 19617
rect 4944 19552 4952 19616
rect 5016 19552 5032 19616
rect 5096 19552 5112 19616
rect 5176 19552 5192 19616
rect 5256 19552 5264 19616
rect 4944 19551 5264 19552
rect 12944 19616 13264 19617
rect 12944 19552 12952 19616
rect 13016 19552 13032 19616
rect 13096 19552 13112 19616
rect 13176 19552 13192 19616
rect 13256 19552 13264 19616
rect 12944 19551 13264 19552
rect 20944 19616 21264 19617
rect 20944 19552 20952 19616
rect 21016 19552 21032 19616
rect 21096 19552 21112 19616
rect 21176 19552 21192 19616
rect 21256 19552 21264 19616
rect 20944 19551 21264 19552
rect 1301 19274 1367 19277
rect 62 19272 1367 19274
rect 62 19216 1306 19272
rect 1362 19216 1367 19272
rect 62 19214 1367 19216
rect 1301 19211 1367 19214
rect 8944 19072 9264 19073
rect 8944 19008 8952 19072
rect 9016 19008 9032 19072
rect 9096 19008 9112 19072
rect 9176 19008 9192 19072
rect 9256 19008 9264 19072
rect 8944 19007 9264 19008
rect 16944 19072 17264 19073
rect 16944 19008 16952 19072
rect 17016 19008 17032 19072
rect 17096 19008 17112 19072
rect 17176 19008 17192 19072
rect 17256 19008 17264 19072
rect 16944 19007 17264 19008
rect 23520 18640 24000 18760
rect 4944 18528 5264 18529
rect 4944 18464 4952 18528
rect 5016 18464 5032 18528
rect 5096 18464 5112 18528
rect 5176 18464 5192 18528
rect 5256 18464 5264 18528
rect 4944 18463 5264 18464
rect 12944 18528 13264 18529
rect 12944 18464 12952 18528
rect 13016 18464 13032 18528
rect 13096 18464 13112 18528
rect 13176 18464 13192 18528
rect 13256 18464 13264 18528
rect 12944 18463 13264 18464
rect 20944 18528 21264 18529
rect 20944 18464 20952 18528
rect 21016 18464 21032 18528
rect 21096 18464 21112 18528
rect 21176 18464 21192 18528
rect 21256 18464 21264 18528
rect 20944 18463 21264 18464
rect 0 18232 480 18352
rect 62 17778 122 18232
rect 21081 18186 21147 18189
rect 23614 18186 23674 18640
rect 21081 18184 23674 18186
rect 21081 18128 21086 18184
rect 21142 18128 23674 18184
rect 21081 18126 23674 18128
rect 21081 18123 21147 18126
rect 8944 17984 9264 17985
rect 8944 17920 8952 17984
rect 9016 17920 9032 17984
rect 9096 17920 9112 17984
rect 9176 17920 9192 17984
rect 9256 17920 9264 17984
rect 8944 17919 9264 17920
rect 16944 17984 17264 17985
rect 16944 17920 16952 17984
rect 17016 17920 17032 17984
rect 17096 17920 17112 17984
rect 17176 17920 17192 17984
rect 17256 17920 17264 17984
rect 16944 17919 17264 17920
rect 1301 17778 1367 17781
rect 62 17776 1367 17778
rect 62 17720 1306 17776
rect 1362 17720 1367 17776
rect 62 17718 1367 17720
rect 1301 17715 1367 17718
rect 9857 17642 9923 17645
rect 17861 17642 17927 17645
rect 18873 17642 18939 17645
rect 9857 17640 18939 17642
rect 9857 17584 9862 17640
rect 9918 17584 17866 17640
rect 17922 17584 18878 17640
rect 18934 17584 18939 17640
rect 9857 17582 18939 17584
rect 9857 17579 9923 17582
rect 17861 17579 17927 17582
rect 18873 17579 18939 17582
rect 4944 17440 5264 17441
rect 4944 17376 4952 17440
rect 5016 17376 5032 17440
rect 5096 17376 5112 17440
rect 5176 17376 5192 17440
rect 5256 17376 5264 17440
rect 4944 17375 5264 17376
rect 12944 17440 13264 17441
rect 12944 17376 12952 17440
rect 13016 17376 13032 17440
rect 13096 17376 13112 17440
rect 13176 17376 13192 17440
rect 13256 17376 13264 17440
rect 12944 17375 13264 17376
rect 20944 17440 21264 17441
rect 20944 17376 20952 17440
rect 21016 17376 21032 17440
rect 21096 17376 21112 17440
rect 21176 17376 21192 17440
rect 21256 17376 21264 17440
rect 20944 17375 21264 17376
rect 23520 17144 24000 17264
rect 11789 16962 11855 16965
rect 12617 16962 12683 16965
rect 11789 16960 12683 16962
rect 11789 16904 11794 16960
rect 11850 16904 12622 16960
rect 12678 16904 12683 16960
rect 11789 16902 12683 16904
rect 11789 16899 11855 16902
rect 12617 16899 12683 16902
rect 8944 16896 9264 16897
rect 8944 16832 8952 16896
rect 9016 16832 9032 16896
rect 9096 16832 9112 16896
rect 9176 16832 9192 16896
rect 9256 16832 9264 16896
rect 8944 16831 9264 16832
rect 16944 16896 17264 16897
rect 16944 16832 16952 16896
rect 17016 16832 17032 16896
rect 17096 16832 17112 16896
rect 17176 16832 17192 16896
rect 17256 16832 17264 16896
rect 16944 16831 17264 16832
rect 0 16600 480 16720
rect 21081 16690 21147 16693
rect 23614 16690 23674 17144
rect 21081 16688 23674 16690
rect 21081 16632 21086 16688
rect 21142 16632 23674 16688
rect 21081 16630 23674 16632
rect 21081 16627 21147 16630
rect 62 16282 122 16600
rect 4944 16352 5264 16353
rect 4944 16288 4952 16352
rect 5016 16288 5032 16352
rect 5096 16288 5112 16352
rect 5176 16288 5192 16352
rect 5256 16288 5264 16352
rect 4944 16287 5264 16288
rect 12944 16352 13264 16353
rect 12944 16288 12952 16352
rect 13016 16288 13032 16352
rect 13096 16288 13112 16352
rect 13176 16288 13192 16352
rect 13256 16288 13264 16352
rect 12944 16287 13264 16288
rect 20944 16352 21264 16353
rect 20944 16288 20952 16352
rect 21016 16288 21032 16352
rect 21096 16288 21112 16352
rect 21176 16288 21192 16352
rect 21256 16288 21264 16352
rect 20944 16287 21264 16288
rect 1577 16282 1643 16285
rect 62 16280 1643 16282
rect 62 16224 1582 16280
rect 1638 16224 1643 16280
rect 62 16222 1643 16224
rect 1577 16219 1643 16222
rect 8944 15808 9264 15809
rect 8944 15744 8952 15808
rect 9016 15744 9032 15808
rect 9096 15744 9112 15808
rect 9176 15744 9192 15808
rect 9256 15744 9264 15808
rect 8944 15743 9264 15744
rect 16944 15808 17264 15809
rect 16944 15744 16952 15808
rect 17016 15744 17032 15808
rect 17096 15744 17112 15808
rect 17176 15744 17192 15808
rect 17256 15744 17264 15808
rect 16944 15743 17264 15744
rect 23520 15648 24000 15768
rect 4944 15264 5264 15265
rect 4944 15200 4952 15264
rect 5016 15200 5032 15264
rect 5096 15200 5112 15264
rect 5176 15200 5192 15264
rect 5256 15200 5264 15264
rect 4944 15199 5264 15200
rect 12944 15264 13264 15265
rect 12944 15200 12952 15264
rect 13016 15200 13032 15264
rect 13096 15200 13112 15264
rect 13176 15200 13192 15264
rect 13256 15200 13264 15264
rect 12944 15199 13264 15200
rect 20944 15264 21264 15265
rect 20944 15200 20952 15264
rect 21016 15200 21032 15264
rect 21096 15200 21112 15264
rect 21176 15200 21192 15264
rect 21256 15200 21264 15264
rect 20944 15199 21264 15200
rect 21909 15194 21975 15197
rect 23614 15194 23674 15648
rect 21909 15192 23674 15194
rect 21909 15136 21914 15192
rect 21970 15136 23674 15192
rect 21909 15134 23674 15136
rect 21909 15131 21975 15134
rect 0 14968 480 15088
rect 62 14514 122 14968
rect 8944 14720 9264 14721
rect 8944 14656 8952 14720
rect 9016 14656 9032 14720
rect 9096 14656 9112 14720
rect 9176 14656 9192 14720
rect 9256 14656 9264 14720
rect 8944 14655 9264 14656
rect 16944 14720 17264 14721
rect 16944 14656 16952 14720
rect 17016 14656 17032 14720
rect 17096 14656 17112 14720
rect 17176 14656 17192 14720
rect 17256 14656 17264 14720
rect 16944 14655 17264 14656
rect 4705 14514 4771 14517
rect 62 14512 4771 14514
rect 62 14456 4710 14512
rect 4766 14456 4771 14512
rect 62 14454 4771 14456
rect 4705 14451 4771 14454
rect 4944 14176 5264 14177
rect 4944 14112 4952 14176
rect 5016 14112 5032 14176
rect 5096 14112 5112 14176
rect 5176 14112 5192 14176
rect 5256 14112 5264 14176
rect 4944 14111 5264 14112
rect 12944 14176 13264 14177
rect 12944 14112 12952 14176
rect 13016 14112 13032 14176
rect 13096 14112 13112 14176
rect 13176 14112 13192 14176
rect 13256 14112 13264 14176
rect 12944 14111 13264 14112
rect 20944 14176 21264 14177
rect 20944 14112 20952 14176
rect 21016 14112 21032 14176
rect 21096 14112 21112 14176
rect 21176 14112 21192 14176
rect 21256 14112 21264 14176
rect 23520 14152 24000 14272
rect 20944 14111 21264 14112
rect 20345 13970 20411 13973
rect 23614 13970 23674 14152
rect 20345 13968 23674 13970
rect 20345 13912 20350 13968
rect 20406 13912 23674 13968
rect 20345 13910 23674 13912
rect 20345 13907 20411 13910
rect 11237 13834 11303 13837
rect 11237 13832 17418 13834
rect 11237 13776 11242 13832
rect 11298 13776 17418 13832
rect 11237 13774 17418 13776
rect 11237 13771 11303 13774
rect 17358 13698 17418 13774
rect 21909 13698 21975 13701
rect 17358 13696 21975 13698
rect 17358 13640 21914 13696
rect 21970 13640 21975 13696
rect 17358 13638 21975 13640
rect 21909 13635 21975 13638
rect 8944 13632 9264 13633
rect 8944 13568 8952 13632
rect 9016 13568 9032 13632
rect 9096 13568 9112 13632
rect 9176 13568 9192 13632
rect 9256 13568 9264 13632
rect 8944 13567 9264 13568
rect 16944 13632 17264 13633
rect 16944 13568 16952 13632
rect 17016 13568 17032 13632
rect 17096 13568 17112 13632
rect 17176 13568 17192 13632
rect 17256 13568 17264 13632
rect 16944 13567 17264 13568
rect 0 13424 480 13456
rect 0 13368 18 13424
rect 74 13368 480 13424
rect 0 13336 480 13368
rect 4705 13290 4771 13293
rect 12341 13290 12407 13293
rect 4705 13288 12407 13290
rect 4705 13232 4710 13288
rect 4766 13232 12346 13288
rect 12402 13232 12407 13288
rect 4705 13230 12407 13232
rect 4705 13227 4771 13230
rect 12341 13227 12407 13230
rect 4944 13088 5264 13089
rect 4944 13024 4952 13088
rect 5016 13024 5032 13088
rect 5096 13024 5112 13088
rect 5176 13024 5192 13088
rect 5256 13024 5264 13088
rect 4944 13023 5264 13024
rect 12944 13088 13264 13089
rect 12944 13024 12952 13088
rect 13016 13024 13032 13088
rect 13096 13024 13112 13088
rect 13176 13024 13192 13088
rect 13256 13024 13264 13088
rect 12944 13023 13264 13024
rect 20944 13088 21264 13089
rect 20944 13024 20952 13088
rect 21016 13024 21032 13088
rect 21096 13024 21112 13088
rect 21176 13024 21192 13088
rect 21256 13024 21264 13088
rect 20944 13023 21264 13024
rect 23520 12746 24000 12776
rect 23484 12744 24000 12746
rect 23484 12688 23570 12744
rect 23626 12688 24000 12744
rect 23484 12686 24000 12688
rect 23520 12656 24000 12686
rect 8944 12544 9264 12545
rect 8944 12480 8952 12544
rect 9016 12480 9032 12544
rect 9096 12480 9112 12544
rect 9176 12480 9192 12544
rect 9256 12480 9264 12544
rect 8944 12479 9264 12480
rect 16944 12544 17264 12545
rect 16944 12480 16952 12544
rect 17016 12480 17032 12544
rect 17096 12480 17112 12544
rect 17176 12480 17192 12544
rect 17256 12480 17264 12544
rect 16944 12479 17264 12480
rect 13486 12276 13492 12340
rect 13556 12338 13562 12340
rect 15101 12338 15167 12341
rect 13556 12336 15167 12338
rect 13556 12280 15106 12336
rect 15162 12280 15167 12336
rect 13556 12278 15167 12280
rect 13556 12276 13562 12278
rect 15101 12275 15167 12278
rect 1761 12202 1827 12205
rect 10409 12202 10475 12205
rect 1761 12200 10475 12202
rect 1761 12144 1766 12200
rect 1822 12144 10414 12200
rect 10470 12144 10475 12200
rect 1761 12142 10475 12144
rect 1761 12139 1827 12142
rect 10409 12139 10475 12142
rect 4944 12000 5264 12001
rect 0 11932 480 11960
rect 4944 11936 4952 12000
rect 5016 11936 5032 12000
rect 5096 11936 5112 12000
rect 5176 11936 5192 12000
rect 5256 11936 5264 12000
rect 4944 11935 5264 11936
rect 12944 12000 13264 12001
rect 12944 11936 12952 12000
rect 13016 11936 13032 12000
rect 13096 11936 13112 12000
rect 13176 11936 13192 12000
rect 13256 11936 13264 12000
rect 12944 11935 13264 11936
rect 20944 12000 21264 12001
rect 20944 11936 20952 12000
rect 21016 11936 21032 12000
rect 21096 11936 21112 12000
rect 21176 11936 21192 12000
rect 21256 11936 21264 12000
rect 20944 11935 21264 11936
rect 0 11868 60 11932
rect 124 11868 480 11932
rect 0 11840 480 11868
rect 9949 11794 10015 11797
rect 12065 11794 12131 11797
rect 20713 11794 20779 11797
rect 9949 11792 20779 11794
rect 9949 11736 9954 11792
rect 10010 11736 12070 11792
rect 12126 11736 20718 11792
rect 20774 11736 20779 11792
rect 9949 11734 20779 11736
rect 9949 11731 10015 11734
rect 12065 11731 12131 11734
rect 20713 11731 20779 11734
rect 54 11596 60 11660
rect 124 11658 130 11660
rect 4797 11658 4863 11661
rect 124 11656 4863 11658
rect 124 11600 4802 11656
rect 4858 11600 4863 11656
rect 124 11598 4863 11600
rect 124 11596 130 11598
rect 4797 11595 4863 11598
rect 8944 11456 9264 11457
rect 8944 11392 8952 11456
rect 9016 11392 9032 11456
rect 9096 11392 9112 11456
rect 9176 11392 9192 11456
rect 9256 11392 9264 11456
rect 8944 11391 9264 11392
rect 16944 11456 17264 11457
rect 16944 11392 16952 11456
rect 17016 11392 17032 11456
rect 17096 11392 17112 11456
rect 17176 11392 17192 11456
rect 17256 11392 17264 11456
rect 16944 11391 17264 11392
rect 21265 11250 21331 11253
rect 23520 11250 24000 11280
rect 21265 11248 24000 11250
rect 21265 11192 21270 11248
rect 21326 11192 24000 11248
rect 21265 11190 24000 11192
rect 21265 11187 21331 11190
rect 23520 11160 24000 11190
rect 4944 10912 5264 10913
rect 4944 10848 4952 10912
rect 5016 10848 5032 10912
rect 5096 10848 5112 10912
rect 5176 10848 5192 10912
rect 5256 10848 5264 10912
rect 4944 10847 5264 10848
rect 12944 10912 13264 10913
rect 12944 10848 12952 10912
rect 13016 10848 13032 10912
rect 13096 10848 13112 10912
rect 13176 10848 13192 10912
rect 13256 10848 13264 10912
rect 12944 10847 13264 10848
rect 20944 10912 21264 10913
rect 20944 10848 20952 10912
rect 21016 10848 21032 10912
rect 21096 10848 21112 10912
rect 21176 10848 21192 10912
rect 21256 10848 21264 10912
rect 20944 10847 21264 10848
rect 8944 10368 9264 10369
rect 0 10296 480 10328
rect 8944 10304 8952 10368
rect 9016 10304 9032 10368
rect 9096 10304 9112 10368
rect 9176 10304 9192 10368
rect 9256 10304 9264 10368
rect 8944 10303 9264 10304
rect 16944 10368 17264 10369
rect 16944 10304 16952 10368
rect 17016 10304 17032 10368
rect 17096 10304 17112 10368
rect 17176 10304 17192 10368
rect 17256 10304 17264 10368
rect 16944 10303 17264 10304
rect 0 10240 110 10296
rect 166 10240 480 10296
rect 0 10208 480 10240
rect 1853 10298 1919 10301
rect 8477 10298 8543 10301
rect 1853 10296 8543 10298
rect 1853 10240 1858 10296
rect 1914 10240 8482 10296
rect 8538 10240 8543 10296
rect 1853 10238 8543 10240
rect 1853 10235 1919 10238
rect 8477 10235 8543 10238
rect 4944 9824 5264 9825
rect 4944 9760 4952 9824
rect 5016 9760 5032 9824
rect 5096 9760 5112 9824
rect 5176 9760 5192 9824
rect 5256 9760 5264 9824
rect 4944 9759 5264 9760
rect 12944 9824 13264 9825
rect 12944 9760 12952 9824
rect 13016 9760 13032 9824
rect 13096 9760 13112 9824
rect 13176 9760 13192 9824
rect 13256 9760 13264 9824
rect 12944 9759 13264 9760
rect 20944 9824 21264 9825
rect 20944 9760 20952 9824
rect 21016 9760 21032 9824
rect 21096 9760 21112 9824
rect 21176 9760 21192 9824
rect 21256 9760 21264 9824
rect 20944 9759 21264 9760
rect 13445 9754 13511 9757
rect 15469 9754 15535 9757
rect 13445 9752 15535 9754
rect 13445 9696 13450 9752
rect 13506 9696 15474 9752
rect 15530 9696 15535 9752
rect 13445 9694 15535 9696
rect 13445 9691 13511 9694
rect 15469 9691 15535 9694
rect 21357 9754 21423 9757
rect 23520 9754 24000 9784
rect 21357 9752 24000 9754
rect 21357 9696 21362 9752
rect 21418 9696 24000 9752
rect 21357 9694 24000 9696
rect 21357 9691 21423 9694
rect 23520 9664 24000 9694
rect 105 9618 171 9621
rect 9949 9618 10015 9621
rect 105 9616 10015 9618
rect 105 9560 110 9616
rect 166 9560 9954 9616
rect 10010 9560 10015 9616
rect 105 9558 10015 9560
rect 105 9555 171 9558
rect 9949 9555 10015 9558
rect 13537 9482 13603 9485
rect 18229 9482 18295 9485
rect 13537 9480 18295 9482
rect 13537 9424 13542 9480
rect 13598 9424 18234 9480
rect 18290 9424 18295 9480
rect 13537 9422 18295 9424
rect 13537 9419 13603 9422
rect 18229 9419 18295 9422
rect 2957 9346 3023 9349
rect 8661 9346 8727 9349
rect 2957 9344 8727 9346
rect 2957 9288 2962 9344
rect 3018 9288 8666 9344
rect 8722 9288 8727 9344
rect 2957 9286 8727 9288
rect 2957 9283 3023 9286
rect 8661 9283 8727 9286
rect 9397 9346 9463 9349
rect 9581 9346 9647 9349
rect 13486 9346 13492 9348
rect 9397 9344 13492 9346
rect 9397 9288 9402 9344
rect 9458 9288 9586 9344
rect 9642 9288 13492 9344
rect 9397 9286 13492 9288
rect 9397 9283 9463 9286
rect 9581 9283 9647 9286
rect 13486 9284 13492 9286
rect 13556 9284 13562 9348
rect 8944 9280 9264 9281
rect 8944 9216 8952 9280
rect 9016 9216 9032 9280
rect 9096 9216 9112 9280
rect 9176 9216 9192 9280
rect 9256 9216 9264 9280
rect 8944 9215 9264 9216
rect 16944 9280 17264 9281
rect 16944 9216 16952 9280
rect 17016 9216 17032 9280
rect 17096 9216 17112 9280
rect 17176 9216 17192 9280
rect 17256 9216 17264 9280
rect 16944 9215 17264 9216
rect 11329 9210 11395 9213
rect 13997 9210 14063 9213
rect 11329 9208 14063 9210
rect 11329 9152 11334 9208
rect 11390 9152 14002 9208
rect 14058 9152 14063 9208
rect 11329 9150 14063 9152
rect 11329 9147 11395 9150
rect 13997 9147 14063 9150
rect 8753 8938 8819 8941
rect 14733 8938 14799 8941
rect 8753 8936 14799 8938
rect 8753 8880 8758 8936
rect 8814 8880 14738 8936
rect 14794 8880 14799 8936
rect 8753 8878 14799 8880
rect 8753 8875 8819 8878
rect 14733 8875 14799 8878
rect 4944 8736 5264 8737
rect 0 8664 480 8696
rect 4944 8672 4952 8736
rect 5016 8672 5032 8736
rect 5096 8672 5112 8736
rect 5176 8672 5192 8736
rect 5256 8672 5264 8736
rect 4944 8671 5264 8672
rect 12944 8736 13264 8737
rect 12944 8672 12952 8736
rect 13016 8672 13032 8736
rect 13096 8672 13112 8736
rect 13176 8672 13192 8736
rect 13256 8672 13264 8736
rect 12944 8671 13264 8672
rect 20944 8736 21264 8737
rect 20944 8672 20952 8736
rect 21016 8672 21032 8736
rect 21096 8672 21112 8736
rect 21176 8672 21192 8736
rect 21256 8672 21264 8736
rect 20944 8671 21264 8672
rect 0 8608 110 8664
rect 166 8608 480 8664
rect 0 8576 480 8608
rect 23520 8258 24000 8288
rect 23484 8256 24000 8258
rect 23484 8200 23570 8256
rect 23626 8200 24000 8256
rect 23484 8198 24000 8200
rect 8944 8192 9264 8193
rect 8944 8128 8952 8192
rect 9016 8128 9032 8192
rect 9096 8128 9112 8192
rect 9176 8128 9192 8192
rect 9256 8128 9264 8192
rect 8944 8127 9264 8128
rect 16944 8192 17264 8193
rect 16944 8128 16952 8192
rect 17016 8128 17032 8192
rect 17096 8128 17112 8192
rect 17176 8128 17192 8192
rect 17256 8128 17264 8192
rect 23520 8168 24000 8198
rect 16944 8127 17264 8128
rect 3785 7986 3851 7989
rect 6729 7986 6795 7989
rect 10501 7986 10567 7989
rect 15929 7986 15995 7989
rect 3785 7984 15995 7986
rect 3785 7928 3790 7984
rect 3846 7928 6734 7984
rect 6790 7928 10506 7984
rect 10562 7928 15934 7984
rect 15990 7928 15995 7984
rect 3785 7926 15995 7928
rect 3785 7923 3851 7926
rect 6729 7923 6795 7926
rect 10501 7923 10567 7926
rect 15929 7923 15995 7926
rect 3141 7850 3207 7853
rect 4102 7850 4108 7852
rect 3141 7848 4108 7850
rect 3141 7792 3146 7848
rect 3202 7792 4108 7848
rect 3141 7790 4108 7792
rect 3141 7787 3207 7790
rect 4102 7788 4108 7790
rect 4172 7788 4178 7852
rect 14222 7788 14228 7852
rect 14292 7850 14298 7852
rect 14457 7850 14523 7853
rect 16481 7850 16547 7853
rect 17953 7850 18019 7853
rect 14292 7848 18019 7850
rect 14292 7792 14462 7848
rect 14518 7792 16486 7848
rect 16542 7792 17958 7848
rect 18014 7792 18019 7848
rect 14292 7790 18019 7792
rect 14292 7788 14298 7790
rect 14457 7787 14523 7790
rect 16481 7787 16547 7790
rect 17953 7787 18019 7790
rect 4944 7648 5264 7649
rect 4944 7584 4952 7648
rect 5016 7584 5032 7648
rect 5096 7584 5112 7648
rect 5176 7584 5192 7648
rect 5256 7584 5264 7648
rect 4944 7583 5264 7584
rect 12944 7648 13264 7649
rect 12944 7584 12952 7648
rect 13016 7584 13032 7648
rect 13096 7584 13112 7648
rect 13176 7584 13192 7648
rect 13256 7584 13264 7648
rect 12944 7583 13264 7584
rect 20944 7648 21264 7649
rect 20944 7584 20952 7648
rect 21016 7584 21032 7648
rect 21096 7584 21112 7648
rect 21176 7584 21192 7648
rect 21256 7584 21264 7648
rect 20944 7583 21264 7584
rect 13353 7442 13419 7445
rect 13486 7442 13492 7444
rect 13353 7440 13492 7442
rect 13353 7384 13358 7440
rect 13414 7384 13492 7440
rect 13353 7382 13492 7384
rect 13353 7379 13419 7382
rect 13486 7380 13492 7382
rect 13556 7380 13562 7444
rect 13261 7306 13327 7309
rect 23565 7306 23631 7309
rect 13261 7304 23631 7306
rect 13261 7248 13266 7304
rect 13322 7248 23570 7304
rect 23626 7248 23631 7304
rect 13261 7246 23631 7248
rect 13261 7243 13327 7246
rect 23565 7243 23631 7246
rect 17493 7170 17559 7173
rect 17493 7168 23674 7170
rect 17493 7112 17498 7168
rect 17554 7112 23674 7168
rect 17493 7110 23674 7112
rect 17493 7107 17559 7110
rect 8944 7104 9264 7105
rect 0 7036 480 7064
rect 8944 7040 8952 7104
rect 9016 7040 9032 7104
rect 9096 7040 9112 7104
rect 9176 7040 9192 7104
rect 9256 7040 9264 7104
rect 8944 7039 9264 7040
rect 16944 7104 17264 7105
rect 16944 7040 16952 7104
rect 17016 7040 17032 7104
rect 17096 7040 17112 7104
rect 17176 7040 17192 7104
rect 17256 7040 17264 7104
rect 16944 7039 17264 7040
rect 0 6972 60 7036
rect 124 6972 480 7036
rect 0 6944 480 6972
rect 3969 6898 4035 6901
rect 12525 6898 12591 6901
rect 3969 6896 12591 6898
rect 3969 6840 3974 6896
rect 4030 6840 12530 6896
rect 12586 6840 12591 6896
rect 3969 6838 12591 6840
rect 3969 6835 4035 6838
rect 12525 6835 12591 6838
rect 54 6700 60 6764
rect 124 6762 130 6764
rect 3972 6762 4032 6835
rect 23614 6792 23674 7110
rect 124 6702 4032 6762
rect 124 6700 130 6702
rect 23520 6672 24000 6792
rect 4944 6560 5264 6561
rect 4944 6496 4952 6560
rect 5016 6496 5032 6560
rect 5096 6496 5112 6560
rect 5176 6496 5192 6560
rect 5256 6496 5264 6560
rect 4944 6495 5264 6496
rect 12944 6560 13264 6561
rect 12944 6496 12952 6560
rect 13016 6496 13032 6560
rect 13096 6496 13112 6560
rect 13176 6496 13192 6560
rect 13256 6496 13264 6560
rect 12944 6495 13264 6496
rect 20944 6560 21264 6561
rect 20944 6496 20952 6560
rect 21016 6496 21032 6560
rect 21096 6496 21112 6560
rect 21176 6496 21192 6560
rect 21256 6496 21264 6560
rect 20944 6495 21264 6496
rect 4613 6354 4679 6357
rect 11697 6354 11763 6357
rect 4613 6352 11763 6354
rect 4613 6296 4618 6352
rect 4674 6296 11702 6352
rect 11758 6296 11763 6352
rect 4613 6294 11763 6296
rect 4613 6291 4679 6294
rect 11697 6291 11763 6294
rect 8944 6016 9264 6017
rect 8944 5952 8952 6016
rect 9016 5952 9032 6016
rect 9096 5952 9112 6016
rect 9176 5952 9192 6016
rect 9256 5952 9264 6016
rect 8944 5951 9264 5952
rect 16944 6016 17264 6017
rect 16944 5952 16952 6016
rect 17016 5952 17032 6016
rect 17096 5952 17112 6016
rect 17176 5952 17192 6016
rect 17256 5952 17264 6016
rect 16944 5951 17264 5952
rect 0 5536 480 5568
rect 0 5480 110 5536
rect 166 5480 480 5536
rect 0 5448 480 5480
rect 4944 5472 5264 5473
rect 4944 5408 4952 5472
rect 5016 5408 5032 5472
rect 5096 5408 5112 5472
rect 5176 5408 5192 5472
rect 5256 5408 5264 5472
rect 4944 5407 5264 5408
rect 12944 5472 13264 5473
rect 12944 5408 12952 5472
rect 13016 5408 13032 5472
rect 13096 5408 13112 5472
rect 13176 5408 13192 5472
rect 13256 5408 13264 5472
rect 12944 5407 13264 5408
rect 20944 5472 21264 5473
rect 20944 5408 20952 5472
rect 21016 5408 21032 5472
rect 21096 5408 21112 5472
rect 21176 5408 21192 5472
rect 21256 5408 21264 5472
rect 20944 5407 21264 5408
rect 23520 5266 24000 5296
rect 23484 5264 24000 5266
rect 23484 5208 23570 5264
rect 23626 5208 24000 5264
rect 23484 5206 24000 5208
rect 23520 5176 24000 5206
rect 3509 5130 3575 5133
rect 5809 5130 5875 5133
rect 11329 5130 11395 5133
rect 11881 5130 11947 5133
rect 3509 5128 11947 5130
rect 3509 5072 3514 5128
rect 3570 5072 5814 5128
rect 5870 5072 11334 5128
rect 11390 5072 11886 5128
rect 11942 5072 11947 5128
rect 3509 5070 11947 5072
rect 3509 5067 3575 5070
rect 5809 5067 5875 5070
rect 11329 5067 11395 5070
rect 11881 5067 11947 5070
rect 8944 4928 9264 4929
rect 8944 4864 8952 4928
rect 9016 4864 9032 4928
rect 9096 4864 9112 4928
rect 9176 4864 9192 4928
rect 9256 4864 9264 4928
rect 8944 4863 9264 4864
rect 16944 4928 17264 4929
rect 16944 4864 16952 4928
rect 17016 4864 17032 4928
rect 17096 4864 17112 4928
rect 17176 4864 17192 4928
rect 17256 4864 17264 4928
rect 16944 4863 17264 4864
rect 4944 4384 5264 4385
rect 4944 4320 4952 4384
rect 5016 4320 5032 4384
rect 5096 4320 5112 4384
rect 5176 4320 5192 4384
rect 5256 4320 5264 4384
rect 4944 4319 5264 4320
rect 12944 4384 13264 4385
rect 12944 4320 12952 4384
rect 13016 4320 13032 4384
rect 13096 4320 13112 4384
rect 13176 4320 13192 4384
rect 13256 4320 13264 4384
rect 12944 4319 13264 4320
rect 20944 4384 21264 4385
rect 20944 4320 20952 4384
rect 21016 4320 21032 4384
rect 21096 4320 21112 4384
rect 21176 4320 21192 4384
rect 21256 4320 21264 4384
rect 20944 4319 21264 4320
rect 13445 4042 13511 4045
rect 23565 4042 23631 4045
rect 13445 4040 23631 4042
rect 13445 3984 13450 4040
rect 13506 3984 23570 4040
rect 23626 3984 23631 4040
rect 13445 3982 23631 3984
rect 13445 3979 13511 3982
rect 23565 3979 23631 3982
rect 0 3904 480 3936
rect 0 3848 110 3904
rect 166 3848 480 3904
rect 0 3816 480 3848
rect 8944 3840 9264 3841
rect 8944 3776 8952 3840
rect 9016 3776 9032 3840
rect 9096 3776 9112 3840
rect 9176 3776 9192 3840
rect 9256 3776 9264 3840
rect 8944 3775 9264 3776
rect 16944 3840 17264 3841
rect 16944 3776 16952 3840
rect 17016 3776 17032 3840
rect 17096 3776 17112 3840
rect 17176 3776 17192 3840
rect 17256 3776 17264 3840
rect 16944 3775 17264 3776
rect 23520 3680 24000 3800
rect 4944 3296 5264 3297
rect 4944 3232 4952 3296
rect 5016 3232 5032 3296
rect 5096 3232 5112 3296
rect 5176 3232 5192 3296
rect 5256 3232 5264 3296
rect 4944 3231 5264 3232
rect 12944 3296 13264 3297
rect 12944 3232 12952 3296
rect 13016 3232 13032 3296
rect 13096 3232 13112 3296
rect 13176 3232 13192 3296
rect 13256 3232 13264 3296
rect 12944 3231 13264 3232
rect 20944 3296 21264 3297
rect 20944 3232 20952 3296
rect 21016 3232 21032 3296
rect 21096 3232 21112 3296
rect 21176 3232 21192 3296
rect 21256 3232 21264 3296
rect 20944 3231 21264 3232
rect 8109 2954 8175 2957
rect 23614 2954 23674 3680
rect 8109 2952 23674 2954
rect 8109 2896 8114 2952
rect 8170 2896 23674 2952
rect 8109 2894 23674 2896
rect 8109 2891 8175 2894
rect 8293 2818 8359 2821
rect 62 2816 8359 2818
rect 62 2760 8298 2816
rect 8354 2760 8359 2816
rect 62 2758 8359 2760
rect 62 2304 122 2758
rect 8293 2755 8359 2758
rect 8944 2752 9264 2753
rect 8944 2688 8952 2752
rect 9016 2688 9032 2752
rect 9096 2688 9112 2752
rect 9176 2688 9192 2752
rect 9256 2688 9264 2752
rect 8944 2687 9264 2688
rect 16944 2752 17264 2753
rect 16944 2688 16952 2752
rect 17016 2688 17032 2752
rect 17096 2688 17112 2752
rect 17176 2688 17192 2752
rect 17256 2688 17264 2752
rect 16944 2687 17264 2688
rect 0 2184 480 2304
rect 4944 2208 5264 2209
rect 4944 2144 4952 2208
rect 5016 2144 5032 2208
rect 5096 2144 5112 2208
rect 5176 2144 5192 2208
rect 5256 2144 5264 2208
rect 4944 2143 5264 2144
rect 12944 2208 13264 2209
rect 12944 2144 12952 2208
rect 13016 2144 13032 2208
rect 13096 2144 13112 2208
rect 13176 2144 13192 2208
rect 13256 2144 13264 2208
rect 12944 2143 13264 2144
rect 20944 2208 21264 2209
rect 20944 2144 20952 2208
rect 21016 2144 21032 2208
rect 21096 2144 21112 2208
rect 21176 2144 21192 2208
rect 21256 2144 21264 2208
rect 23520 2184 24000 2304
rect 20944 2143 21264 2144
rect 9857 1730 9923 1733
rect 23614 1730 23674 2184
rect 9857 1728 23674 1730
rect 9857 1672 9862 1728
rect 9918 1672 23674 1728
rect 9857 1670 23674 1672
rect 9857 1667 9923 1670
rect 8569 1594 8635 1597
rect 17125 1594 17191 1597
rect 8569 1592 17191 1594
rect 8569 1536 8574 1592
rect 8630 1536 17130 1592
rect 17186 1536 17191 1592
rect 8569 1534 17191 1536
rect 8569 1531 8635 1534
rect 17125 1531 17191 1534
rect 4153 1322 4219 1325
rect 62 1320 4219 1322
rect 62 1264 4158 1320
rect 4214 1264 4219 1320
rect 62 1262 4219 1264
rect 62 808 122 1262
rect 4153 1259 4219 1262
rect 5901 1322 5967 1325
rect 21265 1322 21331 1325
rect 5901 1320 21331 1322
rect 5901 1264 5906 1320
rect 5962 1264 21270 1320
rect 21326 1264 21331 1320
rect 5901 1262 21331 1264
rect 5901 1259 5967 1262
rect 21265 1259 21331 1262
rect 0 688 480 808
rect 23520 688 24000 808
rect 5349 234 5415 237
rect 23614 234 23674 688
rect 5349 232 23674 234
rect 5349 176 5354 232
rect 5410 176 23674 232
rect 5349 174 23674 176
rect 5349 171 5415 174
<< via3 >>
rect 4952 21788 5016 21792
rect 4952 21732 4956 21788
rect 4956 21732 5012 21788
rect 5012 21732 5016 21788
rect 4952 21728 5016 21732
rect 5032 21788 5096 21792
rect 5032 21732 5036 21788
rect 5036 21732 5092 21788
rect 5092 21732 5096 21788
rect 5032 21728 5096 21732
rect 5112 21788 5176 21792
rect 5112 21732 5116 21788
rect 5116 21732 5172 21788
rect 5172 21732 5176 21788
rect 5112 21728 5176 21732
rect 5192 21788 5256 21792
rect 5192 21732 5196 21788
rect 5196 21732 5252 21788
rect 5252 21732 5256 21788
rect 5192 21728 5256 21732
rect 12952 21788 13016 21792
rect 12952 21732 12956 21788
rect 12956 21732 13012 21788
rect 13012 21732 13016 21788
rect 12952 21728 13016 21732
rect 13032 21788 13096 21792
rect 13032 21732 13036 21788
rect 13036 21732 13092 21788
rect 13092 21732 13096 21788
rect 13032 21728 13096 21732
rect 13112 21788 13176 21792
rect 13112 21732 13116 21788
rect 13116 21732 13172 21788
rect 13172 21732 13176 21788
rect 13112 21728 13176 21732
rect 13192 21788 13256 21792
rect 13192 21732 13196 21788
rect 13196 21732 13252 21788
rect 13252 21732 13256 21788
rect 13192 21728 13256 21732
rect 20952 21788 21016 21792
rect 20952 21732 20956 21788
rect 20956 21732 21012 21788
rect 21012 21732 21016 21788
rect 20952 21728 21016 21732
rect 21032 21788 21096 21792
rect 21032 21732 21036 21788
rect 21036 21732 21092 21788
rect 21092 21732 21096 21788
rect 21032 21728 21096 21732
rect 21112 21788 21176 21792
rect 21112 21732 21116 21788
rect 21116 21732 21172 21788
rect 21172 21732 21176 21788
rect 21112 21728 21176 21732
rect 21192 21788 21256 21792
rect 21192 21732 21196 21788
rect 21196 21732 21252 21788
rect 21252 21732 21256 21788
rect 21192 21728 21256 21732
rect 8952 21244 9016 21248
rect 8952 21188 8956 21244
rect 8956 21188 9012 21244
rect 9012 21188 9016 21244
rect 8952 21184 9016 21188
rect 9032 21244 9096 21248
rect 9032 21188 9036 21244
rect 9036 21188 9092 21244
rect 9092 21188 9096 21244
rect 9032 21184 9096 21188
rect 9112 21244 9176 21248
rect 9112 21188 9116 21244
rect 9116 21188 9172 21244
rect 9172 21188 9176 21244
rect 9112 21184 9176 21188
rect 9192 21244 9256 21248
rect 9192 21188 9196 21244
rect 9196 21188 9252 21244
rect 9252 21188 9256 21244
rect 9192 21184 9256 21188
rect 16952 21244 17016 21248
rect 16952 21188 16956 21244
rect 16956 21188 17012 21244
rect 17012 21188 17016 21244
rect 16952 21184 17016 21188
rect 17032 21244 17096 21248
rect 17032 21188 17036 21244
rect 17036 21188 17092 21244
rect 17092 21188 17096 21244
rect 17032 21184 17096 21188
rect 17112 21244 17176 21248
rect 17112 21188 17116 21244
rect 17116 21188 17172 21244
rect 17172 21188 17176 21244
rect 17112 21184 17176 21188
rect 17192 21244 17256 21248
rect 17192 21188 17196 21244
rect 17196 21188 17252 21244
rect 17252 21188 17256 21244
rect 17192 21184 17256 21188
rect 4952 20700 5016 20704
rect 4952 20644 4956 20700
rect 4956 20644 5012 20700
rect 5012 20644 5016 20700
rect 4952 20640 5016 20644
rect 5032 20700 5096 20704
rect 5032 20644 5036 20700
rect 5036 20644 5092 20700
rect 5092 20644 5096 20700
rect 5032 20640 5096 20644
rect 5112 20700 5176 20704
rect 5112 20644 5116 20700
rect 5116 20644 5172 20700
rect 5172 20644 5176 20700
rect 5112 20640 5176 20644
rect 5192 20700 5256 20704
rect 5192 20644 5196 20700
rect 5196 20644 5252 20700
rect 5252 20644 5256 20700
rect 5192 20640 5256 20644
rect 12952 20700 13016 20704
rect 12952 20644 12956 20700
rect 12956 20644 13012 20700
rect 13012 20644 13016 20700
rect 12952 20640 13016 20644
rect 13032 20700 13096 20704
rect 13032 20644 13036 20700
rect 13036 20644 13092 20700
rect 13092 20644 13096 20700
rect 13032 20640 13096 20644
rect 13112 20700 13176 20704
rect 13112 20644 13116 20700
rect 13116 20644 13172 20700
rect 13172 20644 13176 20700
rect 13112 20640 13176 20644
rect 13192 20700 13256 20704
rect 13192 20644 13196 20700
rect 13196 20644 13252 20700
rect 13252 20644 13256 20700
rect 13192 20640 13256 20644
rect 20952 20700 21016 20704
rect 20952 20644 20956 20700
rect 20956 20644 21012 20700
rect 21012 20644 21016 20700
rect 20952 20640 21016 20644
rect 21032 20700 21096 20704
rect 21032 20644 21036 20700
rect 21036 20644 21092 20700
rect 21092 20644 21096 20700
rect 21032 20640 21096 20644
rect 21112 20700 21176 20704
rect 21112 20644 21116 20700
rect 21116 20644 21172 20700
rect 21172 20644 21176 20700
rect 21112 20640 21176 20644
rect 21192 20700 21256 20704
rect 21192 20644 21196 20700
rect 21196 20644 21252 20700
rect 21252 20644 21256 20700
rect 21192 20640 21256 20644
rect 8952 20156 9016 20160
rect 8952 20100 8956 20156
rect 8956 20100 9012 20156
rect 9012 20100 9016 20156
rect 8952 20096 9016 20100
rect 9032 20156 9096 20160
rect 9032 20100 9036 20156
rect 9036 20100 9092 20156
rect 9092 20100 9096 20156
rect 9032 20096 9096 20100
rect 9112 20156 9176 20160
rect 9112 20100 9116 20156
rect 9116 20100 9172 20156
rect 9172 20100 9176 20156
rect 9112 20096 9176 20100
rect 9192 20156 9256 20160
rect 9192 20100 9196 20156
rect 9196 20100 9252 20156
rect 9252 20100 9256 20156
rect 9192 20096 9256 20100
rect 16952 20156 17016 20160
rect 16952 20100 16956 20156
rect 16956 20100 17012 20156
rect 17012 20100 17016 20156
rect 16952 20096 17016 20100
rect 17032 20156 17096 20160
rect 17032 20100 17036 20156
rect 17036 20100 17092 20156
rect 17092 20100 17096 20156
rect 17032 20096 17096 20100
rect 17112 20156 17176 20160
rect 17112 20100 17116 20156
rect 17116 20100 17172 20156
rect 17172 20100 17176 20156
rect 17112 20096 17176 20100
rect 17192 20156 17256 20160
rect 17192 20100 17196 20156
rect 17196 20100 17252 20156
rect 17252 20100 17256 20156
rect 17192 20096 17256 20100
rect 4952 19612 5016 19616
rect 4952 19556 4956 19612
rect 4956 19556 5012 19612
rect 5012 19556 5016 19612
rect 4952 19552 5016 19556
rect 5032 19612 5096 19616
rect 5032 19556 5036 19612
rect 5036 19556 5092 19612
rect 5092 19556 5096 19612
rect 5032 19552 5096 19556
rect 5112 19612 5176 19616
rect 5112 19556 5116 19612
rect 5116 19556 5172 19612
rect 5172 19556 5176 19612
rect 5112 19552 5176 19556
rect 5192 19612 5256 19616
rect 5192 19556 5196 19612
rect 5196 19556 5252 19612
rect 5252 19556 5256 19612
rect 5192 19552 5256 19556
rect 12952 19612 13016 19616
rect 12952 19556 12956 19612
rect 12956 19556 13012 19612
rect 13012 19556 13016 19612
rect 12952 19552 13016 19556
rect 13032 19612 13096 19616
rect 13032 19556 13036 19612
rect 13036 19556 13092 19612
rect 13092 19556 13096 19612
rect 13032 19552 13096 19556
rect 13112 19612 13176 19616
rect 13112 19556 13116 19612
rect 13116 19556 13172 19612
rect 13172 19556 13176 19612
rect 13112 19552 13176 19556
rect 13192 19612 13256 19616
rect 13192 19556 13196 19612
rect 13196 19556 13252 19612
rect 13252 19556 13256 19612
rect 13192 19552 13256 19556
rect 20952 19612 21016 19616
rect 20952 19556 20956 19612
rect 20956 19556 21012 19612
rect 21012 19556 21016 19612
rect 20952 19552 21016 19556
rect 21032 19612 21096 19616
rect 21032 19556 21036 19612
rect 21036 19556 21092 19612
rect 21092 19556 21096 19612
rect 21032 19552 21096 19556
rect 21112 19612 21176 19616
rect 21112 19556 21116 19612
rect 21116 19556 21172 19612
rect 21172 19556 21176 19612
rect 21112 19552 21176 19556
rect 21192 19612 21256 19616
rect 21192 19556 21196 19612
rect 21196 19556 21252 19612
rect 21252 19556 21256 19612
rect 21192 19552 21256 19556
rect 8952 19068 9016 19072
rect 8952 19012 8956 19068
rect 8956 19012 9012 19068
rect 9012 19012 9016 19068
rect 8952 19008 9016 19012
rect 9032 19068 9096 19072
rect 9032 19012 9036 19068
rect 9036 19012 9092 19068
rect 9092 19012 9096 19068
rect 9032 19008 9096 19012
rect 9112 19068 9176 19072
rect 9112 19012 9116 19068
rect 9116 19012 9172 19068
rect 9172 19012 9176 19068
rect 9112 19008 9176 19012
rect 9192 19068 9256 19072
rect 9192 19012 9196 19068
rect 9196 19012 9252 19068
rect 9252 19012 9256 19068
rect 9192 19008 9256 19012
rect 16952 19068 17016 19072
rect 16952 19012 16956 19068
rect 16956 19012 17012 19068
rect 17012 19012 17016 19068
rect 16952 19008 17016 19012
rect 17032 19068 17096 19072
rect 17032 19012 17036 19068
rect 17036 19012 17092 19068
rect 17092 19012 17096 19068
rect 17032 19008 17096 19012
rect 17112 19068 17176 19072
rect 17112 19012 17116 19068
rect 17116 19012 17172 19068
rect 17172 19012 17176 19068
rect 17112 19008 17176 19012
rect 17192 19068 17256 19072
rect 17192 19012 17196 19068
rect 17196 19012 17252 19068
rect 17252 19012 17256 19068
rect 17192 19008 17256 19012
rect 4952 18524 5016 18528
rect 4952 18468 4956 18524
rect 4956 18468 5012 18524
rect 5012 18468 5016 18524
rect 4952 18464 5016 18468
rect 5032 18524 5096 18528
rect 5032 18468 5036 18524
rect 5036 18468 5092 18524
rect 5092 18468 5096 18524
rect 5032 18464 5096 18468
rect 5112 18524 5176 18528
rect 5112 18468 5116 18524
rect 5116 18468 5172 18524
rect 5172 18468 5176 18524
rect 5112 18464 5176 18468
rect 5192 18524 5256 18528
rect 5192 18468 5196 18524
rect 5196 18468 5252 18524
rect 5252 18468 5256 18524
rect 5192 18464 5256 18468
rect 12952 18524 13016 18528
rect 12952 18468 12956 18524
rect 12956 18468 13012 18524
rect 13012 18468 13016 18524
rect 12952 18464 13016 18468
rect 13032 18524 13096 18528
rect 13032 18468 13036 18524
rect 13036 18468 13092 18524
rect 13092 18468 13096 18524
rect 13032 18464 13096 18468
rect 13112 18524 13176 18528
rect 13112 18468 13116 18524
rect 13116 18468 13172 18524
rect 13172 18468 13176 18524
rect 13112 18464 13176 18468
rect 13192 18524 13256 18528
rect 13192 18468 13196 18524
rect 13196 18468 13252 18524
rect 13252 18468 13256 18524
rect 13192 18464 13256 18468
rect 20952 18524 21016 18528
rect 20952 18468 20956 18524
rect 20956 18468 21012 18524
rect 21012 18468 21016 18524
rect 20952 18464 21016 18468
rect 21032 18524 21096 18528
rect 21032 18468 21036 18524
rect 21036 18468 21092 18524
rect 21092 18468 21096 18524
rect 21032 18464 21096 18468
rect 21112 18524 21176 18528
rect 21112 18468 21116 18524
rect 21116 18468 21172 18524
rect 21172 18468 21176 18524
rect 21112 18464 21176 18468
rect 21192 18524 21256 18528
rect 21192 18468 21196 18524
rect 21196 18468 21252 18524
rect 21252 18468 21256 18524
rect 21192 18464 21256 18468
rect 8952 17980 9016 17984
rect 8952 17924 8956 17980
rect 8956 17924 9012 17980
rect 9012 17924 9016 17980
rect 8952 17920 9016 17924
rect 9032 17980 9096 17984
rect 9032 17924 9036 17980
rect 9036 17924 9092 17980
rect 9092 17924 9096 17980
rect 9032 17920 9096 17924
rect 9112 17980 9176 17984
rect 9112 17924 9116 17980
rect 9116 17924 9172 17980
rect 9172 17924 9176 17980
rect 9112 17920 9176 17924
rect 9192 17980 9256 17984
rect 9192 17924 9196 17980
rect 9196 17924 9252 17980
rect 9252 17924 9256 17980
rect 9192 17920 9256 17924
rect 16952 17980 17016 17984
rect 16952 17924 16956 17980
rect 16956 17924 17012 17980
rect 17012 17924 17016 17980
rect 16952 17920 17016 17924
rect 17032 17980 17096 17984
rect 17032 17924 17036 17980
rect 17036 17924 17092 17980
rect 17092 17924 17096 17980
rect 17032 17920 17096 17924
rect 17112 17980 17176 17984
rect 17112 17924 17116 17980
rect 17116 17924 17172 17980
rect 17172 17924 17176 17980
rect 17112 17920 17176 17924
rect 17192 17980 17256 17984
rect 17192 17924 17196 17980
rect 17196 17924 17252 17980
rect 17252 17924 17256 17980
rect 17192 17920 17256 17924
rect 4952 17436 5016 17440
rect 4952 17380 4956 17436
rect 4956 17380 5012 17436
rect 5012 17380 5016 17436
rect 4952 17376 5016 17380
rect 5032 17436 5096 17440
rect 5032 17380 5036 17436
rect 5036 17380 5092 17436
rect 5092 17380 5096 17436
rect 5032 17376 5096 17380
rect 5112 17436 5176 17440
rect 5112 17380 5116 17436
rect 5116 17380 5172 17436
rect 5172 17380 5176 17436
rect 5112 17376 5176 17380
rect 5192 17436 5256 17440
rect 5192 17380 5196 17436
rect 5196 17380 5252 17436
rect 5252 17380 5256 17436
rect 5192 17376 5256 17380
rect 12952 17436 13016 17440
rect 12952 17380 12956 17436
rect 12956 17380 13012 17436
rect 13012 17380 13016 17436
rect 12952 17376 13016 17380
rect 13032 17436 13096 17440
rect 13032 17380 13036 17436
rect 13036 17380 13092 17436
rect 13092 17380 13096 17436
rect 13032 17376 13096 17380
rect 13112 17436 13176 17440
rect 13112 17380 13116 17436
rect 13116 17380 13172 17436
rect 13172 17380 13176 17436
rect 13112 17376 13176 17380
rect 13192 17436 13256 17440
rect 13192 17380 13196 17436
rect 13196 17380 13252 17436
rect 13252 17380 13256 17436
rect 13192 17376 13256 17380
rect 20952 17436 21016 17440
rect 20952 17380 20956 17436
rect 20956 17380 21012 17436
rect 21012 17380 21016 17436
rect 20952 17376 21016 17380
rect 21032 17436 21096 17440
rect 21032 17380 21036 17436
rect 21036 17380 21092 17436
rect 21092 17380 21096 17436
rect 21032 17376 21096 17380
rect 21112 17436 21176 17440
rect 21112 17380 21116 17436
rect 21116 17380 21172 17436
rect 21172 17380 21176 17436
rect 21112 17376 21176 17380
rect 21192 17436 21256 17440
rect 21192 17380 21196 17436
rect 21196 17380 21252 17436
rect 21252 17380 21256 17436
rect 21192 17376 21256 17380
rect 8952 16892 9016 16896
rect 8952 16836 8956 16892
rect 8956 16836 9012 16892
rect 9012 16836 9016 16892
rect 8952 16832 9016 16836
rect 9032 16892 9096 16896
rect 9032 16836 9036 16892
rect 9036 16836 9092 16892
rect 9092 16836 9096 16892
rect 9032 16832 9096 16836
rect 9112 16892 9176 16896
rect 9112 16836 9116 16892
rect 9116 16836 9172 16892
rect 9172 16836 9176 16892
rect 9112 16832 9176 16836
rect 9192 16892 9256 16896
rect 9192 16836 9196 16892
rect 9196 16836 9252 16892
rect 9252 16836 9256 16892
rect 9192 16832 9256 16836
rect 16952 16892 17016 16896
rect 16952 16836 16956 16892
rect 16956 16836 17012 16892
rect 17012 16836 17016 16892
rect 16952 16832 17016 16836
rect 17032 16892 17096 16896
rect 17032 16836 17036 16892
rect 17036 16836 17092 16892
rect 17092 16836 17096 16892
rect 17032 16832 17096 16836
rect 17112 16892 17176 16896
rect 17112 16836 17116 16892
rect 17116 16836 17172 16892
rect 17172 16836 17176 16892
rect 17112 16832 17176 16836
rect 17192 16892 17256 16896
rect 17192 16836 17196 16892
rect 17196 16836 17252 16892
rect 17252 16836 17256 16892
rect 17192 16832 17256 16836
rect 4952 16348 5016 16352
rect 4952 16292 4956 16348
rect 4956 16292 5012 16348
rect 5012 16292 5016 16348
rect 4952 16288 5016 16292
rect 5032 16348 5096 16352
rect 5032 16292 5036 16348
rect 5036 16292 5092 16348
rect 5092 16292 5096 16348
rect 5032 16288 5096 16292
rect 5112 16348 5176 16352
rect 5112 16292 5116 16348
rect 5116 16292 5172 16348
rect 5172 16292 5176 16348
rect 5112 16288 5176 16292
rect 5192 16348 5256 16352
rect 5192 16292 5196 16348
rect 5196 16292 5252 16348
rect 5252 16292 5256 16348
rect 5192 16288 5256 16292
rect 12952 16348 13016 16352
rect 12952 16292 12956 16348
rect 12956 16292 13012 16348
rect 13012 16292 13016 16348
rect 12952 16288 13016 16292
rect 13032 16348 13096 16352
rect 13032 16292 13036 16348
rect 13036 16292 13092 16348
rect 13092 16292 13096 16348
rect 13032 16288 13096 16292
rect 13112 16348 13176 16352
rect 13112 16292 13116 16348
rect 13116 16292 13172 16348
rect 13172 16292 13176 16348
rect 13112 16288 13176 16292
rect 13192 16348 13256 16352
rect 13192 16292 13196 16348
rect 13196 16292 13252 16348
rect 13252 16292 13256 16348
rect 13192 16288 13256 16292
rect 20952 16348 21016 16352
rect 20952 16292 20956 16348
rect 20956 16292 21012 16348
rect 21012 16292 21016 16348
rect 20952 16288 21016 16292
rect 21032 16348 21096 16352
rect 21032 16292 21036 16348
rect 21036 16292 21092 16348
rect 21092 16292 21096 16348
rect 21032 16288 21096 16292
rect 21112 16348 21176 16352
rect 21112 16292 21116 16348
rect 21116 16292 21172 16348
rect 21172 16292 21176 16348
rect 21112 16288 21176 16292
rect 21192 16348 21256 16352
rect 21192 16292 21196 16348
rect 21196 16292 21252 16348
rect 21252 16292 21256 16348
rect 21192 16288 21256 16292
rect 8952 15804 9016 15808
rect 8952 15748 8956 15804
rect 8956 15748 9012 15804
rect 9012 15748 9016 15804
rect 8952 15744 9016 15748
rect 9032 15804 9096 15808
rect 9032 15748 9036 15804
rect 9036 15748 9092 15804
rect 9092 15748 9096 15804
rect 9032 15744 9096 15748
rect 9112 15804 9176 15808
rect 9112 15748 9116 15804
rect 9116 15748 9172 15804
rect 9172 15748 9176 15804
rect 9112 15744 9176 15748
rect 9192 15804 9256 15808
rect 9192 15748 9196 15804
rect 9196 15748 9252 15804
rect 9252 15748 9256 15804
rect 9192 15744 9256 15748
rect 16952 15804 17016 15808
rect 16952 15748 16956 15804
rect 16956 15748 17012 15804
rect 17012 15748 17016 15804
rect 16952 15744 17016 15748
rect 17032 15804 17096 15808
rect 17032 15748 17036 15804
rect 17036 15748 17092 15804
rect 17092 15748 17096 15804
rect 17032 15744 17096 15748
rect 17112 15804 17176 15808
rect 17112 15748 17116 15804
rect 17116 15748 17172 15804
rect 17172 15748 17176 15804
rect 17112 15744 17176 15748
rect 17192 15804 17256 15808
rect 17192 15748 17196 15804
rect 17196 15748 17252 15804
rect 17252 15748 17256 15804
rect 17192 15744 17256 15748
rect 4952 15260 5016 15264
rect 4952 15204 4956 15260
rect 4956 15204 5012 15260
rect 5012 15204 5016 15260
rect 4952 15200 5016 15204
rect 5032 15260 5096 15264
rect 5032 15204 5036 15260
rect 5036 15204 5092 15260
rect 5092 15204 5096 15260
rect 5032 15200 5096 15204
rect 5112 15260 5176 15264
rect 5112 15204 5116 15260
rect 5116 15204 5172 15260
rect 5172 15204 5176 15260
rect 5112 15200 5176 15204
rect 5192 15260 5256 15264
rect 5192 15204 5196 15260
rect 5196 15204 5252 15260
rect 5252 15204 5256 15260
rect 5192 15200 5256 15204
rect 12952 15260 13016 15264
rect 12952 15204 12956 15260
rect 12956 15204 13012 15260
rect 13012 15204 13016 15260
rect 12952 15200 13016 15204
rect 13032 15260 13096 15264
rect 13032 15204 13036 15260
rect 13036 15204 13092 15260
rect 13092 15204 13096 15260
rect 13032 15200 13096 15204
rect 13112 15260 13176 15264
rect 13112 15204 13116 15260
rect 13116 15204 13172 15260
rect 13172 15204 13176 15260
rect 13112 15200 13176 15204
rect 13192 15260 13256 15264
rect 13192 15204 13196 15260
rect 13196 15204 13252 15260
rect 13252 15204 13256 15260
rect 13192 15200 13256 15204
rect 20952 15260 21016 15264
rect 20952 15204 20956 15260
rect 20956 15204 21012 15260
rect 21012 15204 21016 15260
rect 20952 15200 21016 15204
rect 21032 15260 21096 15264
rect 21032 15204 21036 15260
rect 21036 15204 21092 15260
rect 21092 15204 21096 15260
rect 21032 15200 21096 15204
rect 21112 15260 21176 15264
rect 21112 15204 21116 15260
rect 21116 15204 21172 15260
rect 21172 15204 21176 15260
rect 21112 15200 21176 15204
rect 21192 15260 21256 15264
rect 21192 15204 21196 15260
rect 21196 15204 21252 15260
rect 21252 15204 21256 15260
rect 21192 15200 21256 15204
rect 8952 14716 9016 14720
rect 8952 14660 8956 14716
rect 8956 14660 9012 14716
rect 9012 14660 9016 14716
rect 8952 14656 9016 14660
rect 9032 14716 9096 14720
rect 9032 14660 9036 14716
rect 9036 14660 9092 14716
rect 9092 14660 9096 14716
rect 9032 14656 9096 14660
rect 9112 14716 9176 14720
rect 9112 14660 9116 14716
rect 9116 14660 9172 14716
rect 9172 14660 9176 14716
rect 9112 14656 9176 14660
rect 9192 14716 9256 14720
rect 9192 14660 9196 14716
rect 9196 14660 9252 14716
rect 9252 14660 9256 14716
rect 9192 14656 9256 14660
rect 16952 14716 17016 14720
rect 16952 14660 16956 14716
rect 16956 14660 17012 14716
rect 17012 14660 17016 14716
rect 16952 14656 17016 14660
rect 17032 14716 17096 14720
rect 17032 14660 17036 14716
rect 17036 14660 17092 14716
rect 17092 14660 17096 14716
rect 17032 14656 17096 14660
rect 17112 14716 17176 14720
rect 17112 14660 17116 14716
rect 17116 14660 17172 14716
rect 17172 14660 17176 14716
rect 17112 14656 17176 14660
rect 17192 14716 17256 14720
rect 17192 14660 17196 14716
rect 17196 14660 17252 14716
rect 17252 14660 17256 14716
rect 17192 14656 17256 14660
rect 4952 14172 5016 14176
rect 4952 14116 4956 14172
rect 4956 14116 5012 14172
rect 5012 14116 5016 14172
rect 4952 14112 5016 14116
rect 5032 14172 5096 14176
rect 5032 14116 5036 14172
rect 5036 14116 5092 14172
rect 5092 14116 5096 14172
rect 5032 14112 5096 14116
rect 5112 14172 5176 14176
rect 5112 14116 5116 14172
rect 5116 14116 5172 14172
rect 5172 14116 5176 14172
rect 5112 14112 5176 14116
rect 5192 14172 5256 14176
rect 5192 14116 5196 14172
rect 5196 14116 5252 14172
rect 5252 14116 5256 14172
rect 5192 14112 5256 14116
rect 12952 14172 13016 14176
rect 12952 14116 12956 14172
rect 12956 14116 13012 14172
rect 13012 14116 13016 14172
rect 12952 14112 13016 14116
rect 13032 14172 13096 14176
rect 13032 14116 13036 14172
rect 13036 14116 13092 14172
rect 13092 14116 13096 14172
rect 13032 14112 13096 14116
rect 13112 14172 13176 14176
rect 13112 14116 13116 14172
rect 13116 14116 13172 14172
rect 13172 14116 13176 14172
rect 13112 14112 13176 14116
rect 13192 14172 13256 14176
rect 13192 14116 13196 14172
rect 13196 14116 13252 14172
rect 13252 14116 13256 14172
rect 13192 14112 13256 14116
rect 20952 14172 21016 14176
rect 20952 14116 20956 14172
rect 20956 14116 21012 14172
rect 21012 14116 21016 14172
rect 20952 14112 21016 14116
rect 21032 14172 21096 14176
rect 21032 14116 21036 14172
rect 21036 14116 21092 14172
rect 21092 14116 21096 14172
rect 21032 14112 21096 14116
rect 21112 14172 21176 14176
rect 21112 14116 21116 14172
rect 21116 14116 21172 14172
rect 21172 14116 21176 14172
rect 21112 14112 21176 14116
rect 21192 14172 21256 14176
rect 21192 14116 21196 14172
rect 21196 14116 21252 14172
rect 21252 14116 21256 14172
rect 21192 14112 21256 14116
rect 8952 13628 9016 13632
rect 8952 13572 8956 13628
rect 8956 13572 9012 13628
rect 9012 13572 9016 13628
rect 8952 13568 9016 13572
rect 9032 13628 9096 13632
rect 9032 13572 9036 13628
rect 9036 13572 9092 13628
rect 9092 13572 9096 13628
rect 9032 13568 9096 13572
rect 9112 13628 9176 13632
rect 9112 13572 9116 13628
rect 9116 13572 9172 13628
rect 9172 13572 9176 13628
rect 9112 13568 9176 13572
rect 9192 13628 9256 13632
rect 9192 13572 9196 13628
rect 9196 13572 9252 13628
rect 9252 13572 9256 13628
rect 9192 13568 9256 13572
rect 16952 13628 17016 13632
rect 16952 13572 16956 13628
rect 16956 13572 17012 13628
rect 17012 13572 17016 13628
rect 16952 13568 17016 13572
rect 17032 13628 17096 13632
rect 17032 13572 17036 13628
rect 17036 13572 17092 13628
rect 17092 13572 17096 13628
rect 17032 13568 17096 13572
rect 17112 13628 17176 13632
rect 17112 13572 17116 13628
rect 17116 13572 17172 13628
rect 17172 13572 17176 13628
rect 17112 13568 17176 13572
rect 17192 13628 17256 13632
rect 17192 13572 17196 13628
rect 17196 13572 17252 13628
rect 17252 13572 17256 13628
rect 17192 13568 17256 13572
rect 4952 13084 5016 13088
rect 4952 13028 4956 13084
rect 4956 13028 5012 13084
rect 5012 13028 5016 13084
rect 4952 13024 5016 13028
rect 5032 13084 5096 13088
rect 5032 13028 5036 13084
rect 5036 13028 5092 13084
rect 5092 13028 5096 13084
rect 5032 13024 5096 13028
rect 5112 13084 5176 13088
rect 5112 13028 5116 13084
rect 5116 13028 5172 13084
rect 5172 13028 5176 13084
rect 5112 13024 5176 13028
rect 5192 13084 5256 13088
rect 5192 13028 5196 13084
rect 5196 13028 5252 13084
rect 5252 13028 5256 13084
rect 5192 13024 5256 13028
rect 12952 13084 13016 13088
rect 12952 13028 12956 13084
rect 12956 13028 13012 13084
rect 13012 13028 13016 13084
rect 12952 13024 13016 13028
rect 13032 13084 13096 13088
rect 13032 13028 13036 13084
rect 13036 13028 13092 13084
rect 13092 13028 13096 13084
rect 13032 13024 13096 13028
rect 13112 13084 13176 13088
rect 13112 13028 13116 13084
rect 13116 13028 13172 13084
rect 13172 13028 13176 13084
rect 13112 13024 13176 13028
rect 13192 13084 13256 13088
rect 13192 13028 13196 13084
rect 13196 13028 13252 13084
rect 13252 13028 13256 13084
rect 13192 13024 13256 13028
rect 20952 13084 21016 13088
rect 20952 13028 20956 13084
rect 20956 13028 21012 13084
rect 21012 13028 21016 13084
rect 20952 13024 21016 13028
rect 21032 13084 21096 13088
rect 21032 13028 21036 13084
rect 21036 13028 21092 13084
rect 21092 13028 21096 13084
rect 21032 13024 21096 13028
rect 21112 13084 21176 13088
rect 21112 13028 21116 13084
rect 21116 13028 21172 13084
rect 21172 13028 21176 13084
rect 21112 13024 21176 13028
rect 21192 13084 21256 13088
rect 21192 13028 21196 13084
rect 21196 13028 21252 13084
rect 21252 13028 21256 13084
rect 21192 13024 21256 13028
rect 8952 12540 9016 12544
rect 8952 12484 8956 12540
rect 8956 12484 9012 12540
rect 9012 12484 9016 12540
rect 8952 12480 9016 12484
rect 9032 12540 9096 12544
rect 9032 12484 9036 12540
rect 9036 12484 9092 12540
rect 9092 12484 9096 12540
rect 9032 12480 9096 12484
rect 9112 12540 9176 12544
rect 9112 12484 9116 12540
rect 9116 12484 9172 12540
rect 9172 12484 9176 12540
rect 9112 12480 9176 12484
rect 9192 12540 9256 12544
rect 9192 12484 9196 12540
rect 9196 12484 9252 12540
rect 9252 12484 9256 12540
rect 9192 12480 9256 12484
rect 16952 12540 17016 12544
rect 16952 12484 16956 12540
rect 16956 12484 17012 12540
rect 17012 12484 17016 12540
rect 16952 12480 17016 12484
rect 17032 12540 17096 12544
rect 17032 12484 17036 12540
rect 17036 12484 17092 12540
rect 17092 12484 17096 12540
rect 17032 12480 17096 12484
rect 17112 12540 17176 12544
rect 17112 12484 17116 12540
rect 17116 12484 17172 12540
rect 17172 12484 17176 12540
rect 17112 12480 17176 12484
rect 17192 12540 17256 12544
rect 17192 12484 17196 12540
rect 17196 12484 17252 12540
rect 17252 12484 17256 12540
rect 17192 12480 17256 12484
rect 13492 12276 13556 12340
rect 4952 11996 5016 12000
rect 4952 11940 4956 11996
rect 4956 11940 5012 11996
rect 5012 11940 5016 11996
rect 4952 11936 5016 11940
rect 5032 11996 5096 12000
rect 5032 11940 5036 11996
rect 5036 11940 5092 11996
rect 5092 11940 5096 11996
rect 5032 11936 5096 11940
rect 5112 11996 5176 12000
rect 5112 11940 5116 11996
rect 5116 11940 5172 11996
rect 5172 11940 5176 11996
rect 5112 11936 5176 11940
rect 5192 11996 5256 12000
rect 5192 11940 5196 11996
rect 5196 11940 5252 11996
rect 5252 11940 5256 11996
rect 5192 11936 5256 11940
rect 12952 11996 13016 12000
rect 12952 11940 12956 11996
rect 12956 11940 13012 11996
rect 13012 11940 13016 11996
rect 12952 11936 13016 11940
rect 13032 11996 13096 12000
rect 13032 11940 13036 11996
rect 13036 11940 13092 11996
rect 13092 11940 13096 11996
rect 13032 11936 13096 11940
rect 13112 11996 13176 12000
rect 13112 11940 13116 11996
rect 13116 11940 13172 11996
rect 13172 11940 13176 11996
rect 13112 11936 13176 11940
rect 13192 11996 13256 12000
rect 13192 11940 13196 11996
rect 13196 11940 13252 11996
rect 13252 11940 13256 11996
rect 13192 11936 13256 11940
rect 20952 11996 21016 12000
rect 20952 11940 20956 11996
rect 20956 11940 21012 11996
rect 21012 11940 21016 11996
rect 20952 11936 21016 11940
rect 21032 11996 21096 12000
rect 21032 11940 21036 11996
rect 21036 11940 21092 11996
rect 21092 11940 21096 11996
rect 21032 11936 21096 11940
rect 21112 11996 21176 12000
rect 21112 11940 21116 11996
rect 21116 11940 21172 11996
rect 21172 11940 21176 11996
rect 21112 11936 21176 11940
rect 21192 11996 21256 12000
rect 21192 11940 21196 11996
rect 21196 11940 21252 11996
rect 21252 11940 21256 11996
rect 21192 11936 21256 11940
rect 60 11868 124 11932
rect 60 11596 124 11660
rect 8952 11452 9016 11456
rect 8952 11396 8956 11452
rect 8956 11396 9012 11452
rect 9012 11396 9016 11452
rect 8952 11392 9016 11396
rect 9032 11452 9096 11456
rect 9032 11396 9036 11452
rect 9036 11396 9092 11452
rect 9092 11396 9096 11452
rect 9032 11392 9096 11396
rect 9112 11452 9176 11456
rect 9112 11396 9116 11452
rect 9116 11396 9172 11452
rect 9172 11396 9176 11452
rect 9112 11392 9176 11396
rect 9192 11452 9256 11456
rect 9192 11396 9196 11452
rect 9196 11396 9252 11452
rect 9252 11396 9256 11452
rect 9192 11392 9256 11396
rect 16952 11452 17016 11456
rect 16952 11396 16956 11452
rect 16956 11396 17012 11452
rect 17012 11396 17016 11452
rect 16952 11392 17016 11396
rect 17032 11452 17096 11456
rect 17032 11396 17036 11452
rect 17036 11396 17092 11452
rect 17092 11396 17096 11452
rect 17032 11392 17096 11396
rect 17112 11452 17176 11456
rect 17112 11396 17116 11452
rect 17116 11396 17172 11452
rect 17172 11396 17176 11452
rect 17112 11392 17176 11396
rect 17192 11452 17256 11456
rect 17192 11396 17196 11452
rect 17196 11396 17252 11452
rect 17252 11396 17256 11452
rect 17192 11392 17256 11396
rect 4952 10908 5016 10912
rect 4952 10852 4956 10908
rect 4956 10852 5012 10908
rect 5012 10852 5016 10908
rect 4952 10848 5016 10852
rect 5032 10908 5096 10912
rect 5032 10852 5036 10908
rect 5036 10852 5092 10908
rect 5092 10852 5096 10908
rect 5032 10848 5096 10852
rect 5112 10908 5176 10912
rect 5112 10852 5116 10908
rect 5116 10852 5172 10908
rect 5172 10852 5176 10908
rect 5112 10848 5176 10852
rect 5192 10908 5256 10912
rect 5192 10852 5196 10908
rect 5196 10852 5252 10908
rect 5252 10852 5256 10908
rect 5192 10848 5256 10852
rect 12952 10908 13016 10912
rect 12952 10852 12956 10908
rect 12956 10852 13012 10908
rect 13012 10852 13016 10908
rect 12952 10848 13016 10852
rect 13032 10908 13096 10912
rect 13032 10852 13036 10908
rect 13036 10852 13092 10908
rect 13092 10852 13096 10908
rect 13032 10848 13096 10852
rect 13112 10908 13176 10912
rect 13112 10852 13116 10908
rect 13116 10852 13172 10908
rect 13172 10852 13176 10908
rect 13112 10848 13176 10852
rect 13192 10908 13256 10912
rect 13192 10852 13196 10908
rect 13196 10852 13252 10908
rect 13252 10852 13256 10908
rect 13192 10848 13256 10852
rect 20952 10908 21016 10912
rect 20952 10852 20956 10908
rect 20956 10852 21012 10908
rect 21012 10852 21016 10908
rect 20952 10848 21016 10852
rect 21032 10908 21096 10912
rect 21032 10852 21036 10908
rect 21036 10852 21092 10908
rect 21092 10852 21096 10908
rect 21032 10848 21096 10852
rect 21112 10908 21176 10912
rect 21112 10852 21116 10908
rect 21116 10852 21172 10908
rect 21172 10852 21176 10908
rect 21112 10848 21176 10852
rect 21192 10908 21256 10912
rect 21192 10852 21196 10908
rect 21196 10852 21252 10908
rect 21252 10852 21256 10908
rect 21192 10848 21256 10852
rect 8952 10364 9016 10368
rect 8952 10308 8956 10364
rect 8956 10308 9012 10364
rect 9012 10308 9016 10364
rect 8952 10304 9016 10308
rect 9032 10364 9096 10368
rect 9032 10308 9036 10364
rect 9036 10308 9092 10364
rect 9092 10308 9096 10364
rect 9032 10304 9096 10308
rect 9112 10364 9176 10368
rect 9112 10308 9116 10364
rect 9116 10308 9172 10364
rect 9172 10308 9176 10364
rect 9112 10304 9176 10308
rect 9192 10364 9256 10368
rect 9192 10308 9196 10364
rect 9196 10308 9252 10364
rect 9252 10308 9256 10364
rect 9192 10304 9256 10308
rect 16952 10364 17016 10368
rect 16952 10308 16956 10364
rect 16956 10308 17012 10364
rect 17012 10308 17016 10364
rect 16952 10304 17016 10308
rect 17032 10364 17096 10368
rect 17032 10308 17036 10364
rect 17036 10308 17092 10364
rect 17092 10308 17096 10364
rect 17032 10304 17096 10308
rect 17112 10364 17176 10368
rect 17112 10308 17116 10364
rect 17116 10308 17172 10364
rect 17172 10308 17176 10364
rect 17112 10304 17176 10308
rect 17192 10364 17256 10368
rect 17192 10308 17196 10364
rect 17196 10308 17252 10364
rect 17252 10308 17256 10364
rect 17192 10304 17256 10308
rect 4952 9820 5016 9824
rect 4952 9764 4956 9820
rect 4956 9764 5012 9820
rect 5012 9764 5016 9820
rect 4952 9760 5016 9764
rect 5032 9820 5096 9824
rect 5032 9764 5036 9820
rect 5036 9764 5092 9820
rect 5092 9764 5096 9820
rect 5032 9760 5096 9764
rect 5112 9820 5176 9824
rect 5112 9764 5116 9820
rect 5116 9764 5172 9820
rect 5172 9764 5176 9820
rect 5112 9760 5176 9764
rect 5192 9820 5256 9824
rect 5192 9764 5196 9820
rect 5196 9764 5252 9820
rect 5252 9764 5256 9820
rect 5192 9760 5256 9764
rect 12952 9820 13016 9824
rect 12952 9764 12956 9820
rect 12956 9764 13012 9820
rect 13012 9764 13016 9820
rect 12952 9760 13016 9764
rect 13032 9820 13096 9824
rect 13032 9764 13036 9820
rect 13036 9764 13092 9820
rect 13092 9764 13096 9820
rect 13032 9760 13096 9764
rect 13112 9820 13176 9824
rect 13112 9764 13116 9820
rect 13116 9764 13172 9820
rect 13172 9764 13176 9820
rect 13112 9760 13176 9764
rect 13192 9820 13256 9824
rect 13192 9764 13196 9820
rect 13196 9764 13252 9820
rect 13252 9764 13256 9820
rect 13192 9760 13256 9764
rect 20952 9820 21016 9824
rect 20952 9764 20956 9820
rect 20956 9764 21012 9820
rect 21012 9764 21016 9820
rect 20952 9760 21016 9764
rect 21032 9820 21096 9824
rect 21032 9764 21036 9820
rect 21036 9764 21092 9820
rect 21092 9764 21096 9820
rect 21032 9760 21096 9764
rect 21112 9820 21176 9824
rect 21112 9764 21116 9820
rect 21116 9764 21172 9820
rect 21172 9764 21176 9820
rect 21112 9760 21176 9764
rect 21192 9820 21256 9824
rect 21192 9764 21196 9820
rect 21196 9764 21252 9820
rect 21252 9764 21256 9820
rect 21192 9760 21256 9764
rect 13492 9284 13556 9348
rect 8952 9276 9016 9280
rect 8952 9220 8956 9276
rect 8956 9220 9012 9276
rect 9012 9220 9016 9276
rect 8952 9216 9016 9220
rect 9032 9276 9096 9280
rect 9032 9220 9036 9276
rect 9036 9220 9092 9276
rect 9092 9220 9096 9276
rect 9032 9216 9096 9220
rect 9112 9276 9176 9280
rect 9112 9220 9116 9276
rect 9116 9220 9172 9276
rect 9172 9220 9176 9276
rect 9112 9216 9176 9220
rect 9192 9276 9256 9280
rect 9192 9220 9196 9276
rect 9196 9220 9252 9276
rect 9252 9220 9256 9276
rect 9192 9216 9256 9220
rect 16952 9276 17016 9280
rect 16952 9220 16956 9276
rect 16956 9220 17012 9276
rect 17012 9220 17016 9276
rect 16952 9216 17016 9220
rect 17032 9276 17096 9280
rect 17032 9220 17036 9276
rect 17036 9220 17092 9276
rect 17092 9220 17096 9276
rect 17032 9216 17096 9220
rect 17112 9276 17176 9280
rect 17112 9220 17116 9276
rect 17116 9220 17172 9276
rect 17172 9220 17176 9276
rect 17112 9216 17176 9220
rect 17192 9276 17256 9280
rect 17192 9220 17196 9276
rect 17196 9220 17252 9276
rect 17252 9220 17256 9276
rect 17192 9216 17256 9220
rect 4952 8732 5016 8736
rect 4952 8676 4956 8732
rect 4956 8676 5012 8732
rect 5012 8676 5016 8732
rect 4952 8672 5016 8676
rect 5032 8732 5096 8736
rect 5032 8676 5036 8732
rect 5036 8676 5092 8732
rect 5092 8676 5096 8732
rect 5032 8672 5096 8676
rect 5112 8732 5176 8736
rect 5112 8676 5116 8732
rect 5116 8676 5172 8732
rect 5172 8676 5176 8732
rect 5112 8672 5176 8676
rect 5192 8732 5256 8736
rect 5192 8676 5196 8732
rect 5196 8676 5252 8732
rect 5252 8676 5256 8732
rect 5192 8672 5256 8676
rect 12952 8732 13016 8736
rect 12952 8676 12956 8732
rect 12956 8676 13012 8732
rect 13012 8676 13016 8732
rect 12952 8672 13016 8676
rect 13032 8732 13096 8736
rect 13032 8676 13036 8732
rect 13036 8676 13092 8732
rect 13092 8676 13096 8732
rect 13032 8672 13096 8676
rect 13112 8732 13176 8736
rect 13112 8676 13116 8732
rect 13116 8676 13172 8732
rect 13172 8676 13176 8732
rect 13112 8672 13176 8676
rect 13192 8732 13256 8736
rect 13192 8676 13196 8732
rect 13196 8676 13252 8732
rect 13252 8676 13256 8732
rect 13192 8672 13256 8676
rect 20952 8732 21016 8736
rect 20952 8676 20956 8732
rect 20956 8676 21012 8732
rect 21012 8676 21016 8732
rect 20952 8672 21016 8676
rect 21032 8732 21096 8736
rect 21032 8676 21036 8732
rect 21036 8676 21092 8732
rect 21092 8676 21096 8732
rect 21032 8672 21096 8676
rect 21112 8732 21176 8736
rect 21112 8676 21116 8732
rect 21116 8676 21172 8732
rect 21172 8676 21176 8732
rect 21112 8672 21176 8676
rect 21192 8732 21256 8736
rect 21192 8676 21196 8732
rect 21196 8676 21252 8732
rect 21252 8676 21256 8732
rect 21192 8672 21256 8676
rect 8952 8188 9016 8192
rect 8952 8132 8956 8188
rect 8956 8132 9012 8188
rect 9012 8132 9016 8188
rect 8952 8128 9016 8132
rect 9032 8188 9096 8192
rect 9032 8132 9036 8188
rect 9036 8132 9092 8188
rect 9092 8132 9096 8188
rect 9032 8128 9096 8132
rect 9112 8188 9176 8192
rect 9112 8132 9116 8188
rect 9116 8132 9172 8188
rect 9172 8132 9176 8188
rect 9112 8128 9176 8132
rect 9192 8188 9256 8192
rect 9192 8132 9196 8188
rect 9196 8132 9252 8188
rect 9252 8132 9256 8188
rect 9192 8128 9256 8132
rect 16952 8188 17016 8192
rect 16952 8132 16956 8188
rect 16956 8132 17012 8188
rect 17012 8132 17016 8188
rect 16952 8128 17016 8132
rect 17032 8188 17096 8192
rect 17032 8132 17036 8188
rect 17036 8132 17092 8188
rect 17092 8132 17096 8188
rect 17032 8128 17096 8132
rect 17112 8188 17176 8192
rect 17112 8132 17116 8188
rect 17116 8132 17172 8188
rect 17172 8132 17176 8188
rect 17112 8128 17176 8132
rect 17192 8188 17256 8192
rect 17192 8132 17196 8188
rect 17196 8132 17252 8188
rect 17252 8132 17256 8188
rect 17192 8128 17256 8132
rect 4108 7788 4172 7852
rect 14228 7788 14292 7852
rect 4952 7644 5016 7648
rect 4952 7588 4956 7644
rect 4956 7588 5012 7644
rect 5012 7588 5016 7644
rect 4952 7584 5016 7588
rect 5032 7644 5096 7648
rect 5032 7588 5036 7644
rect 5036 7588 5092 7644
rect 5092 7588 5096 7644
rect 5032 7584 5096 7588
rect 5112 7644 5176 7648
rect 5112 7588 5116 7644
rect 5116 7588 5172 7644
rect 5172 7588 5176 7644
rect 5112 7584 5176 7588
rect 5192 7644 5256 7648
rect 5192 7588 5196 7644
rect 5196 7588 5252 7644
rect 5252 7588 5256 7644
rect 5192 7584 5256 7588
rect 12952 7644 13016 7648
rect 12952 7588 12956 7644
rect 12956 7588 13012 7644
rect 13012 7588 13016 7644
rect 12952 7584 13016 7588
rect 13032 7644 13096 7648
rect 13032 7588 13036 7644
rect 13036 7588 13092 7644
rect 13092 7588 13096 7644
rect 13032 7584 13096 7588
rect 13112 7644 13176 7648
rect 13112 7588 13116 7644
rect 13116 7588 13172 7644
rect 13172 7588 13176 7644
rect 13112 7584 13176 7588
rect 13192 7644 13256 7648
rect 13192 7588 13196 7644
rect 13196 7588 13252 7644
rect 13252 7588 13256 7644
rect 13192 7584 13256 7588
rect 20952 7644 21016 7648
rect 20952 7588 20956 7644
rect 20956 7588 21012 7644
rect 21012 7588 21016 7644
rect 20952 7584 21016 7588
rect 21032 7644 21096 7648
rect 21032 7588 21036 7644
rect 21036 7588 21092 7644
rect 21092 7588 21096 7644
rect 21032 7584 21096 7588
rect 21112 7644 21176 7648
rect 21112 7588 21116 7644
rect 21116 7588 21172 7644
rect 21172 7588 21176 7644
rect 21112 7584 21176 7588
rect 21192 7644 21256 7648
rect 21192 7588 21196 7644
rect 21196 7588 21252 7644
rect 21252 7588 21256 7644
rect 21192 7584 21256 7588
rect 13492 7380 13556 7444
rect 8952 7100 9016 7104
rect 8952 7044 8956 7100
rect 8956 7044 9012 7100
rect 9012 7044 9016 7100
rect 8952 7040 9016 7044
rect 9032 7100 9096 7104
rect 9032 7044 9036 7100
rect 9036 7044 9092 7100
rect 9092 7044 9096 7100
rect 9032 7040 9096 7044
rect 9112 7100 9176 7104
rect 9112 7044 9116 7100
rect 9116 7044 9172 7100
rect 9172 7044 9176 7100
rect 9112 7040 9176 7044
rect 9192 7100 9256 7104
rect 9192 7044 9196 7100
rect 9196 7044 9252 7100
rect 9252 7044 9256 7100
rect 9192 7040 9256 7044
rect 16952 7100 17016 7104
rect 16952 7044 16956 7100
rect 16956 7044 17012 7100
rect 17012 7044 17016 7100
rect 16952 7040 17016 7044
rect 17032 7100 17096 7104
rect 17032 7044 17036 7100
rect 17036 7044 17092 7100
rect 17092 7044 17096 7100
rect 17032 7040 17096 7044
rect 17112 7100 17176 7104
rect 17112 7044 17116 7100
rect 17116 7044 17172 7100
rect 17172 7044 17176 7100
rect 17112 7040 17176 7044
rect 17192 7100 17256 7104
rect 17192 7044 17196 7100
rect 17196 7044 17252 7100
rect 17252 7044 17256 7100
rect 17192 7040 17256 7044
rect 60 6972 124 7036
rect 60 6700 124 6764
rect 4952 6556 5016 6560
rect 4952 6500 4956 6556
rect 4956 6500 5012 6556
rect 5012 6500 5016 6556
rect 4952 6496 5016 6500
rect 5032 6556 5096 6560
rect 5032 6500 5036 6556
rect 5036 6500 5092 6556
rect 5092 6500 5096 6556
rect 5032 6496 5096 6500
rect 5112 6556 5176 6560
rect 5112 6500 5116 6556
rect 5116 6500 5172 6556
rect 5172 6500 5176 6556
rect 5112 6496 5176 6500
rect 5192 6556 5256 6560
rect 5192 6500 5196 6556
rect 5196 6500 5252 6556
rect 5252 6500 5256 6556
rect 5192 6496 5256 6500
rect 12952 6556 13016 6560
rect 12952 6500 12956 6556
rect 12956 6500 13012 6556
rect 13012 6500 13016 6556
rect 12952 6496 13016 6500
rect 13032 6556 13096 6560
rect 13032 6500 13036 6556
rect 13036 6500 13092 6556
rect 13092 6500 13096 6556
rect 13032 6496 13096 6500
rect 13112 6556 13176 6560
rect 13112 6500 13116 6556
rect 13116 6500 13172 6556
rect 13172 6500 13176 6556
rect 13112 6496 13176 6500
rect 13192 6556 13256 6560
rect 13192 6500 13196 6556
rect 13196 6500 13252 6556
rect 13252 6500 13256 6556
rect 13192 6496 13256 6500
rect 20952 6556 21016 6560
rect 20952 6500 20956 6556
rect 20956 6500 21012 6556
rect 21012 6500 21016 6556
rect 20952 6496 21016 6500
rect 21032 6556 21096 6560
rect 21032 6500 21036 6556
rect 21036 6500 21092 6556
rect 21092 6500 21096 6556
rect 21032 6496 21096 6500
rect 21112 6556 21176 6560
rect 21112 6500 21116 6556
rect 21116 6500 21172 6556
rect 21172 6500 21176 6556
rect 21112 6496 21176 6500
rect 21192 6556 21256 6560
rect 21192 6500 21196 6556
rect 21196 6500 21252 6556
rect 21252 6500 21256 6556
rect 21192 6496 21256 6500
rect 8952 6012 9016 6016
rect 8952 5956 8956 6012
rect 8956 5956 9012 6012
rect 9012 5956 9016 6012
rect 8952 5952 9016 5956
rect 9032 6012 9096 6016
rect 9032 5956 9036 6012
rect 9036 5956 9092 6012
rect 9092 5956 9096 6012
rect 9032 5952 9096 5956
rect 9112 6012 9176 6016
rect 9112 5956 9116 6012
rect 9116 5956 9172 6012
rect 9172 5956 9176 6012
rect 9112 5952 9176 5956
rect 9192 6012 9256 6016
rect 9192 5956 9196 6012
rect 9196 5956 9252 6012
rect 9252 5956 9256 6012
rect 9192 5952 9256 5956
rect 16952 6012 17016 6016
rect 16952 5956 16956 6012
rect 16956 5956 17012 6012
rect 17012 5956 17016 6012
rect 16952 5952 17016 5956
rect 17032 6012 17096 6016
rect 17032 5956 17036 6012
rect 17036 5956 17092 6012
rect 17092 5956 17096 6012
rect 17032 5952 17096 5956
rect 17112 6012 17176 6016
rect 17112 5956 17116 6012
rect 17116 5956 17172 6012
rect 17172 5956 17176 6012
rect 17112 5952 17176 5956
rect 17192 6012 17256 6016
rect 17192 5956 17196 6012
rect 17196 5956 17252 6012
rect 17252 5956 17256 6012
rect 17192 5952 17256 5956
rect 4952 5468 5016 5472
rect 4952 5412 4956 5468
rect 4956 5412 5012 5468
rect 5012 5412 5016 5468
rect 4952 5408 5016 5412
rect 5032 5468 5096 5472
rect 5032 5412 5036 5468
rect 5036 5412 5092 5468
rect 5092 5412 5096 5468
rect 5032 5408 5096 5412
rect 5112 5468 5176 5472
rect 5112 5412 5116 5468
rect 5116 5412 5172 5468
rect 5172 5412 5176 5468
rect 5112 5408 5176 5412
rect 5192 5468 5256 5472
rect 5192 5412 5196 5468
rect 5196 5412 5252 5468
rect 5252 5412 5256 5468
rect 5192 5408 5256 5412
rect 12952 5468 13016 5472
rect 12952 5412 12956 5468
rect 12956 5412 13012 5468
rect 13012 5412 13016 5468
rect 12952 5408 13016 5412
rect 13032 5468 13096 5472
rect 13032 5412 13036 5468
rect 13036 5412 13092 5468
rect 13092 5412 13096 5468
rect 13032 5408 13096 5412
rect 13112 5468 13176 5472
rect 13112 5412 13116 5468
rect 13116 5412 13172 5468
rect 13172 5412 13176 5468
rect 13112 5408 13176 5412
rect 13192 5468 13256 5472
rect 13192 5412 13196 5468
rect 13196 5412 13252 5468
rect 13252 5412 13256 5468
rect 13192 5408 13256 5412
rect 20952 5468 21016 5472
rect 20952 5412 20956 5468
rect 20956 5412 21012 5468
rect 21012 5412 21016 5468
rect 20952 5408 21016 5412
rect 21032 5468 21096 5472
rect 21032 5412 21036 5468
rect 21036 5412 21092 5468
rect 21092 5412 21096 5468
rect 21032 5408 21096 5412
rect 21112 5468 21176 5472
rect 21112 5412 21116 5468
rect 21116 5412 21172 5468
rect 21172 5412 21176 5468
rect 21112 5408 21176 5412
rect 21192 5468 21256 5472
rect 21192 5412 21196 5468
rect 21196 5412 21252 5468
rect 21252 5412 21256 5468
rect 21192 5408 21256 5412
rect 8952 4924 9016 4928
rect 8952 4868 8956 4924
rect 8956 4868 9012 4924
rect 9012 4868 9016 4924
rect 8952 4864 9016 4868
rect 9032 4924 9096 4928
rect 9032 4868 9036 4924
rect 9036 4868 9092 4924
rect 9092 4868 9096 4924
rect 9032 4864 9096 4868
rect 9112 4924 9176 4928
rect 9112 4868 9116 4924
rect 9116 4868 9172 4924
rect 9172 4868 9176 4924
rect 9112 4864 9176 4868
rect 9192 4924 9256 4928
rect 9192 4868 9196 4924
rect 9196 4868 9252 4924
rect 9252 4868 9256 4924
rect 9192 4864 9256 4868
rect 16952 4924 17016 4928
rect 16952 4868 16956 4924
rect 16956 4868 17012 4924
rect 17012 4868 17016 4924
rect 16952 4864 17016 4868
rect 17032 4924 17096 4928
rect 17032 4868 17036 4924
rect 17036 4868 17092 4924
rect 17092 4868 17096 4924
rect 17032 4864 17096 4868
rect 17112 4924 17176 4928
rect 17112 4868 17116 4924
rect 17116 4868 17172 4924
rect 17172 4868 17176 4924
rect 17112 4864 17176 4868
rect 17192 4924 17256 4928
rect 17192 4868 17196 4924
rect 17196 4868 17252 4924
rect 17252 4868 17256 4924
rect 17192 4864 17256 4868
rect 4952 4380 5016 4384
rect 4952 4324 4956 4380
rect 4956 4324 5012 4380
rect 5012 4324 5016 4380
rect 4952 4320 5016 4324
rect 5032 4380 5096 4384
rect 5032 4324 5036 4380
rect 5036 4324 5092 4380
rect 5092 4324 5096 4380
rect 5032 4320 5096 4324
rect 5112 4380 5176 4384
rect 5112 4324 5116 4380
rect 5116 4324 5172 4380
rect 5172 4324 5176 4380
rect 5112 4320 5176 4324
rect 5192 4380 5256 4384
rect 5192 4324 5196 4380
rect 5196 4324 5252 4380
rect 5252 4324 5256 4380
rect 5192 4320 5256 4324
rect 12952 4380 13016 4384
rect 12952 4324 12956 4380
rect 12956 4324 13012 4380
rect 13012 4324 13016 4380
rect 12952 4320 13016 4324
rect 13032 4380 13096 4384
rect 13032 4324 13036 4380
rect 13036 4324 13092 4380
rect 13092 4324 13096 4380
rect 13032 4320 13096 4324
rect 13112 4380 13176 4384
rect 13112 4324 13116 4380
rect 13116 4324 13172 4380
rect 13172 4324 13176 4380
rect 13112 4320 13176 4324
rect 13192 4380 13256 4384
rect 13192 4324 13196 4380
rect 13196 4324 13252 4380
rect 13252 4324 13256 4380
rect 13192 4320 13256 4324
rect 20952 4380 21016 4384
rect 20952 4324 20956 4380
rect 20956 4324 21012 4380
rect 21012 4324 21016 4380
rect 20952 4320 21016 4324
rect 21032 4380 21096 4384
rect 21032 4324 21036 4380
rect 21036 4324 21092 4380
rect 21092 4324 21096 4380
rect 21032 4320 21096 4324
rect 21112 4380 21176 4384
rect 21112 4324 21116 4380
rect 21116 4324 21172 4380
rect 21172 4324 21176 4380
rect 21112 4320 21176 4324
rect 21192 4380 21256 4384
rect 21192 4324 21196 4380
rect 21196 4324 21252 4380
rect 21252 4324 21256 4380
rect 21192 4320 21256 4324
rect 8952 3836 9016 3840
rect 8952 3780 8956 3836
rect 8956 3780 9012 3836
rect 9012 3780 9016 3836
rect 8952 3776 9016 3780
rect 9032 3836 9096 3840
rect 9032 3780 9036 3836
rect 9036 3780 9092 3836
rect 9092 3780 9096 3836
rect 9032 3776 9096 3780
rect 9112 3836 9176 3840
rect 9112 3780 9116 3836
rect 9116 3780 9172 3836
rect 9172 3780 9176 3836
rect 9112 3776 9176 3780
rect 9192 3836 9256 3840
rect 9192 3780 9196 3836
rect 9196 3780 9252 3836
rect 9252 3780 9256 3836
rect 9192 3776 9256 3780
rect 16952 3836 17016 3840
rect 16952 3780 16956 3836
rect 16956 3780 17012 3836
rect 17012 3780 17016 3836
rect 16952 3776 17016 3780
rect 17032 3836 17096 3840
rect 17032 3780 17036 3836
rect 17036 3780 17092 3836
rect 17092 3780 17096 3836
rect 17032 3776 17096 3780
rect 17112 3836 17176 3840
rect 17112 3780 17116 3836
rect 17116 3780 17172 3836
rect 17172 3780 17176 3836
rect 17112 3776 17176 3780
rect 17192 3836 17256 3840
rect 17192 3780 17196 3836
rect 17196 3780 17252 3836
rect 17252 3780 17256 3836
rect 17192 3776 17256 3780
rect 4952 3292 5016 3296
rect 4952 3236 4956 3292
rect 4956 3236 5012 3292
rect 5012 3236 5016 3292
rect 4952 3232 5016 3236
rect 5032 3292 5096 3296
rect 5032 3236 5036 3292
rect 5036 3236 5092 3292
rect 5092 3236 5096 3292
rect 5032 3232 5096 3236
rect 5112 3292 5176 3296
rect 5112 3236 5116 3292
rect 5116 3236 5172 3292
rect 5172 3236 5176 3292
rect 5112 3232 5176 3236
rect 5192 3292 5256 3296
rect 5192 3236 5196 3292
rect 5196 3236 5252 3292
rect 5252 3236 5256 3292
rect 5192 3232 5256 3236
rect 12952 3292 13016 3296
rect 12952 3236 12956 3292
rect 12956 3236 13012 3292
rect 13012 3236 13016 3292
rect 12952 3232 13016 3236
rect 13032 3292 13096 3296
rect 13032 3236 13036 3292
rect 13036 3236 13092 3292
rect 13092 3236 13096 3292
rect 13032 3232 13096 3236
rect 13112 3292 13176 3296
rect 13112 3236 13116 3292
rect 13116 3236 13172 3292
rect 13172 3236 13176 3292
rect 13112 3232 13176 3236
rect 13192 3292 13256 3296
rect 13192 3236 13196 3292
rect 13196 3236 13252 3292
rect 13252 3236 13256 3292
rect 13192 3232 13256 3236
rect 20952 3292 21016 3296
rect 20952 3236 20956 3292
rect 20956 3236 21012 3292
rect 21012 3236 21016 3292
rect 20952 3232 21016 3236
rect 21032 3292 21096 3296
rect 21032 3236 21036 3292
rect 21036 3236 21092 3292
rect 21092 3236 21096 3292
rect 21032 3232 21096 3236
rect 21112 3292 21176 3296
rect 21112 3236 21116 3292
rect 21116 3236 21172 3292
rect 21172 3236 21176 3292
rect 21112 3232 21176 3236
rect 21192 3292 21256 3296
rect 21192 3236 21196 3292
rect 21196 3236 21252 3292
rect 21252 3236 21256 3292
rect 21192 3232 21256 3236
rect 8952 2748 9016 2752
rect 8952 2692 8956 2748
rect 8956 2692 9012 2748
rect 9012 2692 9016 2748
rect 8952 2688 9016 2692
rect 9032 2748 9096 2752
rect 9032 2692 9036 2748
rect 9036 2692 9092 2748
rect 9092 2692 9096 2748
rect 9032 2688 9096 2692
rect 9112 2748 9176 2752
rect 9112 2692 9116 2748
rect 9116 2692 9172 2748
rect 9172 2692 9176 2748
rect 9112 2688 9176 2692
rect 9192 2748 9256 2752
rect 9192 2692 9196 2748
rect 9196 2692 9252 2748
rect 9252 2692 9256 2748
rect 9192 2688 9256 2692
rect 16952 2748 17016 2752
rect 16952 2692 16956 2748
rect 16956 2692 17012 2748
rect 17012 2692 17016 2748
rect 16952 2688 17016 2692
rect 17032 2748 17096 2752
rect 17032 2692 17036 2748
rect 17036 2692 17092 2748
rect 17092 2692 17096 2748
rect 17032 2688 17096 2692
rect 17112 2748 17176 2752
rect 17112 2692 17116 2748
rect 17116 2692 17172 2748
rect 17172 2692 17176 2748
rect 17112 2688 17176 2692
rect 17192 2748 17256 2752
rect 17192 2692 17196 2748
rect 17196 2692 17252 2748
rect 17252 2692 17256 2748
rect 17192 2688 17256 2692
rect 4952 2204 5016 2208
rect 4952 2148 4956 2204
rect 4956 2148 5012 2204
rect 5012 2148 5016 2204
rect 4952 2144 5016 2148
rect 5032 2204 5096 2208
rect 5032 2148 5036 2204
rect 5036 2148 5092 2204
rect 5092 2148 5096 2204
rect 5032 2144 5096 2148
rect 5112 2204 5176 2208
rect 5112 2148 5116 2204
rect 5116 2148 5172 2204
rect 5172 2148 5176 2204
rect 5112 2144 5176 2148
rect 5192 2204 5256 2208
rect 5192 2148 5196 2204
rect 5196 2148 5252 2204
rect 5252 2148 5256 2204
rect 5192 2144 5256 2148
rect 12952 2204 13016 2208
rect 12952 2148 12956 2204
rect 12956 2148 13012 2204
rect 13012 2148 13016 2204
rect 12952 2144 13016 2148
rect 13032 2204 13096 2208
rect 13032 2148 13036 2204
rect 13036 2148 13092 2204
rect 13092 2148 13096 2204
rect 13032 2144 13096 2148
rect 13112 2204 13176 2208
rect 13112 2148 13116 2204
rect 13116 2148 13172 2204
rect 13172 2148 13176 2204
rect 13112 2144 13176 2148
rect 13192 2204 13256 2208
rect 13192 2148 13196 2204
rect 13196 2148 13252 2204
rect 13252 2148 13256 2204
rect 13192 2144 13256 2148
rect 20952 2204 21016 2208
rect 20952 2148 20956 2204
rect 20956 2148 21012 2204
rect 21012 2148 21016 2204
rect 20952 2144 21016 2148
rect 21032 2204 21096 2208
rect 21032 2148 21036 2204
rect 21036 2148 21092 2204
rect 21092 2148 21096 2204
rect 21032 2144 21096 2148
rect 21112 2204 21176 2208
rect 21112 2148 21116 2204
rect 21116 2148 21172 2204
rect 21172 2148 21176 2204
rect 21112 2144 21176 2148
rect 21192 2204 21256 2208
rect 21192 2148 21196 2204
rect 21196 2148 21252 2204
rect 21252 2148 21256 2204
rect 21192 2144 21256 2148
<< metal4 >>
rect 4944 21792 5264 21808
rect 4944 21728 4952 21792
rect 5016 21728 5032 21792
rect 5096 21728 5112 21792
rect 5176 21728 5192 21792
rect 5256 21728 5264 21792
rect 4944 20704 5264 21728
rect 4944 20640 4952 20704
rect 5016 20640 5032 20704
rect 5096 20640 5112 20704
rect 5176 20640 5192 20704
rect 5256 20640 5264 20704
rect 4944 19616 5264 20640
rect 4944 19552 4952 19616
rect 5016 19552 5032 19616
rect 5096 19552 5112 19616
rect 5176 19552 5192 19616
rect 5256 19552 5264 19616
rect 4944 18528 5264 19552
rect 4944 18464 4952 18528
rect 5016 18464 5032 18528
rect 5096 18464 5112 18528
rect 5176 18464 5192 18528
rect 5256 18464 5264 18528
rect 4944 17440 5264 18464
rect 4944 17376 4952 17440
rect 5016 17376 5032 17440
rect 5096 17376 5112 17440
rect 5176 17376 5192 17440
rect 5256 17376 5264 17440
rect 4944 16352 5264 17376
rect 4944 16288 4952 16352
rect 5016 16288 5032 16352
rect 5096 16288 5112 16352
rect 5176 16288 5192 16352
rect 5256 16288 5264 16352
rect 4944 15264 5264 16288
rect 4944 15200 4952 15264
rect 5016 15200 5032 15264
rect 5096 15200 5112 15264
rect 5176 15200 5192 15264
rect 5256 15200 5264 15264
rect 4944 14176 5264 15200
rect 4944 14112 4952 14176
rect 5016 14112 5032 14176
rect 5096 14112 5112 14176
rect 5176 14112 5192 14176
rect 5256 14112 5264 14176
rect 4944 13088 5264 14112
rect 4944 13024 4952 13088
rect 5016 13024 5032 13088
rect 5096 13024 5112 13088
rect 5176 13024 5192 13088
rect 5256 13024 5264 13088
rect 4944 12000 5264 13024
rect 4944 11936 4952 12000
rect 5016 11936 5032 12000
rect 5096 11936 5112 12000
rect 5176 11936 5192 12000
rect 5256 11936 5264 12000
rect 59 11932 125 11933
rect 59 11868 60 11932
rect 124 11868 125 11932
rect 59 11867 125 11868
rect 62 11661 122 11867
rect 59 11660 125 11661
rect 59 11596 60 11660
rect 124 11596 125 11660
rect 59 11595 125 11596
rect 4944 10912 5264 11936
rect 4944 10848 4952 10912
rect 5016 10848 5032 10912
rect 5096 10848 5112 10912
rect 5176 10848 5192 10912
rect 5256 10848 5264 10912
rect 4944 9824 5264 10848
rect 4944 9760 4952 9824
rect 5016 9760 5032 9824
rect 5096 9760 5112 9824
rect 5176 9760 5192 9824
rect 5256 9760 5264 9824
rect 4944 8736 5264 9760
rect 4944 8672 4952 8736
rect 5016 8672 5032 8736
rect 5096 8672 5112 8736
rect 5176 8672 5192 8736
rect 5256 8672 5264 8736
rect 4944 7648 5264 8672
rect 4944 7584 4952 7648
rect 5016 7584 5032 7648
rect 5096 7584 5112 7648
rect 5176 7584 5192 7648
rect 5256 7584 5264 7648
rect 59 7036 125 7037
rect 59 6972 60 7036
rect 124 6972 125 7036
rect 59 6971 125 6972
rect 62 6765 122 6971
rect 59 6764 125 6765
rect 59 6700 60 6764
rect 124 6700 125 6764
rect 59 6699 125 6700
rect 4944 6560 5264 7584
rect 4944 6496 4952 6560
rect 5016 6496 5032 6560
rect 5096 6496 5112 6560
rect 5176 6496 5192 6560
rect 5256 6496 5264 6560
rect 4944 5472 5264 6496
rect 4944 5408 4952 5472
rect 5016 5408 5032 5472
rect 5096 5408 5112 5472
rect 5176 5408 5192 5472
rect 5256 5408 5264 5472
rect 4944 4384 5264 5408
rect 4944 4320 4952 4384
rect 5016 4320 5032 4384
rect 5096 4320 5112 4384
rect 5176 4320 5192 4384
rect 5256 4320 5264 4384
rect 4944 3296 5264 4320
rect 4944 3232 4952 3296
rect 5016 3232 5032 3296
rect 5096 3232 5112 3296
rect 5176 3232 5192 3296
rect 5256 3232 5264 3296
rect 4944 2208 5264 3232
rect 4944 2144 4952 2208
rect 5016 2144 5032 2208
rect 5096 2144 5112 2208
rect 5176 2144 5192 2208
rect 5256 2144 5264 2208
rect 4944 2128 5264 2144
rect 8944 21248 9264 21808
rect 8944 21184 8952 21248
rect 9016 21184 9032 21248
rect 9096 21184 9112 21248
rect 9176 21184 9192 21248
rect 9256 21184 9264 21248
rect 8944 20160 9264 21184
rect 8944 20096 8952 20160
rect 9016 20096 9032 20160
rect 9096 20096 9112 20160
rect 9176 20096 9192 20160
rect 9256 20096 9264 20160
rect 8944 19072 9264 20096
rect 8944 19008 8952 19072
rect 9016 19008 9032 19072
rect 9096 19008 9112 19072
rect 9176 19008 9192 19072
rect 9256 19008 9264 19072
rect 8944 17984 9264 19008
rect 8944 17920 8952 17984
rect 9016 17920 9032 17984
rect 9096 17920 9112 17984
rect 9176 17920 9192 17984
rect 9256 17920 9264 17984
rect 8944 16896 9264 17920
rect 8944 16832 8952 16896
rect 9016 16832 9032 16896
rect 9096 16832 9112 16896
rect 9176 16832 9192 16896
rect 9256 16832 9264 16896
rect 8944 15808 9264 16832
rect 8944 15744 8952 15808
rect 9016 15744 9032 15808
rect 9096 15744 9112 15808
rect 9176 15744 9192 15808
rect 9256 15744 9264 15808
rect 8944 14720 9264 15744
rect 8944 14656 8952 14720
rect 9016 14656 9032 14720
rect 9096 14656 9112 14720
rect 9176 14656 9192 14720
rect 9256 14656 9264 14720
rect 8944 13632 9264 14656
rect 8944 13568 8952 13632
rect 9016 13568 9032 13632
rect 9096 13568 9112 13632
rect 9176 13568 9192 13632
rect 9256 13568 9264 13632
rect 8944 12544 9264 13568
rect 8944 12480 8952 12544
rect 9016 12480 9032 12544
rect 9096 12480 9112 12544
rect 9176 12480 9192 12544
rect 9256 12480 9264 12544
rect 8944 11456 9264 12480
rect 8944 11392 8952 11456
rect 9016 11392 9032 11456
rect 9096 11392 9112 11456
rect 9176 11392 9192 11456
rect 9256 11392 9264 11456
rect 8944 10368 9264 11392
rect 8944 10304 8952 10368
rect 9016 10304 9032 10368
rect 9096 10304 9112 10368
rect 9176 10304 9192 10368
rect 9256 10304 9264 10368
rect 8944 9280 9264 10304
rect 8944 9216 8952 9280
rect 9016 9216 9032 9280
rect 9096 9216 9112 9280
rect 9176 9216 9192 9280
rect 9256 9216 9264 9280
rect 8944 8192 9264 9216
rect 8944 8128 8952 8192
rect 9016 8128 9032 8192
rect 9096 8128 9112 8192
rect 9176 8128 9192 8192
rect 9256 8128 9264 8192
rect 8944 7104 9264 8128
rect 8944 7040 8952 7104
rect 9016 7040 9032 7104
rect 9096 7040 9112 7104
rect 9176 7040 9192 7104
rect 9256 7040 9264 7104
rect 8944 6016 9264 7040
rect 8944 5952 8952 6016
rect 9016 5952 9032 6016
rect 9096 5952 9112 6016
rect 9176 5952 9192 6016
rect 9256 5952 9264 6016
rect 8944 4928 9264 5952
rect 8944 4864 8952 4928
rect 9016 4864 9032 4928
rect 9096 4864 9112 4928
rect 9176 4864 9192 4928
rect 9256 4864 9264 4928
rect 8944 3840 9264 4864
rect 8944 3776 8952 3840
rect 9016 3776 9032 3840
rect 9096 3776 9112 3840
rect 9176 3776 9192 3840
rect 9256 3776 9264 3840
rect 8944 2752 9264 3776
rect 8944 2688 8952 2752
rect 9016 2688 9032 2752
rect 9096 2688 9112 2752
rect 9176 2688 9192 2752
rect 9256 2688 9264 2752
rect 8944 2128 9264 2688
rect 12944 21792 13264 21808
rect 12944 21728 12952 21792
rect 13016 21728 13032 21792
rect 13096 21728 13112 21792
rect 13176 21728 13192 21792
rect 13256 21728 13264 21792
rect 12944 20704 13264 21728
rect 12944 20640 12952 20704
rect 13016 20640 13032 20704
rect 13096 20640 13112 20704
rect 13176 20640 13192 20704
rect 13256 20640 13264 20704
rect 12944 19616 13264 20640
rect 12944 19552 12952 19616
rect 13016 19552 13032 19616
rect 13096 19552 13112 19616
rect 13176 19552 13192 19616
rect 13256 19552 13264 19616
rect 12944 18528 13264 19552
rect 12944 18464 12952 18528
rect 13016 18464 13032 18528
rect 13096 18464 13112 18528
rect 13176 18464 13192 18528
rect 13256 18464 13264 18528
rect 12944 17440 13264 18464
rect 12944 17376 12952 17440
rect 13016 17376 13032 17440
rect 13096 17376 13112 17440
rect 13176 17376 13192 17440
rect 13256 17376 13264 17440
rect 12944 16352 13264 17376
rect 12944 16288 12952 16352
rect 13016 16288 13032 16352
rect 13096 16288 13112 16352
rect 13176 16288 13192 16352
rect 13256 16288 13264 16352
rect 12944 15264 13264 16288
rect 12944 15200 12952 15264
rect 13016 15200 13032 15264
rect 13096 15200 13112 15264
rect 13176 15200 13192 15264
rect 13256 15200 13264 15264
rect 12944 14176 13264 15200
rect 12944 14112 12952 14176
rect 13016 14112 13032 14176
rect 13096 14112 13112 14176
rect 13176 14112 13192 14176
rect 13256 14112 13264 14176
rect 12944 13088 13264 14112
rect 12944 13024 12952 13088
rect 13016 13024 13032 13088
rect 13096 13024 13112 13088
rect 13176 13024 13192 13088
rect 13256 13024 13264 13088
rect 12944 12000 13264 13024
rect 16944 21248 17264 21808
rect 16944 21184 16952 21248
rect 17016 21184 17032 21248
rect 17096 21184 17112 21248
rect 17176 21184 17192 21248
rect 17256 21184 17264 21248
rect 16944 20160 17264 21184
rect 16944 20096 16952 20160
rect 17016 20096 17032 20160
rect 17096 20096 17112 20160
rect 17176 20096 17192 20160
rect 17256 20096 17264 20160
rect 16944 19072 17264 20096
rect 16944 19008 16952 19072
rect 17016 19008 17032 19072
rect 17096 19008 17112 19072
rect 17176 19008 17192 19072
rect 17256 19008 17264 19072
rect 16944 17984 17264 19008
rect 16944 17920 16952 17984
rect 17016 17920 17032 17984
rect 17096 17920 17112 17984
rect 17176 17920 17192 17984
rect 17256 17920 17264 17984
rect 16944 16896 17264 17920
rect 16944 16832 16952 16896
rect 17016 16832 17032 16896
rect 17096 16832 17112 16896
rect 17176 16832 17192 16896
rect 17256 16832 17264 16896
rect 16944 15808 17264 16832
rect 16944 15744 16952 15808
rect 17016 15744 17032 15808
rect 17096 15744 17112 15808
rect 17176 15744 17192 15808
rect 17256 15744 17264 15808
rect 16944 14720 17264 15744
rect 16944 14656 16952 14720
rect 17016 14656 17032 14720
rect 17096 14656 17112 14720
rect 17176 14656 17192 14720
rect 17256 14656 17264 14720
rect 16944 13632 17264 14656
rect 16944 13568 16952 13632
rect 17016 13568 17032 13632
rect 17096 13568 17112 13632
rect 17176 13568 17192 13632
rect 17256 13568 17264 13632
rect 16944 12544 17264 13568
rect 16944 12480 16952 12544
rect 17016 12480 17032 12544
rect 17096 12480 17112 12544
rect 17176 12480 17192 12544
rect 17256 12480 17264 12544
rect 13491 12340 13557 12341
rect 13491 12276 13492 12340
rect 13556 12276 13557 12340
rect 13491 12275 13557 12276
rect 12944 11936 12952 12000
rect 13016 11936 13032 12000
rect 13096 11936 13112 12000
rect 13176 11936 13192 12000
rect 13256 11936 13264 12000
rect 12944 10912 13264 11936
rect 12944 10848 12952 10912
rect 13016 10848 13032 10912
rect 13096 10848 13112 10912
rect 13176 10848 13192 10912
rect 13256 10848 13264 10912
rect 12944 9824 13264 10848
rect 12944 9760 12952 9824
rect 13016 9760 13032 9824
rect 13096 9760 13112 9824
rect 13176 9760 13192 9824
rect 13256 9760 13264 9824
rect 12944 8736 13264 9760
rect 13494 9349 13554 12275
rect 16944 11456 17264 12480
rect 16944 11392 16952 11456
rect 17016 11392 17032 11456
rect 17096 11392 17112 11456
rect 17176 11392 17192 11456
rect 17256 11392 17264 11456
rect 16944 10368 17264 11392
rect 16944 10304 16952 10368
rect 17016 10304 17032 10368
rect 17096 10304 17112 10368
rect 17176 10304 17192 10368
rect 17256 10304 17264 10368
rect 13491 9348 13557 9349
rect 13491 9284 13492 9348
rect 13556 9284 13557 9348
rect 13491 9283 13557 9284
rect 12944 8672 12952 8736
rect 13016 8672 13032 8736
rect 13096 8672 13112 8736
rect 13176 8672 13192 8736
rect 13256 8672 13264 8736
rect 12944 7648 13264 8672
rect 12944 7584 12952 7648
rect 13016 7584 13032 7648
rect 13096 7584 13112 7648
rect 13176 7584 13192 7648
rect 13256 7584 13264 7648
rect 12944 6560 13264 7584
rect 13494 7445 13554 9283
rect 16944 9280 17264 10304
rect 16944 9216 16952 9280
rect 17016 9216 17032 9280
rect 17096 9216 17112 9280
rect 17176 9216 17192 9280
rect 17256 9216 17264 9280
rect 16944 8192 17264 9216
rect 16944 8128 16952 8192
rect 17016 8128 17032 8192
rect 17096 8128 17112 8192
rect 17176 8128 17192 8192
rect 17256 8128 17264 8192
rect 13491 7444 13557 7445
rect 13491 7380 13492 7444
rect 13556 7380 13557 7444
rect 13491 7379 13557 7380
rect 12944 6496 12952 6560
rect 13016 6496 13032 6560
rect 13096 6496 13112 6560
rect 13176 6496 13192 6560
rect 13256 6496 13264 6560
rect 12944 5472 13264 6496
rect 12944 5408 12952 5472
rect 13016 5408 13032 5472
rect 13096 5408 13112 5472
rect 13176 5408 13192 5472
rect 13256 5408 13264 5472
rect 12944 4384 13264 5408
rect 12944 4320 12952 4384
rect 13016 4320 13032 4384
rect 13096 4320 13112 4384
rect 13176 4320 13192 4384
rect 13256 4320 13264 4384
rect 12944 3296 13264 4320
rect 12944 3232 12952 3296
rect 13016 3232 13032 3296
rect 13096 3232 13112 3296
rect 13176 3232 13192 3296
rect 13256 3232 13264 3296
rect 12944 2208 13264 3232
rect 12944 2144 12952 2208
rect 13016 2144 13032 2208
rect 13096 2144 13112 2208
rect 13176 2144 13192 2208
rect 13256 2144 13264 2208
rect 12944 2128 13264 2144
rect 16944 7104 17264 8128
rect 16944 7040 16952 7104
rect 17016 7040 17032 7104
rect 17096 7040 17112 7104
rect 17176 7040 17192 7104
rect 17256 7040 17264 7104
rect 16944 6016 17264 7040
rect 16944 5952 16952 6016
rect 17016 5952 17032 6016
rect 17096 5952 17112 6016
rect 17176 5952 17192 6016
rect 17256 5952 17264 6016
rect 16944 4928 17264 5952
rect 16944 4864 16952 4928
rect 17016 4864 17032 4928
rect 17096 4864 17112 4928
rect 17176 4864 17192 4928
rect 17256 4864 17264 4928
rect 16944 3840 17264 4864
rect 16944 3776 16952 3840
rect 17016 3776 17032 3840
rect 17096 3776 17112 3840
rect 17176 3776 17192 3840
rect 17256 3776 17264 3840
rect 16944 2752 17264 3776
rect 16944 2688 16952 2752
rect 17016 2688 17032 2752
rect 17096 2688 17112 2752
rect 17176 2688 17192 2752
rect 17256 2688 17264 2752
rect 16944 2128 17264 2688
rect 20944 21792 21264 21808
rect 20944 21728 20952 21792
rect 21016 21728 21032 21792
rect 21096 21728 21112 21792
rect 21176 21728 21192 21792
rect 21256 21728 21264 21792
rect 20944 20704 21264 21728
rect 20944 20640 20952 20704
rect 21016 20640 21032 20704
rect 21096 20640 21112 20704
rect 21176 20640 21192 20704
rect 21256 20640 21264 20704
rect 20944 19616 21264 20640
rect 20944 19552 20952 19616
rect 21016 19552 21032 19616
rect 21096 19552 21112 19616
rect 21176 19552 21192 19616
rect 21256 19552 21264 19616
rect 20944 18528 21264 19552
rect 20944 18464 20952 18528
rect 21016 18464 21032 18528
rect 21096 18464 21112 18528
rect 21176 18464 21192 18528
rect 21256 18464 21264 18528
rect 20944 17440 21264 18464
rect 20944 17376 20952 17440
rect 21016 17376 21032 17440
rect 21096 17376 21112 17440
rect 21176 17376 21192 17440
rect 21256 17376 21264 17440
rect 20944 16352 21264 17376
rect 20944 16288 20952 16352
rect 21016 16288 21032 16352
rect 21096 16288 21112 16352
rect 21176 16288 21192 16352
rect 21256 16288 21264 16352
rect 20944 15264 21264 16288
rect 20944 15200 20952 15264
rect 21016 15200 21032 15264
rect 21096 15200 21112 15264
rect 21176 15200 21192 15264
rect 21256 15200 21264 15264
rect 20944 14176 21264 15200
rect 20944 14112 20952 14176
rect 21016 14112 21032 14176
rect 21096 14112 21112 14176
rect 21176 14112 21192 14176
rect 21256 14112 21264 14176
rect 20944 13088 21264 14112
rect 20944 13024 20952 13088
rect 21016 13024 21032 13088
rect 21096 13024 21112 13088
rect 21176 13024 21192 13088
rect 21256 13024 21264 13088
rect 20944 12000 21264 13024
rect 20944 11936 20952 12000
rect 21016 11936 21032 12000
rect 21096 11936 21112 12000
rect 21176 11936 21192 12000
rect 21256 11936 21264 12000
rect 20944 10912 21264 11936
rect 20944 10848 20952 10912
rect 21016 10848 21032 10912
rect 21096 10848 21112 10912
rect 21176 10848 21192 10912
rect 21256 10848 21264 10912
rect 20944 9824 21264 10848
rect 20944 9760 20952 9824
rect 21016 9760 21032 9824
rect 21096 9760 21112 9824
rect 21176 9760 21192 9824
rect 21256 9760 21264 9824
rect 20944 8736 21264 9760
rect 20944 8672 20952 8736
rect 21016 8672 21032 8736
rect 21096 8672 21112 8736
rect 21176 8672 21192 8736
rect 21256 8672 21264 8736
rect 20944 7648 21264 8672
rect 20944 7584 20952 7648
rect 21016 7584 21032 7648
rect 21096 7584 21112 7648
rect 21176 7584 21192 7648
rect 21256 7584 21264 7648
rect 20944 6560 21264 7584
rect 20944 6496 20952 6560
rect 21016 6496 21032 6560
rect 21096 6496 21112 6560
rect 21176 6496 21192 6560
rect 21256 6496 21264 6560
rect 20944 5472 21264 6496
rect 20944 5408 20952 5472
rect 21016 5408 21032 5472
rect 21096 5408 21112 5472
rect 21176 5408 21192 5472
rect 21256 5408 21264 5472
rect 20944 4384 21264 5408
rect 20944 4320 20952 4384
rect 21016 4320 21032 4384
rect 21096 4320 21112 4384
rect 21176 4320 21192 4384
rect 21256 4320 21264 4384
rect 20944 3296 21264 4320
rect 20944 3232 20952 3296
rect 21016 3232 21032 3296
rect 21096 3232 21112 3296
rect 21176 3232 21192 3296
rect 21256 3232 21264 3296
rect 20944 2208 21264 3232
rect 20944 2144 20952 2208
rect 21016 2144 21032 2208
rect 21096 2144 21112 2208
rect 21176 2144 21192 2208
rect 21256 2144 21264 2208
rect 20944 2128 21264 2144
<< via4 >>
rect 4022 7852 4258 7938
rect 4022 7788 4108 7852
rect 4108 7788 4172 7852
rect 4172 7788 4258 7852
rect 4022 7702 4258 7788
rect 14142 7852 14378 7938
rect 14142 7788 14228 7852
rect 14228 7788 14292 7852
rect 14292 7788 14378 7852
rect 14142 7702 14378 7788
<< metal5 >>
rect 3980 7938 14420 7980
rect 3980 7702 4022 7938
rect 4258 7702 14142 7938
rect 14378 7702 14420 7938
rect 3980 7660 14420 7702
use scs8hd_decap_3  PHY_0 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1104 0 -1 2720
box -38 -48 314 592
use scs8hd_decap_3  PHY_2
timestamp 1586364061
transform 1 0 1104 0 1 2720
box -38 -48 314 592
use scs8hd_decap_12  FILLER_0_3 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1380 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_3
timestamp 1586364061
transform 1 0 1380 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_15
timestamp 1586364061
transform 1 0 2484 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_0_27 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 3588 0 -1 2720
box -38 -48 406 592
use scs8hd_decap_12  FILLER_1_15
timestamp 1586364061
transform 1 0 2484 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_1_27
timestamp 1586364061
transform 1 0 3588 0 1 2720
box -38 -48 406 592
use scs8hd_inv_8  _048_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 4692 0 1 2720
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_72 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 3956 0 -1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__042__A tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 4048 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__048__A
timestamp 1586364061
transform 1 0 4508 0 1 2720
box -38 -48 222 592
use scs8hd_decap_12  FILLER_0_32
timestamp 1586364061
transform 1 0 4048 0 -1 2720
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_1_31 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 3956 0 1 2720
box -38 -48 130 592
use scs8hd_decap_3  FILLER_1_34
timestamp 1586364061
transform 1 0 4232 0 1 2720
box -38 -48 314 592
use scs8hd_buf_2  _155_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 5704 0 -1 2720
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__050__A
timestamp 1586364061
transform 1 0 5796 0 1 2720
box -38 -48 222 592
use scs8hd_decap_6  FILLER_0_44 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 5152 0 -1 2720
box -38 -48 590 592
use scs8hd_fill_2  FILLER_0_54 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 6072 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_3  FILLER_1_48
timestamp 1586364061
transform 1 0 5520 0 1 2720
box -38 -48 314 592
use scs8hd_decap_6  FILLER_1_53
timestamp 1586364061
transform 1 0 5980 0 1 2720
box -38 -48 590 592
use scs8hd_decap_3  FILLER_1_62
timestamp 1586364061
transform 1 0 6808 0 1 2720
box -38 -48 314 592
use scs8hd_fill_2  FILLER_0_58
timestamp 1586364061
transform 1 0 6440 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__067__B
timestamp 1586364061
transform 1 0 6532 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__049__A
timestamp 1586364061
transform 1 0 6624 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__155__A
timestamp 1586364061
transform 1 0 6256 0 -1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_79
timestamp 1586364061
transform 1 0 6716 0 1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_73
timestamp 1586364061
transform 1 0 6808 0 -1 2720
box -38 -48 130 592
use scs8hd_fill_2  FILLER_1_67
timestamp 1586364061
transform 1 0 7268 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__067__A
timestamp 1586364061
transform 1 0 7084 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__107__C
timestamp 1586364061
transform 1 0 7452 0 1 2720
box -38 -48 222 592
use scs8hd_inv_8  _049_
timestamp 1586364061
transform 1 0 6900 0 -1 2720
box -38 -48 866 592
use scs8hd_nor3_4  _107_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 7636 0 1 2720
box -38 -48 1234 592
use scs8hd_buf_2  _147_
timestamp 1586364061
transform 1 0 8556 0 -1 2720
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__107__A
timestamp 1586364061
transform 1 0 7912 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__107__B
timestamp 1586364061
transform 1 0 8280 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_72
timestamp 1586364061
transform 1 0 7728 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_76
timestamp 1586364061
transform 1 0 8096 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_1  FILLER_0_80
timestamp 1586364061
transform 1 0 8464 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_4  FILLER_1_84
timestamp 1586364061
transform 1 0 8832 0 1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_0_89
timestamp 1586364061
transform 1 0 9292 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_85
timestamp 1586364061
transform 1 0 8924 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_1.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 9200 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__147__A
timestamp 1586364061
transform 1 0 9108 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_94
timestamp 1586364061
transform 1 0 9752 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_90
timestamp 1586364061
transform 1 0 9384 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 9568 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_1.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 9476 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_1.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 9936 0 1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_74
timestamp 1586364061
transform 1 0 9660 0 -1 2720
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  mem_top_ipin_1.LATCH_0_.latch tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 9752 0 -1 2720
box -38 -48 1050 592
use scs8hd_ebufn_2  mux_top_ipin_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 10396 0 1 2720
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_1.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 10948 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_105
timestamp 1586364061
transform 1 0 10764 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_0_109
timestamp 1586364061
transform 1 0 11132 0 -1 2720
box -38 -48 406 592
use scs8hd_decap_3  FILLER_1_98
timestamp 1586364061
transform 1 0 10120 0 1 2720
box -38 -48 314 592
use scs8hd_fill_2  FILLER_1_110
timestamp 1586364061
transform 1 0 11224 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_114
timestamp 1586364061
transform 1 0 11592 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_116
timestamp 1586364061
transform 1 0 11776 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 11408 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11776 0 1 2720
box -38 -48 222 592
use scs8hd_inv_1  mux_top_ipin_1.INVTX1_0_.scs8hd_inv_1 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 11500 0 -1 2720
box -38 -48 314 592
use scs8hd_fill_2  FILLER_1_118
timestamp 1586364061
transform 1 0 11960 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_120
timestamp 1586364061
transform 1 0 12144 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 12328 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 12144 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_1.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 11960 0 -1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_80
timestamp 1586364061
transform 1 0 12328 0 1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_75
timestamp 1586364061
transform 1 0 12512 0 -1 2720
box -38 -48 130 592
use scs8hd_ebufn_2  mux_top_ipin_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12420 0 1 2720
box -38 -48 866 592
use scs8hd_ebufn_2  mux_top_ipin_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12604 0 -1 2720
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 13616 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 13432 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_1.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 13800 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_134
timestamp 1586364061
transform 1 0 13432 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_0_138
timestamp 1586364061
transform 1 0 13800 0 -1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_1_132
timestamp 1586364061
transform 1 0 13248 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_136
timestamp 1586364061
transform 1 0 13616 0 1 2720
box -38 -48 222 592
use scs8hd_conb_1  _140_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 13984 0 1 2720
box -38 -48 314 592
use scs8hd_buf_2  _145_
timestamp 1586364061
transform 1 0 14168 0 -1 2720
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__145__A
timestamp 1586364061
transform 1 0 14720 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_146
timestamp 1586364061
transform 1 0 14536 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_0_150
timestamp 1586364061
transform 1 0 14904 0 -1 2720
box -38 -48 406 592
use scs8hd_decap_12  FILLER_1_143
timestamp 1586364061
transform 1 0 14260 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_76
timestamp 1586364061
transform 1 0 15364 0 -1 2720
box -38 -48 130 592
use scs8hd_fill_1  FILLER_0_154
timestamp 1586364061
transform 1 0 15272 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_12  FILLER_0_156
timestamp 1586364061
transform 1 0 15456 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_155
timestamp 1586364061
transform 1 0 15364 0 1 2720
box -38 -48 1142 592
use scs8hd_buf_2  _157_
timestamp 1586364061
transform 1 0 17112 0 -1 2720
box -38 -48 406 592
use scs8hd_decap_6  FILLER_0_168
timestamp 1586364061
transform 1 0 16560 0 -1 2720
box -38 -48 590 592
use scs8hd_fill_2  FILLER_0_178
timestamp 1586364061
transform 1 0 17480 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_12  FILLER_1_167
timestamp 1586364061
transform 1 0 16468 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_1_179
timestamp 1586364061
transform 1 0 17572 0 1 2720
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_77
timestamp 1586364061
transform 1 0 18216 0 -1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_81
timestamp 1586364061
transform 1 0 17940 0 1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__157__A
timestamp 1586364061
transform 1 0 17664 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_0_182
timestamp 1586364061
transform 1 0 17848 0 -1 2720
box -38 -48 406 592
use scs8hd_decap_12  FILLER_0_187
timestamp 1586364061
transform 1 0 18308 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_184
timestamp 1586364061
transform 1 0 18032 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_199
timestamp 1586364061
transform 1 0 19412 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_196
timestamp 1586364061
transform 1 0 19136 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_78
timestamp 1586364061
transform 1 0 21068 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_211
timestamp 1586364061
transform 1 0 20516 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_0_218
timestamp 1586364061
transform 1 0 21160 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_208
timestamp 1586364061
transform 1 0 20240 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_220
timestamp 1586364061
transform 1 0 21344 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_3  PHY_1
timestamp 1586364061
transform -1 0 22816 0 -1 2720
box -38 -48 314 592
use scs8hd_decap_3  PHY_3
timestamp 1586364061
transform -1 0 22816 0 1 2720
box -38 -48 314 592
use scs8hd_decap_3  FILLER_0_230
timestamp 1586364061
transform 1 0 22264 0 -1 2720
box -38 -48 314 592
use scs8hd_fill_1  FILLER_1_232
timestamp 1586364061
transform 1 0 22448 0 1 2720
box -38 -48 130 592
use scs8hd_decap_3  PHY_4
timestamp 1586364061
transform 1 0 1104 0 -1 3808
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 1564 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 1932 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_3
timestamp 1586364061
transform 1 0 1380 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_7
timestamp 1586364061
transform 1 0 1748 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_12  FILLER_2_11
timestamp 1586364061
transform 1 0 2116 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_2_23 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 3220 0 -1 3808
box -38 -48 774 592
use scs8hd_inv_8  _042_
timestamp 1586364061
transform 1 0 4048 0 -1 3808
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_82
timestamp 1586364061
transform 1 0 3956 0 -1 3808
box -38 -48 130 592
use scs8hd_fill_2  FILLER_2_41
timestamp 1586364061
transform 1 0 4876 0 -1 3808
box -38 -48 222 592
use scs8hd_inv_8  _050_
timestamp 1586364061
transform 1 0 5796 0 -1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__061__A
timestamp 1586364061
transform 1 0 5520 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__057__B
timestamp 1586364061
transform 1 0 5060 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_3  FILLER_2_45
timestamp 1586364061
transform 1 0 5244 0 -1 3808
box -38 -48 314 592
use scs8hd_fill_1  FILLER_2_50
timestamp 1586364061
transform 1 0 5704 0 -1 3808
box -38 -48 130 592
use scs8hd_nand2_4  _067_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 7360 0 -1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__053__C
timestamp 1586364061
transform 1 0 7084 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_2_60
timestamp 1586364061
transform 1 0 6624 0 -1 3808
box -38 -48 406 592
use scs8hd_fill_1  FILLER_2_64
timestamp 1586364061
transform 1 0 6992 0 -1 3808
box -38 -48 130 592
use scs8hd_fill_1  FILLER_2_67
timestamp 1586364061
transform 1 0 7268 0 -1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__106__C
timestamp 1586364061
transform 1 0 8372 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_77
timestamp 1586364061
transform 1 0 8188 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_8  FILLER_2_81
timestamp 1586364061
transform 1 0 8556 0 -1 3808
box -38 -48 774 592
use scs8hd_lpflow_inputisolatch_1  mem_top_ipin_1.LATCH_1_.latch
timestamp 1586364061
transform 1 0 9936 0 -1 3808
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_83
timestamp 1586364061
transform 1 0 9568 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_3  FILLER_2_89
timestamp 1586364061
transform 1 0 9292 0 -1 3808
box -38 -48 314 592
use scs8hd_decap_3  FILLER_2_93
timestamp 1586364061
transform 1 0 9660 0 -1 3808
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11132 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_107
timestamp 1586364061
transform 1 0 10948 0 -1 3808
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_ipin_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 11684 0 -1 3808
box -38 -48 866 592
use scs8hd_decap_4  FILLER_2_111
timestamp 1586364061
transform 1 0 11316 0 -1 3808
box -38 -48 406 592
use scs8hd_fill_2  FILLER_2_124
timestamp 1586364061
transform 1 0 12512 0 -1 3808
box -38 -48 222 592
use scs8hd_inv_1  mux_top_ipin_1.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 13248 0 -1 3808
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__043__A
timestamp 1586364061
transform 1 0 12696 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_2_128
timestamp 1586364061
transform 1 0 12880 0 -1 3808
box -38 -48 406 592
use scs8hd_decap_12  FILLER_2_135
timestamp 1586364061
transform 1 0 13524 0 -1 3808
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA__119__A
timestamp 1586364061
transform 1 0 14904 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_3  FILLER_2_147
timestamp 1586364061
transform 1 0 14628 0 -1 3808
box -38 -48 314 592
use scs8hd_fill_1  FILLER_2_152
timestamp 1586364061
transform 1 0 15088 0 -1 3808
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_84
timestamp 1586364061
transform 1 0 15180 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_2_154
timestamp 1586364061
transform 1 0 15272 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_166
timestamp 1586364061
transform 1 0 16376 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_2_178
timestamp 1586364061
transform 1 0 17480 0 -1 3808
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA__118__A
timestamp 1586364061
transform 1 0 18032 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_12  FILLER_2_186
timestamp 1586364061
transform 1 0 18216 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_198
timestamp 1586364061
transform 1 0 19320 0 -1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_85
timestamp 1586364061
transform 1 0 20792 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_4  FILLER_2_210
timestamp 1586364061
transform 1 0 20424 0 -1 3808
box -38 -48 406 592
use scs8hd_decap_12  FILLER_2_215
timestamp 1586364061
transform 1 0 20884 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_3  PHY_5
timestamp 1586364061
transform -1 0 22816 0 -1 3808
box -38 -48 314 592
use scs8hd_decap_6  FILLER_2_227
timestamp 1586364061
transform 1 0 21988 0 -1 3808
box -38 -48 590 592
use scs8hd_inv_8  _045_
timestamp 1586364061
transform 1 0 1564 0 1 3808
box -38 -48 866 592
use scs8hd_decap_3  PHY_6
timestamp 1586364061
transform 1 0 1104 0 1 3808
box -38 -48 314 592
use scs8hd_fill_2  FILLER_3_3
timestamp 1586364061
transform 1 0 1380 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__054__B
timestamp 1586364061
transform 1 0 3404 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__045__A
timestamp 1586364061
transform 1 0 2576 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_14
timestamp 1586364061
transform 1 0 2392 0 1 3808
box -38 -48 222 592
use scs8hd_decap_6  FILLER_3_18
timestamp 1586364061
transform 1 0 2760 0 1 3808
box -38 -48 590 592
use scs8hd_fill_1  FILLER_3_24
timestamp 1586364061
transform 1 0 3312 0 1 3808
box -38 -48 130 592
use scs8hd_fill_2  FILLER_3_27
timestamp 1586364061
transform 1 0 3588 0 1 3808
box -38 -48 222 592
use scs8hd_or3_4  _057_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 4692 0 1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__057__C
timestamp 1586364061
transform 1 0 4508 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__057__A
timestamp 1586364061
transform 1 0 4140 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__054__A
timestamp 1586364061
transform 1 0 3772 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_31
timestamp 1586364061
transform 1 0 3956 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_35
timestamp 1586364061
transform 1 0 4324 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__061__C
timestamp 1586364061
transform 1 0 5704 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__061__B
timestamp 1586364061
transform 1 0 6072 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_48
timestamp 1586364061
transform 1 0 5520 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_52
timestamp 1586364061
transform 1 0 5888 0 1 3808
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_86
timestamp 1586364061
transform 1 0 6716 0 1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__053__A
timestamp 1586364061
transform 1 0 7084 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__053__B
timestamp 1586364061
transform 1 0 6532 0 1 3808
box -38 -48 222 592
use scs8hd_decap_3  FILLER_3_56
timestamp 1586364061
transform 1 0 6256 0 1 3808
box -38 -48 314 592
use scs8hd_decap_3  FILLER_3_62
timestamp 1586364061
transform 1 0 6808 0 1 3808
box -38 -48 314 592
use scs8hd_decap_4  FILLER_3_67
timestamp 1586364061
transform 1 0 7268 0 1 3808
box -38 -48 406 592
use scs8hd_nor3_4  _106_
timestamp 1586364061
transform 1 0 7912 0 1 3808
box -38 -48 1234 592
use scs8hd_diode_2  ANTENNA__106__A
timestamp 1586364061
transform 1 0 7728 0 1 3808
box -38 -48 222 592
use scs8hd_fill_1  FILLER_3_71
timestamp 1586364061
transform 1 0 7636 0 1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__052__A
timestamp 1586364061
transform 1 0 9660 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__044__A
timestamp 1586364061
transform 1 0 9292 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_87
timestamp 1586364061
transform 1 0 9108 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_91
timestamp 1586364061
transform 1 0 9476 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_95
timestamp 1586364061
transform 1 0 9844 0 1 3808
box -38 -48 222 592
use scs8hd_inv_8  _044_
timestamp 1586364061
transform 1 0 10028 0 1 3808
box -38 -48 866 592
use scs8hd_decap_6  FILLER_3_106
timestamp 1586364061
transform 1 0 10856 0 1 3808
box -38 -48 590 592
use scs8hd_inv_8  _043_
timestamp 1586364061
transform 1 0 12420 0 1 3808
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_87
timestamp 1586364061
transform 1 0 12328 0 1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__122__B
timestamp 1586364061
transform 1 0 11868 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__122__A
timestamp 1586364061
transform 1 0 11500 0 1 3808
box -38 -48 222 592
use scs8hd_fill_1  FILLER_3_112
timestamp 1586364061
transform 1 0 11408 0 1 3808
box -38 -48 130 592
use scs8hd_fill_2  FILLER_3_115
timestamp 1586364061
transform 1 0 11684 0 1 3808
box -38 -48 222 592
use scs8hd_decap_3  FILLER_3_119
timestamp 1586364061
transform 1 0 12052 0 1 3808
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__117__B
timestamp 1586364061
transform 1 0 13432 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__117__A
timestamp 1586364061
transform 1 0 13800 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_132
timestamp 1586364061
transform 1 0 13248 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_136
timestamp 1586364061
transform 1 0 13616 0 1 3808
box -38 -48 222 592
use scs8hd_nor2_4  _119_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 14904 0 1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__119__B
timestamp 1586364061
transform 1 0 14720 0 1 3808
box -38 -48 222 592
use scs8hd_decap_8  FILLER_3_140
timestamp 1586364061
transform 1 0 13984 0 1 3808
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_1.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 15916 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_1.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 16284 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_159
timestamp 1586364061
transform 1 0 15732 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_163
timestamp 1586364061
transform 1 0 16100 0 1 3808
box -38 -48 222 592
use scs8hd_decap_12  FILLER_3_167
timestamp 1586364061
transform 1 0 16468 0 1 3808
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_3_179
timestamp 1586364061
transform 1 0 17572 0 1 3808
box -38 -48 222 592
use scs8hd_nor2_4  _118_
timestamp 1586364061
transform 1 0 18032 0 1 3808
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_88
timestamp 1586364061
transform 1 0 17940 0 1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__118__B
timestamp 1586364061
transform 1 0 17756 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_193
timestamp 1586364061
transform 1 0 18860 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_1.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 19044 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_1.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 19412 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_197
timestamp 1586364061
transform 1 0 19228 0 1 3808
box -38 -48 222 592
use scs8hd_decap_12  FILLER_3_201
timestamp 1586364061
transform 1 0 19596 0 1 3808
box -38 -48 1142 592
use scs8hd_inv_1  mux_bottom_ipin_1.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 20884 0 1 3808
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 21344 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_213
timestamp 1586364061
transform 1 0 20700 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_218
timestamp 1586364061
transform 1 0 21160 0 1 3808
box -38 -48 222 592
use scs8hd_decap_3  PHY_7
timestamp 1586364061
transform -1 0 22816 0 1 3808
box -38 -48 314 592
use scs8hd_decap_8  FILLER_3_222
timestamp 1586364061
transform 1 0 21528 0 1 3808
box -38 -48 774 592
use scs8hd_decap_3  FILLER_3_230
timestamp 1586364061
transform 1 0 22264 0 1 3808
box -38 -48 314 592
use scs8hd_ebufn_2  mux_top_ipin_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 1380 0 -1 4896
box -38 -48 866 592
use scs8hd_decap_3  PHY_8
timestamp 1586364061
transform 1 0 1104 0 -1 4896
box -38 -48 314 592
use scs8hd_fill_2  FILLER_4_12
timestamp 1586364061
transform 1 0 2208 0 -1 4896
box -38 -48 222 592
use scs8hd_conb_1  _141_
timestamp 1586364061
transform 1 0 2944 0 -1 4896
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 2392 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_4_16
timestamp 1586364061
transform 1 0 2576 0 -1 4896
box -38 -48 406 592
use scs8hd_decap_8  FILLER_4_23
timestamp 1586364061
transform 1 0 3220 0 -1 4896
box -38 -48 774 592
use scs8hd_or2_4  _054_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 4140 0 -1 4896
box -38 -48 682 592
use scs8hd_tapvpwrvgnd_1  PHY_89
timestamp 1586364061
transform 1 0 3956 0 -1 4896
box -38 -48 130 592
use scs8hd_fill_1  FILLER_4_32
timestamp 1586364061
transform 1 0 4048 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_4  FILLER_4_40
timestamp 1586364061
transform 1 0 4784 0 -1 4896
box -38 -48 406 592
use scs8hd_or3_4  _061_
timestamp 1586364061
transform 1 0 5520 0 -1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__063__B
timestamp 1586364061
transform 1 0 5152 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_46
timestamp 1586364061
transform 1 0 5336 0 -1 4896
box -38 -48 222 592
use scs8hd_or3_4  _053_
timestamp 1586364061
transform 1 0 7084 0 -1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__059__C
timestamp 1586364061
transform 1 0 6532 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_57
timestamp 1586364061
transform 1 0 6348 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_4_61
timestamp 1586364061
transform 1 0 6716 0 -1 4896
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__106__B
timestamp 1586364061
transform 1 0 8096 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_74
timestamp 1586364061
transform 1 0 7912 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_12  FILLER_4_78
timestamp 1586364061
transform 1 0 8280 0 -1 4896
box -38 -48 1142 592
use scs8hd_inv_8  _052_
timestamp 1586364061
transform 1 0 9660 0 -1 4896
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_90
timestamp 1586364061
transform 1 0 9568 0 -1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__075__C
timestamp 1586364061
transform 1 0 9384 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_12  FILLER_4_102
timestamp 1586364061
transform 1 0 10488 0 -1 4896
box -38 -48 1142 592
use scs8hd_nor2_4  _122_
timestamp 1586364061
transform 1 0 11868 0 -1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__123__B
timestamp 1586364061
transform 1 0 11592 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_1  FILLER_4_116
timestamp 1586364061
transform 1 0 11776 0 -1 4896
box -38 -48 130 592
use scs8hd_or2_4  _117_
timestamp 1586364061
transform 1 0 13432 0 -1 4896
box -38 -48 682 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 13156 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_4_126
timestamp 1586364061
transform 1 0 12696 0 -1 4896
box -38 -48 406 592
use scs8hd_fill_1  FILLER_4_130
timestamp 1586364061
transform 1 0 13064 0 -1 4896
box -38 -48 130 592
use scs8hd_fill_1  FILLER_4_133
timestamp 1586364061
transform 1 0 13340 0 -1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14260 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_141
timestamp 1586364061
transform 1 0 14076 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_8  FILLER_4_145
timestamp 1586364061
transform 1 0 14444 0 -1 4896
box -38 -48 774 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_1.LATCH_4_.latch
timestamp 1586364061
transform 1 0 15456 0 -1 4896
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_91
timestamp 1586364061
transform 1 0 15180 0 -1 4896
box -38 -48 130 592
use scs8hd_fill_2  FILLER_4_154
timestamp 1586364061
transform 1 0 15272 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 16652 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 17480 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_167
timestamp 1586364061
transform 1 0 16468 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_6  FILLER_4_171
timestamp 1586364061
transform 1 0 16836 0 -1 4896
box -38 -48 590 592
use scs8hd_fill_1  FILLER_4_177
timestamp 1586364061
transform 1 0 17388 0 -1 4896
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_1.LATCH_5_.latch
timestamp 1586364061
transform 1 0 18584 0 -1 4896
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_1.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 18032 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_4_180
timestamp 1586364061
transform 1 0 17664 0 -1 4896
box -38 -48 406 592
use scs8hd_decap_4  FILLER_4_186
timestamp 1586364061
transform 1 0 18216 0 -1 4896
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 19780 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_201
timestamp 1586364061
transform 1 0 19596 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_8  FILLER_4_205
timestamp 1586364061
transform 1 0 19964 0 -1 4896
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_92
timestamp 1586364061
transform 1 0 20792 0 -1 4896
box -38 -48 130 592
use scs8hd_fill_1  FILLER_4_213
timestamp 1586364061
transform 1 0 20700 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_4_215
timestamp 1586364061
transform 1 0 20884 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_3  PHY_9
timestamp 1586364061
transform -1 0 22816 0 -1 4896
box -38 -48 314 592
use scs8hd_decap_6  FILLER_4_227
timestamp 1586364061
transform 1 0 21988 0 -1 4896
box -38 -48 590 592
use scs8hd_lpflow_inputisolatch_1  mem_top_ipin_2.LATCH_1_.latch
timestamp 1586364061
transform 1 0 1932 0 1 4896
box -38 -48 1050 592
use scs8hd_decap_3  PHY_10
timestamp 1586364061
transform 1 0 1104 0 1 4896
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_2.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 1748 0 1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_5_3
timestamp 1586364061
transform 1 0 1380 0 1 4896
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_2.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 3128 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_20
timestamp 1586364061
transform 1 0 2944 0 1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_5_24
timestamp 1586364061
transform 1 0 3312 0 1 4896
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__108__A
timestamp 1586364061
transform 1 0 4048 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__108__B
timestamp 1586364061
transform 1 0 4416 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__108__C
timestamp 1586364061
transform 1 0 3680 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_30
timestamp 1586364061
transform 1 0 3864 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_34
timestamp 1586364061
transform 1 0 4232 0 1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_5_38
timestamp 1586364061
transform 1 0 4600 0 1 4896
box -38 -48 406 592
use scs8hd_or3_4  _063_
timestamp 1586364061
transform 1 0 5152 0 1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__063__A
timestamp 1586364061
transform 1 0 4968 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__059__B
timestamp 1586364061
transform 1 0 6164 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_53
timestamp 1586364061
transform 1 0 5980 0 1 4896
box -38 -48 222 592
use scs8hd_inv_8  _047_
timestamp 1586364061
transform 1 0 6808 0 1 4896
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_93
timestamp 1586364061
transform 1 0 6716 0 1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__047__A
timestamp 1586364061
transform 1 0 6532 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_57
timestamp 1586364061
transform 1 0 6348 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__098__A
timestamp 1586364061
transform 1 0 7820 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__075__A
timestamp 1586364061
transform 1 0 8556 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__098__B
timestamp 1586364061
transform 1 0 8188 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_71
timestamp 1586364061
transform 1 0 7636 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_75
timestamp 1586364061
transform 1 0 8004 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_79
timestamp 1586364061
transform 1 0 8372 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_83
timestamp 1586364061
transform 1 0 8740 0 1 4896
box -38 -48 222 592
use scs8hd_or3_4  _075_
timestamp 1586364061
transform 1 0 9476 0 1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__075__B
timestamp 1586364061
transform 1 0 9292 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__083__A
timestamp 1586364061
transform 1 0 8924 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_87
timestamp 1586364061
transform 1 0 9108 0 1 4896
box -38 -48 222 592
use scs8hd_inv_1  mux_top_ipin_1.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 11040 0 1 4896
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__083__C
timestamp 1586364061
transform 1 0 10488 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__083__B
timestamp 1586364061
transform 1 0 10856 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_100
timestamp 1586364061
transform 1 0 10304 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_104
timestamp 1586364061
transform 1 0 10672 0 1 4896
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_1.LATCH_1_.latch
timestamp 1586364061
transform 1 0 12512 0 1 4896
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_94
timestamp 1586364061
transform 1 0 12328 0 1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_1.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 11500 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_1.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 12144 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_111
timestamp 1586364061
transform 1 0 11316 0 1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_5_115
timestamp 1586364061
transform 1 0 11684 0 1 4896
box -38 -48 406 592
use scs8hd_fill_1  FILLER_5_119
timestamp 1586364061
transform 1 0 12052 0 1 4896
box -38 -48 130 592
use scs8hd_fill_1  FILLER_5_123
timestamp 1586364061
transform 1 0 12420 0 1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 13708 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_135
timestamp 1586364061
transform 1 0 13524 0 1 4896
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_ipin_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 14260 0 1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 14076 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_139
timestamp 1586364061
transform 1 0 13892 0 1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_5_152
timestamp 1586364061
transform 1 0 15088 0 1 4896
box -38 -48 406 592
use scs8hd_ebufn_2  mux_bottom_ipin_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 16192 0 1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__120__B
timestamp 1586364061
transform 1 0 15916 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__120__A
timestamp 1586364061
transform 1 0 15548 0 1 4896
box -38 -48 222 592
use scs8hd_fill_1  FILLER_5_156
timestamp 1586364061
transform 1 0 15456 0 1 4896
box -38 -48 130 592
use scs8hd_fill_2  FILLER_5_159
timestamp 1586364061
transform 1 0 15732 0 1 4896
box -38 -48 222 592
use scs8hd_fill_1  FILLER_5_163
timestamp 1586364061
transform 1 0 16100 0 1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 17388 0 1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_5_173
timestamp 1586364061
transform 1 0 17020 0 1 4896
box -38 -48 406 592
use scs8hd_fill_2  FILLER_5_179
timestamp 1586364061
transform 1 0 17572 0 1 4896
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_1.LATCH_3_.latch
timestamp 1586364061
transform 1 0 18032 0 1 4896
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_95
timestamp 1586364061
transform 1 0 17940 0 1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_1.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 17756 0 1 4896
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_ipin_1.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 19780 0 1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 19596 0 1 4896
box -38 -48 222 592
use scs8hd_decap_6  FILLER_5_195
timestamp 1586364061
transform 1 0 19044 0 1 4896
box -38 -48 590 592
use scs8hd_decap_12  FILLER_5_212
timestamp 1586364061
transform 1 0 20608 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_3  PHY_11
timestamp 1586364061
transform -1 0 22816 0 1 4896
box -38 -48 314 592
use scs8hd_decap_8  FILLER_5_224
timestamp 1586364061
transform 1 0 21712 0 1 4896
box -38 -48 774 592
use scs8hd_fill_1  FILLER_5_232
timestamp 1586364061
transform 1 0 22448 0 1 4896
box -38 -48 130 592
use scs8hd_fill_2  FILLER_7_6
timestamp 1586364061
transform 1 0 1656 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_3
timestamp 1586364061
transform 1 0 1380 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 1564 0 -1 5984
box -38 -48 222 592
use scs8hd_decap_3  PHY_14
timestamp 1586364061
transform 1 0 1104 0 1 5984
box -38 -48 314 592
use scs8hd_decap_3  PHY_12
timestamp 1586364061
transform 1 0 1104 0 -1 5984
box -38 -48 314 592
use scs8hd_inv_1  mux_top_ipin_2.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1380 0 1 5984
box -38 -48 314 592
use scs8hd_fill_2  FILLER_7_10
timestamp 1586364061
transform 1 0 2024 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_2.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 2208 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_2.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 1840 0 1 5984
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_ipin_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 1748 0 -1 5984
box -38 -48 866 592
use scs8hd_fill_1  FILLER_7_18
timestamp 1586364061
transform 1 0 2760 0 1 5984
box -38 -48 130 592
use scs8hd_decap_4  FILLER_7_14
timestamp 1586364061
transform 1 0 2392 0 1 5984
box -38 -48 406 592
use scs8hd_decap_4  FILLER_6_20
timestamp 1586364061
transform 1 0 2944 0 -1 5984
box -38 -48 406 592
use scs8hd_fill_2  FILLER_6_16
timestamp 1586364061
transform 1 0 2576 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_2.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 2760 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__109__B
timestamp 1586364061
transform 1 0 2852 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_21
timestamp 1586364061
transform 1 0 3036 0 1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_6_27
timestamp 1586364061
transform 1 0 3588 0 -1 5984
box -38 -48 406 592
use scs8hd_fill_1  FILLER_6_24
timestamp 1586364061
transform 1 0 3312 0 -1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__109__A
timestamp 1586364061
transform 1 0 3404 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__109__C
timestamp 1586364061
transform 1 0 3220 0 1 5984
box -38 -48 222 592
use scs8hd_nor3_4  _109_
timestamp 1586364061
transform 1 0 3404 0 1 5984
box -38 -48 1234 592
use scs8hd_nor3_4  _108_
timestamp 1586364061
transform 1 0 4048 0 -1 5984
box -38 -48 1234 592
use scs8hd_tapvpwrvgnd_1  PHY_96
timestamp 1586364061
transform 1 0 3956 0 -1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_5.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 4784 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_38
timestamp 1586364061
transform 1 0 4600 0 1 5984
box -38 -48 222 592
use scs8hd_decap_6  FILLER_7_42
timestamp 1586364061
transform 1 0 4968 0 1 5984
box -38 -48 590 592
use scs8hd_fill_2  FILLER_6_45
timestamp 1586364061
transform 1 0 5244 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__063__C
timestamp 1586364061
transform 1 0 5428 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__065__C
timestamp 1586364061
transform 1 0 5520 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_54
timestamp 1586364061
transform 1 0 6072 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_50
timestamp 1586364061
transform 1 0 5704 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_49
timestamp 1586364061
transform 1 0 5612 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__059__A
timestamp 1586364061
transform 1 0 5796 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__065__A
timestamp 1586364061
transform 1 0 5888 0 1 5984
box -38 -48 222 592
use scs8hd_or3_4  _059_
timestamp 1586364061
transform 1 0 5980 0 -1 5984
box -38 -48 866 592
use scs8hd_decap_3  FILLER_7_58
timestamp 1586364061
transform 1 0 6440 0 1 5984
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__065__B
timestamp 1586364061
transform 1 0 6256 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_62
timestamp 1586364061
transform 1 0 6808 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_62
timestamp 1586364061
transform 1 0 6808 0 -1 5984
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_100
timestamp 1586364061
transform 1 0 6716 0 1 5984
box -38 -48 130 592
use scs8hd_fill_2  FILLER_7_66
timestamp 1586364061
transform 1 0 7176 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_66
timestamp 1586364061
transform 1 0 7176 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__110__A
timestamp 1586364061
transform 1 0 6992 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__068__C
timestamp 1586364061
transform 1 0 6992 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__068__D
timestamp 1586364061
transform 1 0 7360 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__110__C
timestamp 1586364061
transform 1 0 7360 0 1 5984
box -38 -48 222 592
use scs8hd_or4_4  _068_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 7544 0 1 5984
box -38 -48 866 592
use scs8hd_or2_4  _098_
timestamp 1586364061
transform 1 0 7544 0 -1 5984
box -38 -48 682 592
use scs8hd_diode_2  ANTENNA__110__B
timestamp 1586364061
transform 1 0 8556 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__068__B
timestamp 1586364061
transform 1 0 8372 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_77
timestamp 1586364061
transform 1 0 8188 0 -1 5984
box -38 -48 222 592
use scs8hd_decap_6  FILLER_6_81
timestamp 1586364061
transform 1 0 8556 0 -1 5984
box -38 -48 590 592
use scs8hd_fill_2  FILLER_7_79
timestamp 1586364061
transform 1 0 8372 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_83
timestamp 1586364061
transform 1 0 8740 0 1 5984
box -38 -48 222 592
use scs8hd_or3_4  _083_
timestamp 1586364061
transform 1 0 9660 0 -1 5984
box -38 -48 866 592
use scs8hd_or4_4  _099_
timestamp 1586364061
transform 1 0 9108 0 1 5984
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_97
timestamp 1586364061
transform 1 0 9568 0 -1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__099__C
timestamp 1586364061
transform 1 0 8924 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__099__B
timestamp 1586364061
transform 1 0 9108 0 -1 5984
box -38 -48 222 592
use scs8hd_decap_3  FILLER_6_89
timestamp 1586364061
transform 1 0 9292 0 -1 5984
box -38 -48 314 592
use scs8hd_fill_2  FILLER_7_96
timestamp 1586364061
transform 1 0 9936 0 1 5984
box -38 -48 222 592
use scs8hd_inv_8  _051_
timestamp 1586364061
transform 1 0 10672 0 1 5984
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__051__A
timestamp 1586364061
transform 1 0 10488 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__099__A
timestamp 1586364061
transform 1 0 10120 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__055__A
timestamp 1586364061
transform 1 0 10672 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__055__C
timestamp 1586364061
transform 1 0 11040 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_102
timestamp 1586364061
transform 1 0 10488 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_106
timestamp 1586364061
transform 1 0 10856 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_110
timestamp 1586364061
transform 1 0 11224 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_100
timestamp 1586364061
transform 1 0 10304 0 1 5984
box -38 -48 222 592
use scs8hd_nor2_4  _123_
timestamp 1586364061
transform 1 0 11592 0 -1 5984
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_101
timestamp 1586364061
transform 1 0 12328 0 1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 11684 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__123__A
timestamp 1586364061
transform 1 0 11408 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_1.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 12144 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_123
timestamp 1586364061
transform 1 0 12420 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_113
timestamp 1586364061
transform 1 0 11500 0 1 5984
box -38 -48 222 592
use scs8hd_decap_3  FILLER_7_117
timestamp 1586364061
transform 1 0 11868 0 1 5984
box -38 -48 314 592
use scs8hd_fill_2  FILLER_7_123
timestamp 1586364061
transform 1 0 12420 0 1 5984
box -38 -48 222 592
use scs8hd_inv_1  mux_bottom_ipin_1.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 12604 0 1 5984
box -38 -48 314 592
use scs8hd_ebufn_2  mux_bottom_ipin_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 13616 0 1 5984
box -38 -48 866 592
use scs8hd_ebufn_2  mux_bottom_ipin_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 13156 0 -1 5984
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 13064 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_1.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 13432 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_1.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 12604 0 -1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_6_127
timestamp 1586364061
transform 1 0 12788 0 -1 5984
box -38 -48 406 592
use scs8hd_fill_2  FILLER_7_128
timestamp 1586364061
transform 1 0 12880 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_132
timestamp 1586364061
transform 1 0 13248 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_1.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 15088 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_1.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 14720 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14168 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_140
timestamp 1586364061
transform 1 0 13984 0 -1 5984
box -38 -48 222 592
use scs8hd_decap_8  FILLER_6_144
timestamp 1586364061
transform 1 0 14352 0 -1 5984
box -38 -48 774 592
use scs8hd_fill_1  FILLER_6_152
timestamp 1586364061
transform 1 0 15088 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_3  FILLER_7_145
timestamp 1586364061
transform 1 0 14444 0 1 5984
box -38 -48 314 592
use scs8hd_fill_2  FILLER_7_150
timestamp 1586364061
transform 1 0 14904 0 1 5984
box -38 -48 222 592
use scs8hd_nor2_4  _120_
timestamp 1586364061
transform 1 0 15916 0 -1 5984
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_1.LATCH_2_.latch
timestamp 1586364061
transform 1 0 15272 0 1 5984
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_98
timestamp 1586364061
transform 1 0 15180 0 -1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 15732 0 -1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_6_154
timestamp 1586364061
transform 1 0 15272 0 -1 5984
box -38 -48 406 592
use scs8hd_fill_1  FILLER_6_158
timestamp 1586364061
transform 1 0 15640 0 -1 5984
box -38 -48 130 592
use scs8hd_fill_2  FILLER_7_165
timestamp 1586364061
transform 1 0 16284 0 1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_7_169
timestamp 1586364061
transform 1 0 16652 0 1 5984
box -38 -48 406 592
use scs8hd_fill_2  FILLER_6_170
timestamp 1586364061
transform 1 0 16744 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 16928 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 16468 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_179
timestamp 1586364061
transform 1 0 17572 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_175
timestamp 1586364061
transform 1 0 17204 0 1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_6_174
timestamp 1586364061
transform 1 0 17112 0 -1 5984
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__094__A
timestamp 1586364061
transform 1 0 17020 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__121__B
timestamp 1586364061
transform 1 0 17388 0 1 5984
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_ipin_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 17480 0 -1 5984
box -38 -48 866 592
use scs8hd_nor2_4  _121_
timestamp 1586364061
transform 1 0 18032 0 1 5984
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_102
timestamp 1586364061
transform 1 0 17940 0 1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__094__B
timestamp 1586364061
transform 1 0 17756 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__121__A
timestamp 1586364061
transform 1 0 18492 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_187
timestamp 1586364061
transform 1 0 18308 0 -1 5984
box -38 -48 222 592
use scs8hd_decap_6  FILLER_6_191
timestamp 1586364061
transform 1 0 18676 0 -1 5984
box -38 -48 590 592
use scs8hd_decap_6  FILLER_7_193
timestamp 1586364061
transform 1 0 18860 0 1 5984
box -38 -48 590 592
use scs8hd_nor2_4  _092_
timestamp 1586364061
transform 1 0 19596 0 1 5984
box -38 -48 866 592
use scs8hd_conb_1  _132_
timestamp 1586364061
transform 1 0 19320 0 -1 5984
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__092__B
timestamp 1586364061
transform 1 0 19412 0 1 5984
box -38 -48 222 592
use scs8hd_fill_1  FILLER_6_197
timestamp 1586364061
transform 1 0 19228 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_201
timestamp 1586364061
transform 1 0 19596 0 -1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_99
timestamp 1586364061
transform 1 0 20792 0 -1 5984
box -38 -48 130 592
use scs8hd_fill_1  FILLER_6_213
timestamp 1586364061
transform 1 0 20700 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_215
timestamp 1586364061
transform 1 0 20884 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_210
timestamp 1586364061
transform 1 0 20424 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_3  PHY_13
timestamp 1586364061
transform -1 0 22816 0 -1 5984
box -38 -48 314 592
use scs8hd_decap_3  PHY_15
timestamp 1586364061
transform -1 0 22816 0 1 5984
box -38 -48 314 592
use scs8hd_decap_6  FILLER_6_227
timestamp 1586364061
transform 1 0 21988 0 -1 5984
box -38 -48 590 592
use scs8hd_decap_8  FILLER_7_222
timestamp 1586364061
transform 1 0 21528 0 1 5984
box -38 -48 774 592
use scs8hd_decap_3  FILLER_7_230
timestamp 1586364061
transform 1 0 22264 0 1 5984
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_top_ipin_2.LATCH_0_.latch
timestamp 1586364061
transform 1 0 1656 0 -1 7072
box -38 -48 1050 592
use scs8hd_decap_3  PHY_16
timestamp 1586364061
transform 1 0 1104 0 -1 7072
box -38 -48 314 592
use scs8hd_decap_3  FILLER_8_3
timestamp 1586364061
transform 1 0 1380 0 -1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__081__B
timestamp 1586364061
transform 1 0 3312 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 2852 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_17
timestamp 1586364061
transform 1 0 2668 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_3  FILLER_8_21
timestamp 1586364061
transform 1 0 3036 0 -1 7072
box -38 -48 314 592
use scs8hd_decap_4  FILLER_8_26
timestamp 1586364061
transform 1 0 3496 0 -1 7072
box -38 -48 406 592
use scs8hd_inv_1  mux_bottom_ipin_5.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 4232 0 -1 7072
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_103
timestamp 1586364061
transform 1 0 3956 0 -1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_5.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 4692 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_1  FILLER_8_30
timestamp 1586364061
transform 1 0 3864 0 -1 7072
box -38 -48 130 592
use scs8hd_fill_2  FILLER_8_32
timestamp 1586364061
transform 1 0 4048 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_37
timestamp 1586364061
transform 1 0 4508 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_3  FILLER_8_41
timestamp 1586364061
transform 1 0 4876 0 -1 7072
box -38 -48 314 592
use scs8hd_or3_4  _065_
timestamp 1586364061
transform 1 0 5520 0 -1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__080__A
timestamp 1586364061
transform 1 0 5152 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_46
timestamp 1586364061
transform 1 0 5336 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__076__B
timestamp 1586364061
transform 1 0 7176 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__068__A
timestamp 1586364061
transform 1 0 6808 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_8_57
timestamp 1586364061
transform 1 0 6348 0 -1 7072
box -38 -48 406 592
use scs8hd_fill_1  FILLER_8_61
timestamp 1586364061
transform 1 0 6716 0 -1 7072
box -38 -48 130 592
use scs8hd_fill_2  FILLER_8_64
timestamp 1586364061
transform 1 0 6992 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_68
timestamp 1586364061
transform 1 0 7360 0 -1 7072
box -38 -48 222 592
use scs8hd_or4_4  _110_
timestamp 1586364061
transform 1 0 7544 0 -1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__110__D
timestamp 1586364061
transform 1 0 8556 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_79
timestamp 1586364061
transform 1 0 8372 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_8_83
timestamp 1586364061
transform 1 0 8740 0 -1 7072
box -38 -48 406 592
use scs8hd_or4_4  _055_
timestamp 1586364061
transform 1 0 9844 0 -1 7072
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_104
timestamp 1586364061
transform 1 0 9568 0 -1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__099__D
timestamp 1586364061
transform 1 0 9108 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_3  FILLER_8_89
timestamp 1586364061
transform 1 0 9292 0 -1 7072
box -38 -48 314 592
use scs8hd_fill_2  FILLER_8_93
timestamp 1586364061
transform 1 0 9660 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__055__B
timestamp 1586364061
transform 1 0 10856 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__055__D
timestamp 1586364061
transform 1 0 11224 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_104
timestamp 1586364061
transform 1 0 10672 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_108
timestamp 1586364061
transform 1 0 11040 0 -1 7072
box -38 -48 222 592
use scs8hd_inv_1  mux_bottom_ipin_1.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 11592 0 -1 7072
box -38 -48 314 592
use scs8hd_fill_2  FILLER_8_112
timestamp 1586364061
transform 1 0 11408 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_8  FILLER_8_117
timestamp 1586364061
transform 1 0 11868 0 -1 7072
box -38 -48 774 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_1.LATCH_0_.latch
timestamp 1586364061
transform 1 0 12604 0 -1 7072
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 13800 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_136
timestamp 1586364061
transform 1 0 13616 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14168 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_140
timestamp 1586364061
transform 1 0 13984 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_8  FILLER_8_144
timestamp 1586364061
transform 1 0 14352 0 -1 7072
box -38 -48 774 592
use scs8hd_fill_1  FILLER_8_152
timestamp 1586364061
transform 1 0 15088 0 -1 7072
box -38 -48 130 592
use scs8hd_ebufn_2  mux_bottom_ipin_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 16008 0 -1 7072
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_105
timestamp 1586364061
transform 1 0 15180 0 -1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 15548 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_3  FILLER_8_154
timestamp 1586364061
transform 1 0 15272 0 -1 7072
box -38 -48 314 592
use scs8hd_decap_3  FILLER_8_159
timestamp 1586364061
transform 1 0 15732 0 -1 7072
box -38 -48 314 592
use scs8hd_decap_12  FILLER_8_171
timestamp 1586364061
transform 1 0 16836 0 -1 7072
box -38 -48 1142 592
use scs8hd_nor2_4  _094_
timestamp 1586364061
transform 1 0 17940 0 -1 7072
box -38 -48 866 592
use scs8hd_fill_2  FILLER_8_192
timestamp 1586364061
transform 1 0 18768 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_7.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 18952 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__092__A
timestamp 1586364061
transform 1 0 19596 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_7.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 19964 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_8_196
timestamp 1586364061
transform 1 0 19136 0 -1 7072
box -38 -48 406 592
use scs8hd_fill_1  FILLER_8_200
timestamp 1586364061
transform 1 0 19504 0 -1 7072
box -38 -48 130 592
use scs8hd_fill_2  FILLER_8_203
timestamp 1586364061
transform 1 0 19780 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_6  FILLER_8_207
timestamp 1586364061
transform 1 0 20148 0 -1 7072
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_106
timestamp 1586364061
transform 1 0 20792 0 -1 7072
box -38 -48 130 592
use scs8hd_fill_1  FILLER_8_213
timestamp 1586364061
transform 1 0 20700 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_8_215
timestamp 1586364061
transform 1 0 20884 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_3  PHY_17
timestamp 1586364061
transform -1 0 22816 0 -1 7072
box -38 -48 314 592
use scs8hd_decap_6  FILLER_8_227
timestamp 1586364061
transform 1 0 21988 0 -1 7072
box -38 -48 590 592
use scs8hd_ebufn_2  mux_top_ipin_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 1748 0 1 7072
box -38 -48 866 592
use scs8hd_decap_3  PHY_18
timestamp 1586364061
transform 1 0 1104 0 1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 1564 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_3
timestamp 1586364061
transform 1 0 1380 0 1 7072
box -38 -48 222 592
use scs8hd_nor2_4  _081_
timestamp 1586364061
transform 1 0 3312 0 1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_2.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 2944 0 1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_9_16
timestamp 1586364061
transform 1 0 2576 0 1 7072
box -38 -48 406 592
use scs8hd_fill_2  FILLER_9_22
timestamp 1586364061
transform 1 0 3128 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_5.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 4324 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_33
timestamp 1586364061
transform 1 0 4140 0 1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_9_37
timestamp 1586364061
transform 1 0 4508 0 1 7072
box -38 -48 406 592
use scs8hd_fill_1  FILLER_9_41
timestamp 1586364061
transform 1 0 4876 0 1 7072
box -38 -48 130 592
use scs8hd_nor2_4  _080_
timestamp 1586364061
transform 1 0 5152 0 1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__080__B
timestamp 1586364061
transform 1 0 4968 0 1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_9_53
timestamp 1586364061
transform 1 0 5980 0 1 7072
box -38 -48 406 592
use scs8hd_or2_4  _076_
timestamp 1586364061
transform 1 0 7176 0 1 7072
box -38 -48 682 592
use scs8hd_tapvpwrvgnd_1  PHY_107
timestamp 1586364061
transform 1 0 6716 0 1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_5.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 6440 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__076__A
timestamp 1586364061
transform 1 0 6992 0 1 7072
box -38 -48 222 592
use scs8hd_fill_1  FILLER_9_57
timestamp 1586364061
transform 1 0 6348 0 1 7072
box -38 -48 130 592
use scs8hd_fill_1  FILLER_9_60
timestamp 1586364061
transform 1 0 6624 0 1 7072
box -38 -48 130 592
use scs8hd_fill_2  FILLER_9_62
timestamp 1586364061
transform 1 0 6808 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_5.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 8188 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__084__B
timestamp 1586364061
transform 1 0 8740 0 1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_9_73
timestamp 1586364061
transform 1 0 7820 0 1 7072
box -38 -48 406 592
use scs8hd_decap_4  FILLER_9_79
timestamp 1586364061
transform 1 0 8372 0 1 7072
box -38 -48 406 592
use scs8hd_or4_4  _091_
timestamp 1586364061
transform 1 0 9660 0 1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__091__D
timestamp 1586364061
transform 1 0 9476 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__084__A
timestamp 1586364061
transform 1 0 9108 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_85
timestamp 1586364061
transform 1 0 8924 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_89
timestamp 1586364061
transform 1 0 9292 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_6.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 11040 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__091__A
timestamp 1586364061
transform 1 0 10672 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_102
timestamp 1586364061
transform 1 0 10488 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_106
timestamp 1586364061
transform 1 0 10856 0 1 7072
box -38 -48 222 592
use scs8hd_fill_1  FILLER_9_110
timestamp 1586364061
transform 1 0 11224 0 1 7072
box -38 -48 130 592
use scs8hd_inv_1  mux_bottom_ipin_6.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 11316 0 1 7072
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_108
timestamp 1586364061
transform 1 0 12328 0 1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_6.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 11776 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__124__A
timestamp 1586364061
transform 1 0 12144 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_114
timestamp 1586364061
transform 1 0 11592 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_118
timestamp 1586364061
transform 1 0 11960 0 1 7072
box -38 -48 222 592
use scs8hd_decap_3  FILLER_9_123
timestamp 1586364061
transform 1 0 12420 0 1 7072
box -38 -48 314 592
use scs8hd_inv_1  mux_bottom_ipin_1.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 12696 0 1 7072
box -38 -48 314 592
use scs8hd_ebufn_2  mux_bottom_ipin_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 13708 0 1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 13156 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__124__B
timestamp 1586364061
transform 1 0 13524 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_129
timestamp 1586364061
transform 1 0 12972 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_133
timestamp 1586364061
transform 1 0 13340 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 14720 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_146
timestamp 1586364061
transform 1 0 14536 0 1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_9_150
timestamp 1586364061
transform 1 0 14904 0 1 7072
box -38 -48 406 592
use scs8hd_ebufn_2  mux_bottom_ipin_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15548 0 1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 15272 0 1 7072
box -38 -48 222 592
use scs8hd_fill_1  FILLER_9_156
timestamp 1586364061
transform 1 0 15456 0 1 7072
box -38 -48 130 592
use scs8hd_fill_2  FILLER_9_166
timestamp 1586364061
transform 1 0 16376 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_7.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 16560 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_7.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 16928 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_170
timestamp 1586364061
transform 1 0 16744 0 1 7072
box -38 -48 222 592
use scs8hd_decap_8  FILLER_9_174
timestamp 1586364061
transform 1 0 17112 0 1 7072
box -38 -48 774 592
use scs8hd_inv_1  mux_bottom_ipin_1.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 18032 0 1 7072
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_109
timestamp 1586364061
transform 1 0 17940 0 1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 18492 0 1 7072
box -38 -48 222 592
use scs8hd_fill_1  FILLER_9_182
timestamp 1586364061
transform 1 0 17848 0 1 7072
box -38 -48 130 592
use scs8hd_fill_2  FILLER_9_187
timestamp 1586364061
transform 1 0 18308 0 1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_9_191
timestamp 1586364061
transform 1 0 18676 0 1 7072
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_7.LATCH_5_.latch
timestamp 1586364061
transform 1 0 19320 0 1 7072
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_7.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 19136 0 1 7072
box -38 -48 222 592
use scs8hd_fill_1  FILLER_9_195
timestamp 1586364061
transform 1 0 19044 0 1 7072
box -38 -48 130 592
use scs8hd_conb_1  _138_
timestamp 1586364061
transform 1 0 21068 0 1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_7.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 20884 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_7.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 20516 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_209
timestamp 1586364061
transform 1 0 20332 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_213
timestamp 1586364061
transform 1 0 20700 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_220
timestamp 1586364061
transform 1 0 21344 0 1 7072
box -38 -48 222 592
use scs8hd_decap_3  PHY_19
timestamp 1586364061
transform -1 0 22816 0 1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_7.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 21528 0 1 7072
box -38 -48 222 592
use scs8hd_decap_8  FILLER_9_224
timestamp 1586364061
transform 1 0 21712 0 1 7072
box -38 -48 774 592
use scs8hd_fill_1  FILLER_9_232
timestamp 1586364061
transform 1 0 22448 0 1 7072
box -38 -48 130 592
use scs8hd_ebufn_2  mux_top_ipin_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 1380 0 -1 8160
box -38 -48 866 592
use scs8hd_decap_3  PHY_20
timestamp 1586364061
transform 1 0 1104 0 -1 8160
box -38 -48 314 592
use scs8hd_fill_2  FILLER_10_12
timestamp 1586364061
transform 1 0 2208 0 -1 8160
box -38 -48 222 592
use scs8hd_inv_1  mux_top_ipin_2.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 2944 0 -1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__081__A
timestamp 1586364061
transform 1 0 3404 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 2392 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 2760 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_16
timestamp 1586364061
transform 1 0 2576 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_23
timestamp 1586364061
transform 1 0 3220 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_10_27
timestamp 1586364061
transform 1 0 3588 0 -1 8160
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_5.LATCH_1_.latch
timestamp 1586364061
transform 1 0 4048 0 -1 8160
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_110
timestamp 1586364061
transform 1 0 3956 0 -1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_5.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 5244 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_43
timestamp 1586364061
transform 1 0 5060 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_8  FILLER_10_47
timestamp 1586364061
transform 1 0 5428 0 -1 8160
box -38 -48 774 592
use scs8hd_fill_1  FILLER_10_55
timestamp 1586364061
transform 1 0 6164 0 -1 8160
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_5.LATCH_2_.latch
timestamp 1586364061
transform 1 0 6440 0 -1 8160
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_5.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 6256 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_69
timestamp 1586364061
transform 1 0 7452 0 -1 8160
box -38 -48 222 592
use scs8hd_inv_1  mux_bottom_ipin_5.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 8188 0 -1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_5.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 7636 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_10_73
timestamp 1586364061
transform 1 0 7820 0 -1 8160
box -38 -48 406 592
use scs8hd_decap_8  FILLER_10_80
timestamp 1586364061
transform 1 0 8464 0 -1 8160
box -38 -48 774 592
use scs8hd_or2_4  _084_
timestamp 1586364061
transform 1 0 9660 0 -1 8160
box -38 -48 682 592
use scs8hd_tapvpwrvgnd_1  PHY_111
timestamp 1586364061
transform 1 0 9568 0 -1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__091__C
timestamp 1586364061
transform 1 0 9384 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_88
timestamp 1586364061
transform 1 0 9200 0 -1 8160
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_6.LATCH_0_.latch
timestamp 1586364061
transform 1 0 11040 0 -1 8160
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA__091__B
timestamp 1586364061
transform 1 0 10488 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_6.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 10856 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_100
timestamp 1586364061
transform 1 0 10304 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_104
timestamp 1586364061
transform 1 0 10672 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_6.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 12236 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_119
timestamp 1586364061
transform 1 0 12052 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_123
timestamp 1586364061
transform 1 0 12420 0 -1 8160
box -38 -48 222 592
use scs8hd_or2_4  _124_
timestamp 1586364061
transform 1 0 12788 0 -1 8160
box -38 -48 682 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 13708 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_6.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 12604 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_3  FILLER_10_134
timestamp 1586364061
transform 1 0 13432 0 -1 8160
box -38 -48 314 592
use scs8hd_inv_1  mux_bottom_ipin_1.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 14168 0 -1 8160
box -38 -48 314 592
use scs8hd_decap_3  FILLER_10_139
timestamp 1586364061
transform 1 0 13892 0 -1 8160
box -38 -48 314 592
use scs8hd_decap_8  FILLER_10_145
timestamp 1586364061
transform 1 0 14444 0 -1 8160
box -38 -48 774 592
use scs8hd_inv_1  mux_bottom_ipin_1.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 15272 0 -1 8160
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_112
timestamp 1586364061
transform 1 0 15180 0 -1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_7.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 15732 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 16100 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_157
timestamp 1586364061
transform 1 0 15548 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_161
timestamp 1586364061
transform 1 0 15916 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_3  FILLER_10_165
timestamp 1586364061
transform 1 0 16284 0 -1 8160
box -38 -48 314 592
use scs8hd_ebufn_2  mux_bottom_ipin_7.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 16560 0 -1 8160
box -38 -48 866 592
use scs8hd_decap_8  FILLER_10_177
timestamp 1586364061
transform 1 0 17388 0 -1 8160
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA__093__A
timestamp 1586364061
transform 1 0 18124 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_6  FILLER_10_187
timestamp 1586364061
transform 1 0 18308 0 -1 8160
box -38 -48 590 592
use scs8hd_fill_1  FILLER_10_193
timestamp 1586364061
transform 1 0 18860 0 -1 8160
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_7.LATCH_3_.latch
timestamp 1586364061
transform 1 0 18952 0 -1 8160
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_7.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 20148 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_205
timestamp 1586364061
transform 1 0 19964 0 -1 8160
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_ipin_7.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 20884 0 -1 8160
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_113
timestamp 1586364061
transform 1 0 20792 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_4  FILLER_10_209
timestamp 1586364061
transform 1 0 20332 0 -1 8160
box -38 -48 406 592
use scs8hd_fill_1  FILLER_10_213
timestamp 1586364061
transform 1 0 20700 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_3  PHY_21
timestamp 1586364061
transform -1 0 22816 0 -1 8160
box -38 -48 314 592
use scs8hd_decap_8  FILLER_10_224
timestamp 1586364061
transform 1 0 21712 0 -1 8160
box -38 -48 774 592
use scs8hd_fill_1  FILLER_10_232
timestamp 1586364061
transform 1 0 22448 0 -1 8160
box -38 -48 130 592
use scs8hd_inv_8  _046_
timestamp 1586364061
transform 1 0 1380 0 1 8160
box -38 -48 866 592
use scs8hd_decap_3  PHY_22
timestamp 1586364061
transform 1 0 1104 0 1 8160
box -38 -48 314 592
use scs8hd_fill_2  FILLER_11_12
timestamp 1586364061
transform 1 0 2208 0 1 8160
box -38 -48 222 592
use scs8hd_inv_1  mux_bottom_ipin_5.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 3404 0 1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__079__B
timestamp 1586364061
transform 1 0 2392 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__079__A
timestamp 1586364061
transform 1 0 2760 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__046__A
timestamp 1586364061
transform 1 0 3128 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_16
timestamp 1586364061
transform 1 0 2576 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_20
timestamp 1586364061
transform 1 0 2944 0 1 8160
box -38 -48 222 592
use scs8hd_fill_1  FILLER_11_24
timestamp 1586364061
transform 1 0 3312 0 1 8160
box -38 -48 130 592
use scs8hd_ebufn_2  mux_bottom_ipin_5.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 4416 0 1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_5.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 3864 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_5.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 4232 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_28
timestamp 1586364061
transform 1 0 3680 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_32
timestamp 1586364061
transform 1 0 4048 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_5.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 5428 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_5.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 6164 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_5.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 5796 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_45
timestamp 1586364061
transform 1 0 5244 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_49
timestamp 1586364061
transform 1 0 5612 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_53
timestamp 1586364061
transform 1 0 5980 0 1 8160
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_ipin_5.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 7452 0 1 8160
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_114
timestamp 1586364061
transform 1 0 6716 0 1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_5.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 7268 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_5.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 6532 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_57
timestamp 1586364061
transform 1 0 6348 0 1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_11_62
timestamp 1586364061
transform 1 0 6808 0 1 8160
box -38 -48 406 592
use scs8hd_fill_1  FILLER_11_66
timestamp 1586364061
transform 1 0 7176 0 1 8160
box -38 -48 130 592
use scs8hd_decap_6  FILLER_11_78
timestamp 1586364061
transform 1 0 8280 0 1 8160
box -38 -48 590 592
use scs8hd_inv_1  mux_bottom_ipin_5.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 9016 0 1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_5.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 9476 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__089__B
timestamp 1586364061
transform 1 0 8832 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_89
timestamp 1586364061
transform 1 0 9292 0 1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_11_93
timestamp 1586364061
transform 1 0 9660 0 1 8160
box -38 -48 406 592
use scs8hd_nor2_4  _090_
timestamp 1586364061
transform 1 0 10212 0 1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__090__B
timestamp 1586364061
transform 1 0 10028 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__089__A
timestamp 1586364061
transform 1 0 11224 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_108
timestamp 1586364061
transform 1 0 11040 0 1 8160
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_ipin_6.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12420 0 1 8160
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_115
timestamp 1586364061
transform 1 0 12328 0 1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_6.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 12144 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_6.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 11776 0 1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_11_112
timestamp 1586364061
transform 1 0 11408 0 1 8160
box -38 -48 406 592
use scs8hd_fill_2  FILLER_11_118
timestamp 1586364061
transform 1 0 11960 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_6.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 13616 0 1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_11_132
timestamp 1586364061
transform 1 0 13248 0 1 8160
box -38 -48 406 592
use scs8hd_fill_2  FILLER_11_138
timestamp 1586364061
transform 1 0 13800 0 1 8160
box -38 -48 222 592
use scs8hd_inv_1  mux_bottom_ipin_6.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 13984 0 1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_6.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 14444 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_7.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 15088 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_143
timestamp 1586364061
transform 1 0 14260 0 1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_11_147
timestamp 1586364061
transform 1 0 14628 0 1 8160
box -38 -48 406 592
use scs8hd_fill_1  FILLER_11_151
timestamp 1586364061
transform 1 0 14996 0 1 8160
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_7.LATCH_0_.latch
timestamp 1586364061
transform 1 0 15272 0 1 8160
box -38 -48 1050 592
use scs8hd_decap_3  FILLER_11_165
timestamp 1586364061
transform 1 0 16284 0 1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_7.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 16560 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_7.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 16928 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_170
timestamp 1586364061
transform 1 0 16744 0 1 8160
box -38 -48 222 592
use scs8hd_decap_6  FILLER_11_174
timestamp 1586364061
transform 1 0 17112 0 1 8160
box -38 -48 590 592
use scs8hd_inv_1  mux_bottom_ipin_7.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 18032 0 1 8160
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_116
timestamp 1586364061
transform 1 0 17940 0 1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_7.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 18492 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_7.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 18860 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__093__B
timestamp 1586364061
transform 1 0 17756 0 1 8160
box -38 -48 222 592
use scs8hd_fill_1  FILLER_11_180
timestamp 1586364061
transform 1 0 17664 0 1 8160
box -38 -48 130 592
use scs8hd_fill_2  FILLER_11_187
timestamp 1586364061
transform 1 0 18308 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_191
timestamp 1586364061
transform 1 0 18676 0 1 8160
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_7.LATCH_4_.latch
timestamp 1586364061
transform 1 0 19044 0 1 8160
box -38 -48 1050 592
use scs8hd_fill_2  FILLER_11_206
timestamp 1586364061
transform 1 0 20056 0 1 8160
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_ipin_7.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 20792 0 1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_7.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 20608 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_7.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 20240 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_210
timestamp 1586364061
transform 1 0 20424 0 1 8160
box -38 -48 222 592
use scs8hd_decap_3  PHY_23
timestamp 1586364061
transform -1 0 22816 0 1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_7.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 21804 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_7.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 22172 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_223
timestamp 1586364061
transform 1 0 21620 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_227
timestamp 1586364061
transform 1 0 21988 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_231
timestamp 1586364061
transform 1 0 22356 0 1 8160
box -38 -48 222 592
use scs8hd_inv_1  mux_top_ipin_2.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1380 0 -1 9248
box -38 -48 314 592
use scs8hd_decap_3  PHY_24
timestamp 1586364061
transform 1 0 1104 0 -1 9248
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_2.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 1840 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__077__B
timestamp 1586364061
transform 1 0 2208 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_6
timestamp 1586364061
transform 1 0 1656 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_10
timestamp 1586364061
transform 1 0 2024 0 -1 9248
box -38 -48 222 592
use scs8hd_nor2_4  _079_
timestamp 1586364061
transform 1 0 2392 0 -1 9248
box -38 -48 866 592
use scs8hd_decap_8  FILLER_12_23
timestamp 1586364061
transform 1 0 3220 0 -1 9248
box -38 -48 774 592
use scs8hd_ebufn_2  mux_bottom_ipin_5.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 4508 0 -1 9248
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_117
timestamp 1586364061
transform 1 0 3956 0 -1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_5.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 4324 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_3  FILLER_12_32
timestamp 1586364061
transform 1 0 4048 0 -1 9248
box -38 -48 314 592
use scs8hd_decap_12  FILLER_12_46
timestamp 1586364061
transform 1 0 5336 0 -1 9248
box -38 -48 1142 592
use scs8hd_ebufn_2  mux_bottom_ipin_5.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 6992 0 -1 9248
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_5.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 6716 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_3  FILLER_12_58
timestamp 1586364061
transform 1 0 6440 0 -1 9248
box -38 -48 314 592
use scs8hd_fill_1  FILLER_12_63
timestamp 1586364061
transform 1 0 6900 0 -1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_5.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 8004 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_73
timestamp 1586364061
transform 1 0 7820 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_12  FILLER_12_77
timestamp 1586364061
transform 1 0 8188 0 -1 9248
box -38 -48 1142 592
use scs8hd_nor2_4  _089_
timestamp 1586364061
transform 1 0 9660 0 -1 9248
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_118
timestamp 1586364061
transform 1 0 9568 0 -1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_6.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 9384 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_1  FILLER_12_89
timestamp 1586364061
transform 1 0 9292 0 -1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__090__A
timestamp 1586364061
transform 1 0 10672 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_102
timestamp 1586364061
transform 1 0 10488 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_8  FILLER_12_106
timestamp 1586364061
transform 1 0 10856 0 -1 9248
box -38 -48 774 592
use scs8hd_ebufn_2  mux_bottom_ipin_6.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12052 0 -1 9248
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_6.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11868 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_3  FILLER_12_114
timestamp 1586364061
transform 1 0 11592 0 -1 9248
box -38 -48 314 592
use scs8hd_inv_1  mux_bottom_ipin_6.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 13616 0 -1 9248
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_6.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 13064 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_128
timestamp 1586364061
transform 1 0 12880 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_12_132
timestamp 1586364061
transform 1 0 13248 0 -1 9248
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__097__A
timestamp 1586364061
transform 1 0 14444 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_6.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14076 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_139
timestamp 1586364061
transform 1 0 13892 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_143
timestamp 1586364061
transform 1 0 14260 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_6  FILLER_12_147
timestamp 1586364061
transform 1 0 14628 0 -1 9248
box -38 -48 590 592
use scs8hd_inv_1  mux_bottom_ipin_7.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 15548 0 -1 9248
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_119
timestamp 1586364061
transform 1 0 15180 0 -1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_7.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 16008 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_7.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 16376 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_3  FILLER_12_154
timestamp 1586364061
transform 1 0 15272 0 -1 9248
box -38 -48 314 592
use scs8hd_fill_2  FILLER_12_160
timestamp 1586364061
transform 1 0 15824 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_164
timestamp 1586364061
transform 1 0 16192 0 -1 9248
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_ipin_7.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 16560 0 -1 9248
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_7.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 17572 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_177
timestamp 1586364061
transform 1 0 17388 0 -1 9248
box -38 -48 222 592
use scs8hd_nor2_4  _093_
timestamp 1586364061
transform 1 0 18124 0 -1 9248
box -38 -48 866 592
use scs8hd_decap_4  FILLER_12_181
timestamp 1586364061
transform 1 0 17756 0 -1 9248
box -38 -48 406 592
use scs8hd_inv_1  mux_bottom_ipin_7.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 19780 0 -1 9248
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_7.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 19136 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_7.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 19504 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_194
timestamp 1586364061
transform 1 0 18952 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_198
timestamp 1586364061
transform 1 0 19320 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_1  FILLER_12_202
timestamp 1586364061
transform 1 0 19688 0 -1 9248
box -38 -48 130 592
use scs8hd_fill_2  FILLER_12_206
timestamp 1586364061
transform 1 0 20056 0 -1 9248
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_ipin_7.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 20884 0 -1 9248
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_120
timestamp 1586364061
transform 1 0 20792 0 -1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_7.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 20240 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_12_210
timestamp 1586364061
transform 1 0 20424 0 -1 9248
box -38 -48 406 592
use scs8hd_decap_3  PHY_25
timestamp 1586364061
transform -1 0 22816 0 -1 9248
box -38 -48 314 592
use scs8hd_decap_8  FILLER_12_224
timestamp 1586364061
transform 1 0 21712 0 -1 9248
box -38 -48 774 592
use scs8hd_fill_1  FILLER_12_232
timestamp 1586364061
transform 1 0 22448 0 -1 9248
box -38 -48 130 592
use scs8hd_nor2_4  _077_
timestamp 1586364061
transform 1 0 1564 0 1 9248
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_5.LATCH_5_.latch
timestamp 1586364061
transform 1 0 1472 0 -1 10336
box -38 -48 1050 592
use scs8hd_decap_3  PHY_26
timestamp 1586364061
transform 1 0 1104 0 1 9248
box -38 -48 314 592
use scs8hd_decap_3  PHY_28
timestamp 1586364061
transform 1 0 1104 0 -1 10336
box -38 -48 314 592
use scs8hd_fill_2  FILLER_13_3
timestamp 1586364061
transform 1 0 1380 0 1 9248
box -38 -48 222 592
use scs8hd_fill_1  FILLER_14_3
timestamp 1586364061
transform 1 0 1380 0 -1 10336
box -38 -48 130 592
use scs8hd_fill_2  FILLER_14_15
timestamp 1586364061
transform 1 0 2484 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_18
timestamp 1586364061
transform 1 0 2760 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_14
timestamp 1586364061
transform 1 0 2392 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_5.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 2668 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__077__A
timestamp 1586364061
transform 1 0 2944 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_5.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 2576 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_26
timestamp 1586364061
transform 1 0 3496 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_22
timestamp 1586364061
transform 1 0 3128 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_5.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 3312 0 1 9248
box -38 -48 222 592
use scs8hd_decap_12  FILLER_14_19
timestamp 1586364061
transform 1 0 2852 0 -1 10336
box -38 -48 1142 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_5.LATCH_4_.latch
timestamp 1586364061
transform 1 0 4048 0 -1 10336
box -38 -48 1050 592
use scs8hd_ebufn_2  mux_bottom_ipin_5.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 4324 0 1 9248
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_124
timestamp 1586364061
transform 1 0 3956 0 -1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_5.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 4048 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_5.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 3680 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_30
timestamp 1586364061
transform 1 0 3864 0 1 9248
box -38 -48 222 592
use scs8hd_fill_1  FILLER_13_34
timestamp 1586364061
transform 1 0 4232 0 1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_5.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 5244 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_5.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 5336 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_44
timestamp 1586364061
transform 1 0 5152 0 1 9248
box -38 -48 222 592
use scs8hd_decap_8  FILLER_13_48
timestamp 1586364061
transform 1 0 5520 0 1 9248
box -38 -48 774 592
use scs8hd_fill_2  FILLER_14_43
timestamp 1586364061
transform 1 0 5060 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_12  FILLER_14_47
timestamp 1586364061
transform 1 0 5428 0 -1 10336
box -38 -48 1142 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_5.LATCH_0_.latch
timestamp 1586364061
transform 1 0 6716 0 -1 10336
box -38 -48 1050 592
use scs8hd_ebufn_2  mux_bottom_ipin_5.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 7268 0 1 9248
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_121
timestamp 1586364061
transform 1 0 6716 0 1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_5.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 6992 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_5.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 6532 0 1 9248
box -38 -48 222 592
use scs8hd_decap_3  FILLER_13_56
timestamp 1586364061
transform 1 0 6256 0 1 9248
box -38 -48 314 592
use scs8hd_fill_2  FILLER_13_62
timestamp 1586364061
transform 1 0 6808 0 1 9248
box -38 -48 222 592
use scs8hd_fill_1  FILLER_13_66
timestamp 1586364061
transform 1 0 7176 0 1 9248
box -38 -48 130 592
use scs8hd_fill_2  FILLER_14_59
timestamp 1586364061
transform 1 0 6532 0 -1 10336
box -38 -48 222 592
use scs8hd_inv_1  mux_bottom_ipin_6.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 8556 0 -1 10336
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_6.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 8556 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_5.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 7912 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_13_76
timestamp 1586364061
transform 1 0 8096 0 1 9248
box -38 -48 406 592
use scs8hd_fill_1  FILLER_13_80
timestamp 1586364061
transform 1 0 8464 0 1 9248
box -38 -48 130 592
use scs8hd_fill_1  FILLER_13_83
timestamp 1586364061
transform 1 0 8740 0 1 9248
box -38 -48 130 592
use scs8hd_fill_2  FILLER_14_72
timestamp 1586364061
transform 1 0 7728 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_14_76
timestamp 1586364061
transform 1 0 8096 0 -1 10336
box -38 -48 406 592
use scs8hd_fill_1  FILLER_14_80
timestamp 1586364061
transform 1 0 8464 0 -1 10336
box -38 -48 130 592
use scs8hd_fill_1  FILLER_14_88
timestamp 1586364061
transform 1 0 9200 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_4  FILLER_14_84
timestamp 1586364061
transform 1 0 8832 0 -1 10336
box -38 -48 406 592
use scs8hd_fill_2  FILLER_13_87
timestamp 1586364061
transform 1 0 9108 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__088__A
timestamp 1586364061
transform 1 0 9292 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_5.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 9292 0 1 9248
box -38 -48 222 592
use scs8hd_inv_1  mux_bottom_ipin_5.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 8832 0 1 9248
box -38 -48 314 592
use scs8hd_fill_2  FILLER_14_93
timestamp 1586364061
transform 1 0 9660 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_1  FILLER_14_91
timestamp 1586364061
transform 1 0 9476 0 -1 10336
box -38 -48 130 592
use scs8hd_fill_2  FILLER_13_91
timestamp 1586364061
transform 1 0 9476 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_6.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 9844 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_6.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 9660 0 1 9248
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_125
timestamp 1586364061
transform 1 0 9568 0 -1 10336
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_6.LATCH_1_.latch
timestamp 1586364061
transform 1 0 9844 0 1 9248
box -38 -48 1050 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_6.LATCH_2_.latch
timestamp 1586364061
transform 1 0 10028 0 -1 10336
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_6.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 11040 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_106
timestamp 1586364061
transform 1 0 10856 0 1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_13_110
timestamp 1586364061
transform 1 0 11224 0 1 9248
box -38 -48 406 592
use scs8hd_decap_8  FILLER_14_108
timestamp 1586364061
transform 1 0 11040 0 -1 10336
box -38 -48 774 592
use scs8hd_ebufn_2  mux_bottom_ipin_6.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12420 0 1 9248
box -38 -48 866 592
use scs8hd_ebufn_2  mux_bottom_ipin_6.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12052 0 -1 10336
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_122
timestamp 1586364061
transform 1 0 12328 0 1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_6.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 12052 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_6.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 11684 0 1 9248
box -38 -48 222 592
use scs8hd_fill_1  FILLER_13_114
timestamp 1586364061
transform 1 0 11592 0 1 9248
box -38 -48 130 592
use scs8hd_fill_2  FILLER_13_117
timestamp 1586364061
transform 1 0 11868 0 1 9248
box -38 -48 222 592
use scs8hd_fill_1  FILLER_13_121
timestamp 1586364061
transform 1 0 12236 0 1 9248
box -38 -48 130 592
use scs8hd_decap_3  FILLER_14_116
timestamp 1586364061
transform 1 0 11776 0 -1 10336
box -38 -48 314 592
use scs8hd_ebufn_2  mux_bottom_ipin_6.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 13616 0 -1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__062__B
timestamp 1586364061
transform 1 0 13432 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_6.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 13616 0 1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_13_132
timestamp 1586364061
transform 1 0 13248 0 1 9248
box -38 -48 406 592
use scs8hd_decap_4  FILLER_13_138
timestamp 1586364061
transform 1 0 13800 0 1 9248
box -38 -48 406 592
use scs8hd_decap_6  FILLER_14_128
timestamp 1586364061
transform 1 0 12880 0 -1 10336
box -38 -48 590 592
use scs8hd_nor2_4  _097_
timestamp 1586364061
transform 1 0 14444 0 1 9248
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__097__B
timestamp 1586364061
transform 1 0 14260 0 1 9248
box -38 -48 222 592
use scs8hd_fill_1  FILLER_13_142
timestamp 1586364061
transform 1 0 14168 0 1 9248
box -38 -48 130 592
use scs8hd_decap_8  FILLER_14_145
timestamp 1586364061
transform 1 0 14444 0 -1 10336
box -38 -48 774 592
use scs8hd_fill_1  FILLER_14_154
timestamp 1586364061
transform 1 0 15272 0 -1 10336
box -38 -48 130 592
use scs8hd_fill_2  FILLER_13_158
timestamp 1586364061
transform 1 0 15640 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_154
timestamp 1586364061
transform 1 0 15272 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_7.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 15456 0 1 9248
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_126
timestamp 1586364061
transform 1 0 15180 0 -1 10336
box -38 -48 130 592
use scs8hd_fill_2  FILLER_13_162
timestamp 1586364061
transform 1 0 16008 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_7.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 15824 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_7.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 16192 0 1 9248
box -38 -48 222 592
use scs8hd_decap_8  FILLER_14_166
timestamp 1586364061
transform 1 0 16376 0 -1 10336
box -38 -48 774 592
use scs8hd_ebufn_2  mux_bottom_ipin_7.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 16376 0 1 9248
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_7.LATCH_2_.latch
timestamp 1586364061
transform 1 0 15364 0 -1 10336
box -38 -48 1050 592
use scs8hd_ebufn_2  mux_bottom_ipin_7.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 17112 0 -1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_7.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 17388 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_175
timestamp 1586364061
transform 1 0 17204 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_179
timestamp 1586364061
transform 1 0 17572 0 1 9248
box -38 -48 222 592
use scs8hd_nor2_4  _096_
timestamp 1586364061
transform 1 0 18032 0 1 9248
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_7.LATCH_1_.latch
timestamp 1586364061
transform 1 0 18676 0 -1 10336
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_123
timestamp 1586364061
transform 1 0 17940 0 1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__096__B
timestamp 1586364061
transform 1 0 17756 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__096__A
timestamp 1586364061
transform 1 0 18124 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_193
timestamp 1586364061
transform 1 0 18860 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_183
timestamp 1586364061
transform 1 0 17940 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_14_187
timestamp 1586364061
transform 1 0 18308 0 -1 10336
box -38 -48 406 592
use scs8hd_ebufn_2  mux_bottom_ipin_7.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 19596 0 1 9248
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_7.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 19044 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_7.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 19412 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_7.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 19872 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_197
timestamp 1586364061
transform 1 0 19228 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_202
timestamp 1586364061
transform 1 0 19688 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_8  FILLER_14_206
timestamp 1586364061
transform 1 0 20056 0 -1 10336
box -38 -48 774 592
use scs8hd_buf_2  _148_
timestamp 1586364061
transform 1 0 21160 0 1 9248
box -38 -48 406 592
use scs8hd_inv_1  mux_bottom_ipin_7.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 20884 0 -1 10336
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_127
timestamp 1586364061
transform 1 0 20792 0 -1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_7.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 20884 0 1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_13_210
timestamp 1586364061
transform 1 0 20424 0 1 9248
box -38 -48 406 592
use scs8hd_fill_1  FILLER_13_214
timestamp 1586364061
transform 1 0 20792 0 1 9248
box -38 -48 130 592
use scs8hd_fill_1  FILLER_13_217
timestamp 1586364061
transform 1 0 21068 0 1 9248
box -38 -48 130 592
use scs8hd_decap_12  FILLER_14_218
timestamp 1586364061
transform 1 0 21160 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_3  PHY_27
timestamp 1586364061
transform -1 0 22816 0 1 9248
box -38 -48 314 592
use scs8hd_decap_3  PHY_29
timestamp 1586364061
transform -1 0 22816 0 -1 10336
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__148__A
timestamp 1586364061
transform 1 0 21712 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_222
timestamp 1586364061
transform 1 0 21528 0 1 9248
box -38 -48 222 592
use scs8hd_decap_6  FILLER_13_226
timestamp 1586364061
transform 1 0 21896 0 1 9248
box -38 -48 590 592
use scs8hd_fill_1  FILLER_13_232
timestamp 1586364061
transform 1 0 22448 0 1 9248
box -38 -48 130 592
use scs8hd_decap_3  FILLER_14_230
timestamp 1586364061
transform 1 0 22264 0 -1 10336
box -38 -48 314 592
use scs8hd_ebufn_2  mux_bottom_ipin_5.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 1656 0 1 10336
box -38 -48 866 592
use scs8hd_decap_3  PHY_30
timestamp 1586364061
transform 1 0 1104 0 1 10336
box -38 -48 314 592
use scs8hd_decap_3  FILLER_15_3
timestamp 1586364061
transform 1 0 1380 0 1 10336
box -38 -48 314 592
use scs8hd_inv_1  mux_bottom_ipin_5.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 3220 0 1 10336
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__078__B
timestamp 1586364061
transform 1 0 2668 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__078__A
timestamp 1586364061
transform 1 0 3036 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_15
timestamp 1586364061
transform 1 0 2484 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_19
timestamp 1586364061
transform 1 0 2852 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_26
timestamp 1586364061
transform 1 0 3496 0 1 10336
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_5.LATCH_3_.latch
timestamp 1586364061
transform 1 0 4232 0 1 10336
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_5.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 4048 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_5.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 3680 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_30
timestamp 1586364061
transform 1 0 3864 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__082__A
timestamp 1586364061
transform 1 0 5980 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_5.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 5428 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_45
timestamp 1586364061
transform 1 0 5244 0 1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_15_49
timestamp 1586364061
transform 1 0 5612 0 1 10336
box -38 -48 406 592
use scs8hd_fill_2  FILLER_15_55
timestamp 1586364061
transform 1 0 6164 0 1 10336
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_ipin_5.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 7084 0 1 10336
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_128
timestamp 1586364061
transform 1 0 6716 0 1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__082__B
timestamp 1586364061
transform 1 0 6348 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_59
timestamp 1586364061
transform 1 0 6532 0 1 10336
box -38 -48 222 592
use scs8hd_decap_3  FILLER_15_62
timestamp 1586364061
transform 1 0 6808 0 1 10336
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_5.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 8096 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_74
timestamp 1586364061
transform 1 0 7912 0 1 10336
box -38 -48 222 592
use scs8hd_decap_8  FILLER_15_78
timestamp 1586364061
transform 1 0 8280 0 1 10336
box -38 -48 774 592
use scs8hd_nor2_4  _088_
timestamp 1586364061
transform 1 0 9292 0 1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__088__B
timestamp 1586364061
transform 1 0 9108 0 1 10336
box -38 -48 222 592
use scs8hd_fill_1  FILLER_15_86
timestamp 1586364061
transform 1 0 9016 0 1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_6.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 11132 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_6.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 10764 0 1 10336
box -38 -48 222 592
use scs8hd_decap_6  FILLER_15_98
timestamp 1586364061
transform 1 0 10120 0 1 10336
box -38 -48 590 592
use scs8hd_fill_1  FILLER_15_104
timestamp 1586364061
transform 1 0 10672 0 1 10336
box -38 -48 130 592
use scs8hd_fill_2  FILLER_15_107
timestamp 1586364061
transform 1 0 10948 0 1 10336
box -38 -48 222 592
use scs8hd_inv_1  mux_bottom_ipin_6.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 11316 0 1 10336
box -38 -48 314 592
use scs8hd_ebufn_2  mux_bottom_ipin_6.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12420 0 1 10336
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_129
timestamp 1586364061
transform 1 0 12328 0 1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_6.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 11776 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_6.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 12144 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_114
timestamp 1586364061
transform 1 0 11592 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_118
timestamp 1586364061
transform 1 0 11960 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__062__A
timestamp 1586364061
transform 1 0 13616 0 1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_15_132
timestamp 1586364061
transform 1 0 13248 0 1 10336
box -38 -48 406 592
use scs8hd_fill_2  FILLER_15_138
timestamp 1586364061
transform 1 0 13800 0 1 10336
box -38 -48 222 592
use scs8hd_nor2_4  _095_
timestamp 1586364061
transform 1 0 14536 0 1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__095__B
timestamp 1586364061
transform 1 0 14352 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__095__A
timestamp 1586364061
transform 1 0 13984 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_142
timestamp 1586364061
transform 1 0 14168 0 1 10336
box -38 -48 222 592
use scs8hd_inv_1  mux_bottom_ipin_7.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 16284 0 1 10336
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_6.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 15548 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_155
timestamp 1586364061
transform 1 0 15364 0 1 10336
box -38 -48 222 592
use scs8hd_decap_6  FILLER_15_159
timestamp 1586364061
transform 1 0 15732 0 1 10336
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_7.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 16744 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_7.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 17112 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_168
timestamp 1586364061
transform 1 0 16560 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_172
timestamp 1586364061
transform 1 0 16928 0 1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_15_176
timestamp 1586364061
transform 1 0 17296 0 1 10336
box -38 -48 406 592
use scs8hd_inv_1  mux_bottom_ipin_3.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 18032 0 1 10336
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_130
timestamp 1586364061
transform 1 0 17940 0 1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_3.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 18492 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__064__A
timestamp 1586364061
transform 1 0 17664 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__064__B
timestamp 1586364061
transform 1 0 18860 0 1 10336
box -38 -48 222 592
use scs8hd_fill_1  FILLER_15_182
timestamp 1586364061
transform 1 0 17848 0 1 10336
box -38 -48 130 592
use scs8hd_fill_2  FILLER_15_187
timestamp 1586364061
transform 1 0 18308 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_191
timestamp 1586364061
transform 1 0 18676 0 1 10336
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_ipin_7.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 19504 0 1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_7.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 19320 0 1 10336
box -38 -48 222 592
use scs8hd_decap_3  FILLER_15_195
timestamp 1586364061
transform 1 0 19044 0 1 10336
box -38 -48 314 592
use scs8hd_buf_2  _143_
timestamp 1586364061
transform 1 0 21068 0 1 10336
box -38 -48 406 592
use scs8hd_decap_8  FILLER_15_209
timestamp 1586364061
transform 1 0 20332 0 1 10336
box -38 -48 774 592
use scs8hd_fill_2  FILLER_15_221
timestamp 1586364061
transform 1 0 21436 0 1 10336
box -38 -48 222 592
use scs8hd_decap_3  PHY_31
timestamp 1586364061
transform -1 0 22816 0 1 10336
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__143__A
timestamp 1586364061
transform 1 0 21620 0 1 10336
box -38 -48 222 592
use scs8hd_decap_8  FILLER_15_225
timestamp 1586364061
transform 1 0 21804 0 1 10336
box -38 -48 774 592
use scs8hd_conb_1  _136_
timestamp 1586364061
transform 1 0 1380 0 -1 11424
box -38 -48 314 592
use scs8hd_decap_3  PHY_32
timestamp 1586364061
transform 1 0 1104 0 -1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__115__A
timestamp 1586364061
transform 1 0 2208 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_5.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 1840 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_6
timestamp 1586364061
transform 1 0 1656 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_10
timestamp 1586364061
transform 1 0 2024 0 -1 11424
box -38 -48 222 592
use scs8hd_nor2_4  _078_
timestamp 1586364061
transform 1 0 2392 0 -1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_0.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 3404 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_23
timestamp 1586364061
transform 1 0 3220 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_16_27
timestamp 1586364061
transform 1 0 3588 0 -1 11424
box -38 -48 406 592
use scs8hd_ebufn_2  mux_bottom_ipin_5.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 4784 0 -1 11424
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_131
timestamp 1586364061
transform 1 0 3956 0 -1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_5.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 4232 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 4600 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_32
timestamp 1586364061
transform 1 0 4048 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_36
timestamp 1586364061
transform 1 0 4416 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 6164 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_6  FILLER_16_49
timestamp 1586364061
transform 1 0 5612 0 -1 11424
box -38 -48 590 592
use scs8hd_nor2_4  _082_
timestamp 1586364061
transform 1 0 6348 0 -1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 7360 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_66
timestamp 1586364061
transform 1 0 7176 0 -1 11424
box -38 -48 222 592
use scs8hd_inv_1  mux_bottom_ipin_5.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 7912 0 -1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_6.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 8648 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_5.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 7728 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_70
timestamp 1586364061
transform 1 0 7544 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_16_77
timestamp 1586364061
transform 1 0 8188 0 -1 11424
box -38 -48 406 592
use scs8hd_fill_1  FILLER_16_81
timestamp 1586364061
transform 1 0 8556 0 -1 11424
box -38 -48 130 592
use scs8hd_conb_1  _137_
timestamp 1586364061
transform 1 0 9660 0 -1 11424
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_132
timestamp 1586364061
transform 1 0 9568 0 -1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_6.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 9384 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_6  FILLER_16_84
timestamp 1586364061
transform 1 0 8832 0 -1 11424
box -38 -48 590 592
use scs8hd_decap_4  FILLER_16_96
timestamp 1586364061
transform 1 0 9936 0 -1 11424
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_6.LATCH_3_.latch
timestamp 1586364061
transform 1 0 11224 0 -1 11424
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA__087__A
timestamp 1586364061
transform 1 0 10396 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_1  FILLER_16_100
timestamp 1586364061
transform 1 0 10304 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_6  FILLER_16_103
timestamp 1586364061
transform 1 0 10580 0 -1 11424
box -38 -48 590 592
use scs8hd_fill_1  FILLER_16_109
timestamp 1586364061
transform 1 0 11132 0 -1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_6.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 12420 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_121
timestamp 1586364061
transform 1 0 12236 0 -1 11424
box -38 -48 222 592
use scs8hd_nor2_4  _062_
timestamp 1586364061
transform 1 0 13616 0 -1 11424
box -38 -48 866 592
use scs8hd_decap_8  FILLER_16_125
timestamp 1586364061
transform 1 0 12604 0 -1 11424
box -38 -48 774 592
use scs8hd_decap_3  FILLER_16_133
timestamp 1586364061
transform 1 0 13340 0 -1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_3.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 14812 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_16_145
timestamp 1586364061
transform 1 0 14444 0 -1 11424
box -38 -48 406 592
use scs8hd_fill_2  FILLER_16_151
timestamp 1586364061
transform 1 0 14996 0 -1 11424
box -38 -48 222 592
use scs8hd_inv_1  mux_bottom_ipin_6.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 15272 0 -1 11424
box -38 -48 314 592
use scs8hd_inv_1  mux_bottom_ipin_7.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 16284 0 -1 11424
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_133
timestamp 1586364061
transform 1 0 15180 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_8  FILLER_16_157
timestamp 1586364061
transform 1 0 15548 0 -1 11424
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_3.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 17480 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_8  FILLER_16_168
timestamp 1586364061
transform 1 0 16560 0 -1 11424
box -38 -48 774 592
use scs8hd_fill_2  FILLER_16_176
timestamp 1586364061
transform 1 0 17296 0 -1 11424
box -38 -48 222 592
use scs8hd_nor2_4  _064_
timestamp 1586364061
transform 1 0 17664 0 -1 11424
box -38 -48 866 592
use scs8hd_decap_8  FILLER_16_189
timestamp 1586364061
transform 1 0 18492 0 -1 11424
box -38 -48 774 592
use scs8hd_inv_1  mux_bottom_ipin_7.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 19320 0 -1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_7.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 19780 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_1  FILLER_16_197
timestamp 1586364061
transform 1 0 19228 0 -1 11424
box -38 -48 130 592
use scs8hd_fill_2  FILLER_16_201
timestamp 1586364061
transform 1 0 19596 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_8  FILLER_16_205
timestamp 1586364061
transform 1 0 19964 0 -1 11424
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_134
timestamp 1586364061
transform 1 0 20792 0 -1 11424
box -38 -48 130 592
use scs8hd_fill_1  FILLER_16_213
timestamp 1586364061
transform 1 0 20700 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_12  FILLER_16_215
timestamp 1586364061
transform 1 0 20884 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_3  PHY_33
timestamp 1586364061
transform -1 0 22816 0 -1 11424
box -38 -48 314 592
use scs8hd_decap_6  FILLER_16_227
timestamp 1586364061
transform 1 0 21988 0 -1 11424
box -38 -48 590 592
use scs8hd_buf_2  _146_
timestamp 1586364061
transform 1 0 1380 0 1 11424
box -38 -48 406 592
use scs8hd_decap_3  PHY_34
timestamp 1586364061
transform 1 0 1104 0 1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__146__A
timestamp 1586364061
transform 1 0 1932 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_7
timestamp 1586364061
transform 1 0 1748 0 1 11424
box -38 -48 222 592
use scs8hd_decap_3  FILLER_17_11
timestamp 1586364061
transform 1 0 2116 0 1 11424
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_0.LATCH_1_.latch
timestamp 1586364061
transform 1 0 3128 0 1 11424
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_0.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 2944 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__115__B
timestamp 1586364061
transform 1 0 2392 0 1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_17_16
timestamp 1586364061
transform 1 0 2576 0 1 11424
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 4324 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_33
timestamp 1586364061
transform 1 0 4140 0 1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_17_37
timestamp 1586364061
transform 1 0 4508 0 1 11424
box -38 -48 406 592
use scs8hd_fill_1  FILLER_17_41
timestamp 1586364061
transform 1 0 4876 0 1 11424
box -38 -48 130 592
use scs8hd_nor2_4  _116_
timestamp 1586364061
transform 1 0 5152 0 1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 6164 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__116__B
timestamp 1586364061
transform 1 0 4968 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_53
timestamp 1586364061
transform 1 0 5980 0 1 11424
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_0.LATCH_0_.latch
timestamp 1586364061
transform 1 0 6808 0 1 11424
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_135
timestamp 1586364061
transform 1 0 6716 0 1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_0.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 6532 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_57
timestamp 1586364061
transform 1 0 6348 0 1 11424
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_6.LATCH_5_.latch
timestamp 1586364061
transform 1 0 8648 0 1 11424
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 8280 0 1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_17_73
timestamp 1586364061
transform 1 0 7820 0 1 11424
box -38 -48 406 592
use scs8hd_fill_1  FILLER_17_77
timestamp 1586364061
transform 1 0 8188 0 1 11424
box -38 -48 130 592
use scs8hd_fill_2  FILLER_17_80
timestamp 1586364061
transform 1 0 8464 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_6.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9844 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_93
timestamp 1586364061
transform 1 0 9660 0 1 11424
box -38 -48 222 592
use scs8hd_nor2_4  _087_
timestamp 1586364061
transform 1 0 10396 0 1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__087__B
timestamp 1586364061
transform 1 0 10212 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_97
timestamp 1586364061
transform 1 0 10028 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_110
timestamp 1586364061
transform 1 0 11224 0 1 11424
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_ipin_6.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12420 0 1 11424
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_136
timestamp 1586364061
transform 1 0 12328 0 1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_6.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 11408 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_6.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 12144 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_6.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 11776 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_114
timestamp 1586364061
transform 1 0 11592 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_118
timestamp 1586364061
transform 1 0 11960 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_6.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 13432 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_6.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 13800 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_132
timestamp 1586364061
transform 1 0 13248 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_136
timestamp 1586364061
transform 1 0 13616 0 1 11424
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_3.LATCH_2_.latch
timestamp 1586364061
transform 1 0 14812 0 1 11424
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_3.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 14628 0 1 11424
box -38 -48 222 592
use scs8hd_decap_6  FILLER_17_140
timestamp 1586364061
transform 1 0 13984 0 1 11424
box -38 -48 590 592
use scs8hd_fill_1  FILLER_17_146
timestamp 1586364061
transform 1 0 14536 0 1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_3.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 16008 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_3.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 16376 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_160
timestamp 1586364061
transform 1 0 15824 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_164
timestamp 1586364061
transform 1 0 16192 0 1 11424
box -38 -48 222 592
use scs8hd_inv_1  mux_bottom_ipin_3.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 16560 0 1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_3.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 17020 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_3.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 17572 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_171
timestamp 1586364061
transform 1 0 16836 0 1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_17_175
timestamp 1586364061
transform 1 0 17204 0 1 11424
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_3.LATCH_1_.latch
timestamp 1586364061
transform 1 0 18492 0 1 11424
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_137
timestamp 1586364061
transform 1 0 17940 0 1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_3.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 18308 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_181
timestamp 1586364061
transform 1 0 17756 0 1 11424
box -38 -48 222 592
use scs8hd_decap_3  FILLER_17_184
timestamp 1586364061
transform 1 0 18032 0 1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_3.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 19688 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_3.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 20056 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_200
timestamp 1586364061
transform 1 0 19504 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_204
timestamp 1586364061
transform 1 0 19872 0 1 11424
box -38 -48 222 592
use scs8hd_inv_1  mux_bottom_ipin_3.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 20240 0 1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_3.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 20700 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_3.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 21068 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_211
timestamp 1586364061
transform 1 0 20516 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_215
timestamp 1586364061
transform 1 0 20884 0 1 11424
box -38 -48 222 592
use scs8hd_decap_12  FILLER_17_219
timestamp 1586364061
transform 1 0 21252 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_3  PHY_35
timestamp 1586364061
transform -1 0 22816 0 1 11424
box -38 -48 314 592
use scs8hd_fill_2  FILLER_17_231
timestamp 1586364061
transform 1 0 22356 0 1 11424
box -38 -48 222 592
use scs8hd_conb_1  _131_
timestamp 1586364061
transform 1 0 1380 0 -1 12512
box -38 -48 314 592
use scs8hd_decap_3  PHY_36
timestamp 1586364061
transform 1 0 1104 0 -1 12512
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_0.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 1840 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__111__A
timestamp 1586364061
transform 1 0 2208 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_6
timestamp 1586364061
transform 1 0 1656 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_10
timestamp 1586364061
transform 1 0 2024 0 -1 12512
box -38 -48 222 592
use scs8hd_nor2_4  _115_
timestamp 1586364061
transform 1 0 2392 0 -1 12512
box -38 -48 866 592
use scs8hd_decap_6  FILLER_18_23
timestamp 1586364061
transform 1 0 3220 0 -1 12512
box -38 -48 590 592
use scs8hd_ebufn_2  mux_bottom_ipin_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 4048 0 -1 12512
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_138
timestamp 1586364061
transform 1 0 3956 0 -1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 3772 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_3  FILLER_18_41
timestamp 1586364061
transform 1 0 4876 0 -1 12512
box -38 -48 314 592
use scs8hd_inv_1  mux_bottom_ipin_0.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 5704 0 -1 12512
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__116__A
timestamp 1586364061
transform 1 0 5152 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 6164 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_18_46
timestamp 1586364061
transform 1 0 5336 0 -1 12512
box -38 -48 406 592
use scs8hd_fill_2  FILLER_18_53
timestamp 1586364061
transform 1 0 5980 0 -1 12512
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_ipin_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 6716 0 -1 12512
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_0.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 6532 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_57
timestamp 1586364061
transform 1 0 6348 0 -1 12512
box -38 -48 222 592
use scs8hd_inv_1  mux_bottom_ipin_0.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 8280 0 -1 12512
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 7728 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_6.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 8740 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_70
timestamp 1586364061
transform 1 0 7544 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_18_74
timestamp 1586364061
transform 1 0 7912 0 -1 12512
box -38 -48 406 592
use scs8hd_fill_2  FILLER_18_81
timestamp 1586364061
transform 1 0 8556 0 -1 12512
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_ipin_6.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9660 0 -1 12512
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_139
timestamp 1586364061
transform 1 0 9568 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_6  FILLER_18_85
timestamp 1586364061
transform 1 0 8924 0 -1 12512
box -38 -48 590 592
use scs8hd_fill_1  FILLER_18_91
timestamp 1586364061
transform 1 0 9476 0 -1 12512
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_6.LATCH_4_.latch
timestamp 1586364061
transform 1 0 11224 0 -1 12512
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA__086__A
timestamp 1586364061
transform 1 0 10672 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_102
timestamp 1586364061
transform 1 0 10488 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_18_106
timestamp 1586364061
transform 1 0 10856 0 -1 12512
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_6.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 12420 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_121
timestamp 1586364061
transform 1 0 12236 0 -1 12512
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_ipin_6.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12972 0 -1 12512
box -38 -48 866 592
use scs8hd_decap_4  FILLER_18_125
timestamp 1586364061
transform 1 0 12604 0 -1 12512
box -38 -48 406 592
use scs8hd_decap_4  FILLER_18_138
timestamp 1586364061
transform 1 0 13800 0 -1 12512
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_3.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 14260 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_1  FILLER_18_142
timestamp 1586364061
transform 1 0 14168 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_8  FILLER_18_145
timestamp 1586364061
transform 1 0 14444 0 -1 12512
box -38 -48 774 592
use scs8hd_ebufn_2  mux_bottom_ipin_3.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 16008 0 -1 12512
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_140
timestamp 1586364061
transform 1 0 15180 0 -1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_3.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 15824 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_6  FILLER_18_154
timestamp 1586364061
transform 1 0 15272 0 -1 12512
box -38 -48 590 592
use scs8hd_ebufn_2  mux_bottom_ipin_3.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 17572 0 -1 12512
box -38 -48 866 592
use scs8hd_decap_8  FILLER_18_171
timestamp 1586364061
transform 1 0 16836 0 -1 12512
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_3.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 18584 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_188
timestamp 1586364061
transform 1 0 18400 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_3  FILLER_18_192
timestamp 1586364061
transform 1 0 18768 0 -1 12512
box -38 -48 314 592
use scs8hd_ebufn_2  mux_bottom_ipin_3.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 19228 0 -1 12512
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_3.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 19044 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_206
timestamp 1586364061
transform 1 0 20056 0 -1 12512
box -38 -48 222 592
use scs8hd_inv_1  mux_bottom_ipin_3.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 20884 0 -1 12512
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_141
timestamp 1586364061
transform 1 0 20792 0 -1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_3.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 20240 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 21344 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_18_210
timestamp 1586364061
transform 1 0 20424 0 -1 12512
box -38 -48 406 592
use scs8hd_fill_2  FILLER_18_218
timestamp 1586364061
transform 1 0 21160 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_3  PHY_37
timestamp 1586364061
transform -1 0 22816 0 -1 12512
box -38 -48 314 592
use scs8hd_decap_8  FILLER_18_222
timestamp 1586364061
transform 1 0 21528 0 -1 12512
box -38 -48 774 592
use scs8hd_decap_3  FILLER_18_230
timestamp 1586364061
transform 1 0 22264 0 -1 12512
box -38 -48 314 592
use scs8hd_nor2_4  _111_
timestamp 1586364061
transform 1 0 1380 0 1 12512
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_0.LATCH_5_.latch
timestamp 1586364061
transform 1 0 1380 0 -1 13600
box -38 -48 1050 592
use scs8hd_decap_3  PHY_38
timestamp 1586364061
transform 1 0 1104 0 1 12512
box -38 -48 314 592
use scs8hd_decap_3  PHY_40
timestamp 1586364061
transform 1 0 1104 0 -1 13600
box -38 -48 314 592
use scs8hd_fill_2  FILLER_19_12
timestamp 1586364061
transform 1 0 2208 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_14
timestamp 1586364061
transform 1 0 2392 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_1  FILLER_19_20
timestamp 1586364061
transform 1 0 2944 0 1 12512
box -38 -48 130 592
use scs8hd_fill_2  FILLER_19_16
timestamp 1586364061
transform 1 0 2576 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_0.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 2760 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 2576 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__111__B
timestamp 1586364061
transform 1 0 2392 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_26
timestamp 1586364061
transform 1 0 3496 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_24
timestamp 1586364061
transform 1 0 3312 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 3496 0 1 12512
box -38 -48 222 592
use scs8hd_inv_1  mux_bottom_ipin_0.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 3036 0 1 12512
box -38 -48 314 592
use scs8hd_decap_8  FILLER_20_18
timestamp 1586364061
transform 1 0 2760 0 -1 13600
box -38 -48 774 592
use scs8hd_ebufn_2  mux_bottom_ipin_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 4048 0 1 12512
box -38 -48 866 592
use scs8hd_ebufn_2  mux_bottom_ipin_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 4324 0 -1 13600
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_145
timestamp 1586364061
transform 1 0 3956 0 -1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 3864 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 3680 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_28
timestamp 1586364061
transform 1 0 3680 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_41
timestamp 1586364061
transform 1 0 4876 0 1 12512
box -38 -48 222 592
use scs8hd_fill_1  FILLER_20_30
timestamp 1586364061
transform 1 0 3864 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_3  FILLER_20_32
timestamp 1586364061
transform 1 0 4048 0 -1 13600
box -38 -48 314 592
use scs8hd_inv_1  mux_bottom_ipin_0.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 5612 0 1 12512
box -38 -48 314 592
use scs8hd_inv_1  mux_bottom_ipin_0.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 5888 0 -1 13600
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 6072 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 5060 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 5428 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_45
timestamp 1586364061
transform 1 0 5244 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_52
timestamp 1586364061
transform 1 0 5888 0 1 12512
box -38 -48 222 592
use scs8hd_decap_8  FILLER_20_44
timestamp 1586364061
transform 1 0 5152 0 -1 13600
box -38 -48 774 592
use scs8hd_fill_2  FILLER_20_55
timestamp 1586364061
transform 1 0 6164 0 -1 13600
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_ipin_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 6808 0 1 12512
box -38 -48 866 592
use scs8hd_ebufn_2  mux_bottom_ipin_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 6900 0 -1 13600
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_142
timestamp 1586364061
transform 1 0 6716 0 1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 6440 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_0.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 6716 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 6348 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_56
timestamp 1586364061
transform 1 0 6256 0 1 12512
box -38 -48 222 592
use scs8hd_fill_1  FILLER_19_60
timestamp 1586364061
transform 1 0 6624 0 1 12512
box -38 -48 130 592
use scs8hd_fill_2  FILLER_20_59
timestamp 1586364061
transform 1 0 6532 0 -1 13600
box -38 -48 222 592
use scs8hd_nor2_4  _085_
timestamp 1586364061
transform 1 0 8556 0 1 12512
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__085__B
timestamp 1586364061
transform 1 0 8372 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__085__A
timestamp 1586364061
transform 1 0 8556 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 7820 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_71
timestamp 1586364061
transform 1 0 7636 0 1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_19_75
timestamp 1586364061
transform 1 0 8004 0 1 12512
box -38 -48 406 592
use scs8hd_decap_8  FILLER_20_72
timestamp 1586364061
transform 1 0 7728 0 -1 13600
box -38 -48 774 592
use scs8hd_fill_1  FILLER_20_80
timestamp 1586364061
transform 1 0 8464 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_8  FILLER_20_83
timestamp 1586364061
transform 1 0 8740 0 -1 13600
box -38 -48 774 592
use scs8hd_nor2_4  _105_
timestamp 1586364061
transform 1 0 9660 0 -1 13600
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_146
timestamp 1586364061
transform 1 0 9568 0 -1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__105__B
timestamp 1586364061
transform 1 0 9660 0 1 12512
box -38 -48 222 592
use scs8hd_decap_3  FILLER_19_90
timestamp 1586364061
transform 1 0 9384 0 1 12512
box -38 -48 314 592
use scs8hd_decap_3  FILLER_19_95
timestamp 1586364061
transform 1 0 9844 0 1 12512
box -38 -48 314 592
use scs8hd_fill_1  FILLER_20_91
timestamp 1586364061
transform 1 0 9476 0 -1 13600
box -38 -48 130 592
use scs8hd_nor2_4  _086_
timestamp 1586364061
transform 1 0 10304 0 1 12512
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__086__B
timestamp 1586364061
transform 1 0 10120 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_0.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 10672 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_109
timestamp 1586364061
transform 1 0 11132 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_102
timestamp 1586364061
transform 1 0 10488 0 -1 13600
box -38 -48 222 592
use scs8hd_decap_8  FILLER_20_106
timestamp 1586364061
transform 1 0 10856 0 -1 13600
box -38 -48 774 592
use scs8hd_decap_3  FILLER_20_114
timestamp 1586364061
transform 1 0 11592 0 -1 13600
box -38 -48 314 592
use scs8hd_decap_4  FILLER_19_113
timestamp 1586364061
transform 1 0 11500 0 1 12512
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__105__A
timestamp 1586364061
transform 1 0 11316 0 1 12512
box -38 -48 222 592
use scs8hd_decap_3  FILLER_20_120
timestamp 1586364061
transform 1 0 12144 0 -1 13600
box -38 -48 314 592
use scs8hd_decap_3  FILLER_19_119
timestamp 1586364061
transform 1 0 12052 0 1 12512
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 11868 0 1 12512
box -38 -48 222 592
use scs8hd_inv_1  mux_top_ipin_0.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 11868 0 -1 13600
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 12420 0 -1 13600
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_143
timestamp 1586364061
transform 1 0 12328 0 1 12512
box -38 -48 130 592
use scs8hd_inv_1  mux_top_ipin_0.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 12420 0 1 12512
box -38 -48 314 592
use scs8hd_decap_6  FILLER_20_129
timestamp 1586364061
transform 1 0 12972 0 -1 13600
box -38 -48 590 592
use scs8hd_fill_2  FILLER_20_125
timestamp 1586364061
transform 1 0 12604 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_130
timestamp 1586364061
transform 1 0 13064 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_126
timestamp 1586364061
transform 1 0 12696 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 12788 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 12880 0 1 12512
box -38 -48 222 592
use scs8hd_fill_1  FILLER_20_135
timestamp 1586364061
transform 1 0 13524 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_3  FILLER_19_138
timestamp 1586364061
transform 1 0 13800 0 1 12512
box -38 -48 314 592
use scs8hd_fill_2  FILLER_19_134
timestamp 1586364061
transform 1 0 13432 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__066__B
timestamp 1586364061
transform 1 0 13248 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__066__A
timestamp 1586364061
transform 1 0 13616 0 1 12512
box -38 -48 222 592
use scs8hd_nor2_4  _066_
timestamp 1586364061
transform 1 0 13616 0 -1 13600
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_3.LATCH_0_.latch
timestamp 1586364061
transform 1 0 14260 0 1 12512
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_3.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 14076 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__130__A
timestamp 1586364061
transform 1 0 14720 0 -1 13600
box -38 -48 222 592
use scs8hd_decap_3  FILLER_20_145
timestamp 1586364061
transform 1 0 14444 0 -1 13600
box -38 -48 314 592
use scs8hd_decap_3  FILLER_20_150
timestamp 1586364061
transform 1 0 14904 0 -1 13600
box -38 -48 314 592
use scs8hd_ebufn_2  mux_bottom_ipin_3.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15824 0 -1 13600
box -38 -48 866 592
use scs8hd_ebufn_2  mux_bottom_ipin_3.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 16008 0 1 12512
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_147
timestamp 1586364061
transform 1 0 15180 0 -1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_3.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 15824 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_3.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 15456 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_154
timestamp 1586364061
transform 1 0 15272 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_158
timestamp 1586364061
transform 1 0 15640 0 1 12512
box -38 -48 222 592
use scs8hd_decap_6  FILLER_20_154
timestamp 1586364061
transform 1 0 15272 0 -1 13600
box -38 -48 590 592
use scs8hd_fill_2  FILLER_20_169
timestamp 1586364061
transform 1 0 16652 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_171
timestamp 1586364061
transform 1 0 16836 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_3.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 16836 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_1  FILLER_20_177
timestamp 1586364061
transform 1 0 17388 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_4  FILLER_20_173
timestamp 1586364061
transform 1 0 17020 0 -1 13600
box -38 -48 406 592
use scs8hd_fill_2  FILLER_19_179
timestamp 1586364061
transform 1 0 17572 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_175
timestamp 1586364061
transform 1 0 17204 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__058__B
timestamp 1586364061
transform 1 0 17020 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__058__A
timestamp 1586364061
transform 1 0 17388 0 1 12512
box -38 -48 222 592
use scs8hd_nor2_4  _058_
timestamp 1586364061
transform 1 0 17480 0 -1 13600
box -38 -48 866 592
use scs8hd_nor2_4  _060_
timestamp 1586364061
transform 1 0 18032 0 1 12512
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_144
timestamp 1586364061
transform 1 0 17940 0 1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__060__A
timestamp 1586364061
transform 1 0 17756 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__060__B
timestamp 1586364061
transform 1 0 18492 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_193
timestamp 1586364061
transform 1 0 18860 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_187
timestamp 1586364061
transform 1 0 18308 0 -1 13600
box -38 -48 222 592
use scs8hd_decap_4  FILLER_20_191
timestamp 1586364061
transform 1 0 18676 0 -1 13600
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_3.LATCH_4_.latch
timestamp 1586364061
transform 1 0 19044 0 -1 13600
box -38 -48 1050 592
use scs8hd_ebufn_2  mux_bottom_ipin_3.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 19688 0 1 12512
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_3.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 19044 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_3.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 19504 0 1 12512
box -38 -48 222 592
use scs8hd_decap_3  FILLER_19_197
timestamp 1586364061
transform 1 0 19228 0 1 12512
box -38 -48 314 592
use scs8hd_decap_6  FILLER_20_206
timestamp 1586364061
transform 1 0 20056 0 -1 13600
box -38 -48 590 592
use scs8hd_buf_2  _142_
timestamp 1586364061
transform 1 0 21252 0 1 12512
box -38 -48 406 592
use scs8hd_ebufn_2  mux_bottom_ipin_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 20884 0 -1 13600
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_148
timestamp 1586364061
transform 1 0 20792 0 -1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 20884 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_3.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 20608 0 -1 13600
box -38 -48 222 592
use scs8hd_decap_4  FILLER_19_211
timestamp 1586364061
transform 1 0 20516 0 1 12512
box -38 -48 406 592
use scs8hd_fill_2  FILLER_19_217
timestamp 1586364061
transform 1 0 21068 0 1 12512
box -38 -48 222 592
use scs8hd_decap_3  PHY_39
timestamp 1586364061
transform -1 0 22816 0 1 12512
box -38 -48 314 592
use scs8hd_decap_3  PHY_41
timestamp 1586364061
transform -1 0 22816 0 -1 13600
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__142__A
timestamp 1586364061
transform 1 0 21804 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_223
timestamp 1586364061
transform 1 0 21620 0 1 12512
box -38 -48 222 592
use scs8hd_decap_6  FILLER_19_227
timestamp 1586364061
transform 1 0 21988 0 1 12512
box -38 -48 590 592
use scs8hd_decap_8  FILLER_20_224
timestamp 1586364061
transform 1 0 21712 0 -1 13600
box -38 -48 774 592
use scs8hd_fill_1  FILLER_20_232
timestamp 1586364061
transform 1 0 22448 0 -1 13600
box -38 -48 130 592
use scs8hd_ebufn_2  mux_bottom_ipin_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 1472 0 1 13600
box -38 -48 866 592
use scs8hd_decap_3  PHY_42
timestamp 1586364061
transform 1 0 1104 0 1 13600
box -38 -48 314 592
use scs8hd_fill_1  FILLER_21_3
timestamp 1586364061
transform 1 0 1380 0 1 13600
box -38 -48 130 592
use scs8hd_fill_2  FILLER_21_13
timestamp 1586364061
transform 1 0 2300 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_0.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 2484 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_0.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 3496 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_0.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 2852 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_17
timestamp 1586364061
transform 1 0 2668 0 1 13600
box -38 -48 222 592
use scs8hd_decap_4  FILLER_21_21
timestamp 1586364061
transform 1 0 3036 0 1 13600
box -38 -48 406 592
use scs8hd_fill_1  FILLER_21_25
timestamp 1586364061
transform 1 0 3404 0 1 13600
box -38 -48 130 592
use scs8hd_ebufn_2  mux_bottom_ipin_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 3680 0 1 13600
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_0.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 4692 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_37
timestamp 1586364061
transform 1 0 4508 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_41
timestamp 1586364061
transform 1 0 4876 0 1 13600
box -38 -48 222 592
use scs8hd_inv_1  mux_bottom_ipin_0.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 5704 0 1 13600
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 6164 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 5060 0 1 13600
box -38 -48 222 592
use scs8hd_decap_4  FILLER_21_45
timestamp 1586364061
transform 1 0 5244 0 1 13600
box -38 -48 406 592
use scs8hd_fill_1  FILLER_21_49
timestamp 1586364061
transform 1 0 5612 0 1 13600
box -38 -48 130 592
use scs8hd_fill_2  FILLER_21_53
timestamp 1586364061
transform 1 0 5980 0 1 13600
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_0.LATCH_2_.latch
timestamp 1586364061
transform 1 0 6808 0 1 13600
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_149
timestamp 1586364061
transform 1 0 6716 0 1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_0.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 6532 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_57
timestamp 1586364061
transform 1 0 6348 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_4.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 8556 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 8004 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_73
timestamp 1586364061
transform 1 0 7820 0 1 13600
box -38 -48 222 592
use scs8hd_decap_4  FILLER_21_77
timestamp 1586364061
transform 1 0 8188 0 1 13600
box -38 -48 406 592
use scs8hd_decap_8  FILLER_21_83
timestamp 1586364061
transform 1 0 8740 0 1 13600
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_0.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 9844 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_0.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 9476 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_93
timestamp 1586364061
transform 1 0 9660 0 1 13600
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_top_ipin_0.LATCH_0_.latch
timestamp 1586364061
transform 1 0 10396 0 1 13600
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_0.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 10212 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_97
timestamp 1586364061
transform 1 0 10028 0 1 13600
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_ipin_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12420 0 1 13600
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_150
timestamp 1586364061
transform 1 0 12328 0 1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 12144 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 11776 0 1 13600
box -38 -48 222 592
use scs8hd_decap_4  FILLER_21_112
timestamp 1586364061
transform 1 0 11408 0 1 13600
box -38 -48 406 592
use scs8hd_fill_2  FILLER_21_118
timestamp 1586364061
transform 1 0 11960 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 13616 0 1 13600
box -38 -48 222 592
use scs8hd_decap_4  FILLER_21_132
timestamp 1586364061
transform 1 0 13248 0 1 13600
box -38 -48 406 592
use scs8hd_fill_2  FILLER_21_138
timestamp 1586364061
transform 1 0 13800 0 1 13600
box -38 -48 222 592
use scs8hd_nor2_4  _130_
timestamp 1586364061
transform 1 0 14720 0 1 13600
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__130__B
timestamp 1586364061
transform 1 0 14536 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 13984 0 1 13600
box -38 -48 222 592
use scs8hd_decap_4  FILLER_21_142
timestamp 1586364061
transform 1 0 14168 0 1 13600
box -38 -48 406 592
use scs8hd_inv_1  mux_bottom_ipin_2.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 16284 0 1 13600
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 15732 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 16100 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_157
timestamp 1586364061
transform 1 0 15548 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_161
timestamp 1586364061
transform 1 0 15916 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 16744 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__056__B
timestamp 1586364061
transform 1 0 17388 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_168
timestamp 1586364061
transform 1 0 16560 0 1 13600
box -38 -48 222 592
use scs8hd_decap_4  FILLER_21_172
timestamp 1586364061
transform 1 0 16928 0 1 13600
box -38 -48 406 592
use scs8hd_fill_1  FILLER_21_176
timestamp 1586364061
transform 1 0 17296 0 1 13600
box -38 -48 130 592
use scs8hd_fill_2  FILLER_21_179
timestamp 1586364061
transform 1 0 17572 0 1 13600
box -38 -48 222 592
use scs8hd_inv_1  mux_bottom_ipin_3.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 18032 0 1 13600
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_151
timestamp 1586364061
transform 1 0 17940 0 1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_3.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 18492 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_3.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 18860 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__056__A
timestamp 1586364061
transform 1 0 17756 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_187
timestamp 1586364061
transform 1 0 18308 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_191
timestamp 1586364061
transform 1 0 18676 0 1 13600
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_3.LATCH_3_.latch
timestamp 1586364061
transform 1 0 19044 0 1 13600
box -38 -48 1050 592
use scs8hd_fill_2  FILLER_21_206
timestamp 1586364061
transform 1 0 20056 0 1 13600
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_ipin_3.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 20792 0 1 13600
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 20240 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_3.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 20608 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_210
timestamp 1586364061
transform 1 0 20424 0 1 13600
box -38 -48 222 592
use scs8hd_decap_3  PHY_43
timestamp 1586364061
transform -1 0 22816 0 1 13600
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_3.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 21804 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_3.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 22172 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_223
timestamp 1586364061
transform 1 0 21620 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_227
timestamp 1586364061
transform 1 0 21988 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_231
timestamp 1586364061
transform 1 0 22356 0 1 13600
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_0.LATCH_4_.latch
timestamp 1586364061
transform 1 0 2208 0 -1 14688
box -38 -48 1050 592
use scs8hd_decap_3  PHY_44
timestamp 1586364061
transform 1 0 1104 0 -1 14688
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__112__A
timestamp 1586364061
transform 1 0 2024 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 1564 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_3
timestamp 1586364061
transform 1 0 1380 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_3  FILLER_22_7
timestamp 1586364061
transform 1 0 1748 0 -1 14688
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__113__A
timestamp 1586364061
transform 1 0 3588 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_22_23
timestamp 1586364061
transform 1 0 3220 0 -1 14688
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_0.LATCH_3_.latch
timestamp 1586364061
transform 1 0 4048 0 -1 14688
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_152
timestamp 1586364061
transform 1 0 3956 0 -1 14688
box -38 -48 130 592
use scs8hd_fill_2  FILLER_22_29
timestamp 1586364061
transform 1 0 3772 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__072__A
timestamp 1586364061
transform 1 0 5244 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_43
timestamp 1586364061
transform 1 0 5060 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_12  FILLER_22_47
timestamp 1586364061
transform 1 0 5428 0 -1 14688
box -38 -48 1142 592
use scs8hd_ebufn_2  mux_bottom_ipin_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 6808 0 -1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 6624 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_1  FILLER_22_59
timestamp 1586364061
transform 1 0 6532 0 -1 14688
box -38 -48 130 592
use scs8hd_inv_1  mux_bottom_ipin_4.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 8556 0 -1 14688
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_4.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 7820 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_71
timestamp 1586364061
transform 1 0 7636 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_6  FILLER_22_75
timestamp 1586364061
transform 1 0 8004 0 -1 14688
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_153
timestamp 1586364061
transform 1 0 9568 0 -1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__101__A
timestamp 1586364061
transform 1 0 9936 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_8  FILLER_22_84
timestamp 1586364061
transform 1 0 8832 0 -1 14688
box -38 -48 774 592
use scs8hd_decap_3  FILLER_22_93
timestamp 1586364061
transform 1 0 9660 0 -1 14688
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_top_ipin_0.LATCH_2_.latch
timestamp 1586364061
transform 1 0 10212 0 -1 14688
box -38 -48 1050 592
use scs8hd_fill_1  FILLER_22_98
timestamp 1586364061
transform 1 0 10120 0 -1 14688
box -38 -48 130 592
use scs8hd_decap_8  FILLER_22_110
timestamp 1586364061
transform 1 0 11224 0 -1 14688
box -38 -48 774 592
use scs8hd_ebufn_2  mux_top_ipin_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12052 0 -1 14688
box -38 -48 866 592
use scs8hd_fill_1  FILLER_22_118
timestamp 1586364061
transform 1 0 11960 0 -1 14688
box -38 -48 130 592
use scs8hd_ebufn_2  mux_top_ipin_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 13616 0 -1 14688
box -38 -48 866 592
use scs8hd_decap_8  FILLER_22_128
timestamp 1586364061
transform 1 0 12880 0 -1 14688
box -38 -48 774 592
use scs8hd_decap_8  FILLER_22_145
timestamp 1586364061
transform 1 0 14444 0 -1 14688
box -38 -48 774 592
use scs8hd_ebufn_2  mux_bottom_ipin_2.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15640 0 -1 14688
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_154
timestamp 1586364061
transform 1 0 15180 0 -1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_2.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 15456 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_154
timestamp 1586364061
transform 1 0 15272 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_12  FILLER_22_167
timestamp 1586364061
transform 1 0 16468 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_22_179
timestamp 1586364061
transform 1 0 17572 0 -1 14688
box -38 -48 314 592
use scs8hd_nor2_4  _056_
timestamp 1586364061
transform 1 0 17848 0 -1 14688
box -38 -48 866 592
use scs8hd_decap_4  FILLER_22_191
timestamp 1586364061
transform 1 0 18676 0 -1 14688
box -38 -48 406 592
use scs8hd_inv_1  mux_bottom_ipin_2.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 19412 0 -1 14688
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_3.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 19044 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_197
timestamp 1586364061
transform 1 0 19228 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_12  FILLER_22_202
timestamp 1586364061
transform 1 0 19688 0 -1 14688
box -38 -48 1142 592
use scs8hd_ebufn_2  mux_bottom_ipin_3.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 20884 0 -1 14688
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_155
timestamp 1586364061
transform 1 0 20792 0 -1 14688
box -38 -48 130 592
use scs8hd_decap_3  PHY_45
timestamp 1586364061
transform -1 0 22816 0 -1 14688
box -38 -48 314 592
use scs8hd_decap_8  FILLER_22_224
timestamp 1586364061
transform 1 0 21712 0 -1 14688
box -38 -48 774 592
use scs8hd_fill_1  FILLER_22_232
timestamp 1586364061
transform 1 0 22448 0 -1 14688
box -38 -48 130 592
use scs8hd_nor2_4  _112_
timestamp 1586364061
transform 1 0 2024 0 1 14688
box -38 -48 866 592
use scs8hd_decap_3  PHY_46
timestamp 1586364061
transform 1 0 1104 0 1 14688
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__112__B
timestamp 1586364061
transform 1 0 1840 0 1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_23_3
timestamp 1586364061
transform 1 0 1380 0 1 14688
box -38 -48 406 592
use scs8hd_fill_1  FILLER_23_7
timestamp 1586364061
transform 1 0 1748 0 1 14688
box -38 -48 130 592
use scs8hd_nor2_4  _113_
timestamp 1586364061
transform 1 0 3588 0 1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__113__B
timestamp 1586364061
transform 1 0 3404 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 3036 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_19
timestamp 1586364061
transform 1 0 2852 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_23
timestamp 1586364061
transform 1 0 3220 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_4.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 4692 0 1 14688
box -38 -48 222 592
use scs8hd_decap_3  FILLER_23_36
timestamp 1586364061
transform 1 0 4416 0 1 14688
box -38 -48 314 592
use scs8hd_decap_3  FILLER_23_41
timestamp 1586364061
transform 1 0 4876 0 1 14688
box -38 -48 314 592
use scs8hd_nor2_4  _072_
timestamp 1586364061
transform 1 0 5152 0 1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__114__B
timestamp 1586364061
transform 1 0 6164 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_53
timestamp 1586364061
transform 1 0 5980 0 1 14688
box -38 -48 222 592
use scs8hd_nor2_4  _074_
timestamp 1586364061
transform 1 0 7452 0 1 14688
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_156
timestamp 1586364061
transform 1 0 6716 0 1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__074__B
timestamp 1586364061
transform 1 0 7268 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__114__A
timestamp 1586364061
transform 1 0 6532 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_57
timestamp 1586364061
transform 1 0 6348 0 1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_23_62
timestamp 1586364061
transform 1 0 6808 0 1 14688
box -38 -48 406 592
use scs8hd_fill_1  FILLER_23_66
timestamp 1586364061
transform 1 0 7176 0 1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_4.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 8464 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_78
timestamp 1586364061
transform 1 0 8280 0 1 14688
box -38 -48 222 592
use scs8hd_decap_3  FILLER_23_82
timestamp 1586364061
transform 1 0 8648 0 1 14688
box -38 -48 314 592
use scs8hd_nor2_4  _103_
timestamp 1586364061
transform 1 0 9476 0 1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__103__B
timestamp 1586364061
transform 1 0 9292 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__103__A
timestamp 1586364061
transform 1 0 8924 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_87
timestamp 1586364061
transform 1 0 9108 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 11132 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__101__B
timestamp 1586364061
transform 1 0 10488 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_100
timestamp 1586364061
transform 1 0 10304 0 1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_23_104
timestamp 1586364061
transform 1 0 10672 0 1 14688
box -38 -48 406 592
use scs8hd_fill_1  FILLER_23_108
timestamp 1586364061
transform 1 0 11040 0 1 14688
box -38 -48 130 592
use scs8hd_inv_1  mux_top_ipin_0.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 11316 0 1 14688
box -38 -48 314 592
use scs8hd_ebufn_2  mux_top_ipin_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12420 0 1 14688
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_157
timestamp 1586364061
transform 1 0 12328 0 1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 11868 0 1 14688
box -38 -48 222 592
use scs8hd_decap_3  FILLER_23_114
timestamp 1586364061
transform 1 0 11592 0 1 14688
box -38 -48 314 592
use scs8hd_decap_3  FILLER_23_119
timestamp 1586364061
transform 1 0 12052 0 1 14688
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_3.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 13432 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__128__B
timestamp 1586364061
transform 1 0 13800 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_132
timestamp 1586364061
transform 1 0 13248 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_136
timestamp 1586364061
transform 1 0 13616 0 1 14688
box -38 -48 222 592
use scs8hd_nor2_4  _128_
timestamp 1586364061
transform 1 0 13984 0 1 14688
box -38 -48 866 592
use scs8hd_decap_4  FILLER_23_149
timestamp 1586364061
transform 1 0 14812 0 1 14688
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_2.LATCH_0_.latch
timestamp 1586364061
transform 1 0 16008 0 1 14688
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_2.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 15272 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_2.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 15824 0 1 14688
box -38 -48 222 592
use scs8hd_fill_1  FILLER_23_153
timestamp 1586364061
transform 1 0 15180 0 1 14688
box -38 -48 130 592
use scs8hd_decap_4  FILLER_23_156
timestamp 1586364061
transform 1 0 15456 0 1 14688
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 17204 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_173
timestamp 1586364061
transform 1 0 17020 0 1 14688
box -38 -48 222 592
use scs8hd_decap_6  FILLER_23_177
timestamp 1586364061
transform 1 0 17388 0 1 14688
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_158
timestamp 1586364061
transform 1 0 17940 0 1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 18216 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 18584 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_184
timestamp 1586364061
transform 1 0 18032 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_188
timestamp 1586364061
transform 1 0 18400 0 1 14688
box -38 -48 222 592
use scs8hd_decap_6  FILLER_23_192
timestamp 1586364061
transform 1 0 18768 0 1 14688
box -38 -48 590 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_3.LATCH_5_.latch
timestamp 1586364061
transform 1 0 19504 0 1 14688
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_3.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 19320 0 1 14688
box -38 -48 222 592
use scs8hd_conb_1  _134_
timestamp 1586364061
transform 1 0 21252 0 1 14688
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_3.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 20884 0 1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_23_211
timestamp 1586364061
transform 1 0 20516 0 1 14688
box -38 -48 406 592
use scs8hd_fill_2  FILLER_23_217
timestamp 1586364061
transform 1 0 21068 0 1 14688
box -38 -48 222 592
use scs8hd_decap_3  PHY_47
timestamp 1586364061
transform -1 0 22816 0 1 14688
box -38 -48 314 592
use scs8hd_decap_8  FILLER_23_222
timestamp 1586364061
transform 1 0 21528 0 1 14688
box -38 -48 774 592
use scs8hd_decap_3  FILLER_23_230
timestamp 1586364061
transform 1 0 22264 0 1 14688
box -38 -48 314 592
use scs8hd_inv_1  mux_bottom_ipin_0.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1380 0 -1 15776
box -38 -48 314 592
use scs8hd_decap_3  PHY_48
timestamp 1586364061
transform 1 0 1104 0 -1 15776
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__069__B
timestamp 1586364061
transform 1 0 1840 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__069__A
timestamp 1586364061
transform 1 0 2208 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_6
timestamp 1586364061
transform 1 0 1656 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_10
timestamp 1586364061
transform 1 0 2024 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__070__A
timestamp 1586364061
transform 1 0 2576 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_14
timestamp 1586364061
transform 1 0 2392 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_12  FILLER_24_18
timestamp 1586364061
transform 1 0 2760 0 -1 15776
box -38 -48 1142 592
use scs8hd_inv_1  mux_bottom_ipin_4.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 4692 0 -1 15776
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_159
timestamp 1586364061
transform 1 0 3956 0 -1 15776
box -38 -48 130 592
use scs8hd_fill_1  FILLER_24_30
timestamp 1586364061
transform 1 0 3864 0 -1 15776
box -38 -48 130 592
use scs8hd_decap_6  FILLER_24_32
timestamp 1586364061
transform 1 0 4048 0 -1 15776
box -38 -48 590 592
use scs8hd_fill_1  FILLER_24_38
timestamp 1586364061
transform 1 0 4600 0 -1 15776
box -38 -48 130 592
use scs8hd_nor2_4  _114_
timestamp 1586364061
transform 1 0 5704 0 -1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__072__B
timestamp 1586364061
transform 1 0 5152 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_42
timestamp 1586364061
transform 1 0 4968 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_24_46
timestamp 1586364061
transform 1 0 5336 0 -1 15776
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__074__A
timestamp 1586364061
transform 1 0 7452 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_4.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 7084 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_6  FILLER_24_59
timestamp 1586364061
transform 1 0 6532 0 -1 15776
box -38 -48 590 592
use scs8hd_fill_2  FILLER_24_67
timestamp 1586364061
transform 1 0 7268 0 -1 15776
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_4.LATCH_0_.latch
timestamp 1586364061
transform 1 0 7820 0 -1 15776
box -38 -48 1050 592
use scs8hd_fill_2  FILLER_24_71
timestamp 1586364061
transform 1 0 7636 0 -1 15776
box -38 -48 222 592
use scs8hd_nor2_4  _101_
timestamp 1586364061
transform 1 0 9936 0 -1 15776
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_160
timestamp 1586364061
transform 1 0 9568 0 -1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_4.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9016 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_84
timestamp 1586364061
transform 1 0 8832 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_24_88
timestamp 1586364061
transform 1 0 9200 0 -1 15776
box -38 -48 406 592
use scs8hd_decap_3  FILLER_24_93
timestamp 1586364061
transform 1 0 9660 0 -1 15776
box -38 -48 314 592
use scs8hd_decap_12  FILLER_24_105
timestamp 1586364061
transform 1 0 10764 0 -1 15776
box -38 -48 1142 592
use scs8hd_inv_1  mux_top_ipin_0.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 11868 0 -1 15776
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 12420 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_3  FILLER_24_120
timestamp 1586364061
transform 1 0 12144 0 -1 15776
box -38 -48 314 592
use scs8hd_inv_1  mux_bottom_ipin_3.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 13432 0 -1 15776
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 12788 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_125
timestamp 1586364061
transform 1 0 12604 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_24_129
timestamp 1586364061
transform 1 0 12972 0 -1 15776
box -38 -48 406 592
use scs8hd_fill_1  FILLER_24_133
timestamp 1586364061
transform 1 0 13340 0 -1 15776
box -38 -48 130 592
use scs8hd_decap_3  FILLER_24_137
timestamp 1586364061
transform 1 0 13708 0 -1 15776
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__128__A
timestamp 1586364061
transform 1 0 13984 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_8  FILLER_24_142
timestamp 1586364061
transform 1 0 14168 0 -1 15776
box -38 -48 774 592
use scs8hd_decap_3  FILLER_24_150
timestamp 1586364061
transform 1 0 14904 0 -1 15776
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_2.LATCH_2_.latch
timestamp 1586364061
transform 1 0 15272 0 -1 15776
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_161
timestamp 1586364061
transform 1 0 15180 0 -1 15776
box -38 -48 130 592
use scs8hd_fill_2  FILLER_24_165
timestamp 1586364061
transform 1 0 16284 0 -1 15776
box -38 -48 222 592
use scs8hd_inv_1  mux_bottom_ipin_2.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 17020 0 -1 15776
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_2.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 16468 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_24_169
timestamp 1586364061
transform 1 0 16652 0 -1 15776
box -38 -48 406 592
use scs8hd_decap_8  FILLER_24_176
timestamp 1586364061
transform 1 0 17296 0 -1 15776
box -38 -48 774 592
use scs8hd_ebufn_2  mux_bottom_ipin_2.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18124 0 -1 15776
box -38 -48 866 592
use scs8hd_fill_1  FILLER_24_184
timestamp 1586364061
transform 1 0 18032 0 -1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_3.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 19504 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_6  FILLER_24_194
timestamp 1586364061
transform 1 0 18952 0 -1 15776
box -38 -48 590 592
use scs8hd_decap_12  FILLER_24_202
timestamp 1586364061
transform 1 0 19688 0 -1 15776
box -38 -48 1142 592
use scs8hd_inv_1  mux_bottom_ipin_3.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 20884 0 -1 15776
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_162
timestamp 1586364061
transform 1 0 20792 0 -1 15776
box -38 -48 130 592
use scs8hd_decap_12  FILLER_24_218
timestamp 1586364061
transform 1 0 21160 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_3  PHY_49
timestamp 1586364061
transform -1 0 22816 0 -1 15776
box -38 -48 314 592
use scs8hd_decap_3  FILLER_24_230
timestamp 1586364061
transform 1 0 22264 0 -1 15776
box -38 -48 314 592
use scs8hd_buf_2  _151_
timestamp 1586364061
transform 1 0 1380 0 1 15776
box -38 -48 406 592
use scs8hd_decap_3  PHY_50
timestamp 1586364061
transform 1 0 1104 0 1 15776
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__151__A
timestamp 1586364061
transform 1 0 1932 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_7
timestamp 1586364061
transform 1 0 1748 0 1 15776
box -38 -48 222 592
use scs8hd_decap_3  FILLER_25_11
timestamp 1586364061
transform 1 0 2116 0 1 15776
box -38 -48 314 592
use scs8hd_nor2_4  _070_
timestamp 1586364061
transform 1 0 2576 0 1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__070__B
timestamp 1586364061
transform 1 0 2392 0 1 15776
box -38 -48 222 592
use scs8hd_decap_3  FILLER_25_25
timestamp 1586364061
transform 1 0 3404 0 1 15776
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_4.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 4048 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_4.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 4784 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_4.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 4416 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_4.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 3680 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_30
timestamp 1586364061
transform 1 0 3864 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_34
timestamp 1586364061
transform 1 0 4232 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_38
timestamp 1586364061
transform 1 0 4600 0 1 15776
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_4.LATCH_2_.latch
timestamp 1586364061
transform 1 0 4968 0 1 15776
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_4.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 6164 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_53
timestamp 1586364061
transform 1 0 5980 0 1 15776
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_ipin_4.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 6808 0 1 15776
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_163
timestamp 1586364061
transform 1 0 6716 0 1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_4.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 6532 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_57
timestamp 1586364061
transform 1 0 6348 0 1 15776
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_ipin_4.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 8372 0 1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_4.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 8188 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_4.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 7820 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_71
timestamp 1586364061
transform 1 0 7636 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_75
timestamp 1586364061
transform 1 0 8004 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_4.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 9660 0 1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_25_88
timestamp 1586364061
transform 1 0 9200 0 1 15776
box -38 -48 406 592
use scs8hd_fill_1  FILLER_25_92
timestamp 1586364061
transform 1 0 9568 0 1 15776
box -38 -48 130 592
use scs8hd_fill_2  FILLER_25_95
timestamp 1586364061
transform 1 0 9844 0 1 15776
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_top_ipin_0.LATCH_4_.latch
timestamp 1586364061
transform 1 0 10580 0 1 15776
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_0.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 10396 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_0.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 10028 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_99
timestamp 1586364061
transform 1 0 10212 0 1 15776
box -38 -48 222 592
use scs8hd_inv_1  mux_top_ipin_0.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 12420 0 1 15776
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_164
timestamp 1586364061
transform 1 0 12328 0 1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_0.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 11776 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_0.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 12144 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_114
timestamp 1586364061
transform 1 0 11592 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_118
timestamp 1586364061
transform 1 0 11960 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 12880 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 13248 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 13616 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_126
timestamp 1586364061
transform 1 0 12696 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_130
timestamp 1586364061
transform 1 0 13064 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_134
timestamp 1586364061
transform 1 0 13432 0 1 15776
box -38 -48 222 592
use scs8hd_decap_8  FILLER_25_138
timestamp 1586364061
transform 1 0 13800 0 1 15776
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 15088 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14720 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_146
timestamp 1586364061
transform 1 0 14536 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_150
timestamp 1586364061
transform 1 0 14904 0 1 15776
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_ipin_2.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15732 0 1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 15456 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_154
timestamp 1586364061
transform 1 0 15272 0 1 15776
box -38 -48 222 592
use scs8hd_fill_1  FILLER_25_158
timestamp 1586364061
transform 1 0 15640 0 1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__126__B
timestamp 1586364061
transform 1 0 16928 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__126__A
timestamp 1586364061
transform 1 0 17296 0 1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_25_168
timestamp 1586364061
transform 1 0 16560 0 1 15776
box -38 -48 406 592
use scs8hd_fill_2  FILLER_25_174
timestamp 1586364061
transform 1 0 17112 0 1 15776
box -38 -48 222 592
use scs8hd_decap_3  FILLER_25_178
timestamp 1586364061
transform 1 0 17480 0 1 15776
box -38 -48 314 592
use scs8hd_ebufn_2  mux_bottom_ipin_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18032 0 1 15776
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_165
timestamp 1586364061
transform 1 0 17940 0 1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 17756 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_193
timestamp 1586364061
transform 1 0 18860 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_2.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 19044 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_2.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 19412 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_197
timestamp 1586364061
transform 1 0 19228 0 1 15776
box -38 -48 222 592
use scs8hd_decap_12  FILLER_25_201
timestamp 1586364061
transform 1 0 19596 0 1 15776
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA__158__A
timestamp 1586364061
transform 1 0 20884 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_213
timestamp 1586364061
transform 1 0 20700 0 1 15776
box -38 -48 222 592
use scs8hd_decap_12  FILLER_25_217
timestamp 1586364061
transform 1 0 21068 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_3  PHY_51
timestamp 1586364061
transform -1 0 22816 0 1 15776
box -38 -48 314 592
use scs8hd_decap_4  FILLER_25_229
timestamp 1586364061
transform 1 0 22172 0 1 15776
box -38 -48 406 592
use scs8hd_nor2_4  _069_
timestamp 1586364061
transform 1 0 1748 0 -1 16864
box -38 -48 866 592
use scs8hd_ebufn_2  mux_bottom_ipin_4.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 2208 0 1 16864
box -38 -48 866 592
use scs8hd_decap_3  PHY_52
timestamp 1586364061
transform 1 0 1104 0 -1 16864
box -38 -48 314 592
use scs8hd_decap_3  PHY_54
timestamp 1586364061
transform 1 0 1104 0 1 16864
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_4.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 1840 0 1 16864
box -38 -48 222 592
use scs8hd_decap_4  FILLER_26_3
timestamp 1586364061
transform 1 0 1380 0 -1 16864
box -38 -48 406 592
use scs8hd_decap_4  FILLER_27_3
timestamp 1586364061
transform 1 0 1380 0 1 16864
box -38 -48 406 592
use scs8hd_fill_1  FILLER_27_7
timestamp 1586364061
transform 1 0 1748 0 1 16864
box -38 -48 130 592
use scs8hd_fill_2  FILLER_27_10
timestamp 1586364061
transform 1 0 2024 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_4.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 3220 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_4.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 2760 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_16
timestamp 1586364061
transform 1 0 2576 0 -1 16864
box -38 -48 222 592
use scs8hd_decap_8  FILLER_26_20
timestamp 1586364061
transform 1 0 2944 0 -1 16864
box -38 -48 774 592
use scs8hd_fill_2  FILLER_27_21
timestamp 1586364061
transform 1 0 3036 0 1 16864
box -38 -48 222 592
use scs8hd_decap_4  FILLER_27_25
timestamp 1586364061
transform 1 0 3404 0 1 16864
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_4.LATCH_4_.latch
timestamp 1586364061
transform 1 0 4048 0 -1 16864
box -38 -48 1050 592
use scs8hd_ebufn_2  mux_bottom_ipin_4.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 4324 0 1 16864
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_166
timestamp 1586364061
transform 1 0 3956 0 -1 16864
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_4.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 4140 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_4.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 3772 0 1 16864
box -38 -48 222 592
use scs8hd_decap_3  FILLER_26_28
timestamp 1586364061
transform 1 0 3680 0 -1 16864
box -38 -48 314 592
use scs8hd_fill_2  FILLER_27_31
timestamp 1586364061
transform 1 0 3956 0 1 16864
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_ipin_4.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 5796 0 -1 16864
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_4.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 5980 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_4.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 5336 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_4.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 5612 0 -1 16864
box -38 -48 222 592
use scs8hd_decap_6  FILLER_26_43
timestamp 1586364061
transform 1 0 5060 0 -1 16864
box -38 -48 590 592
use scs8hd_fill_2  FILLER_27_44
timestamp 1586364061
transform 1 0 5152 0 1 16864
box -38 -48 222 592
use scs8hd_decap_4  FILLER_27_48
timestamp 1586364061
transform 1 0 5520 0 1 16864
box -38 -48 406 592
use scs8hd_fill_1  FILLER_27_52
timestamp 1586364061
transform 1 0 5888 0 1 16864
box -38 -48 130 592
use scs8hd_decap_6  FILLER_27_55
timestamp 1586364061
transform 1 0 6164 0 1 16864
box -38 -48 590 592
use scs8hd_fill_2  FILLER_26_60
timestamp 1586364061
transform 1 0 6624 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_65
timestamp 1586364061
transform 1 0 7084 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_64
timestamp 1586364061
transform 1 0 6992 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_4.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 6808 0 -1 16864
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_170
timestamp 1586364061
transform 1 0 6716 0 1 16864
box -38 -48 130 592
use scs8hd_inv_1  mux_bottom_ipin_4.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 6808 0 1 16864
box -38 -48 314 592
use scs8hd_fill_2  FILLER_27_69
timestamp 1586364061
transform 1 0 7452 0 1 16864
box -38 -48 222 592
use scs8hd_decap_4  FILLER_26_68
timestamp 1586364061
transform 1 0 7360 0 -1 16864
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_4.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 7176 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_4.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 7268 0 1 16864
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_ipin_4.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 8004 0 -1 16864
box -38 -48 866 592
use scs8hd_ebufn_2  mux_bottom_ipin_4.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 7820 0 1 16864
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_4.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 7636 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_4.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 7820 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_1  FILLER_26_72
timestamp 1586364061
transform 1 0 7728 0 -1 16864
box -38 -48 130 592
use scs8hd_fill_2  FILLER_27_82
timestamp 1586364061
transform 1 0 8648 0 1 16864
box -38 -48 222 592
use scs8hd_inv_1  mux_bottom_ipin_4.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 9384 0 1 16864
box -38 -48 314 592
use scs8hd_inv_1  mux_bottom_ipin_4.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 9660 0 -1 16864
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_167
timestamp 1586364061
transform 1 0 9568 0 -1 16864
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_4.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 9844 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_4.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 8832 0 1 16864
box -38 -48 222 592
use scs8hd_decap_8  FILLER_26_84
timestamp 1586364061
transform 1 0 8832 0 -1 16864
box -38 -48 774 592
use scs8hd_decap_6  FILLER_26_96
timestamp 1586364061
transform 1 0 9936 0 -1 16864
box -38 -48 590 592
use scs8hd_decap_4  FILLER_27_86
timestamp 1586364061
transform 1 0 9016 0 1 16864
box -38 -48 406 592
use scs8hd_fill_2  FILLER_27_93
timestamp 1586364061
transform 1 0 9660 0 1 16864
box -38 -48 222 592
use scs8hd_nor2_4  _104_
timestamp 1586364061
transform 1 0 10396 0 1 16864
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__104__B
timestamp 1586364061
transform 1 0 10212 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__102__A
timestamp 1586364061
transform 1 0 10580 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_1  FILLER_26_102
timestamp 1586364061
transform 1 0 10488 0 -1 16864
box -38 -48 130 592
use scs8hd_decap_6  FILLER_26_105
timestamp 1586364061
transform 1 0 10764 0 -1 16864
box -38 -48 590 592
use scs8hd_fill_2  FILLER_27_97
timestamp 1586364061
transform 1 0 10028 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_110
timestamp 1586364061
transform 1 0 11224 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_114
timestamp 1586364061
transform 1 0 11592 0 1 16864
box -38 -48 222 592
use scs8hd_fill_1  FILLER_26_111
timestamp 1586364061
transform 1 0 11316 0 -1 16864
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 11776 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__102__B
timestamp 1586364061
transform 1 0 11408 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_118
timestamp 1586364061
transform 1 0 11960 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_123
timestamp 1586364061
transform 1 0 12420 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 12144 0 1 16864
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_171
timestamp 1586364061
transform 1 0 12328 0 1 16864
box -38 -48 130 592
use scs8hd_ebufn_2  mux_top_ipin_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12420 0 1 16864
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  mem_top_ipin_0.LATCH_1_.latch
timestamp 1586364061
transform 1 0 11408 0 -1 16864
box -38 -48 1050 592
use scs8hd_ebufn_2  mux_top_ipin_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 13156 0 -1 16864
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__129__B
timestamp 1586364061
transform 1 0 13524 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 12604 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 12972 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_127
timestamp 1586364061
transform 1 0 12788 0 -1 16864
box -38 -48 222 592
use scs8hd_decap_3  FILLER_27_132
timestamp 1586364061
transform 1 0 13248 0 1 16864
box -38 -48 314 592
use scs8hd_fill_2  FILLER_27_137
timestamp 1586364061
transform 1 0 13708 0 1 16864
box -38 -48 222 592
use scs8hd_nor2_4  _129_
timestamp 1586364061
transform 1 0 14076 0 1 16864
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 13892 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__129__A
timestamp 1586364061
transform 1 0 14168 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_140
timestamp 1586364061
transform 1 0 13984 0 -1 16864
box -38 -48 222 592
use scs8hd_decap_8  FILLER_26_144
timestamp 1586364061
transform 1 0 14352 0 -1 16864
box -38 -48 774 592
use scs8hd_fill_1  FILLER_26_152
timestamp 1586364061
transform 1 0 15088 0 -1 16864
box -38 -48 130 592
use scs8hd_decap_4  FILLER_27_150
timestamp 1586364061
transform 1 0 14904 0 1 16864
box -38 -48 406 592
use scs8hd_fill_2  FILLER_27_156
timestamp 1586364061
transform 1 0 15456 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_159
timestamp 1586364061
transform 1 0 15732 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_154
timestamp 1586364061
transform 1 0 15272 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_2.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 15272 0 1 16864
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_168
timestamp 1586364061
transform 1 0 15180 0 -1 16864
box -38 -48 130 592
use scs8hd_inv_1  mux_bottom_ipin_2.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 15456 0 -1 16864
box -38 -48 314 592
use scs8hd_fill_2  FILLER_26_163
timestamp 1586364061
transform 1 0 16100 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 16284 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 15916 0 -1 16864
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_ipin_2.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15640 0 1 16864
box -38 -48 866 592
use scs8hd_nor2_4  _126_
timestamp 1586364061
transform 1 0 16928 0 -1 16864
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_2.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 17112 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_2.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 16652 0 1 16864
box -38 -48 222 592
use scs8hd_decap_4  FILLER_26_167
timestamp 1586364061
transform 1 0 16468 0 -1 16864
box -38 -48 406 592
use scs8hd_fill_1  FILLER_26_171
timestamp 1586364061
transform 1 0 16836 0 -1 16864
box -38 -48 130 592
use scs8hd_fill_2  FILLER_27_167
timestamp 1586364061
transform 1 0 16468 0 1 16864
box -38 -48 222 592
use scs8hd_decap_3  FILLER_27_171
timestamp 1586364061
transform 1 0 16836 0 1 16864
box -38 -48 314 592
use scs8hd_decap_4  FILLER_27_176
timestamp 1586364061
transform 1 0 17296 0 1 16864
box -38 -48 406 592
use scs8hd_fill_1  FILLER_27_180
timestamp 1586364061
transform 1 0 17664 0 1 16864
box -38 -48 130 592
use scs8hd_fill_2  FILLER_26_185
timestamp 1586364061
transform 1 0 18124 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_181
timestamp 1586364061
transform 1 0 17756 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_2.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 17940 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 17756 0 1 16864
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_172
timestamp 1586364061
transform 1 0 17940 0 1 16864
box -38 -48 130 592
use scs8hd_fill_2  FILLER_27_193
timestamp 1586364061
transform 1 0 18860 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 18308 0 -1 16864
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_ipin_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18032 0 1 16864
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_2.LATCH_4_.latch
timestamp 1586364061
transform 1 0 18492 0 -1 16864
box -38 -48 1050 592
use scs8hd_ebufn_2  mux_bottom_ipin_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 19596 0 1 16864
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__125__B
timestamp 1586364061
transform 1 0 19044 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__125__A
timestamp 1586364061
transform 1 0 19412 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 19688 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_200
timestamp 1586364061
transform 1 0 19504 0 -1 16864
box -38 -48 222 592
use scs8hd_decap_8  FILLER_26_204
timestamp 1586364061
transform 1 0 19872 0 -1 16864
box -38 -48 774 592
use scs8hd_fill_2  FILLER_27_197
timestamp 1586364061
transform 1 0 19228 0 1 16864
box -38 -48 222 592
use scs8hd_buf_2  _158_
timestamp 1586364061
transform 1 0 20884 0 -1 16864
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_169
timestamp 1586364061
transform 1 0 20792 0 -1 16864
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__153__A
timestamp 1586364061
transform 1 0 20884 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_212
timestamp 1586364061
transform 1 0 20608 0 -1 16864
box -38 -48 222 592
use scs8hd_decap_12  FILLER_26_219
timestamp 1586364061
transform 1 0 21252 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_27_210
timestamp 1586364061
transform 1 0 20424 0 1 16864
box -38 -48 406 592
use scs8hd_fill_1  FILLER_27_214
timestamp 1586364061
transform 1 0 20792 0 1 16864
box -38 -48 130 592
use scs8hd_decap_12  FILLER_27_217
timestamp 1586364061
transform 1 0 21068 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_3  PHY_53
timestamp 1586364061
transform -1 0 22816 0 -1 16864
box -38 -48 314 592
use scs8hd_decap_3  PHY_55
timestamp 1586364061
transform -1 0 22816 0 1 16864
box -38 -48 314 592
use scs8hd_fill_2  FILLER_26_231
timestamp 1586364061
transform 1 0 22356 0 -1 16864
box -38 -48 222 592
use scs8hd_decap_4  FILLER_27_229
timestamp 1586364061
transform 1 0 22172 0 1 16864
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_4.LATCH_5_.latch
timestamp 1586364061
transform 1 0 1840 0 -1 17952
box -38 -48 1050 592
use scs8hd_decap_3  PHY_56
timestamp 1586364061
transform 1 0 1104 0 -1 17952
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_4.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 1656 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_3  FILLER_28_3
timestamp 1586364061
transform 1 0 1380 0 -1 17952
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__071__A
timestamp 1586364061
transform 1 0 3312 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_4  FILLER_28_19
timestamp 1586364061
transform 1 0 2852 0 -1 17952
box -38 -48 406 592
use scs8hd_fill_1  FILLER_28_23
timestamp 1586364061
transform 1 0 3220 0 -1 17952
box -38 -48 130 592
use scs8hd_decap_4  FILLER_28_26
timestamp 1586364061
transform 1 0 3496 0 -1 17952
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_4.LATCH_3_.latch
timestamp 1586364061
transform 1 0 4232 0 -1 17952
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_173
timestamp 1586364061
transform 1 0 3956 0 -1 17952
box -38 -48 130 592
use scs8hd_fill_1  FILLER_28_30
timestamp 1586364061
transform 1 0 3864 0 -1 17952
box -38 -48 130 592
use scs8hd_fill_2  FILLER_28_32
timestamp 1586364061
transform 1 0 4048 0 -1 17952
box -38 -48 222 592
use scs8hd_inv_1  mux_bottom_ipin_4.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 5980 0 -1 17952
box -38 -48 314 592
use scs8hd_decap_8  FILLER_28_45
timestamp 1586364061
transform 1 0 5244 0 -1 17952
box -38 -48 774 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_4.LATCH_1_.latch
timestamp 1586364061
transform 1 0 7176 0 -1 17952
box -38 -48 1050 592
use scs8hd_decap_8  FILLER_28_56
timestamp 1586364061
transform 1 0 6256 0 -1 17952
box -38 -48 774 592
use scs8hd_fill_2  FILLER_28_64
timestamp 1586364061
transform 1 0 6992 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_12  FILLER_28_77
timestamp 1586364061
transform 1 0 8188 0 -1 17952
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_174
timestamp 1586364061
transform 1 0 9568 0 -1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__100__A
timestamp 1586364061
transform 1 0 9844 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_3  FILLER_28_89
timestamp 1586364061
transform 1 0 9292 0 -1 17952
box -38 -48 314 592
use scs8hd_fill_2  FILLER_28_93
timestamp 1586364061
transform 1 0 9660 0 -1 17952
box -38 -48 222 592
use scs8hd_nor2_4  _102_
timestamp 1586364061
transform 1 0 10580 0 -1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__104__A
timestamp 1586364061
transform 1 0 10396 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_4  FILLER_28_97
timestamp 1586364061
transform 1 0 10028 0 -1 17952
box -38 -48 406 592
use scs8hd_ebufn_2  mux_top_ipin_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12420 0 -1 17952
box -38 -48 866 592
use scs8hd_decap_8  FILLER_28_112
timestamp 1586364061
transform 1 0 11408 0 -1 17952
box -38 -48 774 592
use scs8hd_decap_3  FILLER_28_120
timestamp 1586364061
transform 1 0 12144 0 -1 17952
box -38 -48 314 592
use scs8hd_decap_8  FILLER_28_132
timestamp 1586364061
transform 1 0 13248 0 -1 17952
box -38 -48 774 592
use scs8hd_inv_1  mux_top_ipin_0.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 13984 0 -1 17952
box -38 -48 314 592
use scs8hd_decap_8  FILLER_28_143
timestamp 1586364061
transform 1 0 14260 0 -1 17952
box -38 -48 774 592
use scs8hd_fill_2  FILLER_28_151
timestamp 1586364061
transform 1 0 14996 0 -1 17952
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_2.LATCH_1_.latch
timestamp 1586364061
transform 1 0 15272 0 -1 17952
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_175
timestamp 1586364061
transform 1 0 15180 0 -1 17952
box -38 -48 130 592
use scs8hd_decap_8  FILLER_28_165
timestamp 1586364061
transform 1 0 16284 0 -1 17952
box -38 -48 774 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_2.LATCH_3_.latch
timestamp 1586364061
transform 1 0 17112 0 -1 17952
box -38 -48 1050 592
use scs8hd_fill_1  FILLER_28_173
timestamp 1586364061
transform 1 0 17020 0 -1 17952
box -38 -48 130 592
use scs8hd_nor2_4  _125_
timestamp 1586364061
transform 1 0 18860 0 -1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 18308 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_185
timestamp 1586364061
transform 1 0 18124 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_4  FILLER_28_189
timestamp 1586364061
transform 1 0 18492 0 -1 17952
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 19872 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_202
timestamp 1586364061
transform 1 0 19688 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_4  FILLER_28_206
timestamp 1586364061
transform 1 0 20056 0 -1 17952
box -38 -48 406 592
use scs8hd_buf_2  _153_
timestamp 1586364061
transform 1 0 20884 0 -1 17952
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_176
timestamp 1586364061
transform 1 0 20792 0 -1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 20516 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_1  FILLER_28_210
timestamp 1586364061
transform 1 0 20424 0 -1 17952
box -38 -48 130 592
use scs8hd_fill_1  FILLER_28_213
timestamp 1586364061
transform 1 0 20700 0 -1 17952
box -38 -48 130 592
use scs8hd_decap_12  FILLER_28_219
timestamp 1586364061
transform 1 0 21252 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_3  PHY_57
timestamp 1586364061
transform -1 0 22816 0 -1 17952
box -38 -48 314 592
use scs8hd_fill_2  FILLER_28_231
timestamp 1586364061
transform 1 0 22356 0 -1 17952
box -38 -48 222 592
use scs8hd_conb_1  _135_
timestamp 1586364061
transform 1 0 1932 0 1 17952
box -38 -48 314 592
use scs8hd_decap_3  PHY_58
timestamp 1586364061
transform 1 0 1104 0 1 17952
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_4.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 1564 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_3
timestamp 1586364061
transform 1 0 1380 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_7
timestamp 1586364061
transform 1 0 1748 0 1 17952
box -38 -48 222 592
use scs8hd_decap_8  FILLER_29_12
timestamp 1586364061
transform 1 0 2208 0 1 17952
box -38 -48 774 592
use scs8hd_nor2_4  _071_
timestamp 1586364061
transform 1 0 3312 0 1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__071__B
timestamp 1586364061
transform 1 0 3128 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_20
timestamp 1586364061
transform 1 0 2944 0 1 17952
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_ipin_4.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 4876 0 1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_4.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 4692 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_4.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 4324 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_33
timestamp 1586364061
transform 1 0 4140 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_37
timestamp 1586364061
transform 1 0 4508 0 1 17952
box -38 -48 222 592
use scs8hd_decap_8  FILLER_29_50
timestamp 1586364061
transform 1 0 5704 0 1 17952
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_177
timestamp 1586364061
transform 1 0 6716 0 1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__073__B
timestamp 1586364061
transform 1 0 6992 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__073__A
timestamp 1586364061
transform 1 0 7360 0 1 17952
box -38 -48 222 592
use scs8hd_decap_3  FILLER_29_58
timestamp 1586364061
transform 1 0 6440 0 1 17952
box -38 -48 314 592
use scs8hd_fill_2  FILLER_29_62
timestamp 1586364061
transform 1 0 6808 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_66
timestamp 1586364061
transform 1 0 7176 0 1 17952
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_ipin_4.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 8188 0 1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_4.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 8004 0 1 17952
box -38 -48 222 592
use scs8hd_decap_4  FILLER_29_70
timestamp 1586364061
transform 1 0 7544 0 1 17952
box -38 -48 406 592
use scs8hd_fill_1  FILLER_29_74
timestamp 1586364061
transform 1 0 7912 0 1 17952
box -38 -48 130 592
use scs8hd_nor2_4  _100_
timestamp 1586364061
transform 1 0 9752 0 1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_0.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 9568 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__100__B
timestamp 1586364061
transform 1 0 9200 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_86
timestamp 1586364061
transform 1 0 9016 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_90
timestamp 1586364061
transform 1 0 9384 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_0.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 10764 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_103
timestamp 1586364061
transform 1 0 10580 0 1 17952
box -38 -48 222 592
use scs8hd_decap_4  FILLER_29_107
timestamp 1586364061
transform 1 0 10948 0 1 17952
box -38 -48 406 592
use scs8hd_ebufn_2  mux_top_ipin_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12420 0 1 17952
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_178
timestamp 1586364061
transform 1 0 12328 0 1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_0.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 11408 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 12144 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_0.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 11776 0 1 17952
box -38 -48 222 592
use scs8hd_fill_1  FILLER_29_111
timestamp 1586364061
transform 1 0 11316 0 1 17952
box -38 -48 130 592
use scs8hd_fill_2  FILLER_29_114
timestamp 1586364061
transform 1 0 11592 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_118
timestamp 1586364061
transform 1 0 11960 0 1 17952
box -38 -48 222 592
use scs8hd_decap_8  FILLER_29_132
timestamp 1586364061
transform 1 0 13248 0 1 17952
box -38 -48 774 592
use scs8hd_inv_1  mux_bottom_ipin_2.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 14168 0 1 17952
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 15088 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 14628 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_140
timestamp 1586364061
transform 1 0 13984 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_145
timestamp 1586364061
transform 1 0 14444 0 1 17952
box -38 -48 222 592
use scs8hd_decap_3  FILLER_29_149
timestamp 1586364061
transform 1 0 14812 0 1 17952
box -38 -48 314 592
use scs8hd_ebufn_2  mux_bottom_ipin_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15272 0 1 17952
box -38 -48 866 592
use scs8hd_decap_4  FILLER_29_163
timestamp 1586364061
transform 1 0 16100 0 1 17952
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__127__B
timestamp 1586364061
transform 1 0 16560 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__127__A
timestamp 1586364061
transform 1 0 16928 0 1 17952
box -38 -48 222 592
use scs8hd_fill_1  FILLER_29_167
timestamp 1586364061
transform 1 0 16468 0 1 17952
box -38 -48 130 592
use scs8hd_fill_2  FILLER_29_170
timestamp 1586364061
transform 1 0 16744 0 1 17952
box -38 -48 222 592
use scs8hd_decap_8  FILLER_29_174
timestamp 1586364061
transform 1 0 17112 0 1 17952
box -38 -48 774 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_2.LATCH_5_.latch
timestamp 1586364061
transform 1 0 18768 0 1 17952
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_179
timestamp 1586364061
transform 1 0 17940 0 1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_2.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 18584 0 1 17952
box -38 -48 222 592
use scs8hd_fill_1  FILLER_29_182
timestamp 1586364061
transform 1 0 17848 0 1 17952
box -38 -48 130 592
use scs8hd_decap_6  FILLER_29_184
timestamp 1586364061
transform 1 0 18032 0 1 17952
box -38 -48 590 592
use scs8hd_decap_6  FILLER_29_203
timestamp 1586364061
transform 1 0 19780 0 1 17952
box -38 -48 590 592
use scs8hd_ebufn_2  mux_bottom_ipin_2.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 20516 0 1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 20332 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_220
timestamp 1586364061
transform 1 0 21344 0 1 17952
box -38 -48 222 592
use scs8hd_decap_3  PHY_59
timestamp 1586364061
transform -1 0 22816 0 1 17952
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__152__A
timestamp 1586364061
transform 1 0 21528 0 1 17952
box -38 -48 222 592
use scs8hd_decap_8  FILLER_29_224
timestamp 1586364061
transform 1 0 21712 0 1 17952
box -38 -48 774 592
use scs8hd_fill_1  FILLER_29_232
timestamp 1586364061
transform 1 0 22448 0 1 17952
box -38 -48 130 592
use scs8hd_inv_1  mux_bottom_ipin_4.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1380 0 -1 19040
box -38 -48 314 592
use scs8hd_decap_3  PHY_60
timestamp 1586364061
transform 1 0 1104 0 -1 19040
box -38 -48 314 592
use scs8hd_decap_12  FILLER_30_6
timestamp 1586364061
transform 1 0 1656 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_18
timestamp 1586364061
transform 1 0 2760 0 -1 19040
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_180
timestamp 1586364061
transform 1 0 3956 0 -1 19040
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_4.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 4876 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_1  FILLER_30_30
timestamp 1586364061
transform 1 0 3864 0 -1 19040
box -38 -48 130 592
use scs8hd_decap_8  FILLER_30_32
timestamp 1586364061
transform 1 0 4048 0 -1 19040
box -38 -48 774 592
use scs8hd_fill_1  FILLER_30_40
timestamp 1586364061
transform 1 0 4784 0 -1 19040
box -38 -48 130 592
use scs8hd_decap_12  FILLER_30_43
timestamp 1586364061
transform 1 0 5060 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_30_55
timestamp 1586364061
transform 1 0 6164 0 -1 19040
box -38 -48 406 592
use scs8hd_nor2_4  _073_
timestamp 1586364061
transform 1 0 6624 0 -1 19040
box -38 -48 866 592
use scs8hd_fill_1  FILLER_30_59
timestamp 1586364061
transform 1 0 6532 0 -1 19040
box -38 -48 130 592
use scs8hd_decap_8  FILLER_30_69
timestamp 1586364061
transform 1 0 7452 0 -1 19040
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_4.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 8188 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_12  FILLER_30_79
timestamp 1586364061
transform 1 0 8372 0 -1 19040
box -38 -48 1142 592
use scs8hd_lpflow_inputisolatch_1  mem_top_ipin_0.LATCH_5_.latch
timestamp 1586364061
transform 1 0 9660 0 -1 19040
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_181
timestamp 1586364061
transform 1 0 9568 0 -1 19040
box -38 -48 130 592
use scs8hd_fill_1  FILLER_30_91
timestamp 1586364061
transform 1 0 9476 0 -1 19040
box -38 -48 130 592
use scs8hd_decap_8  FILLER_30_104
timestamp 1586364061
transform 1 0 10672 0 -1 19040
box -38 -48 774 592
use scs8hd_lpflow_inputisolatch_1  mem_top_ipin_0.LATCH_3_.latch
timestamp 1586364061
transform 1 0 11408 0 -1 19040
box -38 -48 1050 592
use scs8hd_fill_2  FILLER_30_123
timestamp 1586364061
transform 1 0 12420 0 -1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 12604 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_12  FILLER_30_127
timestamp 1586364061
transform 1 0 12788 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_139
timestamp 1586364061
transform 1 0 13892 0 -1 19040
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_30_151
timestamp 1586364061
transform 1 0 14996 0 -1 19040
box -38 -48 222 592
use scs8hd_inv_1  mux_bottom_ipin_2.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 15272 0 -1 19040
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_182
timestamp 1586364061
transform 1 0 15180 0 -1 19040
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 15732 0 -1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 16100 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_157
timestamp 1586364061
transform 1 0 15548 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_161
timestamp 1586364061
transform 1 0 15916 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_3  FILLER_30_165
timestamp 1586364061
transform 1 0 16284 0 -1 19040
box -38 -48 314 592
use scs8hd_nor2_4  _127_
timestamp 1586364061
transform 1 0 16560 0 -1 19040
box -38 -48 866 592
use scs8hd_decap_12  FILLER_30_177
timestamp 1586364061
transform 1 0 17388 0 -1 19040
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_2.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 18768 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_3  FILLER_30_189
timestamp 1586364061
transform 1 0 18492 0 -1 19040
box -38 -48 314 592
use scs8hd_conb_1  _133_
timestamp 1586364061
transform 1 0 19412 0 -1 19040
box -38 -48 314 592
use scs8hd_decap_4  FILLER_30_194
timestamp 1586364061
transform 1 0 18952 0 -1 19040
box -38 -48 406 592
use scs8hd_fill_1  FILLER_30_198
timestamp 1586364061
transform 1 0 19320 0 -1 19040
box -38 -48 130 592
use scs8hd_decap_12  FILLER_30_202
timestamp 1586364061
transform 1 0 19688 0 -1 19040
box -38 -48 1142 592
use scs8hd_buf_2  _152_
timestamp 1586364061
transform 1 0 20884 0 -1 19040
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_183
timestamp 1586364061
transform 1 0 20792 0 -1 19040
box -38 -48 130 592
use scs8hd_decap_12  FILLER_30_219
timestamp 1586364061
transform 1 0 21252 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_3  PHY_61
timestamp 1586364061
transform -1 0 22816 0 -1 19040
box -38 -48 314 592
use scs8hd_fill_2  FILLER_30_231
timestamp 1586364061
transform 1 0 22356 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_3  PHY_62
timestamp 1586364061
transform 1 0 1104 0 1 19040
box -38 -48 314 592
use scs8hd_decap_12  FILLER_31_3
timestamp 1586364061
transform 1 0 1380 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_15
timestamp 1586364061
transform 1 0 2484 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_27
timestamp 1586364061
transform 1 0 3588 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_39
timestamp 1586364061
transform 1 0 4692 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_31_51
timestamp 1586364061
transform 1 0 5796 0 1 19040
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_184
timestamp 1586364061
transform 1 0 6716 0 1 19040
box -38 -48 130 592
use scs8hd_fill_2  FILLER_31_59
timestamp 1586364061
transform 1 0 6532 0 1 19040
box -38 -48 222 592
use scs8hd_decap_12  FILLER_31_62
timestamp 1586364061
transform 1 0 6808 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_31_74
timestamp 1586364061
transform 1 0 7912 0 1 19040
box -38 -48 774 592
use scs8hd_fill_2  FILLER_31_82
timestamp 1586364061
transform 1 0 8648 0 1 19040
box -38 -48 222 592
use scs8hd_conb_1  _139_
timestamp 1586364061
transform 1 0 8832 0 1 19040
box -38 -48 314 592
use scs8hd_ebufn_2  mux_top_ipin_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9844 0 1 19040
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9660 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 9292 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_87
timestamp 1586364061
transform 1 0 9108 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_91
timestamp 1586364061
transform 1 0 9476 0 1 19040
box -38 -48 222 592
use scs8hd_decap_12  FILLER_31_104
timestamp 1586364061
transform 1 0 10672 0 1 19040
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_185
timestamp 1586364061
transform 1 0 12328 0 1 19040
box -38 -48 130 592
use scs8hd_decap_6  FILLER_31_116
timestamp 1586364061
transform 1 0 11776 0 1 19040
box -38 -48 590 592
use scs8hd_decap_12  FILLER_31_123
timestamp 1586364061
transform 1 0 12420 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_135
timestamp 1586364061
transform 1 0 13524 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_147
timestamp 1586364061
transform 1 0 14628 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_159
timestamp 1586364061
transform 1 0 15732 0 1 19040
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA__156__A
timestamp 1586364061
transform 1 0 17112 0 1 19040
box -38 -48 222 592
use scs8hd_decap_3  FILLER_31_171
timestamp 1586364061
transform 1 0 16836 0 1 19040
box -38 -48 314 592
use scs8hd_decap_6  FILLER_31_176
timestamp 1586364061
transform 1 0 17296 0 1 19040
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_186
timestamp 1586364061
transform 1 0 17940 0 1 19040
box -38 -48 130 592
use scs8hd_fill_1  FILLER_31_182
timestamp 1586364061
transform 1 0 17848 0 1 19040
box -38 -48 130 592
use scs8hd_decap_12  FILLER_31_184
timestamp 1586364061
transform 1 0 18032 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_196
timestamp 1586364061
transform 1 0 19136 0 1 19040
box -38 -48 1142 592
use scs8hd_inv_1  mux_bottom_ipin_2.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 20884 0 1 19040
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 21344 0 1 19040
box -38 -48 222 592
use scs8hd_decap_6  FILLER_31_208
timestamp 1586364061
transform 1 0 20240 0 1 19040
box -38 -48 590 592
use scs8hd_fill_1  FILLER_31_214
timestamp 1586364061
transform 1 0 20792 0 1 19040
box -38 -48 130 592
use scs8hd_fill_2  FILLER_31_218
timestamp 1586364061
transform 1 0 21160 0 1 19040
box -38 -48 222 592
use scs8hd_decap_3  PHY_63
timestamp 1586364061
transform -1 0 22816 0 1 19040
box -38 -48 314 592
use scs8hd_decap_8  FILLER_31_222
timestamp 1586364061
transform 1 0 21528 0 1 19040
box -38 -48 774 592
use scs8hd_decap_3  FILLER_31_230
timestamp 1586364061
transform 1 0 22264 0 1 19040
box -38 -48 314 592
use scs8hd_decap_3  PHY_64
timestamp 1586364061
transform 1 0 1104 0 -1 20128
box -38 -48 314 592
use scs8hd_decap_12  FILLER_32_3
timestamp 1586364061
transform 1 0 1380 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_15
timestamp 1586364061
transform 1 0 2484 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_32_27
timestamp 1586364061
transform 1 0 3588 0 -1 20128
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_187
timestamp 1586364061
transform 1 0 3956 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_12  FILLER_32_32
timestamp 1586364061
transform 1 0 4048 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_44
timestamp 1586364061
transform 1 0 5152 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_56
timestamp 1586364061
transform 1 0 6256 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_68
timestamp 1586364061
transform 1 0 7360 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_80
timestamp 1586364061
transform 1 0 8464 0 -1 20128
box -38 -48 1142 592
use scs8hd_inv_1  mux_top_ipin_0.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 9660 0 -1 20128
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_188
timestamp 1586364061
transform 1 0 9568 0 -1 20128
box -38 -48 130 592
use scs8hd_fill_2  FILLER_32_96
timestamp 1586364061
transform 1 0 9936 0 -1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 10120 0 -1 20128
box -38 -48 222 592
use scs8hd_decap_12  FILLER_32_100
timestamp 1586364061
transform 1 0 10304 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_112
timestamp 1586364061
transform 1 0 11408 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_124
timestamp 1586364061
transform 1 0 12512 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_136
timestamp 1586364061
transform 1 0 13616 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_32_148
timestamp 1586364061
transform 1 0 14720 0 -1 20128
box -38 -48 406 592
use scs8hd_fill_1  FILLER_32_152
timestamp 1586364061
transform 1 0 15088 0 -1 20128
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_189
timestamp 1586364061
transform 1 0 15180 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_12  FILLER_32_154
timestamp 1586364061
transform 1 0 15272 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_32_166
timestamp 1586364061
transform 1 0 16376 0 -1 20128
box -38 -48 774 592
use scs8hd_buf_2  _156_
timestamp 1586364061
transform 1 0 17112 0 -1 20128
box -38 -48 406 592
use scs8hd_decap_12  FILLER_32_178
timestamp 1586364061
transform 1 0 17480 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_190
timestamp 1586364061
transform 1 0 18584 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_202
timestamp 1586364061
transform 1 0 19688 0 -1 20128
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_190
timestamp 1586364061
transform 1 0 20792 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_12  FILLER_32_215
timestamp 1586364061
transform 1 0 20884 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_3  PHY_65
timestamp 1586364061
transform -1 0 22816 0 -1 20128
box -38 -48 314 592
use scs8hd_decap_6  FILLER_32_227
timestamp 1586364061
transform 1 0 21988 0 -1 20128
box -38 -48 590 592
use scs8hd_inv_1  mux_bottom_ipin_6.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1380 0 1 20128
box -38 -48 314 592
use scs8hd_decap_3  PHY_66
timestamp 1586364061
transform 1 0 1104 0 1 20128
box -38 -48 314 592
use scs8hd_decap_3  PHY_68
timestamp 1586364061
transform 1 0 1104 0 -1 21216
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_6.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 1840 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_6
timestamp 1586364061
transform 1 0 1656 0 1 20128
box -38 -48 222 592
use scs8hd_decap_12  FILLER_33_10
timestamp 1586364061
transform 1 0 2024 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_3
timestamp 1586364061
transform 1 0 1380 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_22
timestamp 1586364061
transform 1 0 3128 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_15
timestamp 1586364061
transform 1 0 2484 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_34_27
timestamp 1586364061
transform 1 0 3588 0 -1 21216
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_194
timestamp 1586364061
transform 1 0 3956 0 -1 21216
box -38 -48 130 592
use scs8hd_decap_12  FILLER_33_34
timestamp 1586364061
transform 1 0 4232 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_32
timestamp 1586364061
transform 1 0 4048 0 -1 21216
box -38 -48 1142 592
use scs8hd_buf_2  _150_
timestamp 1586364061
transform 1 0 5612 0 1 20128
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__150__A
timestamp 1586364061
transform 1 0 6164 0 1 20128
box -38 -48 222 592
use scs8hd_decap_3  FILLER_33_46
timestamp 1586364061
transform 1 0 5336 0 1 20128
box -38 -48 314 592
use scs8hd_fill_2  FILLER_33_53
timestamp 1586364061
transform 1 0 5980 0 1 20128
box -38 -48 222 592
use scs8hd_decap_12  FILLER_34_44
timestamp 1586364061
transform 1 0 5152 0 -1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_191
timestamp 1586364061
transform 1 0 6716 0 1 20128
box -38 -48 130 592
use scs8hd_decap_4  FILLER_33_57
timestamp 1586364061
transform 1 0 6348 0 1 20128
box -38 -48 406 592
use scs8hd_decap_12  FILLER_33_62
timestamp 1586364061
transform 1 0 6808 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_56
timestamp 1586364061
transform 1 0 6256 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_68
timestamp 1586364061
transform 1 0 7360 0 -1 21216
box -38 -48 1142 592
use scs8hd_buf_2  _149_
timestamp 1586364061
transform 1 0 7912 0 1 20128
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__149__A
timestamp 1586364061
transform 1 0 8464 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_78
timestamp 1586364061
transform 1 0 8280 0 1 20128
box -38 -48 222 592
use scs8hd_decap_12  FILLER_33_82
timestamp 1586364061
transform 1 0 8648 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_80
timestamp 1586364061
transform 1 0 8464 0 -1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_195
timestamp 1586364061
transform 1 0 9568 0 -1 21216
box -38 -48 130 592
use scs8hd_decap_8  FILLER_33_94
timestamp 1586364061
transform 1 0 9752 0 1 20128
box -38 -48 774 592
use scs8hd_decap_12  FILLER_34_93
timestamp 1586364061
transform 1 0 9660 0 -1 21216
box -38 -48 1142 592
use scs8hd_buf_2  _144_
timestamp 1586364061
transform 1 0 10672 0 1 20128
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__144__A
timestamp 1586364061
transform 1 0 11224 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_102
timestamp 1586364061
transform 1 0 10488 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_108
timestamp 1586364061
transform 1 0 11040 0 1 20128
box -38 -48 222 592
use scs8hd_decap_12  FILLER_34_105
timestamp 1586364061
transform 1 0 10764 0 -1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_192
timestamp 1586364061
transform 1 0 12328 0 1 20128
box -38 -48 130 592
use scs8hd_decap_8  FILLER_33_112
timestamp 1586364061
transform 1 0 11408 0 1 20128
box -38 -48 774 592
use scs8hd_fill_2  FILLER_33_120
timestamp 1586364061
transform 1 0 12144 0 1 20128
box -38 -48 222 592
use scs8hd_decap_12  FILLER_33_123
timestamp 1586364061
transform 1 0 12420 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_117
timestamp 1586364061
transform 1 0 11868 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_135
timestamp 1586364061
transform 1 0 13524 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_129
timestamp 1586364061
transform 1 0 12972 0 -1 21216
box -38 -48 1142 592
use scs8hd_buf_2  _159_
timestamp 1586364061
transform 1 0 15088 0 1 20128
box -38 -48 406 592
use scs8hd_decap_4  FILLER_33_147
timestamp 1586364061
transform 1 0 14628 0 1 20128
box -38 -48 406 592
use scs8hd_fill_1  FILLER_33_151
timestamp 1586364061
transform 1 0 14996 0 1 20128
box -38 -48 130 592
use scs8hd_decap_12  FILLER_34_141
timestamp 1586364061
transform 1 0 14076 0 -1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_196
timestamp 1586364061
transform 1 0 15180 0 -1 21216
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__159__A
timestamp 1586364061
transform 1 0 15640 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_156
timestamp 1586364061
transform 1 0 15456 0 1 20128
box -38 -48 222 592
use scs8hd_decap_12  FILLER_33_160
timestamp 1586364061
transform 1 0 15824 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_154
timestamp 1586364061
transform 1 0 15272 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_166
timestamp 1586364061
transform 1 0 16376 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_33_172
timestamp 1586364061
transform 1 0 16928 0 1 20128
box -38 -48 774 592
use scs8hd_decap_12  FILLER_34_178
timestamp 1586364061
transform 1 0 17480 0 -1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_193
timestamp 1586364061
transform 1 0 17940 0 1 20128
box -38 -48 130 592
use scs8hd_decap_3  FILLER_33_180
timestamp 1586364061
transform 1 0 17664 0 1 20128
box -38 -48 314 592
use scs8hd_decap_12  FILLER_33_184
timestamp 1586364061
transform 1 0 18032 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_190
timestamp 1586364061
transform 1 0 18584 0 -1 21216
box -38 -48 1142 592
use scs8hd_buf_2  _154_
timestamp 1586364061
transform 1 0 19228 0 1 20128
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__154__A
timestamp 1586364061
transform 1 0 19780 0 1 20128
box -38 -48 222 592
use scs8hd_fill_1  FILLER_33_196
timestamp 1586364061
transform 1 0 19136 0 1 20128
box -38 -48 130 592
use scs8hd_fill_2  FILLER_33_201
timestamp 1586364061
transform 1 0 19596 0 1 20128
box -38 -48 222 592
use scs8hd_decap_12  FILLER_33_205
timestamp 1586364061
transform 1 0 19964 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_202
timestamp 1586364061
transform 1 0 19688 0 -1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_197
timestamp 1586364061
transform 1 0 20792 0 -1 21216
box -38 -48 130 592
use scs8hd_decap_12  FILLER_33_217
timestamp 1586364061
transform 1 0 21068 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_215
timestamp 1586364061
transform 1 0 20884 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_3  PHY_67
timestamp 1586364061
transform -1 0 22816 0 1 20128
box -38 -48 314 592
use scs8hd_decap_3  PHY_69
timestamp 1586364061
transform -1 0 22816 0 -1 21216
box -38 -48 314 592
use scs8hd_decap_4  FILLER_33_229
timestamp 1586364061
transform 1 0 22172 0 1 20128
box -38 -48 406 592
use scs8hd_decap_6  FILLER_34_227
timestamp 1586364061
transform 1 0 21988 0 -1 21216
box -38 -48 590 592
use scs8hd_decap_3  PHY_70
timestamp 1586364061
transform 1 0 1104 0 1 21216
box -38 -48 314 592
use scs8hd_decap_12  FILLER_35_3
timestamp 1586364061
transform 1 0 1380 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_15
timestamp 1586364061
transform 1 0 2484 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_35_27
timestamp 1586364061
transform 1 0 3588 0 1 21216
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_198
timestamp 1586364061
transform 1 0 3956 0 1 21216
box -38 -48 130 592
use scs8hd_decap_12  FILLER_35_32
timestamp 1586364061
transform 1 0 4048 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_44
timestamp 1586364061
transform 1 0 5152 0 1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_199
timestamp 1586364061
transform 1 0 6808 0 1 21216
box -38 -48 130 592
use scs8hd_decap_6  FILLER_35_56
timestamp 1586364061
transform 1 0 6256 0 1 21216
box -38 -48 590 592
use scs8hd_decap_12  FILLER_35_63
timestamp 1586364061
transform 1 0 6900 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_75
timestamp 1586364061
transform 1 0 8004 0 1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_200
timestamp 1586364061
transform 1 0 9660 0 1 21216
box -38 -48 130 592
use scs8hd_decap_6  FILLER_35_87
timestamp 1586364061
transform 1 0 9108 0 1 21216
box -38 -48 590 592
use scs8hd_decap_12  FILLER_35_94
timestamp 1586364061
transform 1 0 9752 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_106
timestamp 1586364061
transform 1 0 10856 0 1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_201
timestamp 1586364061
transform 1 0 12512 0 1 21216
box -38 -48 130 592
use scs8hd_decap_6  FILLER_35_118
timestamp 1586364061
transform 1 0 11960 0 1 21216
box -38 -48 590 592
use scs8hd_decap_12  FILLER_35_125
timestamp 1586364061
transform 1 0 12604 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_137
timestamp 1586364061
transform 1 0 13708 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_35_149
timestamp 1586364061
transform 1 0 14812 0 1 21216
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_202
timestamp 1586364061
transform 1 0 15364 0 1 21216
box -38 -48 130 592
use scs8hd_decap_12  FILLER_35_156
timestamp 1586364061
transform 1 0 15456 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_168
timestamp 1586364061
transform 1 0 16560 0 1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_203
timestamp 1586364061
transform 1 0 18216 0 1 21216
box -38 -48 130 592
use scs8hd_decap_6  FILLER_35_180
timestamp 1586364061
transform 1 0 17664 0 1 21216
box -38 -48 590 592
use scs8hd_decap_12  FILLER_35_187
timestamp 1586364061
transform 1 0 18308 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_199
timestamp 1586364061
transform 1 0 19412 0 1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_204
timestamp 1586364061
transform 1 0 21068 0 1 21216
box -38 -48 130 592
use scs8hd_decap_6  FILLER_35_211
timestamp 1586364061
transform 1 0 20516 0 1 21216
box -38 -48 590 592
use scs8hd_decap_12  FILLER_35_218
timestamp 1586364061
transform 1 0 21160 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_3  PHY_71
timestamp 1586364061
transform -1 0 22816 0 1 21216
box -38 -48 314 592
use scs8hd_decap_3  FILLER_35_230
timestamp 1586364061
transform 1 0 22264 0 1 21216
box -38 -48 314 592
<< labels >>
rlabel metal2 s 4618 0 4674 480 6 address[0]
port 0 nsew default input
rlabel metal3 s 0 688 480 808 6 address[1]
port 1 nsew default input
rlabel metal3 s 23520 688 24000 808 6 address[2]
port 2 nsew default input
rlabel metal3 s 23520 2184 24000 2304 6 address[3]
port 3 nsew default input
rlabel metal3 s 0 2184 480 2304 6 address[4]
port 4 nsew default input
rlabel metal3 s 23520 3680 24000 3800 6 address[5]
port 5 nsew default input
rlabel metal3 s 0 3816 480 3936 6 address[6]
port 6 nsew default input
rlabel metal2 s 938 23520 994 24000 6 bottom_grid_pin_0_
port 7 nsew default tristate
rlabel metal3 s 23520 5176 24000 5296 6 bottom_grid_pin_4_
port 8 nsew default tristate
rlabel metal3 s 0 5448 480 5568 6 bottom_grid_pin_8_
port 9 nsew default tristate
rlabel metal2 s 6458 0 6514 480 6 chanx_left_in[0]
port 10 nsew default input
rlabel metal2 s 2870 23520 2926 24000 6 chanx_left_in[1]
port 11 nsew default input
rlabel metal2 s 8298 0 8354 480 6 chanx_left_in[2]
port 12 nsew default input
rlabel metal2 s 10138 0 10194 480 6 chanx_left_in[3]
port 13 nsew default input
rlabel metal2 s 4894 23520 4950 24000 6 chanx_left_in[4]
port 14 nsew default input
rlabel metal3 s 0 6944 480 7064 6 chanx_left_in[5]
port 15 nsew default input
rlabel metal3 s 23520 6672 24000 6792 6 chanx_left_in[6]
port 16 nsew default input
rlabel metal3 s 0 8576 480 8696 6 chanx_left_in[7]
port 17 nsew default input
rlabel metal3 s 23520 8168 24000 8288 6 chanx_left_in[8]
port 18 nsew default input
rlabel metal2 s 6918 23520 6974 24000 6 chanx_left_out[0]
port 19 nsew default tristate
rlabel metal2 s 8942 23520 8998 24000 6 chanx_left_out[1]
port 20 nsew default tristate
rlabel metal3 s 23520 9664 24000 9784 6 chanx_left_out[2]
port 21 nsew default tristate
rlabel metal2 s 11978 0 12034 480 6 chanx_left_out[3]
port 22 nsew default tristate
rlabel metal3 s 0 10208 480 10328 6 chanx_left_out[4]
port 23 nsew default tristate
rlabel metal2 s 13818 0 13874 480 6 chanx_left_out[5]
port 24 nsew default tristate
rlabel metal2 s 10874 23520 10930 24000 6 chanx_left_out[6]
port 25 nsew default tristate
rlabel metal3 s 23520 11160 24000 11280 6 chanx_left_out[7]
port 26 nsew default tristate
rlabel metal3 s 23520 12656 24000 12776 6 chanx_left_out[8]
port 27 nsew default tristate
rlabel metal3 s 0 11840 480 11960 6 chanx_right_in[0]
port 28 nsew default input
rlabel metal3 s 0 13336 480 13456 6 chanx_right_in[1]
port 29 nsew default input
rlabel metal3 s 23520 14152 24000 14272 6 chanx_right_in[2]
port 30 nsew default input
rlabel metal2 s 12898 23520 12954 24000 6 chanx_right_in[3]
port 31 nsew default input
rlabel metal2 s 14922 23520 14978 24000 6 chanx_right_in[4]
port 32 nsew default input
rlabel metal2 s 15658 0 15714 480 6 chanx_right_in[5]
port 33 nsew default input
rlabel metal2 s 17498 0 17554 480 6 chanx_right_in[6]
port 34 nsew default input
rlabel metal3 s 0 14968 480 15088 6 chanx_right_in[7]
port 35 nsew default input
rlabel metal3 s 23520 15648 24000 15768 6 chanx_right_in[8]
port 36 nsew default input
rlabel metal2 s 16946 23520 17002 24000 6 chanx_right_out[0]
port 37 nsew default tristate
rlabel metal3 s 23520 17144 24000 17264 6 chanx_right_out[1]
port 38 nsew default tristate
rlabel metal2 s 19338 0 19394 480 6 chanx_right_out[2]
port 39 nsew default tristate
rlabel metal2 s 18878 23520 18934 24000 6 chanx_right_out[3]
port 40 nsew default tristate
rlabel metal2 s 21178 0 21234 480 6 chanx_right_out[4]
port 41 nsew default tristate
rlabel metal2 s 20902 23520 20958 24000 6 chanx_right_out[5]
port 42 nsew default tristate
rlabel metal3 s 23520 18640 24000 18760 6 chanx_right_out[6]
port 43 nsew default tristate
rlabel metal3 s 23520 20136 24000 20256 6 chanx_right_out[7]
port 44 nsew default tristate
rlabel metal3 s 0 16600 480 16720 6 chanx_right_out[8]
port 45 nsew default tristate
rlabel metal2 s 2778 0 2834 480 6 data_in
port 46 nsew default input
rlabel metal2 s 938 0 994 480 6 enable
port 47 nsew default input
rlabel metal3 s 0 18232 480 18352 6 top_grid_pin_0_
port 48 nsew default tristate
rlabel metal3 s 0 21360 480 21480 6 top_grid_pin_10_
port 49 nsew default tristate
rlabel metal3 s 0 22992 480 23112 6 top_grid_pin_12_
port 50 nsew default tristate
rlabel metal3 s 23520 23128 24000 23248 6 top_grid_pin_14_
port 51 nsew default tristate
rlabel metal2 s 23018 0 23074 480 6 top_grid_pin_2_
port 52 nsew default tristate
rlabel metal2 s 22926 23520 22982 24000 6 top_grid_pin_4_
port 53 nsew default tristate
rlabel metal3 s 23520 21632 24000 21752 6 top_grid_pin_6_
port 54 nsew default tristate
rlabel metal3 s 0 19728 480 19848 6 top_grid_pin_8_
port 55 nsew default tristate
rlabel metal4 s 4944 2128 5264 21808 6 vpwr
port 56 nsew default input
rlabel metal4 s 8944 2128 9264 21808 6 vgnd
port 57 nsew default input
<< end >>
