VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO cby_1__1_
  CLASS BLOCK ;
  FOREIGN cby_1__1_ ;
  ORIGIN 0.000 0.000 ;
  SIZE 80.000 BY 200.000 ;
  PIN ccff_head
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 78.750 197.600 79.030 200.000 ;
    END
  END ccff_head
  PIN ccff_tail
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 193.160 2.400 193.760 ;
    END
  END ccff_tail
  PIN chany_bottom_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1.010 0.000 1.290 2.400 ;
    END
  END chany_bottom_in[0]
  PIN chany_bottom_in[10]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 20.790 0.000 21.070 2.400 ;
    END
  END chany_bottom_in[10]
  PIN chany_bottom_in[11]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 22.630 0.000 22.910 2.400 ;
    END
  END chany_bottom_in[11]
  PIN chany_bottom_in[12]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 24.930 0.000 25.210 2.400 ;
    END
  END chany_bottom_in[12]
  PIN chany_bottom_in[13]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 26.770 0.000 27.050 2.400 ;
    END
  END chany_bottom_in[13]
  PIN chany_bottom_in[14]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 28.610 0.000 28.890 2.400 ;
    END
  END chany_bottom_in[14]
  PIN chany_bottom_in[15]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 30.910 0.000 31.190 2.400 ;
    END
  END chany_bottom_in[15]
  PIN chany_bottom_in[16]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 32.750 0.000 33.030 2.400 ;
    END
  END chany_bottom_in[16]
  PIN chany_bottom_in[17]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 34.590 0.000 34.870 2.400 ;
    END
  END chany_bottom_in[17]
  PIN chany_bottom_in[18]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 36.890 0.000 37.170 2.400 ;
    END
  END chany_bottom_in[18]
  PIN chany_bottom_in[19]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 38.730 0.000 39.010 2.400 ;
    END
  END chany_bottom_in[19]
  PIN chany_bottom_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2.850 0.000 3.130 2.400 ;
    END
  END chany_bottom_in[1]
  PIN chany_bottom_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 4.690 0.000 4.970 2.400 ;
    END
  END chany_bottom_in[2]
  PIN chany_bottom_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 6.990 0.000 7.270 2.400 ;
    END
  END chany_bottom_in[3]
  PIN chany_bottom_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 8.830 0.000 9.110 2.400 ;
    END
  END chany_bottom_in[4]
  PIN chany_bottom_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 10.670 0.000 10.950 2.400 ;
    END
  END chany_bottom_in[5]
  PIN chany_bottom_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 12.970 0.000 13.250 2.400 ;
    END
  END chany_bottom_in[6]
  PIN chany_bottom_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 14.810 0.000 15.090 2.400 ;
    END
  END chany_bottom_in[7]
  PIN chany_bottom_in[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 16.650 0.000 16.930 2.400 ;
    END
  END chany_bottom_in[8]
  PIN chany_bottom_in[9]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 18.950 0.000 19.230 2.400 ;
    END
  END chany_bottom_in[9]
  PIN chany_bottom_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 41.030 0.000 41.310 2.400 ;
    END
  END chany_bottom_out[0]
  PIN chany_bottom_out[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 60.810 0.000 61.090 2.400 ;
    END
  END chany_bottom_out[10]
  PIN chany_bottom_out[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 62.650 0.000 62.930 2.400 ;
    END
  END chany_bottom_out[11]
  PIN chany_bottom_out[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 64.950 0.000 65.230 2.400 ;
    END
  END chany_bottom_out[12]
  PIN chany_bottom_out[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 66.790 0.000 67.070 2.400 ;
    END
  END chany_bottom_out[13]
  PIN chany_bottom_out[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 68.630 0.000 68.910 2.400 ;
    END
  END chany_bottom_out[14]
  PIN chany_bottom_out[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 70.930 0.000 71.210 2.400 ;
    END
  END chany_bottom_out[15]
  PIN chany_bottom_out[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 72.770 0.000 73.050 2.400 ;
    END
  END chany_bottom_out[16]
  PIN chany_bottom_out[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 74.610 0.000 74.890 2.400 ;
    END
  END chany_bottom_out[17]
  PIN chany_bottom_out[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 76.910 0.000 77.190 2.400 ;
    END
  END chany_bottom_out[18]
  PIN chany_bottom_out[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 78.750 0.000 79.030 2.400 ;
    END
  END chany_bottom_out[19]
  PIN chany_bottom_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 42.870 0.000 43.150 2.400 ;
    END
  END chany_bottom_out[1]
  PIN chany_bottom_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 44.710 0.000 44.990 2.400 ;
    END
  END chany_bottom_out[2]
  PIN chany_bottom_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 47.010 0.000 47.290 2.400 ;
    END
  END chany_bottom_out[3]
  PIN chany_bottom_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 48.850 0.000 49.130 2.400 ;
    END
  END chany_bottom_out[4]
  PIN chany_bottom_out[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 50.690 0.000 50.970 2.400 ;
    END
  END chany_bottom_out[5]
  PIN chany_bottom_out[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 52.990 0.000 53.270 2.400 ;
    END
  END chany_bottom_out[6]
  PIN chany_bottom_out[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 54.830 0.000 55.110 2.400 ;
    END
  END chany_bottom_out[7]
  PIN chany_bottom_out[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 56.670 0.000 56.950 2.400 ;
    END
  END chany_bottom_out[8]
  PIN chany_bottom_out[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 58.970 0.000 59.250 2.400 ;
    END
  END chany_bottom_out[9]
  PIN chany_top_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1.010 197.600 1.290 200.000 ;
    END
  END chany_top_in[0]
  PIN chany_top_in[10]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 20.330 197.600 20.610 200.000 ;
    END
  END chany_top_in[10]
  PIN chany_top_in[11]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 22.170 197.600 22.450 200.000 ;
    END
  END chany_top_in[11]
  PIN chany_top_in[12]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 24.010 197.600 24.290 200.000 ;
    END
  END chany_top_in[12]
  PIN chany_top_in[13]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 26.310 197.600 26.590 200.000 ;
    END
  END chany_top_in[13]
  PIN chany_top_in[14]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 28.150 197.600 28.430 200.000 ;
    END
  END chany_top_in[14]
  PIN chany_top_in[15]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 29.990 197.600 30.270 200.000 ;
    END
  END chany_top_in[15]
  PIN chany_top_in[16]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 31.830 197.600 32.110 200.000 ;
    END
  END chany_top_in[16]
  PIN chany_top_in[17]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 34.130 197.600 34.410 200.000 ;
    END
  END chany_top_in[17]
  PIN chany_top_in[18]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 35.970 197.600 36.250 200.000 ;
    END
  END chany_top_in[18]
  PIN chany_top_in[19]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 37.810 197.600 38.090 200.000 ;
    END
  END chany_top_in[19]
  PIN chany_top_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2.850 197.600 3.130 200.000 ;
    END
  END chany_top_in[1]
  PIN chany_top_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 4.690 197.600 4.970 200.000 ;
    END
  END chany_top_in[2]
  PIN chany_top_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 6.530 197.600 6.810 200.000 ;
    END
  END chany_top_in[3]
  PIN chany_top_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 8.370 197.600 8.650 200.000 ;
    END
  END chany_top_in[4]
  PIN chany_top_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 10.670 197.600 10.950 200.000 ;
    END
  END chany_top_in[5]
  PIN chany_top_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 12.510 197.600 12.790 200.000 ;
    END
  END chany_top_in[6]
  PIN chany_top_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 14.350 197.600 14.630 200.000 ;
    END
  END chany_top_in[7]
  PIN chany_top_in[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 16.190 197.600 16.470 200.000 ;
    END
  END chany_top_in[8]
  PIN chany_top_in[9]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 18.490 197.600 18.770 200.000 ;
    END
  END chany_top_in[9]
  PIN chany_top_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 39.650 197.600 39.930 200.000 ;
    END
  END chany_top_out[0]
  PIN chany_top_out[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 59.430 197.600 59.710 200.000 ;
    END
  END chany_top_out[10]
  PIN chany_top_out[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 61.270 197.600 61.550 200.000 ;
    END
  END chany_top_out[11]
  PIN chany_top_out[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 63.110 197.600 63.390 200.000 ;
    END
  END chany_top_out[12]
  PIN chany_top_out[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 65.410 197.600 65.690 200.000 ;
    END
  END chany_top_out[13]
  PIN chany_top_out[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 67.250 197.600 67.530 200.000 ;
    END
  END chany_top_out[14]
  PIN chany_top_out[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 69.090 197.600 69.370 200.000 ;
    END
  END chany_top_out[15]
  PIN chany_top_out[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 70.930 197.600 71.210 200.000 ;
    END
  END chany_top_out[16]
  PIN chany_top_out[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 73.230 197.600 73.510 200.000 ;
    END
  END chany_top_out[17]
  PIN chany_top_out[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 75.070 197.600 75.350 200.000 ;
    END
  END chany_top_out[18]
  PIN chany_top_out[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 76.910 197.600 77.190 200.000 ;
    END
  END chany_top_out[19]
  PIN chany_top_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 41.950 197.600 42.230 200.000 ;
    END
  END chany_top_out[1]
  PIN chany_top_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 43.790 197.600 44.070 200.000 ;
    END
  END chany_top_out[2]
  PIN chany_top_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 45.630 197.600 45.910 200.000 ;
    END
  END chany_top_out[3]
  PIN chany_top_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 47.470 197.600 47.750 200.000 ;
    END
  END chany_top_out[4]
  PIN chany_top_out[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 49.770 197.600 50.050 200.000 ;
    END
  END chany_top_out[5]
  PIN chany_top_out[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 51.610 197.600 51.890 200.000 ;
    END
  END chany_top_out[6]
  PIN chany_top_out[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 53.450 197.600 53.730 200.000 ;
    END
  END chany_top_out[7]
  PIN chany_top_out[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 55.290 197.600 55.570 200.000 ;
    END
  END chany_top_out[8]
  PIN chany_top_out[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 57.590 197.600 57.870 200.000 ;
    END
  END chany_top_out[9]
  PIN left_grid_pin_0_
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 5.480 2.400 6.080 ;
    END
  END left_grid_pin_0_
  PIN left_grid_pin_10_
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 122.440 2.400 123.040 ;
    END
  END left_grid_pin_10_
  PIN left_grid_pin_11_
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 134.680 2.400 135.280 ;
    END
  END left_grid_pin_11_
  PIN left_grid_pin_12_
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 146.240 2.400 146.840 ;
    END
  END left_grid_pin_12_
  PIN left_grid_pin_13_
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 157.800 2.400 158.400 ;
    END
  END left_grid_pin_13_
  PIN left_grid_pin_14_
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 170.040 2.400 170.640 ;
    END
  END left_grid_pin_14_
  PIN left_grid_pin_15_
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 181.600 2.400 182.200 ;
    END
  END left_grid_pin_15_
  PIN left_grid_pin_1_
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 17.040 2.400 17.640 ;
    END
  END left_grid_pin_1_
  PIN left_grid_pin_2_
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 28.600 2.400 29.200 ;
    END
  END left_grid_pin_2_
  PIN left_grid_pin_3_
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 40.160 2.400 40.760 ;
    END
  END left_grid_pin_3_
  PIN left_grid_pin_4_
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 52.400 2.400 53.000 ;
    END
  END left_grid_pin_4_
  PIN left_grid_pin_5_
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 63.960 2.400 64.560 ;
    END
  END left_grid_pin_5_
  PIN left_grid_pin_6_
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 75.520 2.400 76.120 ;
    END
  END left_grid_pin_6_
  PIN left_grid_pin_7_
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 87.760 2.400 88.360 ;
    END
  END left_grid_pin_7_
  PIN left_grid_pin_8_
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 99.320 2.400 99.920 ;
    END
  END left_grid_pin_8_
  PIN left_grid_pin_9_
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 110.880 2.400 111.480 ;
    END
  END left_grid_pin_9_
  PIN prog_clk
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 77.600 149.640 80.000 150.240 ;
    END
  END prog_clk
  PIN right_grid_pin_52_
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 77.600 49.680 80.000 50.280 ;
    END
  END right_grid_pin_52_
  PIN vpwr
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT 18.055 10.640 19.655 187.920 ;
    END
  END vpwr
  PIN vgnd
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT 31.385 10.640 32.985 187.920 ;
    END
  END vgnd
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 74.060 187.765 ;
      LAYER met1 ;
        RECT 0.990 6.840 79.050 188.660 ;
      LAYER met2 ;
        RECT 1.570 197.320 2.570 197.600 ;
        RECT 3.410 197.320 4.410 197.600 ;
        RECT 5.250 197.320 6.250 197.600 ;
        RECT 7.090 197.320 8.090 197.600 ;
        RECT 8.930 197.320 10.390 197.600 ;
        RECT 11.230 197.320 12.230 197.600 ;
        RECT 13.070 197.320 14.070 197.600 ;
        RECT 14.910 197.320 15.910 197.600 ;
        RECT 16.750 197.320 18.210 197.600 ;
        RECT 19.050 197.320 20.050 197.600 ;
        RECT 20.890 197.320 21.890 197.600 ;
        RECT 22.730 197.320 23.730 197.600 ;
        RECT 24.570 197.320 26.030 197.600 ;
        RECT 26.870 197.320 27.870 197.600 ;
        RECT 28.710 197.320 29.710 197.600 ;
        RECT 30.550 197.320 31.550 197.600 ;
        RECT 32.390 197.320 33.850 197.600 ;
        RECT 34.690 197.320 35.690 197.600 ;
        RECT 36.530 197.320 37.530 197.600 ;
        RECT 38.370 197.320 39.370 197.600 ;
        RECT 40.210 197.320 41.670 197.600 ;
        RECT 42.510 197.320 43.510 197.600 ;
        RECT 44.350 197.320 45.350 197.600 ;
        RECT 46.190 197.320 47.190 197.600 ;
        RECT 48.030 197.320 49.490 197.600 ;
        RECT 50.330 197.320 51.330 197.600 ;
        RECT 52.170 197.320 53.170 197.600 ;
        RECT 54.010 197.320 55.010 197.600 ;
        RECT 55.850 197.320 57.310 197.600 ;
        RECT 58.150 197.320 59.150 197.600 ;
        RECT 59.990 197.320 60.990 197.600 ;
        RECT 61.830 197.320 62.830 197.600 ;
        RECT 63.670 197.320 65.130 197.600 ;
        RECT 65.970 197.320 66.970 197.600 ;
        RECT 67.810 197.320 68.810 197.600 ;
        RECT 69.650 197.320 70.650 197.600 ;
        RECT 71.490 197.320 72.950 197.600 ;
        RECT 73.790 197.320 74.790 197.600 ;
        RECT 75.630 197.320 76.630 197.600 ;
        RECT 77.470 197.320 78.470 197.600 ;
        RECT 1.010 2.680 79.030 197.320 ;
        RECT 1.570 2.400 2.570 2.680 ;
        RECT 3.410 2.400 4.410 2.680 ;
        RECT 5.250 2.400 6.710 2.680 ;
        RECT 7.550 2.400 8.550 2.680 ;
        RECT 9.390 2.400 10.390 2.680 ;
        RECT 11.230 2.400 12.690 2.680 ;
        RECT 13.530 2.400 14.530 2.680 ;
        RECT 15.370 2.400 16.370 2.680 ;
        RECT 17.210 2.400 18.670 2.680 ;
        RECT 19.510 2.400 20.510 2.680 ;
        RECT 21.350 2.400 22.350 2.680 ;
        RECT 23.190 2.400 24.650 2.680 ;
        RECT 25.490 2.400 26.490 2.680 ;
        RECT 27.330 2.400 28.330 2.680 ;
        RECT 29.170 2.400 30.630 2.680 ;
        RECT 31.470 2.400 32.470 2.680 ;
        RECT 33.310 2.400 34.310 2.680 ;
        RECT 35.150 2.400 36.610 2.680 ;
        RECT 37.450 2.400 38.450 2.680 ;
        RECT 39.290 2.400 40.750 2.680 ;
        RECT 41.590 2.400 42.590 2.680 ;
        RECT 43.430 2.400 44.430 2.680 ;
        RECT 45.270 2.400 46.730 2.680 ;
        RECT 47.570 2.400 48.570 2.680 ;
        RECT 49.410 2.400 50.410 2.680 ;
        RECT 51.250 2.400 52.710 2.680 ;
        RECT 53.550 2.400 54.550 2.680 ;
        RECT 55.390 2.400 56.390 2.680 ;
        RECT 57.230 2.400 58.690 2.680 ;
        RECT 59.530 2.400 60.530 2.680 ;
        RECT 61.370 2.400 62.370 2.680 ;
        RECT 63.210 2.400 64.670 2.680 ;
        RECT 65.510 2.400 66.510 2.680 ;
        RECT 67.350 2.400 68.350 2.680 ;
        RECT 69.190 2.400 70.650 2.680 ;
        RECT 71.490 2.400 72.490 2.680 ;
        RECT 73.330 2.400 74.330 2.680 ;
        RECT 75.170 2.400 76.630 2.680 ;
        RECT 77.470 2.400 78.470 2.680 ;
      LAYER met3 ;
        RECT 2.800 192.760 79.055 193.625 ;
        RECT 0.985 182.600 79.055 192.760 ;
        RECT 2.800 181.200 79.055 182.600 ;
        RECT 0.985 171.040 79.055 181.200 ;
        RECT 2.800 169.640 79.055 171.040 ;
        RECT 0.985 158.800 79.055 169.640 ;
        RECT 2.800 157.400 79.055 158.800 ;
        RECT 0.985 150.640 79.055 157.400 ;
        RECT 0.985 149.240 77.200 150.640 ;
        RECT 0.985 147.240 79.055 149.240 ;
        RECT 2.800 145.840 79.055 147.240 ;
        RECT 0.985 135.680 79.055 145.840 ;
        RECT 2.800 134.280 79.055 135.680 ;
        RECT 0.985 123.440 79.055 134.280 ;
        RECT 2.800 122.040 79.055 123.440 ;
        RECT 0.985 111.880 79.055 122.040 ;
        RECT 2.800 110.480 79.055 111.880 ;
        RECT 0.985 100.320 79.055 110.480 ;
        RECT 2.800 98.920 79.055 100.320 ;
        RECT 0.985 88.760 79.055 98.920 ;
        RECT 2.800 87.360 79.055 88.760 ;
        RECT 0.985 76.520 79.055 87.360 ;
        RECT 2.800 75.120 79.055 76.520 ;
        RECT 0.985 64.960 79.055 75.120 ;
        RECT 2.800 63.560 79.055 64.960 ;
        RECT 0.985 53.400 79.055 63.560 ;
        RECT 2.800 52.000 79.055 53.400 ;
        RECT 0.985 50.680 79.055 52.000 ;
        RECT 0.985 49.280 77.200 50.680 ;
        RECT 0.985 41.160 79.055 49.280 ;
        RECT 2.800 39.760 79.055 41.160 ;
        RECT 0.985 29.600 79.055 39.760 ;
        RECT 2.800 28.200 79.055 29.600 ;
        RECT 0.985 18.040 79.055 28.200 ;
        RECT 2.800 16.640 79.055 18.040 ;
        RECT 0.985 6.480 79.055 16.640 ;
        RECT 2.800 5.615 79.055 6.480 ;
      LAYER met4 ;
        RECT 15.935 10.640 17.655 187.920 ;
        RECT 20.055 10.640 30.985 187.920 ;
        RECT 33.385 10.640 72.985 187.920 ;
  END
END cby_1__1_
END LIBRARY

