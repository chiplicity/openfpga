* NGSPICE file created from cbx_1__0_.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_1 abstract view
.subckt sky130_fd_sc_hd__dfxtp_1 D Q CLK VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S X VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A X VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_12 abstract view
.subckt sky130_fd_sc_hd__decap_12 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A X VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A X VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
.subckt sky130_fd_sc_hd__conb_1 HI LO VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A X VGND VNB VPB VPWR
.ends

.subckt cbx_1__0_ bottom_grid_pin_0_ bottom_grid_pin_10_ bottom_grid_pin_12_ bottom_grid_pin_14_
+ bottom_grid_pin_16_ bottom_grid_pin_2_ bottom_grid_pin_4_ bottom_grid_pin_6_ bottom_grid_pin_8_
+ ccff_head ccff_tail chanx_left_in[0] chanx_left_in[10] chanx_left_in[11] chanx_left_in[12]
+ chanx_left_in[13] chanx_left_in[14] chanx_left_in[15] chanx_left_in[16] chanx_left_in[17]
+ chanx_left_in[18] chanx_left_in[19] chanx_left_in[1] chanx_left_in[2] chanx_left_in[3]
+ chanx_left_in[4] chanx_left_in[5] chanx_left_in[6] chanx_left_in[7] chanx_left_in[8]
+ chanx_left_in[9] chanx_left_out[0] chanx_left_out[10] chanx_left_out[11] chanx_left_out[12]
+ chanx_left_out[13] chanx_left_out[14] chanx_left_out[15] chanx_left_out[16] chanx_left_out[17]
+ chanx_left_out[18] chanx_left_out[19] chanx_left_out[1] chanx_left_out[2] chanx_left_out[3]
+ chanx_left_out[4] chanx_left_out[5] chanx_left_out[6] chanx_left_out[7] chanx_left_out[8]
+ chanx_left_out[9] chanx_right_in[0] chanx_right_in[10] chanx_right_in[11] chanx_right_in[12]
+ chanx_right_in[13] chanx_right_in[14] chanx_right_in[15] chanx_right_in[16] chanx_right_in[17]
+ chanx_right_in[18] chanx_right_in[19] chanx_right_in[1] chanx_right_in[2] chanx_right_in[3]
+ chanx_right_in[4] chanx_right_in[5] chanx_right_in[6] chanx_right_in[7] chanx_right_in[8]
+ chanx_right_in[9] chanx_right_out[0] chanx_right_out[10] chanx_right_out[11] chanx_right_out[12]
+ chanx_right_out[13] chanx_right_out[14] chanx_right_out[15] chanx_right_out[16]
+ chanx_right_out[17] chanx_right_out[18] chanx_right_out[19] chanx_right_out[1] chanx_right_out[2]
+ chanx_right_out[3] chanx_right_out[4] chanx_right_out[5] chanx_right_out[6] chanx_right_out[7]
+ chanx_right_out[8] chanx_right_out[9] prog_clk VPWR VGND
Xmem_top_ipin_8.sky130_fd_sc_hd__dfxtp_1_0_ mux_top_ipin_7.mux_l4_in_0_/S mux_top_ipin_8.mux_l1_in_1_/S
+ clkbuf_2_3_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
Xmux_top_ipin_1.mux_l1_in_1_ chanx_right_in[3] chanx_left_in[3] mux_top_ipin_1.mux_l1_in_2_/S
+ mux_top_ipin_1.mux_l1_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_3_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_top_ipin_6.mux_l2_in_0_ mux_top_ipin_6.mux_l1_in_1_/X mux_top_ipin_6.mux_l1_in_0_/X
+ mux_top_ipin_6.mux_l2_in_0_/S mux_top_ipin_6.mux_l2_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_49_ chanx_left_in[0] chanx_right_out[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_18_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_top_ipin_6.mux_l1_in_1_ chanx_right_in[2] chanx_left_in[2] mux_top_ipin_6.mux_l1_in_0_/S
+ mux_top_ipin_6.mux_l1_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_20_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_top_ipin_1.mux_l1_in_0_ chanx_right_in[1] chanx_left_in[1] mux_top_ipin_1.mux_l1_in_2_/S
+ mux_top_ipin_1.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_3_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_48_ chanx_left_in[1] chanx_right_out[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_18_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_top_ipin_6.mux_l1_in_0_ chanx_right_in[0] chanx_left_in[0] mux_top_ipin_6.mux_l1_in_0_/S
+ mux_top_ipin_6.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_20_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_top_ipin_4.sky130_fd_sc_hd__buf_4_0_ mux_top_ipin_4.mux_l4_in_0_/X bottom_grid_pin_8_
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_4
XFILLER_3_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_47_ chanx_left_in[2] chanx_right_out[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_9_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_2_1_0_prog_clk clkbuf_2_1_0_prog_clk/A clkbuf_2_1_0_prog_clk/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_8_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_46_ chanx_left_in[3] chanx_right_out[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_18_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_29_ chanx_right_in[0] chanx_left_out[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_20_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_top_ipin_2.mux_l2_in_3_ _11_/HI chanx_right_in[18] mux_top_ipin_2.mux_l2_in_2_/S
+ mux_top_ipin_2.mux_l2_in_3_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_8_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_45_ chanx_left_in[4] chanx_right_out[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
Xmux_top_ipin_2.mux_l4_in_0_ mux_top_ipin_2.mux_l3_in_1_/X mux_top_ipin_2.mux_l3_in_0_/X
+ mux_top_ipin_2.mux_l4_in_0_/S mux_top_ipin_2.mux_l4_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XFILLER_1_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28_ chanx_right_in[1] chanx_left_out[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
Xmux_top_ipin_7.mux_l2_in_3_ _16_/HI chanx_right_in[17] mux_top_ipin_7.mux_l2_in_1_/S
+ mux_top_ipin_7.mux_l2_in_3_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_19_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_top_ipin_2.mux_l3_in_1_ mux_top_ipin_2.mux_l2_in_3_/X mux_top_ipin_2.mux_l2_in_2_/X
+ mux_top_ipin_2.mux_l3_in_1_/S mux_top_ipin_2.mux_l3_in_1_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XFILLER_6_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_top_ipin_2.mux_l2_in_2_ chanx_left_in[18] chanx_right_in[12] mux_top_ipin_2.mux_l2_in_2_/S
+ mux_top_ipin_2.mux_l2_in_2_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
Xmux_top_ipin_7.mux_l4_in_0_ mux_top_ipin_7.mux_l3_in_1_/X mux_top_ipin_7.mux_l3_in_0_/X
+ mux_top_ipin_7.mux_l4_in_0_/S mux_top_ipin_7.mux_l4_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XFILLER_12_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_top_ipin_7.mux_l3_in_1_ mux_top_ipin_7.mux_l2_in_3_/X mux_top_ipin_7.mux_l2_in_2_/X
+ mux_top_ipin_7.mux_l3_in_1_/S mux_top_ipin_7.mux_l3_in_1_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XFILLER_13_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_44_ chanx_left_in[5] chanx_right_out[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_1_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27_ chanx_right_in[2] chanx_left_out[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_20_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_top_ipin_7.mux_l2_in_2_ chanx_left_in[17] chanx_right_in[11] mux_top_ipin_7.mux_l2_in_1_/S
+ mux_top_ipin_7.mux_l2_in_2_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
Xmux_top_ipin_2.mux_l3_in_0_ mux_top_ipin_2.mux_l2_in_1_/X mux_top_ipin_2.mux_l2_in_0_/X
+ mux_top_ipin_2.mux_l3_in_1_/S mux_top_ipin_2.mux_l3_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XFILLER_10_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_0 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_top_ipin_2.mux_l2_in_1_ chanx_left_in[12] mux_top_ipin_2.mux_l1_in_2_/X mux_top_ipin_2.mux_l2_in_2_/S
+ mux_top_ipin_2.mux_l2_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_8_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_2_0_0_prog_clk clkbuf_2_1_0_prog_clk/A clkbuf_2_0_0_prog_clk/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__clkbuf_1
Xmux_top_ipin_2.mux_l1_in_2_ chanx_right_in[6] chanx_left_in[6] mux_top_ipin_2.mux_l1_in_2_/S
+ mux_top_ipin_2.mux_l1_in_2_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
Xmux_top_ipin_7.mux_l3_in_0_ mux_top_ipin_7.mux_l2_in_1_/X mux_top_ipin_7.mux_l2_in_0_/X
+ mux_top_ipin_7.mux_l3_in_1_/S mux_top_ipin_7.mux_l3_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XFILLER_2_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_43_ chanx_left_in[6] chanx_right_out[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
Xmux_top_ipin_7.sky130_fd_sc_hd__buf_4_0_ mux_top_ipin_7.mux_l4_in_0_/X bottom_grid_pin_14_
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_4
XFILLER_18_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_top_ipin_7.mux_l2_in_1_ chanx_left_in[11] mux_top_ipin_7.mux_l1_in_2_/X mux_top_ipin_7.mux_l2_in_1_/S
+ mux_top_ipin_7.mux_l2_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_1_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_26_ chanx_right_in[3] chanx_left_out[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_19_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09_ _09_/HI _09_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XFILLER_22_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmux_top_ipin_7.mux_l1_in_2_ chanx_right_in[7] chanx_left_in[7] mux_top_ipin_7.mux_l1_in_2_/S
+ mux_top_ipin_7.mux_l1_in_2_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XPHY_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_top_ipin_2.mux_l2_in_0_ mux_top_ipin_2.mux_l1_in_1_/X mux_top_ipin_2.mux_l1_in_0_/X
+ mux_top_ipin_2.mux_l2_in_2_/S mux_top_ipin_2.mux_l2_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XFILLER_8_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_top_ipin_2.mux_l1_in_1_ chanx_right_in[2] chanx_left_in[2] mux_top_ipin_2.mux_l1_in_2_/S
+ mux_top_ipin_2.mux_l1_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_2_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmem_top_ipin_1.sky130_fd_sc_hd__dfxtp_1_3_ mux_top_ipin_1.mux_l3_in_1_/S mux_top_ipin_1.mux_l4_in_0_/S
+ clkbuf_2_0_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
X_42_ chanx_left_in[7] chanx_right_out[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_18_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_top_ipin_7.mux_l2_in_0_ mux_top_ipin_7.mux_l1_in_1_/X mux_top_ipin_7.mux_l1_in_0_/X
+ mux_top_ipin_7.mux_l2_in_1_/S mux_top_ipin_7.mux_l2_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
X_25_ chanx_right_in[4] chanx_left_out[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_19_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_top_ipin_7.mux_l1_in_1_ chanx_right_in[3] chanx_left_in[3] mux_top_ipin_7.mux_l1_in_2_/S
+ mux_top_ipin_7.mux_l1_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XPHY_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmem_top_ipin_4.sky130_fd_sc_hd__dfxtp_1_3_ mux_top_ipin_4.mux_l3_in_1_/S mux_top_ipin_4.mux_l4_in_0_/S
+ clkbuf_2_1_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_12_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmux_top_ipin_2.mux_l1_in_0_ chanx_right_in[0] chanx_left_in[0] mux_top_ipin_2.mux_l1_in_2_/S
+ mux_top_ipin_2.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
Xmem_top_ipin_1.sky130_fd_sc_hd__dfxtp_1_2_ mux_top_ipin_1.mux_l2_in_3_/S mux_top_ipin_1.mux_l3_in_1_/S
+ clkbuf_2_0_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
X_41_ chanx_left_in[8] chanx_right_out[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
X_24_ chanx_right_in[5] chanx_left_out[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_19_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmem_top_ipin_7.sky130_fd_sc_hd__dfxtp_1_3_ mux_top_ipin_7.mux_l3_in_1_/S mux_top_ipin_7.mux_l4_in_0_/S
+ clkbuf_2_3_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
Xmux_top_ipin_0.sky130_fd_sc_hd__buf_4_0_ mux_top_ipin_0.mux_l4_in_0_/X bottom_grid_pin_0_
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_4
XPHY_101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmux_top_ipin_7.mux_l1_in_0_ chanx_right_in[1] chanx_left_in[1] mux_top_ipin_7.mux_l1_in_2_/S
+ mux_top_ipin_7.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XPHY_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmem_top_ipin_4.sky130_fd_sc_hd__dfxtp_1_2_ mux_top_ipin_4.mux_l2_in_3_/S mux_top_ipin_4.mux_l3_in_1_/S
+ clkbuf_2_1_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_12_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmem_top_ipin_1.sky130_fd_sc_hd__dfxtp_1_1_ mux_top_ipin_1.mux_l1_in_2_/S mux_top_ipin_1.mux_l2_in_3_/S
+ clkbuf_2_0_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_4_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_40_ chanx_left_in[9] chanx_right_out[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
X_23_ chanx_right_in[6] chanx_left_out[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_19_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmem_top_ipin_7.sky130_fd_sc_hd__dfxtp_1_2_ mux_top_ipin_7.mux_l2_in_1_/S mux_top_ipin_7.mux_l3_in_1_/S
+ clkbuf_2_3_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XPHY_102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmem_top_ipin_4.sky130_fd_sc_hd__dfxtp_1_1_ mux_top_ipin_4.mux_l1_in_2_/S mux_top_ipin_4.mux_l2_in_3_/S
+ clkbuf_2_1_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
Xmem_top_ipin_1.sky130_fd_sc_hd__dfxtp_1_0_ mux_top_ipin_0.mux_l4_in_0_/S mux_top_ipin_1.mux_l1_in_2_/S
+ clkbuf_2_0_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_1_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22_ chanx_right_in[7] chanx_left_out[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_1_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmem_top_ipin_7.sky130_fd_sc_hd__dfxtp_1_1_ mux_top_ipin_7.mux_l1_in_2_/S mux_top_ipin_7.mux_l2_in_1_/S
+ clkbuf_2_3_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_18_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmem_top_ipin_4.sky130_fd_sc_hd__dfxtp_1_0_ mux_top_ipin_3.mux_l4_in_0_/S mux_top_ipin_4.mux_l1_in_2_/S
+ clkbuf_2_1_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_12_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmux_top_ipin_3.mux_l2_in_3_ _12_/HI chanx_right_in[19] mux_top_ipin_3.mux_l2_in_1_/S
+ mux_top_ipin_3.mux_l2_in_3_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_1_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21_ chanx_right_in[8] chanx_left_out[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_1_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmem_top_ipin_7.sky130_fd_sc_hd__dfxtp_1_0_ mux_top_ipin_6.mux_l4_in_0_/S mux_top_ipin_7.mux_l1_in_2_/S
+ clkbuf_2_3_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_10_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_top_ipin_3.mux_l4_in_0_ mux_top_ipin_3.mux_l3_in_1_/X mux_top_ipin_3.mux_l3_in_0_/X
+ mux_top_ipin_3.mux_l4_in_0_/S mux_top_ipin_3.mux_l4_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XPHY_104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_top_ipin_8.mux_l2_in_3_ _17_/HI chanx_right_in[18] mux_top_ipin_8.mux_l2_in_2_/S
+ mux_top_ipin_8.mux_l2_in_3_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
Xmux_top_ipin_3.mux_l3_in_1_ mux_top_ipin_3.mux_l2_in_3_/X mux_top_ipin_3.mux_l2_in_2_/X
+ mux_top_ipin_3.mux_l3_in_1_/S mux_top_ipin_3.mux_l3_in_1_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XFILLER_12_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_top_ipin_3.mux_l2_in_2_ chanx_left_in[19] chanx_right_in[13] mux_top_ipin_3.mux_l2_in_1_/S
+ mux_top_ipin_3.mux_l2_in_2_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_1_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmux_top_ipin_8.mux_l4_in_0_ mux_top_ipin_8.mux_l3_in_1_/X mux_top_ipin_8.mux_l3_in_0_/X
+ ccff_tail mux_top_ipin_8.mux_l4_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_1_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20_ chanx_right_in[9] chanx_left_out[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
Xmux_top_ipin_8.mux_l3_in_1_ mux_top_ipin_8.mux_l2_in_3_/X mux_top_ipin_8.mux_l2_in_2_/X
+ mux_top_ipin_8.mux_l3_in_0_/S mux_top_ipin_8.mux_l3_in_1_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
Xclkbuf_0_prog_clk prog_clk clkbuf_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__clkbuf_16
XFILLER_10_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_top_ipin_3.sky130_fd_sc_hd__buf_4_0_ mux_top_ipin_3.mux_l4_in_0_/X bottom_grid_pin_6_
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_4
XFILLER_7_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_top_ipin_8.mux_l2_in_2_ chanx_left_in[18] chanx_right_in[12] mux_top_ipin_8.mux_l2_in_2_/S
+ mux_top_ipin_8.mux_l2_in_2_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
Xmux_top_ipin_3.mux_l3_in_0_ mux_top_ipin_3.mux_l2_in_1_/X mux_top_ipin_3.mux_l2_in_0_/X
+ mux_top_ipin_3.mux_l3_in_1_/S mux_top_ipin_3.mux_l3_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XFILLER_16_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_top_ipin_3.mux_l2_in_1_ chanx_left_in[13] mux_top_ipin_3.mux_l1_in_2_/X mux_top_ipin_3.mux_l2_in_1_/S
+ mux_top_ipin_3.mux_l2_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_1_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_top_ipin_3.mux_l1_in_2_ chanx_right_in[7] chanx_left_in[7] mux_top_ipin_3.mux_l1_in_2_/S
+ mux_top_ipin_3.mux_l1_in_2_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
Xmux_top_ipin_8.mux_l3_in_0_ mux_top_ipin_8.mux_l2_in_1_/X mux_top_ipin_8.mux_l2_in_0_/X
+ mux_top_ipin_8.mux_l3_in_0_/S mux_top_ipin_8.mux_l3_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XFILLER_10_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_top_ipin_8.mux_l2_in_1_ chanx_left_in[12] mux_top_ipin_8.mux_l1_in_2_/X mux_top_ipin_8.mux_l2_in_2_/S
+ mux_top_ipin_8.mux_l2_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_21_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmux_top_ipin_8.mux_l1_in_2_ chanx_right_in[8] chanx_left_in[8] mux_top_ipin_8.mux_l1_in_1_/S
+ mux_top_ipin_8.mux_l1_in_2_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
Xmux_top_ipin_3.mux_l2_in_0_ mux_top_ipin_3.mux_l1_in_1_/X mux_top_ipin_3.mux_l1_in_0_/X
+ mux_top_ipin_3.mux_l2_in_1_/S mux_top_ipin_3.mux_l2_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XFILLER_13_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_top_ipin_3.mux_l1_in_1_ chanx_right_in[3] chanx_left_in[3] mux_top_ipin_3.mux_l1_in_2_/S
+ mux_top_ipin_3.mux_l1_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_10_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_top_ipin_8.mux_l2_in_0_ mux_top_ipin_8.mux_l1_in_1_/X mux_top_ipin_8.mux_l1_in_0_/X
+ mux_top_ipin_8.mux_l2_in_2_/S mux_top_ipin_8.mux_l2_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XFILLER_21_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_top_ipin_8.mux_l1_in_1_ chanx_right_in[2] chanx_left_in[2] mux_top_ipin_8.mux_l1_in_1_/S
+ mux_top_ipin_8.mux_l1_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_13_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_top_ipin_3.mux_l1_in_0_ chanx_right_in[1] chanx_left_in[1] mux_top_ipin_3.mux_l1_in_2_/S
+ mux_top_ipin_3.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_10_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmux_top_ipin_8.mux_l1_in_0_ chanx_right_in[0] chanx_left_in[0] mux_top_ipin_8.mux_l1_in_1_/S
+ mux_top_ipin_8.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_13_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmux_top_ipin_6.sky130_fd_sc_hd__buf_4_0_ mux_top_ipin_6.mux_l4_in_0_/X bottom_grid_pin_12_
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_4
XFILLER_14_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_90 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmux_top_ipin_4.mux_l2_in_3_ _13_/HI chanx_right_in[14] mux_top_ipin_4.mux_l2_in_3_/S
+ mux_top_ipin_4.mux_l2_in_3_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_19_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_91 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_80 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_57_ chanx_right_in[12] chanx_left_out[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_15_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_top_ipin_4.mux_l4_in_0_ mux_top_ipin_4.mux_l3_in_1_/X mux_top_ipin_4.mux_l3_in_0_/X
+ mux_top_ipin_4.mux_l4_in_0_/S mux_top_ipin_4.mux_l4_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
Xmem_top_ipin_0.sky130_fd_sc_hd__dfxtp_1_3_ mux_top_ipin_0.mux_l3_in_1_/S mux_top_ipin_0.mux_l4_in_0_/S
+ clkbuf_2_0_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_7_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_top_ipin_4.mux_l3_in_1_ mux_top_ipin_4.mux_l2_in_3_/X mux_top_ipin_4.mux_l2_in_2_/X
+ mux_top_ipin_4.mux_l3_in_1_/S mux_top_ipin_4.mux_l3_in_1_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_top_ipin_4.mux_l2_in_2_ chanx_left_in[14] chanx_right_in[8] mux_top_ipin_4.mux_l2_in_3_/S
+ mux_top_ipin_4.mux_l2_in_2_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_14_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_92 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmem_top_ipin_3.sky130_fd_sc_hd__dfxtp_1_3_ mux_top_ipin_3.mux_l3_in_1_/S mux_top_ipin_3.mux_l4_in_0_/S
+ clkbuf_2_1_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XPHY_81 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_70 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_56_ chanx_right_in[13] chanx_left_out[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
X_39_ chanx_left_in[10] chanx_right_out[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
Xmem_top_ipin_0.sky130_fd_sc_hd__dfxtp_1_2_ mux_top_ipin_0.mux_l2_in_2_/S mux_top_ipin_0.mux_l3_in_1_/S
+ clkbuf_2_0_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_11_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_top_ipin_4.mux_l3_in_0_ mux_top_ipin_4.mux_l2_in_1_/X mux_top_ipin_4.mux_l2_in_0_/X
+ mux_top_ipin_4.mux_l3_in_1_/S mux_top_ipin_4.mux_l3_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
Xmem_top_ipin_6.sky130_fd_sc_hd__dfxtp_1_3_ mux_top_ipin_6.mux_l3_in_1_/S mux_top_ipin_6.mux_l4_in_0_/S
+ clkbuf_2_2_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_19_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_top_ipin_4.mux_l2_in_1_ chanx_left_in[8] mux_top_ipin_4.mux_l1_in_2_/X mux_top_ipin_4.mux_l2_in_3_/S
+ mux_top_ipin_4.mux_l2_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XPHY_93 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_82 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_60 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_71 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmem_top_ipin_3.sky130_fd_sc_hd__dfxtp_1_2_ mux_top_ipin_3.mux_l2_in_1_/S mux_top_ipin_3.mux_l3_in_1_/S
+ clkbuf_2_1_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_2_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_55_ chanx_right_in[14] chanx_left_out[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_15_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_top_ipin_4.mux_l1_in_2_ chanx_right_in[4] chanx_left_in[4] mux_top_ipin_4.mux_l1_in_2_/S
+ mux_top_ipin_4.mux_l1_in_2_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_20_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_38_ chanx_left_in[11] chanx_right_out[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_22_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmem_top_ipin_0.sky130_fd_sc_hd__dfxtp_1_1_ mux_top_ipin_0.mux_l1_in_1_/S mux_top_ipin_0.mux_l2_in_2_/S
+ clkbuf_2_2_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_11_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmem_top_ipin_6.sky130_fd_sc_hd__dfxtp_1_2_ mux_top_ipin_6.mux_l2_in_0_/S mux_top_ipin_6.mux_l3_in_1_/S
+ clkbuf_2_2_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
Xmux_top_ipin_4.mux_l2_in_0_ mux_top_ipin_4.mux_l1_in_1_/X mux_top_ipin_4.mux_l1_in_0_/X
+ mux_top_ipin_4.mux_l2_in_3_/S mux_top_ipin_4.mux_l2_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XFILLER_18_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_94 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_83 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_50 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_61 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_72 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmem_top_ipin_3.sky130_fd_sc_hd__dfxtp_1_1_ mux_top_ipin_3.mux_l1_in_2_/S mux_top_ipin_3.mux_l2_in_1_/S
+ clkbuf_2_1_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
X_54_ chanx_right_in[15] chanx_left_out[15] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_2_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_top_ipin_4.mux_l1_in_1_ chanx_right_in[2] chanx_left_in[2] mux_top_ipin_4.mux_l1_in_2_/S
+ mux_top_ipin_4.mux_l1_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_2_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_37_ chanx_left_in[12] chanx_right_out[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
Xmem_top_ipin_0.sky130_fd_sc_hd__dfxtp_1_0_ ccff_head mux_top_ipin_0.mux_l1_in_1_/S
+ clkbuf_2_2_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_8_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmem_top_ipin_6.sky130_fd_sc_hd__dfxtp_1_1_ mux_top_ipin_6.mux_l1_in_0_/S mux_top_ipin_6.mux_l2_in_0_/S
+ clkbuf_2_2_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_14_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_95 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_84 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_51 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_62 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_73 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmem_top_ipin_3.sky130_fd_sc_hd__dfxtp_1_0_ mux_top_ipin_2.mux_l4_in_0_/S mux_top_ipin_3.mux_l1_in_2_/S
+ clkbuf_2_1_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
X_53_ chanx_right_in[16] chanx_left_out[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_14_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_top_ipin_4.mux_l1_in_0_ chanx_right_in[0] chanx_left_in[0] mux_top_ipin_4.mux_l1_in_2_/S
+ mux_top_ipin_4.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
X_36_ chanx_left_in[13] chanx_right_out[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_22_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19_ chanx_right_in[10] chanx_left_out[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_17_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmem_top_ipin_6.sky130_fd_sc_hd__dfxtp_1_0_ mux_top_ipin_5.mux_l4_in_0_/S mux_top_ipin_6.mux_l1_in_0_/S
+ clkbuf_2_2_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_10_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_top_ipin_2.sky130_fd_sc_hd__buf_4_0_ mux_top_ipin_2.mux_l4_in_0_/X bottom_grid_pin_4_
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_4
XPHY_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_96 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_85 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_52 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_63 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_52_ chanx_right_in[17] chanx_left_out[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XPHY_74 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_35_ chanx_left_in[14] chanx_right_out[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_22_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18_ chanx_right_in[11] chanx_left_out[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_3_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_97 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_86 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_53 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_64 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_75 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_51_ chanx_right_in[18] chanx_left_out[18] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_11_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_34_ chanx_left_in[15] chanx_right_out[15] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_22_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17_ _17_/HI _17_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XFILLER_3_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_top_ipin_0.mux_l2_in_3_ _09_/HI chanx_right_in[16] mux_top_ipin_0.mux_l2_in_2_/S
+ mux_top_ipin_0.mux_l2_in_3_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_5_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_98 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_87 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_54 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmux_top_ipin_0.mux_l4_in_0_ mux_top_ipin_0.mux_l3_in_1_/X mux_top_ipin_0.mux_l3_in_0_/X
+ mux_top_ipin_0.mux_l4_in_0_/S mux_top_ipin_0.mux_l4_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XPHY_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_65 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_76 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_50_ chanx_right_in[19] chanx_left_out[19] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_2_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_33_ chanx_left_in[16] chanx_right_out[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
Xmux_top_ipin_5.mux_l2_in_3_ _14_/HI chanx_right_in[15] mux_top_ipin_5.mux_l2_in_1_/S
+ mux_top_ipin_5.mux_l2_in_3_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_22_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_top_ipin_0.mux_l3_in_1_ mux_top_ipin_0.mux_l2_in_3_/X mux_top_ipin_0.mux_l2_in_2_/X
+ mux_top_ipin_0.mux_l3_in_1_/S mux_top_ipin_0.mux_l3_in_1_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XFILLER_7_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16_ _16_/HI _16_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XFILLER_17_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_top_ipin_5.mux_l4_in_0_ mux_top_ipin_5.mux_l3_in_1_/X mux_top_ipin_5.mux_l3_in_0_/X
+ mux_top_ipin_5.mux_l4_in_0_/S mux_top_ipin_5.mux_l4_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
Xmux_top_ipin_0.mux_l2_in_2_ chanx_left_in[16] chanx_right_in[10] mux_top_ipin_0.mux_l2_in_2_/S
+ mux_top_ipin_0.mux_l2_in_2_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_0_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_top_ipin_5.mux_l3_in_1_ mux_top_ipin_5.mux_l2_in_3_/X mux_top_ipin_5.mux_l2_in_2_/X
+ mux_top_ipin_5.mux_l3_in_0_/S mux_top_ipin_5.mux_l3_in_1_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XPHY_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_99 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_88 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_55 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_66 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_77 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_32_ chanx_left_in[17] chanx_right_out[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
Xmux_top_ipin_5.mux_l2_in_2_ chanx_left_in[15] chanx_right_in[9] mux_top_ipin_5.mux_l2_in_1_/S
+ mux_top_ipin_5.mux_l2_in_2_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_22_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmux_top_ipin_0.mux_l3_in_0_ mux_top_ipin_0.mux_l2_in_1_/X mux_top_ipin_0.mux_l2_in_0_/X
+ mux_top_ipin_0.mux_l3_in_1_/S mux_top_ipin_0.mux_l3_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XFILLER_19_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15_ _15_/HI _15_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XFILLER_6_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_top_ipin_0.mux_l2_in_1_ chanx_left_in[10] mux_top_ipin_0.mux_l1_in_2_/X mux_top_ipin_0.mux_l2_in_2_/S
+ mux_top_ipin_0.mux_l2_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_0_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmux_top_ipin_0.mux_l1_in_2_ chanx_right_in[4] chanx_left_in[4] mux_top_ipin_0.mux_l1_in_1_/S
+ mux_top_ipin_0.mux_l1_in_2_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XPHY_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_top_ipin_5.mux_l3_in_0_ mux_top_ipin_5.mux_l2_in_1_/X mux_top_ipin_5.mux_l2_in_0_/X
+ mux_top_ipin_5.mux_l3_in_0_/S mux_top_ipin_5.mux_l3_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
Xmux_top_ipin_5.sky130_fd_sc_hd__buf_4_0_ mux_top_ipin_5.mux_l4_in_0_/X bottom_grid_pin_10_
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_4
XPHY_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_89 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_56 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_67 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_78 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_31_ chanx_left_in[18] chanx_right_out[18] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
Xmux_top_ipin_5.mux_l2_in_1_ chanx_left_in[9] mux_top_ipin_5.mux_l1_in_2_/X mux_top_ipin_5.mux_l2_in_1_/S
+ mux_top_ipin_5.mux_l2_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_11_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14_ _14_/HI _14_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
Xmux_top_ipin_5.mux_l1_in_2_ chanx_right_in[5] chanx_left_in[5] mux_top_ipin_5.mux_l1_in_0_/S
+ mux_top_ipin_5.mux_l1_in_2_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
Xmux_top_ipin_0.mux_l2_in_0_ mux_top_ipin_0.mux_l1_in_1_/X mux_top_ipin_0.mux_l1_in_0_/X
+ mux_top_ipin_0.mux_l2_in_2_/S mux_top_ipin_0.mux_l2_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
Xmux_top_ipin_0.mux_l1_in_1_ chanx_right_in[2] chanx_left_in[2] mux_top_ipin_0.mux_l1_in_1_/S
+ mux_top_ipin_0.mux_l1_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XPHY_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_79 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_46 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_57 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_68 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_30_ chanx_left_in[19] chanx_right_out[19] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_9_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmux_top_ipin_5.mux_l2_in_0_ mux_top_ipin_5.mux_l1_in_1_/X mux_top_ipin_5.mux_l1_in_0_/X
+ mux_top_ipin_5.mux_l2_in_1_/S mux_top_ipin_5.mux_l2_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XFILLER_12_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13_ _13_/HI _13_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XFILLER_17_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_top_ipin_5.mux_l1_in_1_ chanx_right_in[3] chanx_left_in[3] mux_top_ipin_5.mux_l1_in_0_/S
+ mux_top_ipin_5.mux_l1_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_0_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_top_ipin_0.mux_l1_in_0_ chanx_right_in[0] chanx_left_in[0] mux_top_ipin_0.mux_l1_in_1_/S
+ mux_top_ipin_0.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_20_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_47 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_58 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_69 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12_ _12_/HI _12_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XFILLER_10_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_top_ipin_5.mux_l1_in_0_ chanx_right_in[1] chanx_left_in[1] mux_top_ipin_5.mux_l1_in_0_/S
+ mux_top_ipin_5.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_3_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_48 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_59 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11_ _11_/HI _11_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XFILLER_10_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_1_1_0_prog_clk clkbuf_0_prog_clk/X clkbuf_2_3_0_prog_clk/A VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__clkbuf_1
Xmem_top_ipin_2.sky130_fd_sc_hd__dfxtp_1_3_ mux_top_ipin_2.mux_l3_in_1_/S mux_top_ipin_2.mux_l4_in_0_/S
+ clkbuf_2_1_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_20_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_49 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_top_ipin_8.sky130_fd_sc_hd__buf_4_0_ mux_top_ipin_8.mux_l4_in_0_/X bottom_grid_pin_16_
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_4
XFILLER_7_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10_ _10_/HI _10_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
Xmem_top_ipin_5.sky130_fd_sc_hd__dfxtp_1_3_ mux_top_ipin_5.mux_l3_in_0_/S mux_top_ipin_5.mux_l4_in_0_/S
+ clkbuf_2_2_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
Xclkbuf_2_3_0_prog_clk clkbuf_2_3_0_prog_clk/A clkbuf_2_3_0_prog_clk/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_18_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmem_top_ipin_2.sky130_fd_sc_hd__dfxtp_1_2_ mux_top_ipin_2.mux_l2_in_2_/S mux_top_ipin_2.mux_l3_in_1_/S
+ clkbuf_2_1_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XPHY_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_top_ipin_1.mux_l2_in_3_ _10_/HI chanx_right_in[17] mux_top_ipin_1.mux_l2_in_3_/S
+ mux_top_ipin_1.mux_l2_in_3_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XPHY_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmem_top_ipin_8.sky130_fd_sc_hd__dfxtp_1_3_ mux_top_ipin_8.mux_l3_in_0_/S ccff_tail
+ clkbuf_2_2_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
Xmux_top_ipin_1.mux_l4_in_0_ mux_top_ipin_1.mux_l3_in_1_/X mux_top_ipin_1.mux_l3_in_0_/X
+ mux_top_ipin_1.mux_l4_in_0_/S mux_top_ipin_1.mux_l4_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XFILLER_6_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmem_top_ipin_5.sky130_fd_sc_hd__dfxtp_1_2_ mux_top_ipin_5.mux_l2_in_1_/S mux_top_ipin_5.mux_l3_in_0_/S
+ clkbuf_2_3_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_0_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmux_top_ipin_6.mux_l2_in_3_ _15_/HI chanx_right_in[16] mux_top_ipin_6.mux_l2_in_0_/S
+ mux_top_ipin_6.mux_l2_in_3_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
Xmux_top_ipin_1.mux_l3_in_1_ mux_top_ipin_1.mux_l2_in_3_/X mux_top_ipin_1.mux_l2_in_2_/X
+ mux_top_ipin_1.mux_l3_in_1_/S mux_top_ipin_1.mux_l3_in_1_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XFILLER_15_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmem_top_ipin_2.sky130_fd_sc_hd__dfxtp_1_1_ mux_top_ipin_2.mux_l1_in_2_/S mux_top_ipin_2.mux_l2_in_2_/S
+ clkbuf_2_0_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_6_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_top_ipin_1.mux_l2_in_2_ chanx_left_in[17] chanx_right_in[11] mux_top_ipin_1.mux_l2_in_3_/S
+ mux_top_ipin_1.mux_l2_in_2_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XPHY_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_top_ipin_6.mux_l4_in_0_ mux_top_ipin_6.mux_l3_in_1_/X mux_top_ipin_6.mux_l3_in_0_/X
+ mux_top_ipin_6.mux_l4_in_0_/S mux_top_ipin_6.mux_l4_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XPHY_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmem_top_ipin_8.sky130_fd_sc_hd__dfxtp_1_2_ mux_top_ipin_8.mux_l2_in_2_/S mux_top_ipin_8.mux_l3_in_0_/S
+ clkbuf_2_3_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_3_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_top_ipin_6.mux_l3_in_1_ mux_top_ipin_6.mux_l2_in_3_/X mux_top_ipin_6.mux_l2_in_2_/X
+ mux_top_ipin_6.mux_l3_in_1_/S mux_top_ipin_6.mux_l3_in_1_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XFILLER_12_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_top_ipin_1.sky130_fd_sc_hd__buf_4_0_ mux_top_ipin_1.mux_l4_in_0_/X bottom_grid_pin_2_
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_4
Xmem_top_ipin_5.sky130_fd_sc_hd__dfxtp_1_1_ mux_top_ipin_5.mux_l1_in_0_/S mux_top_ipin_5.mux_l2_in_1_/S
+ clkbuf_2_3_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
Xmux_top_ipin_6.mux_l2_in_2_ chanx_left_in[16] chanx_right_in[10] mux_top_ipin_6.mux_l2_in_0_/S
+ mux_top_ipin_6.mux_l2_in_2_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_0_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_top_ipin_1.mux_l3_in_0_ mux_top_ipin_1.mux_l2_in_1_/X mux_top_ipin_1.mux_l2_in_0_/X
+ mux_top_ipin_1.mux_l3_in_1_/S mux_top_ipin_1.mux_l3_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XFILLER_9_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmem_top_ipin_2.sky130_fd_sc_hd__dfxtp_1_0_ mux_top_ipin_1.mux_l4_in_0_/S mux_top_ipin_2.mux_l1_in_2_/S
+ clkbuf_2_0_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
Xmux_top_ipin_1.mux_l2_in_1_ chanx_left_in[11] mux_top_ipin_1.mux_l1_in_2_/X mux_top_ipin_1.mux_l2_in_3_/S
+ mux_top_ipin_1.mux_l2_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_6_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_1_0_0_prog_clk clkbuf_0_prog_clk/X clkbuf_2_1_0_prog_clk/A VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__clkbuf_1
Xmux_top_ipin_1.mux_l1_in_2_ chanx_right_in[5] chanx_left_in[5] mux_top_ipin_1.mux_l1_in_2_/S
+ mux_top_ipin_1.mux_l1_in_2_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
Xmem_top_ipin_8.sky130_fd_sc_hd__dfxtp_1_1_ mux_top_ipin_8.mux_l1_in_1_/S mux_top_ipin_8.mux_l2_in_2_/S
+ clkbuf_2_3_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_13_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_top_ipin_6.mux_l3_in_0_ mux_top_ipin_6.mux_l2_in_1_/X mux_top_ipin_6.mux_l2_in_0_/X
+ mux_top_ipin_6.mux_l3_in_1_/S mux_top_ipin_6.mux_l3_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XFILLER_12_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmem_top_ipin_5.sky130_fd_sc_hd__dfxtp_1_0_ mux_top_ipin_4.mux_l4_in_0_/S mux_top_ipin_5.mux_l1_in_0_/S
+ clkbuf_2_3_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_2_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_top_ipin_6.mux_l2_in_1_ chanx_left_in[10] mux_top_ipin_6.mux_l1_in_2_/X mux_top_ipin_6.mux_l2_in_0_/S
+ mux_top_ipin_6.mux_l2_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_0_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_top_ipin_6.mux_l1_in_2_ chanx_right_in[6] chanx_left_in[6] mux_top_ipin_6.mux_l1_in_0_/S
+ mux_top_ipin_6.mux_l1_in_2_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
Xmux_top_ipin_1.mux_l2_in_0_ mux_top_ipin_1.mux_l1_in_1_/X mux_top_ipin_1.mux_l1_in_0_/X
+ mux_top_ipin_1.mux_l2_in_3_/S mux_top_ipin_1.mux_l2_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
Xclkbuf_2_2_0_prog_clk clkbuf_2_3_0_prog_clk/A clkbuf_2_2_0_prog_clk/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_20_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
.ends

