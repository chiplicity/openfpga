* NGSPICE file created from cby_1__1_.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_1 abstract view
.subckt sky130_fd_sc_hd__dfxtp_1 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_8 abstract view
.subckt sky130_fd_sc_hd__buf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
.subckt sky130_fd_sc_hd__conb_1 VGND VNB VPB VPWR HI LO
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_12 abstract view
.subckt sky130_fd_sc_hd__decap_12 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

.subckt cby_1__1_ Test_en_E_in Test_en_E_out Test_en_N_out Test_en_S_in Test_en_W_in
+ Test_en_W_out ccff_head ccff_tail chany_bottom_in[0] chany_bottom_in[10] chany_bottom_in[11]
+ chany_bottom_in[12] chany_bottom_in[13] chany_bottom_in[14] chany_bottom_in[15]
+ chany_bottom_in[16] chany_bottom_in[17] chany_bottom_in[18] chany_bottom_in[19]
+ chany_bottom_in[1] chany_bottom_in[2] chany_bottom_in[3] chany_bottom_in[4] chany_bottom_in[5]
+ chany_bottom_in[6] chany_bottom_in[7] chany_bottom_in[8] chany_bottom_in[9] chany_bottom_out[0]
+ chany_bottom_out[10] chany_bottom_out[11] chany_bottom_out[12] chany_bottom_out[13]
+ chany_bottom_out[14] chany_bottom_out[15] chany_bottom_out[16] chany_bottom_out[17]
+ chany_bottom_out[18] chany_bottom_out[19] chany_bottom_out[1] chany_bottom_out[2]
+ chany_bottom_out[3] chany_bottom_out[4] chany_bottom_out[5] chany_bottom_out[6]
+ chany_bottom_out[7] chany_bottom_out[8] chany_bottom_out[9] chany_top_in[0] chany_top_in[10]
+ chany_top_in[11] chany_top_in[12] chany_top_in[13] chany_top_in[14] chany_top_in[15]
+ chany_top_in[16] chany_top_in[17] chany_top_in[18] chany_top_in[19] chany_top_in[1]
+ chany_top_in[2] chany_top_in[3] chany_top_in[4] chany_top_in[5] chany_top_in[6]
+ chany_top_in[7] chany_top_in[8] chany_top_in[9] chany_top_out[0] chany_top_out[10]
+ chany_top_out[11] chany_top_out[12] chany_top_out[13] chany_top_out[14] chany_top_out[15]
+ chany_top_out[16] chany_top_out[17] chany_top_out[18] chany_top_out[19] chany_top_out[1]
+ chany_top_out[2] chany_top_out[3] chany_top_out[4] chany_top_out[5] chany_top_out[6]
+ chany_top_out[7] chany_top_out[8] chany_top_out[9] clk_2_N_in clk_2_N_out clk_2_S_in
+ clk_2_S_out clk_3_N_in clk_3_N_out clk_3_S_in clk_3_S_out left_grid_pin_16_ left_grid_pin_17_
+ left_grid_pin_18_ left_grid_pin_19_ left_grid_pin_20_ left_grid_pin_21_ left_grid_pin_22_
+ left_grid_pin_23_ left_grid_pin_24_ left_grid_pin_25_ left_grid_pin_26_ left_grid_pin_27_
+ left_grid_pin_28_ left_grid_pin_29_ left_grid_pin_30_ left_grid_pin_31_ prog_clk_0_N_out
+ prog_clk_0_S_out prog_clk_0_W_in prog_clk_2_N_in prog_clk_2_N_out prog_clk_2_S_in
+ prog_clk_2_S_out prog_clk_3_N_in prog_clk_3_N_out prog_clk_3_S_in prog_clk_3_S_out
+ VPWR VGND
XFILLER_22_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_right_ipin_11.mux_l2_in_0_ mux_right_ipin_11.mux_l1_in_1_/X mux_right_ipin_11.mux_l1_in_0_/X
+ mux_right_ipin_11.mux_l2_in_0_/S VGND VGND VPWR VPWR mux_right_ipin_11.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_12_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_66_ chany_bottom_in[7] VGND VGND VPWR VPWR chany_top_out[7] sky130_fd_sc_hd__buf_2
Xmem_right_ipin_15.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_6_0_mem_right_ipin_0.prog_clk/X
+ mux_right_ipin_15.mux_l1_in_0_/S VGND VGND VPWR VPWR mux_right_ipin_15.mux_l2_in_2_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_2_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_right_ipin_11.mux_l1_in_1_ chany_top_in[3] chany_bottom_in[3] mux_right_ipin_11.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_right_ipin_11.mux_l1_in_1_/X sky130_fd_sc_hd__mux2_1
X_49_ chany_top_in[4] VGND VGND VPWR VPWR chany_bottom_out[4] sky130_fd_sc_hd__buf_2
XFILLER_22_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmem_right_ipin_12.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_7_0_mem_right_ipin_0.prog_clk/X
+ mux_right_ipin_11.mux_l4_in_0_/S VGND VGND VPWR VPWR mux_right_ipin_12.mux_l1_in_2_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_20_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_65_ chany_bottom_in[8] VGND VGND VPWR VPWR chany_top_out[8] sky130_fd_sc_hd__buf_2
Xmux_right_ipin_8.sky130_fd_sc_hd__buf_4_0_ mux_right_ipin_8.mux_l4_in_0_/X VGND VGND
+ VPWR VPWR left_grid_pin_24_ sky130_fd_sc_hd__buf_4
Xmem_right_ipin_15.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_7_0_mem_right_ipin_0.prog_clk/X
+ mux_right_ipin_14.mux_l4_in_0_/S VGND VGND VPWR VPWR mux_right_ipin_15.mux_l1_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_right_ipin_11.mux_l1_in_0_ chany_top_in[1] chany_bottom_in[1] mux_right_ipin_11.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_right_ipin_11.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
X_48_ chany_top_in[5] VGND VGND VPWR VPWR chany_bottom_out[5] sky130_fd_sc_hd__buf_2
XFILLER_18_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_64_ chany_bottom_in[9] VGND VGND VPWR VPWR chany_top_out[9] sky130_fd_sc_hd__buf_2
XFILLER_5_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_right_ipin_3.mux_l2_in_3_ _29_/HI chany_top_in[19] mux_right_ipin_3.mux_l2_in_2_/S
+ VGND VGND VPWR VPWR mux_right_ipin_3.mux_l2_in_3_/X sky130_fd_sc_hd__mux2_1
XFILLER_3_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_47_ chany_top_in[6] VGND VGND VPWR VPWR chany_bottom_out[6] sky130_fd_sc_hd__buf_2
XFILLER_9_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_right_ipin_3.mux_l4_in_0_ mux_right_ipin_3.mux_l3_in_1_/X mux_right_ipin_3.mux_l3_in_0_/X
+ mux_right_ipin_3.mux_l4_in_0_/S VGND VGND VPWR VPWR mux_right_ipin_3.mux_l4_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_25_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmux_right_ipin_8.mux_l2_in_3_ _18_/HI chany_top_in[18] mux_right_ipin_8.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_right_ipin_8.mux_l2_in_3_/X sky130_fd_sc_hd__mux2_1
XFILLER_26_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_right_ipin_3.mux_l3_in_1_ mux_right_ipin_3.mux_l2_in_3_/X mux_right_ipin_3.mux_l2_in_2_/X
+ mux_right_ipin_3.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_right_ipin_3.mux_l3_in_1_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_9_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_63_ chany_bottom_in[10] VGND VGND VPWR VPWR chany_top_out[10] sky130_fd_sc_hd__buf_2
Xmux_right_ipin_3.mux_l2_in_2_ chany_bottom_in[19] chany_top_in[13] mux_right_ipin_3.mux_l2_in_2_/S
+ VGND VGND VPWR VPWR mux_right_ipin_3.mux_l2_in_2_/X sky130_fd_sc_hd__mux2_1
XFILLER_23_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xprog_clk_0_FTB00 prog_clk_0_W_in VGND VGND VPWR VPWR prog_clk_0_FTB00/X sky130_fd_sc_hd__buf_8
Xmux_right_ipin_8.mux_l4_in_0_ mux_right_ipin_8.mux_l3_in_1_/X mux_right_ipin_8.mux_l3_in_0_/X
+ mux_right_ipin_8.mux_l4_in_0_/S VGND VGND VPWR VPWR mux_right_ipin_8.mux_l4_in_0_/X
+ sky130_fd_sc_hd__mux2_1
X_46_ chany_top_in[7] VGND VGND VPWR VPWR chany_bottom_out[7] sky130_fd_sc_hd__buf_2
Xclkbuf_1_0_0_mem_right_ipin_0.prog_clk clkbuf_0_mem_right_ipin_0.prog_clk/X VGND
+ VGND VPWR VPWR clkbuf_2_1_0_mem_right_ipin_0.prog_clk/A sky130_fd_sc_hd__clkbuf_1
Xmux_right_ipin_1.sky130_fd_sc_hd__buf_4_0_ mux_right_ipin_1.mux_l4_in_0_/X VGND VGND
+ VPWR VPWR left_grid_pin_17_ sky130_fd_sc_hd__buf_4
X_29_ VGND VGND VPWR VPWR _29_/HI _29_/LO sky130_fd_sc_hd__conb_1
Xmux_right_ipin_8.mux_l3_in_1_ mux_right_ipin_8.mux_l2_in_3_/X mux_right_ipin_8.mux_l2_in_2_/X
+ mux_right_ipin_8.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_right_ipin_8.mux_l3_in_1_/X
+ sky130_fd_sc_hd__mux2_1
Xprog_clk_3_N_FTB01 prog_clk_3_N_in VGND VGND VPWR VPWR prog_clk_3_N_out sky130_fd_sc_hd__buf_4
XFILLER_19_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_right_ipin_8.mux_l2_in_2_ chany_bottom_in[18] chany_top_in[12] mux_right_ipin_8.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_right_ipin_8.mux_l2_in_2_/X sky130_fd_sc_hd__mux2_1
XFILLER_11_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_right_ipin_3.mux_l3_in_0_ mux_right_ipin_3.mux_l2_in_1_/X mux_right_ipin_3.mux_l2_in_0_/X
+ mux_right_ipin_3.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_right_ipin_3.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_8_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_62_ chany_bottom_in[11] VGND VGND VPWR VPWR chany_top_out[11] sky130_fd_sc_hd__buf_2
Xmux_right_ipin_3.mux_l2_in_1_ chany_bottom_in[13] mux_right_ipin_3.mux_l1_in_2_/X
+ mux_right_ipin_3.mux_l2_in_2_/S VGND VGND VPWR VPWR mux_right_ipin_3.mux_l2_in_1_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_23_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_45_ chany_top_in[8] VGND VGND VPWR VPWR chany_bottom_out[8] sky130_fd_sc_hd__buf_2
Xmux_right_ipin_12.mux_l2_in_3_ _24_/HI chany_top_in[16] mux_right_ipin_12.mux_l2_in_2_/S
+ VGND VGND VPWR VPWR mux_right_ipin_12.mux_l2_in_3_/X sky130_fd_sc_hd__mux2_1
Xmux_right_ipin_3.mux_l1_in_2_ chany_top_in[7] chany_bottom_in[7] mux_right_ipin_3.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR mux_right_ipin_3.mux_l1_in_2_/X sky130_fd_sc_hd__mux2_1
X_28_ VGND VGND VPWR VPWR _28_/HI _28_/LO sky130_fd_sc_hd__conb_1
Xmux_right_ipin_8.mux_l3_in_0_ mux_right_ipin_8.mux_l2_in_1_/X mux_right_ipin_8.mux_l2_in_0_/X
+ mux_right_ipin_8.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_right_ipin_8.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_20_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_right_ipin_8.mux_l2_in_1_ chany_bottom_in[12] mux_right_ipin_8.mux_l1_in_2_/X
+ mux_right_ipin_8.mux_l2_in_3_/S VGND VGND VPWR VPWR mux_right_ipin_8.mux_l2_in_1_/X
+ sky130_fd_sc_hd__mux2_1
Xmux_right_ipin_12.mux_l4_in_0_ mux_right_ipin_12.mux_l3_in_1_/X mux_right_ipin_12.mux_l3_in_0_/X
+ mux_right_ipin_12.mux_l4_in_0_/S VGND VGND VPWR VPWR mux_right_ipin_12.mux_l4_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_26_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_right_ipin_8.mux_l1_in_2_ chany_top_in[8] chany_bottom_in[8] mux_right_ipin_8.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR mux_right_ipin_8.mux_l1_in_2_/X sky130_fd_sc_hd__mux2_1
X_61_ chany_bottom_in[12] VGND VGND VPWR VPWR chany_top_out[12] sky130_fd_sc_hd__buf_2
Xmux_right_ipin_12.mux_l3_in_1_ mux_right_ipin_12.mux_l2_in_3_/X mux_right_ipin_12.mux_l2_in_2_/X
+ mux_right_ipin_12.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_right_ipin_12.mux_l3_in_1_/X
+ sky130_fd_sc_hd__mux2_1
Xmux_right_ipin_3.mux_l2_in_0_ mux_right_ipin_3.mux_l1_in_1_/X mux_right_ipin_3.mux_l1_in_0_/X
+ mux_right_ipin_3.mux_l2_in_2_/S VGND VGND VPWR VPWR mux_right_ipin_3.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_5_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_44_ chany_top_in[9] VGND VGND VPWR VPWR chany_bottom_out[9] sky130_fd_sc_hd__buf_2
Xmux_right_ipin_12.mux_l2_in_2_ chany_bottom_in[16] chany_top_in[12] mux_right_ipin_12.mux_l2_in_2_/S
+ VGND VGND VPWR VPWR mux_right_ipin_12.mux_l2_in_2_/X sky130_fd_sc_hd__mux2_1
XFILLER_18_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_right_ipin_3.mux_l1_in_1_ chany_top_in[3] chany_bottom_in[3] mux_right_ipin_3.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR mux_right_ipin_3.mux_l1_in_1_/X sky130_fd_sc_hd__mux2_1
X_27_ VGND VGND VPWR VPWR _27_/HI _27_/LO sky130_fd_sc_hd__conb_1
XFILLER_19_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmux_right_ipin_8.mux_l2_in_0_ mux_right_ipin_8.mux_l1_in_1_/X mux_right_ipin_8.mux_l1_in_0_/X
+ mux_right_ipin_8.mux_l2_in_3_/S VGND VGND VPWR VPWR mux_right_ipin_8.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XPHY_0 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_right_ipin_8.mux_l1_in_1_ chany_top_in[2] chany_bottom_in[2] mux_right_ipin_8.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR mux_right_ipin_8.mux_l1_in_1_/X sky130_fd_sc_hd__mux2_1
XFILLER_12_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_60_ chany_bottom_in[13] VGND VGND VPWR VPWR chany_top_out[13] sky130_fd_sc_hd__buf_2
Xmux_right_ipin_12.mux_l3_in_0_ mux_right_ipin_12.mux_l2_in_1_/X mux_right_ipin_12.mux_l2_in_0_/X
+ mux_right_ipin_12.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_right_ipin_12.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_23_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_43_ chany_top_in[10] VGND VGND VPWR VPWR chany_bottom_out[10] sky130_fd_sc_hd__buf_2
Xmux_right_ipin_12.mux_l2_in_1_ chany_bottom_in[12] mux_right_ipin_12.mux_l1_in_2_/X
+ mux_right_ipin_12.mux_l2_in_2_/S VGND VGND VPWR VPWR mux_right_ipin_12.mux_l2_in_1_/X
+ sky130_fd_sc_hd__mux2_1
Xprog_clk_2_S_FTB01 prog_clk_2_N_in VGND VGND VPWR VPWR prog_clk_2_S_out sky130_fd_sc_hd__buf_4
Xmux_right_ipin_3.mux_l1_in_0_ chany_top_in[1] chany_bottom_in[1] mux_right_ipin_3.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR mux_right_ipin_3.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_27_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_3_2_0_mem_right_ipin_0.prog_clk clkbuf_3_3_0_mem_right_ipin_0.prog_clk/A VGND
+ VGND VPWR VPWR clkbuf_3_2_0_mem_right_ipin_0.prog_clk/X sky130_fd_sc_hd__clkbuf_1
X_26_ VGND VGND VPWR VPWR _26_/HI _26_/LO sky130_fd_sc_hd__conb_1
XFILLER_20_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_right_ipin_12.mux_l1_in_2_ chany_top_in[6] chany_bottom_in[6] mux_right_ipin_12.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR mux_right_ipin_12.mux_l1_in_2_/X sky130_fd_sc_hd__mux2_1
XPHY_121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmem_right_ipin_0.sky130_fd_sc_hd__dfxtp_1_3_ clkbuf_3_0_0_mem_right_ipin_0.prog_clk/X
+ mux_right_ipin_0.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_right_ipin_0.mux_l4_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
Xmux_right_ipin_8.mux_l1_in_0_ chany_top_in[0] chany_bottom_in[0] mux_right_ipin_8.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR mux_right_ipin_8.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
Xclkbuf_3_5_0_mem_right_ipin_0.prog_clk clkbuf_3_5_0_mem_right_ipin_0.prog_clk/A VGND
+ VGND VPWR VPWR clkbuf_3_5_0_mem_right_ipin_0.prog_clk/X sky130_fd_sc_hd__clkbuf_1
XFILLER_23_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_42_ chany_top_in[11] VGND VGND VPWR VPWR chany_bottom_out[11] sky130_fd_sc_hd__buf_2
Xmux_right_ipin_12.mux_l2_in_0_ mux_right_ipin_12.mux_l1_in_1_/X mux_right_ipin_12.mux_l1_in_0_/X
+ mux_right_ipin_12.mux_l2_in_2_/S VGND VGND VPWR VPWR mux_right_ipin_12.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_18_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25_ VGND VGND VPWR VPWR _25_/HI _25_/LO sky130_fd_sc_hd__conb_1
Xmux_right_ipin_12.sky130_fd_sc_hd__buf_4_0_ mux_right_ipin_12.mux_l4_in_0_/X VGND
+ VGND VPWR VPWR left_grid_pin_28_ sky130_fd_sc_hd__buf_4
XFILLER_25_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_right_ipin_12.mux_l1_in_1_ chany_top_in[2] chany_bottom_in[2] mux_right_ipin_12.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR mux_right_ipin_12.mux_l1_in_1_/X sky130_fd_sc_hd__mux2_1
Xmux_right_ipin_4.sky130_fd_sc_hd__buf_4_0_ mux_right_ipin_4.mux_l4_in_0_/X VGND VGND
+ VPWR VPWR left_grid_pin_20_ sky130_fd_sc_hd__buf_4
Xmem_right_ipin_3.sky130_fd_sc_hd__dfxtp_1_3_ clkbuf_3_1_0_mem_right_ipin_0.prog_clk/X
+ mux_right_ipin_3.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_right_ipin_3.mux_l4_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_25_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmem_right_ipin_0.sky130_fd_sc_hd__dfxtp_1_2_ clkbuf_3_0_0_mem_right_ipin_0.prog_clk/X
+ mux_right_ipin_0.mux_l2_in_3_/S VGND VGND VPWR VPWR mux_right_ipin_0.mux_l3_in_1_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_12_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_41_ chany_top_in[12] VGND VGND VPWR VPWR chany_bottom_out[12] sky130_fd_sc_hd__buf_2
Xmem_right_ipin_6.sky130_fd_sc_hd__dfxtp_1_3_ clkbuf_3_3_0_mem_right_ipin_0.prog_clk/X
+ mux_right_ipin_6.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_right_ipin_6.mux_l4_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
X_24_ VGND VGND VPWR VPWR _24_/HI _24_/LO sky130_fd_sc_hd__conb_1
Xmem_right_ipin_3.sky130_fd_sc_hd__dfxtp_1_2_ clkbuf_3_3_0_mem_right_ipin_0.prog_clk/X
+ mux_right_ipin_3.mux_l2_in_2_/S VGND VGND VPWR VPWR mux_right_ipin_3.mux_l3_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
Xmux_right_ipin_12.mux_l1_in_0_ chany_top_in[0] chany_bottom_in[0] mux_right_ipin_12.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR mux_right_ipin_12.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XPHY_123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmem_right_ipin_0.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_2_0_mem_right_ipin_0.prog_clk/X
+ mux_right_ipin_0.mux_l1_in_2_/S VGND VGND VPWR VPWR mux_right_ipin_0.mux_l2_in_3_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_8_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmem_right_ipin_9.sky130_fd_sc_hd__dfxtp_1_3_ clkbuf_3_4_0_mem_right_ipin_0.prog_clk/X
+ mux_right_ipin_9.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_right_ipin_9.mux_l4_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
Xmem_right_ipin_11.sky130_fd_sc_hd__dfxtp_1_3_ clkbuf_3_5_0_mem_right_ipin_0.prog_clk/X
+ mux_right_ipin_11.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_right_ipin_11.mux_l4_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
X_40_ chany_top_in[13] VGND VGND VPWR VPWR chany_bottom_out[13] sky130_fd_sc_hd__buf_2
Xmem_right_ipin_6.sky130_fd_sc_hd__dfxtp_1_2_ clkbuf_3_1_0_mem_right_ipin_0.prog_clk/X
+ mux_right_ipin_6.mux_l2_in_1_/S VGND VGND VPWR VPWR mux_right_ipin_6.mux_l3_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
X_23_ VGND VGND VPWR VPWR _23_/HI _23_/LO sky130_fd_sc_hd__conb_1
Xmux_right_ipin_4.mux_l2_in_3_ _30_/HI chany_top_in[14] mux_right_ipin_4.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_right_ipin_4.mux_l2_in_3_/X sky130_fd_sc_hd__mux2_1
XTest_en_E_FTB01 Test_en_E_in VGND VGND VPWR VPWR Test_en_E_out sky130_fd_sc_hd__buf_4
Xmem_right_ipin_3.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_2_0_mem_right_ipin_0.prog_clk/X
+ mux_right_ipin_3.mux_l1_in_2_/S VGND VGND VPWR VPWR mux_right_ipin_3.mux_l2_in_2_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_25_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmux_right_ipin_4.mux_l4_in_0_ mux_right_ipin_4.mux_l3_in_1_/X mux_right_ipin_4.mux_l3_in_0_/X
+ mux_right_ipin_4.mux_l4_in_0_/S VGND VGND VPWR VPWR mux_right_ipin_4.mux_l4_in_0_/X
+ sky130_fd_sc_hd__mux2_1
Xmem_right_ipin_0.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_0_0_mem_right_ipin_0.prog_clk/X
+ ccff_head VGND VGND VPWR VPWR mux_right_ipin_0.mux_l1_in_2_/S sky130_fd_sc_hd__dfxtp_1
Xmem_right_ipin_14.sky130_fd_sc_hd__dfxtp_1_3_ clkbuf_3_5_0_mem_right_ipin_0.prog_clk/X
+ mux_right_ipin_14.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_right_ipin_14.mux_l4_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_12_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmem_right_ipin_9.sky130_fd_sc_hd__dfxtp_1_2_ clkbuf_3_1_0_mem_right_ipin_0.prog_clk/X
+ mux_right_ipin_9.mux_l2_in_1_/S VGND VGND VPWR VPWR mux_right_ipin_9.mux_l3_in_1_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_27_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_right_ipin_9.mux_l2_in_3_ _19_/HI chany_top_in[13] mux_right_ipin_9.mux_l2_in_1_/S
+ VGND VGND VPWR VPWR mux_right_ipin_9.mux_l2_in_3_/X sky130_fd_sc_hd__mux2_1
Xmux_right_ipin_4.mux_l3_in_1_ mux_right_ipin_4.mux_l2_in_3_/X mux_right_ipin_4.mux_l2_in_2_/X
+ mux_right_ipin_4.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_right_ipin_4.mux_l3_in_1_/X
+ sky130_fd_sc_hd__mux2_1
Xmem_right_ipin_11.sky130_fd_sc_hd__dfxtp_1_2_ clkbuf_3_7_0_mem_right_ipin_0.prog_clk/X
+ mux_right_ipin_11.mux_l2_in_0_/S VGND VGND VPWR VPWR mux_right_ipin_11.mux_l3_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_1_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmem_right_ipin_6.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_3_0_mem_right_ipin_0.prog_clk/X
+ mux_right_ipin_6.mux_l1_in_0_/S VGND VGND VPWR VPWR mux_right_ipin_6.mux_l2_in_1_/S
+ sky130_fd_sc_hd__dfxtp_1
X_22_ VGND VGND VPWR VPWR _22_/HI _22_/LO sky130_fd_sc_hd__conb_1
XFILLER_1_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_right_ipin_4.mux_l2_in_2_ chany_bottom_in[14] chany_top_in[8] mux_right_ipin_4.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_right_ipin_4.mux_l2_in_2_/X sky130_fd_sc_hd__mux2_1
Xmux_right_ipin_9.mux_l4_in_0_ mux_right_ipin_9.mux_l3_in_1_/X mux_right_ipin_9.mux_l3_in_0_/X
+ mux_right_ipin_9.mux_l4_in_0_/S VGND VGND VPWR VPWR mux_right_ipin_9.mux_l4_in_0_/X
+ sky130_fd_sc_hd__mux2_1
Xmem_right_ipin_3.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_0_0_mem_right_ipin_0.prog_clk/X
+ mux_right_ipin_2.mux_l4_in_0_/S VGND VGND VPWR VPWR mux_right_ipin_3.mux_l1_in_2_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_18_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_right_ipin_9.mux_l3_in_1_ mux_right_ipin_9.mux_l2_in_3_/X mux_right_ipin_9.mux_l2_in_2_/X
+ mux_right_ipin_9.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_right_ipin_9.mux_l3_in_1_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_21_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmem_right_ipin_14.sky130_fd_sc_hd__dfxtp_1_2_ clkbuf_3_5_0_mem_right_ipin_0.prog_clk/X
+ mux_right_ipin_14.mux_l2_in_3_/S VGND VGND VPWR VPWR mux_right_ipin_14.mux_l3_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_8_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmem_right_ipin_9.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_6_0_mem_right_ipin_0.prog_clk/X
+ mux_right_ipin_9.mux_l1_in_0_/S VGND VGND VPWR VPWR mux_right_ipin_9.mux_l2_in_1_/S
+ sky130_fd_sc_hd__dfxtp_1
Xclkbuf_2_2_0_mem_right_ipin_0.prog_clk clkbuf_2_2_0_mem_right_ipin_0.prog_clk/A VGND
+ VGND VPWR VPWR clkbuf_3_5_0_mem_right_ipin_0.prog_clk/A sky130_fd_sc_hd__clkbuf_1
Xmux_right_ipin_9.mux_l2_in_2_ chany_bottom_in[13] chany_top_in[5] mux_right_ipin_9.mux_l2_in_1_/S
+ VGND VGND VPWR VPWR mux_right_ipin_9.mux_l2_in_2_/X sky130_fd_sc_hd__mux2_1
XFILLER_5_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_right_ipin_4.mux_l3_in_0_ mux_right_ipin_4.mux_l2_in_1_/X mux_right_ipin_4.mux_l2_in_0_/X
+ mux_right_ipin_4.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_right_ipin_4.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
Xmem_right_ipin_11.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_7_0_mem_right_ipin_0.prog_clk/X
+ mux_right_ipin_11.mux_l1_in_0_/S VGND VGND VPWR VPWR mux_right_ipin_11.mux_l2_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
Xclk_3_S_FTB01 clk_3_N_in VGND VGND VPWR VPWR clk_3_S_out sky130_fd_sc_hd__buf_4
XFILLER_1_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmem_right_ipin_6.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_1_0_mem_right_ipin_0.prog_clk/X
+ mux_right_ipin_5.mux_l4_in_0_/S VGND VGND VPWR VPWR mux_right_ipin_6.mux_l1_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
X_21_ VGND VGND VPWR VPWR _21_/HI _21_/LO sky130_fd_sc_hd__conb_1
Xmux_right_ipin_4.mux_l2_in_1_ chany_bottom_in[8] mux_right_ipin_4.mux_l1_in_2_/X
+ mux_right_ipin_4.mux_l2_in_3_/S VGND VGND VPWR VPWR mux_right_ipin_4.mux_l2_in_1_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_1_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_right_ipin_15.sky130_fd_sc_hd__buf_4_0_ mux_right_ipin_15.mux_l4_in_0_/X VGND
+ VGND VPWR VPWR left_grid_pin_31_ sky130_fd_sc_hd__buf_4
Xmux_right_ipin_13.mux_l2_in_3_ _25_/HI chany_top_in[17] mux_right_ipin_13.mux_l2_in_2_/S
+ VGND VGND VPWR VPWR mux_right_ipin_13.mux_l2_in_3_/X sky130_fd_sc_hd__mux2_1
XPHY_126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmux_right_ipin_4.mux_l1_in_2_ chany_top_in[4] chany_bottom_in[4] mux_right_ipin_4.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_right_ipin_4.mux_l1_in_2_/X sky130_fd_sc_hd__mux2_1
Xmux_right_ipin_7.sky130_fd_sc_hd__buf_4_0_ mux_right_ipin_7.mux_l4_in_0_/X VGND VGND
+ VPWR VPWR left_grid_pin_23_ sky130_fd_sc_hd__buf_4
XFILLER_15_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_right_ipin_9.mux_l3_in_0_ mux_right_ipin_9.mux_l2_in_1_/X mux_right_ipin_9.mux_l2_in_0_/X
+ mux_right_ipin_9.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_right_ipin_9.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
Xmem_right_ipin_14.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_6_0_mem_right_ipin_0.prog_clk/X
+ mux_right_ipin_14.mux_l1_in_0_/S VGND VGND VPWR VPWR mux_right_ipin_14.mux_l2_in_3_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_8_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmem_right_ipin_9.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_6_0_mem_right_ipin_0.prog_clk/X
+ mux_right_ipin_8.mux_l4_in_0_/S VGND VGND VPWR VPWR mux_right_ipin_9.mux_l1_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
Xmux_right_ipin_9.mux_l2_in_1_ chany_bottom_in[5] chany_top_in[3] mux_right_ipin_9.mux_l2_in_1_/S
+ VGND VGND VPWR VPWR mux_right_ipin_9.mux_l2_in_1_/X sky130_fd_sc_hd__mux2_1
XFILLER_27_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_right_ipin_13.mux_l4_in_0_ mux_right_ipin_13.mux_l3_in_1_/X mux_right_ipin_13.mux_l3_in_0_/X
+ mux_right_ipin_13.mux_l4_in_0_/S VGND VGND VPWR VPWR mux_right_ipin_13.mux_l4_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_4_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmem_right_ipin_11.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_5_0_mem_right_ipin_0.prog_clk/X
+ mux_right_ipin_10.mux_l4_in_0_/S VGND VGND VPWR VPWR mux_right_ipin_11.mux_l1_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
Xmux_right_ipin_13.mux_l3_in_1_ mux_right_ipin_13.mux_l2_in_3_/X mux_right_ipin_13.mux_l2_in_2_/X
+ mux_right_ipin_13.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_right_ipin_13.mux_l3_in_1_/X
+ sky130_fd_sc_hd__mux2_1
Xmux_right_ipin_4.mux_l2_in_0_ mux_right_ipin_4.mux_l1_in_1_/X mux_right_ipin_4.mux_l1_in_0_/X
+ mux_right_ipin_4.mux_l2_in_3_/S VGND VGND VPWR VPWR mux_right_ipin_4.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_1_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20_ VGND VGND VPWR VPWR _20_/HI _20_/LO sky130_fd_sc_hd__conb_1
XFILLER_19_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_right_ipin_13.mux_l2_in_2_ chany_bottom_in[17] chany_top_in[9] mux_right_ipin_13.mux_l2_in_2_/S
+ VGND VGND VPWR VPWR mux_right_ipin_13.mux_l2_in_2_/X sky130_fd_sc_hd__mux2_1
XFILLER_24_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmux_right_ipin_4.mux_l1_in_1_ chany_top_in[2] chany_bottom_in[2] mux_right_ipin_4.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_right_ipin_4.mux_l1_in_1_/X sky130_fd_sc_hd__mux2_1
XPHY_127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xprog_clk_2_N_FTB01 prog_clk_2_N_in VGND VGND VPWR VPWR prog_clk_2_N_out sky130_fd_sc_hd__buf_4
XFILLER_24_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmem_right_ipin_14.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_6_0_mem_right_ipin_0.prog_clk/X
+ mux_right_ipin_13.mux_l4_in_0_/S VGND VGND VPWR VPWR mux_right_ipin_14.mux_l1_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_16_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_right_ipin_9.mux_l2_in_0_ chany_bottom_in[3] mux_right_ipin_9.mux_l1_in_0_/X
+ mux_right_ipin_9.mux_l2_in_1_/S VGND VGND VPWR VPWR mux_right_ipin_9.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_27_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_right_ipin_13.mux_l3_in_0_ mux_right_ipin_13.mux_l2_in_1_/X mux_right_ipin_13.mux_l2_in_0_/X
+ mux_right_ipin_13.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_right_ipin_13.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_24_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_right_ipin_13.mux_l2_in_1_ chany_bottom_in[9] chany_top_in[3] mux_right_ipin_13.mux_l2_in_2_/S
+ VGND VGND VPWR VPWR mux_right_ipin_13.mux_l2_in_1_/X sky130_fd_sc_hd__mux2_1
XFILLER_18_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_right_ipin_4.mux_l1_in_0_ chany_top_in[0] chany_bottom_in[0] mux_right_ipin_4.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_right_ipin_4.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XPHY_128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_right_ipin_0.sky130_fd_sc_hd__buf_4_0_ mux_right_ipin_0.mux_l4_in_0_/X VGND VGND
+ VPWR VPWR left_grid_pin_16_ sky130_fd_sc_hd__buf_4
XFILLER_4_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_right_ipin_9.mux_l1_in_0_ chany_top_in[1] chany_bottom_in[1] mux_right_ipin_9.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_right_ipin_9.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_24_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmux_right_ipin_13.mux_l2_in_0_ chany_bottom_in[3] mux_right_ipin_13.mux_l1_in_0_/X
+ mux_right_ipin_13.mux_l2_in_2_/S VGND VGND VPWR VPWR mux_right_ipin_13.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XPHY_118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_77_ prog_clk_3_N_in VGND VGND VPWR VPWR prog_clk_3_S_in sky130_fd_sc_hd__buf_2
XFILLER_19_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_right_ipin_13.mux_l1_in_0_ chany_top_in[1] chany_bottom_in[1] mux_right_ipin_13.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_right_ipin_13.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_21_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_right_ipin_0.mux_l2_in_3_ _20_/HI chany_top_in[16] mux_right_ipin_0.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_right_ipin_0.mux_l2_in_3_/X sky130_fd_sc_hd__mux2_1
XFILLER_1_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_76_ prog_clk_2_N_in VGND VGND VPWR VPWR prog_clk_2_S_in sky130_fd_sc_hd__buf_2
XFILLER_14_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_right_ipin_0.mux_l4_in_0_ mux_right_ipin_0.mux_l3_in_1_/X mux_right_ipin_0.mux_l3_in_0_/X
+ mux_right_ipin_0.mux_l4_in_0_/S VGND VGND VPWR VPWR mux_right_ipin_0.mux_l4_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_10_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_59_ chany_bottom_in[14] VGND VGND VPWR VPWR chany_top_out[14] sky130_fd_sc_hd__buf_2
XPHY_109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmux_right_ipin_5.mux_l2_in_3_ _31_/HI chany_top_in[17] mux_right_ipin_5.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_right_ipin_5.mux_l2_in_3_/X sky130_fd_sc_hd__mux2_1
XFILLER_11_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_right_ipin_0.mux_l3_in_1_ mux_right_ipin_0.mux_l2_in_3_/X mux_right_ipin_0.mux_l2_in_2_/X
+ mux_right_ipin_0.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_right_ipin_0.mux_l3_in_1_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_16_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_right_ipin_0.mux_l2_in_2_ chany_bottom_in[16] chany_top_in[10] mux_right_ipin_0.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_right_ipin_0.mux_l2_in_2_/X sky130_fd_sc_hd__mux2_1
XFILLER_4_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_right_ipin_5.mux_l4_in_0_ mux_right_ipin_5.mux_l3_in_1_/X mux_right_ipin_5.mux_l3_in_0_/X
+ mux_right_ipin_5.mux_l4_in_0_/S VGND VGND VPWR VPWR mux_right_ipin_5.mux_l4_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_24_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_right_ipin_5.mux_l3_in_1_ mux_right_ipin_5.mux_l2_in_3_/X mux_right_ipin_5.mux_l2_in_2_/X
+ mux_right_ipin_5.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_right_ipin_5.mux_l3_in_1_/X
+ sky130_fd_sc_hd__mux2_1
X_75_ clk_3_N_in VGND VGND VPWR VPWR clk_3_S_in sky130_fd_sc_hd__buf_2
XFILLER_10_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_58_ chany_bottom_in[15] VGND VGND VPWR VPWR chany_top_out[15] sky130_fd_sc_hd__buf_2
XFILLER_24_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_90 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclk_3_N_FTB01 clk_3_N_in VGND VGND VPWR VPWR clk_3_N_out sky130_fd_sc_hd__buf_4
XFILLER_21_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_right_ipin_5.mux_l2_in_2_ chany_bottom_in[17] chany_top_in[9] mux_right_ipin_5.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_right_ipin_5.mux_l2_in_2_/X sky130_fd_sc_hd__mux2_1
XFILLER_21_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_right_ipin_0.mux_l3_in_0_ mux_right_ipin_0.mux_l2_in_1_/X mux_right_ipin_0.mux_l2_in_0_/X
+ mux_right_ipin_0.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_right_ipin_0.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_7_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_right_ipin_11.sky130_fd_sc_hd__buf_4_0_ mux_right_ipin_11.mux_l4_in_0_/X VGND
+ VGND VPWR VPWR left_grid_pin_27_ sky130_fd_sc_hd__buf_4
Xmux_right_ipin_0.mux_l2_in_1_ chany_bottom_in[10] mux_right_ipin_0.mux_l1_in_2_/X
+ mux_right_ipin_0.mux_l2_in_3_/S VGND VGND VPWR VPWR mux_right_ipin_0.mux_l2_in_1_/X
+ sky130_fd_sc_hd__mux2_1
Xclkbuf_3_1_0_mem_right_ipin_0.prog_clk clkbuf_3_1_0_mem_right_ipin_0.prog_clk/A VGND
+ VGND VPWR VPWR clkbuf_3_1_0_mem_right_ipin_0.prog_clk/X sky130_fd_sc_hd__clkbuf_1
Xmux_right_ipin_3.sky130_fd_sc_hd__buf_4_0_ mux_right_ipin_3.mux_l4_in_0_/X VGND VGND
+ VPWR VPWR left_grid_pin_19_ sky130_fd_sc_hd__buf_4
XFILLER_1_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_right_ipin_0.mux_l1_in_2_ chany_top_in[4] chany_bottom_in[4] mux_right_ipin_0.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR mux_right_ipin_0.mux_l1_in_2_/X sky130_fd_sc_hd__mux2_1
Xmux_right_ipin_5.mux_l3_in_0_ mux_right_ipin_5.mux_l2_in_1_/X mux_right_ipin_5.mux_l2_in_0_/X
+ mux_right_ipin_5.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_right_ipin_5.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
X_74_ clk_2_N_in VGND VGND VPWR VPWR clk_2_S_in sky130_fd_sc_hd__buf_2
XFILLER_19_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_91 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_80 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_57_ chany_bottom_in[16] VGND VGND VPWR VPWR chany_top_out[16] sky130_fd_sc_hd__buf_2
Xmux_right_ipin_5.mux_l2_in_1_ chany_bottom_in[9] chany_top_in[3] mux_right_ipin_5.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_right_ipin_5.mux_l2_in_1_/X sky130_fd_sc_hd__mux2_1
Xclkbuf_3_4_0_mem_right_ipin_0.prog_clk clkbuf_3_5_0_mem_right_ipin_0.prog_clk/A VGND
+ VGND VPWR VPWR clkbuf_3_4_0_mem_right_ipin_0.prog_clk/X sky130_fd_sc_hd__clkbuf_1
XFILLER_16_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_right_ipin_14.mux_l2_in_3_ _26_/HI chany_top_in[18] mux_right_ipin_14.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_right_ipin_14.mux_l2_in_3_/X sky130_fd_sc_hd__mux2_1
Xmux_right_ipin_0.mux_l2_in_0_ mux_right_ipin_0.mux_l1_in_1_/X mux_right_ipin_0.mux_l1_in_0_/X
+ mux_right_ipin_0.mux_l2_in_3_/S VGND VGND VPWR VPWR mux_right_ipin_0.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_4_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmem_right_ipin_2.sky130_fd_sc_hd__dfxtp_1_3_ clkbuf_3_0_0_mem_right_ipin_0.prog_clk/X
+ mux_right_ipin_2.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_right_ipin_2.mux_l4_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
Xmux_right_ipin_14.mux_l4_in_0_ mux_right_ipin_14.mux_l3_in_1_/X mux_right_ipin_14.mux_l3_in_0_/X
+ mux_right_ipin_14.mux_l4_in_0_/S VGND VGND VPWR VPWR mux_right_ipin_14.mux_l4_in_0_/X
+ sky130_fd_sc_hd__mux2_1
Xmux_right_ipin_0.mux_l1_in_1_ chany_top_in[2] chany_bottom_in[2] mux_right_ipin_0.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR mux_right_ipin_0.mux_l1_in_1_/X sky130_fd_sc_hd__mux2_1
XFILLER_6_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_73_ chany_bottom_in[0] VGND VGND VPWR VPWR chany_top_out[0] sky130_fd_sc_hd__buf_2
XFILLER_27_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_3_7_0_mem_right_ipin_0.prog_clk clkbuf_3_7_0_mem_right_ipin_0.prog_clk/A VGND
+ VGND VPWR VPWR clkbuf_3_7_0_mem_right_ipin_0.prog_clk/X sky130_fd_sc_hd__clkbuf_1
XPHY_92 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_70 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_81 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_56_ chany_bottom_in[17] VGND VGND VPWR VPWR chany_top_out[17] sky130_fd_sc_hd__buf_2
Xmux_right_ipin_14.mux_l3_in_1_ mux_right_ipin_14.mux_l2_in_3_/X mux_right_ipin_14.mux_l2_in_2_/X
+ mux_right_ipin_14.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_right_ipin_14.mux_l3_in_1_/X
+ sky130_fd_sc_hd__mux2_1
Xmux_right_ipin_5.mux_l2_in_0_ chany_bottom_in[3] mux_right_ipin_5.mux_l1_in_0_/X
+ mux_right_ipin_5.mux_l2_in_3_/S VGND VGND VPWR VPWR mux_right_ipin_5.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_15_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_39_ chany_top_in[14] VGND VGND VPWR VPWR chany_bottom_out[14] sky130_fd_sc_hd__buf_2
Xmux_right_ipin_14.mux_l2_in_2_ chany_bottom_in[18] chany_top_in[10] mux_right_ipin_14.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_right_ipin_14.mux_l2_in_2_/X sky130_fd_sc_hd__mux2_1
XFILLER_11_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmem_right_ipin_5.sky130_fd_sc_hd__dfxtp_1_3_ clkbuf_3_1_0_mem_right_ipin_0.prog_clk/X
+ mux_right_ipin_5.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_right_ipin_5.mux_l4_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_4_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_right_ipin_2.sky130_fd_sc_hd__dfxtp_1_2_ clkbuf_3_2_0_mem_right_ipin_0.prog_clk/X
+ mux_right_ipin_2.mux_l2_in_2_/S VGND VGND VPWR VPWR mux_right_ipin_2.mux_l3_in_1_/S
+ sky130_fd_sc_hd__dfxtp_1
Xmux_right_ipin_0.mux_l1_in_0_ chany_top_in[0] chany_bottom_in[0] mux_right_ipin_0.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR mux_right_ipin_0.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
X_72_ chany_bottom_in[1] VGND VGND VPWR VPWR chany_top_out[1] sky130_fd_sc_hd__buf_2
Xclk_2_S_FTB01 clk_2_N_in VGND VGND VPWR VPWR clk_2_S_out sky130_fd_sc_hd__buf_4
XFILLER_14_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_60 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_71 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_82 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_93 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_55_ chany_bottom_in[18] VGND VGND VPWR VPWR chany_top_out[18] sky130_fd_sc_hd__buf_2
XFILLER_24_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmux_right_ipin_14.mux_l3_in_0_ mux_right_ipin_14.mux_l2_in_1_/X mux_right_ipin_14.mux_l2_in_0_/X
+ mux_right_ipin_14.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_right_ipin_14.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_23_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmem_right_ipin_8.sky130_fd_sc_hd__dfxtp_1_3_ clkbuf_3_1_0_mem_right_ipin_0.prog_clk/X
+ mux_right_ipin_8.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_right_ipin_8.mux_l4_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_20_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_38_ chany_top_in[15] VGND VGND VPWR VPWR chany_bottom_out[15] sky130_fd_sc_hd__buf_2
Xmem_right_ipin_10.sky130_fd_sc_hd__dfxtp_1_3_ clkbuf_3_4_0_mem_right_ipin_0.prog_clk/X
+ mux_right_ipin_10.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_right_ipin_10.mux_l4_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_11_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_right_ipin_14.mux_l2_in_1_ chany_bottom_in[10] chany_top_in[2] mux_right_ipin_14.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_right_ipin_14.mux_l2_in_1_/X sky130_fd_sc_hd__mux2_1
Xmux_right_ipin_5.mux_l1_in_0_ chany_top_in[1] chany_bottom_in[1] mux_right_ipin_5.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_right_ipin_5.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
Xmem_right_ipin_5.sky130_fd_sc_hd__dfxtp_1_2_ clkbuf_3_3_0_mem_right_ipin_0.prog_clk/X
+ mux_right_ipin_5.mux_l2_in_3_/S VGND VGND VPWR VPWR mux_right_ipin_5.mux_l3_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_4_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmem_right_ipin_2.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_2_0_mem_right_ipin_0.prog_clk/X
+ mux_right_ipin_2.mux_l1_in_0_/S VGND VGND VPWR VPWR mux_right_ipin_2.mux_l2_in_2_/S
+ sky130_fd_sc_hd__dfxtp_1
X_71_ chany_bottom_in[2] VGND VGND VPWR VPWR chany_top_out[2] sky130_fd_sc_hd__buf_2
XFILLER_27_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_94 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_61 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_72 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_83 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_54_ chany_bottom_in[19] VGND VGND VPWR VPWR chany_top_out[19] sky130_fd_sc_hd__buf_2
Xmem_right_ipin_13.sky130_fd_sc_hd__dfxtp_1_3_ clkbuf_3_5_0_mem_right_ipin_0.prog_clk/X
+ mux_right_ipin_13.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_right_ipin_13.mux_l4_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_2_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmem_right_ipin_8.sky130_fd_sc_hd__dfxtp_1_2_ clkbuf_3_3_0_mem_right_ipin_0.prog_clk/X
+ mux_right_ipin_8.mux_l2_in_3_/S VGND VGND VPWR VPWR mux_right_ipin_8.mux_l3_in_1_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_14_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_37_ chany_top_in[16] VGND VGND VPWR VPWR chany_bottom_out[16] sky130_fd_sc_hd__buf_2
Xmem_right_ipin_10.sky130_fd_sc_hd__dfxtp_1_2_ clkbuf_3_4_0_mem_right_ipin_0.prog_clk/X
+ mux_right_ipin_10.mux_l2_in_0_/S VGND VGND VPWR VPWR mux_right_ipin_10.mux_l3_in_1_/S
+ sky130_fd_sc_hd__dfxtp_1
Xmux_right_ipin_14.mux_l2_in_0_ chany_bottom_in[2] mux_right_ipin_14.mux_l1_in_0_/X
+ mux_right_ipin_14.mux_l2_in_3_/S VGND VGND VPWR VPWR mux_right_ipin_14.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
Xmem_right_ipin_5.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_2_0_mem_right_ipin_0.prog_clk/X
+ mux_right_ipin_5.mux_l1_in_0_/S VGND VGND VPWR VPWR mux_right_ipin_5.mux_l2_in_3_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_8_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmux_right_ipin_14.sky130_fd_sc_hd__buf_4_0_ mux_right_ipin_14.mux_l4_in_0_/X VGND
+ VGND VPWR VPWR left_grid_pin_30_ sky130_fd_sc_hd__buf_4
Xmux_right_ipin_6.sky130_fd_sc_hd__buf_4_0_ mux_right_ipin_6.mux_l4_in_0_/X VGND VGND
+ VPWR VPWR left_grid_pin_22_ sky130_fd_sc_hd__buf_4
XFILLER_0_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmem_right_ipin_2.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_0_0_mem_right_ipin_0.prog_clk/X
+ mux_right_ipin_1.mux_l4_in_0_/S VGND VGND VPWR VPWR mux_right_ipin_2.mux_l1_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_5_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_70_ chany_bottom_in[3] VGND VGND VPWR VPWR chany_top_out[3] sky130_fd_sc_hd__buf_2
XTest_en_W_FTB01 Test_en_E_in VGND VGND VPWR VPWR Test_en_W_out sky130_fd_sc_hd__buf_4
XFILLER_18_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmem_right_ipin_13.sky130_fd_sc_hd__dfxtp_1_2_ clkbuf_3_7_0_mem_right_ipin_0.prog_clk/X
+ mux_right_ipin_13.mux_l2_in_2_/S VGND VGND VPWR VPWR mux_right_ipin_13.mux_l3_in_1_/S
+ sky130_fd_sc_hd__dfxtp_1
XPHY_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_95 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_62 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_53_ chany_top_in[0] VGND VGND VPWR VPWR chany_bottom_out[0] sky130_fd_sc_hd__buf_2
XPHY_73 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_84 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmem_right_ipin_8.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_3_0_mem_right_ipin_0.prog_clk/X
+ mux_right_ipin_8.mux_l1_in_2_/S VGND VGND VPWR VPWR mux_right_ipin_8.mux_l2_in_3_/S
+ sky130_fd_sc_hd__dfxtp_1
Xclkbuf_2_1_0_mem_right_ipin_0.prog_clk clkbuf_2_1_0_mem_right_ipin_0.prog_clk/A VGND
+ VGND VPWR VPWR clkbuf_3_3_0_mem_right_ipin_0.prog_clk/A sky130_fd_sc_hd__clkbuf_1
XFILLER_20_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_36_ chany_top_in[17] VGND VGND VPWR VPWR chany_bottom_out[17] sky130_fd_sc_hd__buf_2
XFILLER_22_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmem_right_ipin_10.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_4_0_mem_right_ipin_0.prog_clk/X
+ mux_right_ipin_10.mux_l1_in_0_/S VGND VGND VPWR VPWR mux_right_ipin_10.mux_l2_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_11_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19_ VGND VGND VPWR VPWR _19_/HI _19_/LO sky130_fd_sc_hd__conb_1
Xmem_right_ipin_5.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_0_0_mem_right_ipin_0.prog_clk/X
+ mux_right_ipin_4.mux_l4_in_0_/S VGND VGND VPWR VPWR mux_right_ipin_5.mux_l1_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
Xmux_right_ipin_14.mux_l1_in_0_ chany_top_in[0] chany_bottom_in[0] mux_right_ipin_14.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_right_ipin_14.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_10_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_right_ipin_1.mux_l2_in_3_ _21_/HI chany_top_in[13] mux_right_ipin_1.mux_l2_in_1_/S
+ VGND VGND VPWR VPWR mux_right_ipin_1.mux_l2_in_3_/X sky130_fd_sc_hd__mux2_1
XFILLER_27_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmem_right_ipin_13.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_7_0_mem_right_ipin_0.prog_clk/X
+ mux_right_ipin_13.mux_l1_in_0_/S VGND VGND VPWR VPWR mux_right_ipin_13.mux_l2_in_2_/S
+ sky130_fd_sc_hd__dfxtp_1
XPHY_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_96 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_63 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_52_ chany_top_in[1] VGND VGND VPWR VPWR chany_bottom_out[1] sky130_fd_sc_hd__buf_2
XPHY_74 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_85 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmem_right_ipin_8.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_3_0_mem_right_ipin_0.prog_clk/X
+ mux_right_ipin_7.mux_l4_in_0_/S VGND VGND VPWR VPWR mux_right_ipin_8.mux_l1_in_2_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_23_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_35_ chany_top_in[18] VGND VGND VPWR VPWR chany_bottom_out[18] sky130_fd_sc_hd__buf_2
Xmux_right_ipin_1.mux_l4_in_0_ mux_right_ipin_1.mux_l3_in_1_/X mux_right_ipin_1.mux_l3_in_0_/X
+ mux_right_ipin_1.mux_l4_in_0_/S VGND VGND VPWR VPWR mux_right_ipin_1.mux_l4_in_0_/X
+ sky130_fd_sc_hd__mux2_1
Xmem_right_ipin_10.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_4_0_mem_right_ipin_0.prog_clk/X
+ mux_right_ipin_9.mux_l4_in_0_/S VGND VGND VPWR VPWR mux_right_ipin_10.mux_l1_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_8_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18_ VGND VGND VPWR VPWR _18_/HI _18_/LO sky130_fd_sc_hd__conb_1
Xmux_right_ipin_6.mux_l2_in_3_ _16_/HI chany_top_in[18] mux_right_ipin_6.mux_l2_in_1_/S
+ VGND VGND VPWR VPWR mux_right_ipin_6.mux_l2_in_3_/X sky130_fd_sc_hd__mux2_1
XFILLER_17_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_right_ipin_1.mux_l3_in_1_ mux_right_ipin_1.mux_l2_in_3_/X mux_right_ipin_1.mux_l2_in_2_/X
+ mux_right_ipin_1.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_right_ipin_1.mux_l3_in_1_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_right_ipin_1.mux_l2_in_2_ chany_bottom_in[13] chany_top_in[5] mux_right_ipin_1.mux_l2_in_1_/S
+ VGND VGND VPWR VPWR mux_right_ipin_1.mux_l2_in_2_/X sky130_fd_sc_hd__mux2_1
XFILLER_14_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_right_ipin_6.mux_l4_in_0_ mux_right_ipin_6.mux_l3_in_1_/X mux_right_ipin_6.mux_l3_in_0_/X
+ mux_right_ipin_6.mux_l4_in_0_/S VGND VGND VPWR VPWR mux_right_ipin_6.mux_l4_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XPHY_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmem_right_ipin_13.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_5_0_mem_right_ipin_0.prog_clk/X
+ mux_right_ipin_12.mux_l4_in_0_/S VGND VGND VPWR VPWR mux_right_ipin_13.mux_l1_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XPHY_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_97 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_64 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_75 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_86 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_51_ chany_top_in[2] VGND VGND VPWR VPWR chany_bottom_out[2] sky130_fd_sc_hd__buf_2
XFILLER_23_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xprog_clk_0_S_FTB01 prog_clk_0_W_in VGND VGND VPWR VPWR prog_clk_0_S_out sky130_fd_sc_hd__buf_4
Xmux_right_ipin_6.mux_l3_in_1_ mux_right_ipin_6.mux_l2_in_3_/X mux_right_ipin_6.mux_l2_in_2_/X
+ mux_right_ipin_6.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_right_ipin_6.mux_l3_in_1_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_11_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_34_ chany_top_in[19] VGND VGND VPWR VPWR chany_bottom_out[19] sky130_fd_sc_hd__buf_2
XFILLER_22_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_right_ipin_6.mux_l2_in_2_ chany_bottom_in[18] chany_top_in[10] mux_right_ipin_6.mux_l2_in_1_/S
+ VGND VGND VPWR VPWR mux_right_ipin_6.mux_l2_in_2_/X sky130_fd_sc_hd__mux2_1
X_17_ VGND VGND VPWR VPWR _17_/HI _17_/LO sky130_fd_sc_hd__conb_1
Xmux_right_ipin_1.mux_l3_in_0_ mux_right_ipin_1.mux_l2_in_1_/X mux_right_ipin_1.mux_l2_in_0_/X
+ mux_right_ipin_1.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_right_ipin_1.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_3_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_right_ipin_1.mux_l2_in_1_ chany_bottom_in[5] chany_top_in[3] mux_right_ipin_1.mux_l2_in_1_/S
+ VGND VGND VPWR VPWR mux_right_ipin_1.mux_l2_in_1_/X sky130_fd_sc_hd__mux2_1
XPHY_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_98 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_65 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_76 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_87 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_50_ chany_top_in[3] VGND VGND VPWR VPWR chany_bottom_out[3] sky130_fd_sc_hd__buf_2
Xmux_right_ipin_10.mux_l2_in_3_ _22_/HI chany_top_in[14] mux_right_ipin_10.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR mux_right_ipin_10.mux_l2_in_3_/X sky130_fd_sc_hd__mux2_1
Xmux_right_ipin_6.mux_l3_in_0_ mux_right_ipin_6.mux_l2_in_1_/X mux_right_ipin_6.mux_l2_in_0_/X
+ mux_right_ipin_6.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_right_ipin_6.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_11_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_33_ Test_en_E_in VGND VGND VPWR VPWR Test_en_W_in sky130_fd_sc_hd__buf_2
XFILLER_11_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_right_ipin_6.mux_l2_in_1_ chany_bottom_in[10] chany_top_in[2] mux_right_ipin_6.mux_l2_in_1_/S
+ VGND VGND VPWR VPWR mux_right_ipin_6.mux_l2_in_1_/X sky130_fd_sc_hd__mux2_1
X_16_ VGND VGND VPWR VPWR _16_/HI _16_/LO sky130_fd_sc_hd__conb_1
XFILLER_6_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_right_ipin_10.mux_l4_in_0_ mux_right_ipin_10.mux_l3_in_1_/X mux_right_ipin_10.mux_l3_in_0_/X
+ mux_right_ipin_10.mux_l4_in_0_/S VGND VGND VPWR VPWR mux_right_ipin_10.mux_l4_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_right_ipin_15.mux_l2_in_3_ _27_/HI chany_top_in[19] mux_right_ipin_15.mux_l2_in_2_/S
+ VGND VGND VPWR VPWR mux_right_ipin_15.mux_l2_in_3_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_right_ipin_10.mux_l3_in_1_ mux_right_ipin_10.mux_l2_in_3_/X mux_right_ipin_10.mux_l2_in_2_/X
+ mux_right_ipin_10.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_right_ipin_10.mux_l3_in_1_/X
+ sky130_fd_sc_hd__mux2_1
Xmux_right_ipin_9.sky130_fd_sc_hd__buf_4_0_ mux_right_ipin_9.mux_l4_in_0_/X VGND VGND
+ VPWR VPWR left_grid_pin_25_ sky130_fd_sc_hd__buf_4
Xmux_right_ipin_1.mux_l2_in_0_ chany_bottom_in[3] mux_right_ipin_1.mux_l1_in_0_/X
+ mux_right_ipin_1.mux_l2_in_1_/S VGND VGND VPWR VPWR mux_right_ipin_1.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_26_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_99 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_66 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_77 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_88 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_right_ipin_10.mux_l2_in_2_ chany_bottom_in[14] chany_top_in[6] mux_right_ipin_10.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR mux_right_ipin_10.mux_l2_in_2_/X sky130_fd_sc_hd__mux2_1
XFILLER_11_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_right_ipin_15.mux_l4_in_0_ mux_right_ipin_15.mux_l3_in_1_/X mux_right_ipin_15.mux_l3_in_0_/X
+ ccff_tail VGND VGND VPWR VPWR mux_right_ipin_15.mux_l4_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_14_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_32_ Test_en_E_in VGND VGND VPWR VPWR Test_en_S_in sky130_fd_sc_hd__buf_2
Xclk_2_N_FTB01 clk_2_N_in VGND VGND VPWR VPWR clk_2_N_out sky130_fd_sc_hd__buf_4
XFILLER_22_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_right_ipin_15.mux_l3_in_1_ mux_right_ipin_15.mux_l2_in_3_/X mux_right_ipin_15.mux_l2_in_2_/X
+ mux_right_ipin_15.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_right_ipin_15.mux_l3_in_1_/X
+ sky130_fd_sc_hd__mux2_1
Xmux_right_ipin_6.mux_l2_in_0_ chany_bottom_in[2] mux_right_ipin_6.mux_l1_in_0_/X
+ mux_right_ipin_6.mux_l2_in_1_/S VGND VGND VPWR VPWR mux_right_ipin_6.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_3_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_right_ipin_15.mux_l2_in_2_ chany_bottom_in[19] chany_top_in[15] mux_right_ipin_15.mux_l2_in_2_/S
+ VGND VGND VPWR VPWR mux_right_ipin_15.mux_l2_in_2_/X sky130_fd_sc_hd__mux2_1
Xclkbuf_1_1_0_mem_right_ipin_0.prog_clk clkbuf_0_mem_right_ipin_0.prog_clk/X VGND
+ VGND VPWR VPWR clkbuf_2_2_0_mem_right_ipin_0.prog_clk/A sky130_fd_sc_hd__clkbuf_1
Xmux_right_ipin_10.mux_l3_in_0_ mux_right_ipin_10.mux_l2_in_1_/X mux_right_ipin_10.mux_l2_in_0_/X
+ mux_right_ipin_10.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_right_ipin_10.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XPHY_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_56 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_67 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_78 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_89 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmux_right_ipin_10.mux_l2_in_1_ chany_bottom_in[6] chany_top_in[2] mux_right_ipin_10.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR mux_right_ipin_10.mux_l2_in_1_/X sky130_fd_sc_hd__mux2_1
Xmux_right_ipin_1.mux_l1_in_0_ chany_top_in[1] chany_bottom_in[1] mux_right_ipin_1.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_right_ipin_1.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
X_31_ VGND VGND VPWR VPWR _31_/HI _31_/LO sky130_fd_sc_hd__conb_1
XFILLER_11_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_right_ipin_15.mux_l3_in_0_ mux_right_ipin_15.mux_l2_in_1_/X mux_right_ipin_15.mux_l2_in_0_/X
+ mux_right_ipin_15.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_right_ipin_15.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_17_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_right_ipin_6.mux_l1_in_0_ chany_top_in[0] chany_bottom_in[0] mux_right_ipin_6.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_right_ipin_6.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
Xmux_right_ipin_15.mux_l2_in_1_ chany_bottom_in[15] mux_right_ipin_15.mux_l1_in_2_/X
+ mux_right_ipin_15.mux_l2_in_2_/S VGND VGND VPWR VPWR mux_right_ipin_15.mux_l2_in_1_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_14_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_right_ipin_15.mux_l1_in_2_ chany_top_in[9] chany_bottom_in[9] mux_right_ipin_15.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_right_ipin_15.mux_l1_in_2_/X sky130_fd_sc_hd__mux2_1
XPHY_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_57 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_68 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_79 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_right_ipin_10.sky130_fd_sc_hd__buf_4_0_ mux_right_ipin_10.mux_l4_in_0_/X VGND
+ VGND VPWR VPWR left_grid_pin_26_ sky130_fd_sc_hd__buf_4
Xmux_right_ipin_10.mux_l2_in_0_ chany_bottom_in[2] mux_right_ipin_10.mux_l1_in_0_/X
+ mux_right_ipin_10.mux_l2_in_0_/S VGND VGND VPWR VPWR mux_right_ipin_10.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_17_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_30_ VGND VGND VPWR VPWR _30_/HI _30_/LO sky130_fd_sc_hd__conb_1
Xmux_right_ipin_2.sky130_fd_sc_hd__buf_4_0_ mux_right_ipin_2.mux_l4_in_0_/X VGND VGND
+ VPWR VPWR left_grid_pin_18_ sky130_fd_sc_hd__buf_4
XFILLER_22_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_right_ipin_15.mux_l2_in_0_ mux_right_ipin_15.mux_l1_in_1_/X mux_right_ipin_15.mux_l1_in_0_/X
+ mux_right_ipin_15.mux_l2_in_2_/S VGND VGND VPWR VPWR mux_right_ipin_15.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_5_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_right_ipin_15.mux_l1_in_1_ chany_top_in[3] chany_bottom_in[3] mux_right_ipin_15.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_right_ipin_15.mux_l1_in_1_/X sky130_fd_sc_hd__mux2_1
XPHY_58 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_69 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_3_0_0_mem_right_ipin_0.prog_clk clkbuf_3_1_0_mem_right_ipin_0.prog_clk/A VGND
+ VGND VPWR VPWR clkbuf_3_0_0_mem_right_ipin_0.prog_clk/X sky130_fd_sc_hd__clkbuf_1
XFILLER_9_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_right_ipin_10.mux_l1_in_0_ chany_top_in[0] chany_bottom_in[0] mux_right_ipin_10.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_right_ipin_10.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_10_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_3_3_0_mem_right_ipin_0.prog_clk clkbuf_3_3_0_mem_right_ipin_0.prog_clk/A VGND
+ VGND VPWR VPWR clkbuf_3_3_0_mem_right_ipin_0.prog_clk/X sky130_fd_sc_hd__clkbuf_1
XPHY_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_right_ipin_15.mux_l1_in_0_ chany_top_in[1] chany_bottom_in[1] mux_right_ipin_15.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_right_ipin_15.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XPHY_59 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_right_ipin_2.mux_l2_in_3_ _28_/HI chany_top_in[14] mux_right_ipin_2.mux_l2_in_2_/S
+ VGND VGND VPWR VPWR mux_right_ipin_2.mux_l2_in_3_/X sky130_fd_sc_hd__mux2_1
XFILLER_14_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmem_right_ipin_1.sky130_fd_sc_hd__dfxtp_1_3_ clkbuf_3_0_0_mem_right_ipin_0.prog_clk/X
+ mux_right_ipin_1.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_right_ipin_1.mux_l4_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
Xprog_clk_0_N_FTB01 prog_clk_0_W_in VGND VGND VPWR VPWR prog_clk_0_N_out sky130_fd_sc_hd__buf_4
Xmux_right_ipin_2.mux_l4_in_0_ mux_right_ipin_2.mux_l3_in_1_/X mux_right_ipin_2.mux_l3_in_0_/X
+ mux_right_ipin_2.mux_l4_in_0_/S VGND VGND VPWR VPWR mux_right_ipin_2.mux_l4_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_3_6_0_mem_right_ipin_0.prog_clk clkbuf_3_7_0_mem_right_ipin_0.prog_clk/A VGND
+ VGND VPWR VPWR clkbuf_3_6_0_mem_right_ipin_0.prog_clk/X sky130_fd_sc_hd__clkbuf_1
Xmux_right_ipin_7.mux_l2_in_3_ _17_/HI chany_top_in[17] mux_right_ipin_7.mux_l2_in_1_/S
+ VGND VGND VPWR VPWR mux_right_ipin_7.mux_l2_in_3_/X sky130_fd_sc_hd__mux2_1
Xmux_right_ipin_2.mux_l3_in_1_ mux_right_ipin_2.mux_l2_in_3_/X mux_right_ipin_2.mux_l2_in_2_/X
+ mux_right_ipin_2.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_right_ipin_2.mux_l3_in_1_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_20_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_0 _28_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_right_ipin_2.mux_l2_in_2_ chany_bottom_in[14] chany_top_in[6] mux_right_ipin_2.mux_l2_in_2_/S
+ VGND VGND VPWR VPWR mux_right_ipin_2.mux_l2_in_2_/X sky130_fd_sc_hd__mux2_1
Xmem_right_ipin_4.sky130_fd_sc_hd__dfxtp_1_3_ clkbuf_3_1_0_mem_right_ipin_0.prog_clk/X
+ mux_right_ipin_4.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_right_ipin_4.mux_l4_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_7_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_right_ipin_7.mux_l4_in_0_ mux_right_ipin_7.mux_l3_in_1_/X mux_right_ipin_7.mux_l3_in_0_/X
+ mux_right_ipin_7.mux_l4_in_0_/S VGND VGND VPWR VPWR mux_right_ipin_7.mux_l4_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_9_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_right_ipin_7.mux_l3_in_1_ mux_right_ipin_7.mux_l2_in_3_/X mux_right_ipin_7.mux_l2_in_2_/X
+ mux_right_ipin_7.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_right_ipin_7.mux_l3_in_1_/X
+ sky130_fd_sc_hd__mux2_1
Xmem_right_ipin_1.sky130_fd_sc_hd__dfxtp_1_2_ clkbuf_3_2_0_mem_right_ipin_0.prog_clk/X
+ mux_right_ipin_1.mux_l2_in_1_/S VGND VGND VPWR VPWR mux_right_ipin_1.mux_l3_in_1_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_3_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_right_ipin_7.mux_l2_in_2_ chany_bottom_in[17] chany_top_in[11] mux_right_ipin_7.mux_l2_in_1_/S
+ VGND VGND VPWR VPWR mux_right_ipin_7.mux_l2_in_2_/X sky130_fd_sc_hd__mux2_1
XFILLER_22_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_right_ipin_2.mux_l3_in_0_ mux_right_ipin_2.mux_l2_in_1_/X mux_right_ipin_2.mux_l2_in_0_/X
+ mux_right_ipin_2.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_right_ipin_2.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
Xmem_right_ipin_7.sky130_fd_sc_hd__dfxtp_1_3_ clkbuf_3_1_0_mem_right_ipin_0.prog_clk/X
+ mux_right_ipin_7.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_right_ipin_7.mux_l4_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_26_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_1 _28_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_right_ipin_2.mux_l2_in_1_ chany_bottom_in[6] chany_top_in[2] mux_right_ipin_2.mux_l2_in_2_/S
+ VGND VGND VPWR VPWR mux_right_ipin_2.mux_l2_in_1_/X sky130_fd_sc_hd__mux2_1
Xmux_right_ipin_13.sky130_fd_sc_hd__buf_4_0_ mux_right_ipin_13.mux_l4_in_0_/X VGND
+ VGND VPWR VPWR left_grid_pin_29_ sky130_fd_sc_hd__buf_4
Xmem_right_ipin_4.sky130_fd_sc_hd__dfxtp_1_2_ clkbuf_3_0_0_mem_right_ipin_0.prog_clk/X
+ mux_right_ipin_4.mux_l2_in_3_/S VGND VGND VPWR VPWR mux_right_ipin_4.mux_l3_in_1_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_9_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_right_ipin_5.sky130_fd_sc_hd__buf_4_0_ mux_right_ipin_5.mux_l4_in_0_/X VGND VGND
+ VPWR VPWR left_grid_pin_21_ sky130_fd_sc_hd__buf_4
XFILLER_6_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_right_ipin_11.mux_l2_in_3_ _23_/HI chany_top_in[15] mux_right_ipin_11.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR mux_right_ipin_11.mux_l2_in_3_/X sky130_fd_sc_hd__mux2_1
X_69_ chany_bottom_in[4] VGND VGND VPWR VPWR chany_top_out[4] sky130_fd_sc_hd__buf_2
Xprog_clk_3_S_FTB01 prog_clk_3_N_in VGND VGND VPWR VPWR prog_clk_3_S_out sky130_fd_sc_hd__buf_4
Xmem_right_ipin_1.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_3_0_mem_right_ipin_0.prog_clk/X
+ mux_right_ipin_1.mux_l1_in_0_/S VGND VGND VPWR VPWR mux_right_ipin_1.mux_l2_in_1_/S
+ sky130_fd_sc_hd__dfxtp_1
Xmux_right_ipin_7.mux_l3_in_0_ mux_right_ipin_7.mux_l2_in_1_/X mux_right_ipin_7.mux_l2_in_0_/X
+ mux_right_ipin_7.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_right_ipin_7.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
Xmem_right_ipin_12.sky130_fd_sc_hd__dfxtp_1_3_ clkbuf_3_5_0_mem_right_ipin_0.prog_clk/X
+ mux_right_ipin_12.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_right_ipin_12.mux_l4_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_15_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_right_ipin_7.mux_l2_in_1_ chany_bottom_in[11] mux_right_ipin_7.mux_l1_in_2_/X
+ mux_right_ipin_7.mux_l2_in_1_/S VGND VGND VPWR VPWR mux_right_ipin_7.mux_l2_in_1_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_20_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_right_ipin_11.mux_l4_in_0_ mux_right_ipin_11.mux_l3_in_1_/X mux_right_ipin_11.mux_l3_in_0_/X
+ mux_right_ipin_11.mux_l4_in_0_/S VGND VGND VPWR VPWR mux_right_ipin_11.mux_l4_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_2 _30_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_right_ipin_7.sky130_fd_sc_hd__dfxtp_1_2_ clkbuf_3_3_0_mem_right_ipin_0.prog_clk/X
+ mux_right_ipin_7.mux_l2_in_1_/S VGND VGND VPWR VPWR mux_right_ipin_7.mux_l3_in_1_/S
+ sky130_fd_sc_hd__dfxtp_1
XPHY_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_right_ipin_7.mux_l1_in_2_ chany_top_in[7] chany_bottom_in[7] mux_right_ipin_7.mux_l1_in_1_/S
+ VGND VGND VPWR VPWR mux_right_ipin_7.mux_l1_in_2_/X sky130_fd_sc_hd__mux2_1
Xmux_right_ipin_11.mux_l3_in_1_ mux_right_ipin_11.mux_l2_in_3_/X mux_right_ipin_11.mux_l2_in_2_/X
+ mux_right_ipin_11.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_right_ipin_11.mux_l3_in_1_/X
+ sky130_fd_sc_hd__mux2_1
Xmux_right_ipin_2.mux_l2_in_0_ chany_bottom_in[2] mux_right_ipin_2.mux_l1_in_0_/X
+ mux_right_ipin_2.mux_l2_in_2_/S VGND VGND VPWR VPWR mux_right_ipin_2.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_13_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmem_right_ipin_4.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_2_0_mem_right_ipin_0.prog_clk/X
+ mux_right_ipin_4.mux_l1_in_0_/S VGND VGND VPWR VPWR mux_right_ipin_4.mux_l2_in_3_/S
+ sky130_fd_sc_hd__dfxtp_1
XTest_en_N_FTB01 Test_en_E_in VGND VGND VPWR VPWR Test_en_N_out sky130_fd_sc_hd__buf_4
Xmux_right_ipin_11.mux_l2_in_2_ chany_bottom_in[15] chany_top_in[11] mux_right_ipin_11.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR mux_right_ipin_11.mux_l2_in_2_/X sky130_fd_sc_hd__mux2_1
X_68_ chany_bottom_in[5] VGND VGND VPWR VPWR chany_top_out[5] sky130_fd_sc_hd__buf_2
Xmem_right_ipin_15.sky130_fd_sc_hd__dfxtp_1_3_ clkbuf_3_6_0_mem_right_ipin_0.prog_clk/X
+ mux_right_ipin_15.mux_l3_in_0_/S VGND VGND VPWR VPWR ccff_tail sky130_fd_sc_hd__dfxtp_1
Xmem_right_ipin_1.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_0_0_mem_right_ipin_0.prog_clk/X
+ mux_right_ipin_0.mux_l4_in_0_/S VGND VGND VPWR VPWR mux_right_ipin_1.mux_l1_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_2_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmem_right_ipin_12.sky130_fd_sc_hd__dfxtp_1_2_ clkbuf_3_6_0_mem_right_ipin_0.prog_clk/X
+ mux_right_ipin_12.mux_l2_in_2_/S VGND VGND VPWR VPWR mux_right_ipin_12.mux_l3_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
Xmux_right_ipin_7.mux_l2_in_0_ mux_right_ipin_7.mux_l1_in_1_/X mux_right_ipin_7.mux_l1_in_0_/X
+ mux_right_ipin_7.mux_l2_in_1_/S VGND VGND VPWR VPWR mux_right_ipin_7.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
Xclkbuf_0_mem_right_ipin_0.prog_clk prog_clk_0_FTB00/X VGND VGND VPWR VPWR clkbuf_0_mem_right_ipin_0.prog_clk/X
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA_3 _30_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_right_ipin_7.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_1_0_mem_right_ipin_0.prog_clk/X
+ mux_right_ipin_7.mux_l1_in_1_/S VGND VGND VPWR VPWR mux_right_ipin_7.mux_l2_in_1_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_6_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_2_0_0_mem_right_ipin_0.prog_clk clkbuf_2_1_0_mem_right_ipin_0.prog_clk/A VGND
+ VGND VPWR VPWR clkbuf_3_1_0_mem_right_ipin_0.prog_clk/A sky130_fd_sc_hd__clkbuf_1
XPHY_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_right_ipin_7.mux_l1_in_1_ chany_top_in[3] chany_bottom_in[3] mux_right_ipin_7.mux_l1_in_1_/S
+ VGND VGND VPWR VPWR mux_right_ipin_7.mux_l1_in_1_/X sky130_fd_sc_hd__mux2_1
Xmux_right_ipin_11.mux_l3_in_0_ mux_right_ipin_11.mux_l2_in_1_/X mux_right_ipin_11.mux_l2_in_0_/X
+ mux_right_ipin_11.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_right_ipin_11.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_26_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmem_right_ipin_4.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_2_0_mem_right_ipin_0.prog_clk/X
+ mux_right_ipin_3.mux_l4_in_0_/S VGND VGND VPWR VPWR mux_right_ipin_4.mux_l1_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_13_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_right_ipin_11.mux_l2_in_1_ chany_bottom_in[11] mux_right_ipin_11.mux_l1_in_2_/X
+ mux_right_ipin_11.mux_l2_in_0_/S VGND VGND VPWR VPWR mux_right_ipin_11.mux_l2_in_1_/X
+ sky130_fd_sc_hd__mux2_1
Xmux_right_ipin_2.mux_l1_in_0_ chany_top_in[0] chany_bottom_in[0] mux_right_ipin_2.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_right_ipin_2.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_5_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_67_ chany_bottom_in[6] VGND VGND VPWR VPWR chany_top_out[6] sky130_fd_sc_hd__buf_2
Xmem_right_ipin_15.sky130_fd_sc_hd__dfxtp_1_2_ clkbuf_3_6_0_mem_right_ipin_0.prog_clk/X
+ mux_right_ipin_15.mux_l2_in_2_/S VGND VGND VPWR VPWR mux_right_ipin_15.mux_l3_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_24_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_2_3_0_mem_right_ipin_0.prog_clk clkbuf_2_2_0_mem_right_ipin_0.prog_clk/A VGND
+ VGND VPWR VPWR clkbuf_3_7_0_mem_right_ipin_0.prog_clk/A sky130_fd_sc_hd__clkbuf_1
XFILLER_9_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_right_ipin_11.mux_l1_in_2_ chany_top_in[5] chany_bottom_in[5] mux_right_ipin_11.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_right_ipin_11.mux_l1_in_2_/X sky130_fd_sc_hd__mux2_1
Xmem_right_ipin_12.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_7_0_mem_right_ipin_0.prog_clk/X
+ mux_right_ipin_12.mux_l1_in_2_/S VGND VGND VPWR VPWR mux_right_ipin_12.mux_l2_in_2_/S
+ sky130_fd_sc_hd__dfxtp_1
Xmem_right_ipin_7.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_1_0_mem_right_ipin_0.prog_clk/X
+ mux_right_ipin_6.mux_l4_in_0_/S VGND VGND VPWR VPWR mux_right_ipin_7.mux_l1_in_1_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_20_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_right_ipin_7.mux_l1_in_0_ chany_top_in[1] chany_bottom_in[1] mux_right_ipin_7.mux_l1_in_1_/S
+ VGND VGND VPWR VPWR mux_right_ipin_7.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_16_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
.ends

