magic
tech sky130A
magscale 1 2
timestamp 1608228718
<< checkpaint >>
rect -1260 -1260 25660 25660
<< locali >>
rect 11713 21879 11747 21981
rect 12357 21947 12391 22117
rect 19257 21947 19291 22117
rect 5917 21471 5951 21641
rect 17325 21403 17359 21641
rect 20913 21403 20947 21641
rect 14565 20859 14599 21029
rect 4997 20383 5031 20553
rect 3157 19703 3191 19873
rect 5273 19839 5307 19941
rect 19073 19839 19107 19941
rect 9689 17663 9723 17833
rect 2237 16983 2271 17085
rect 9597 16983 9631 17153
rect 17325 16983 17359 17153
rect 8585 16643 8619 16745
rect 9137 16439 9171 16609
rect 12173 16575 12207 16745
rect 17785 16031 17819 16201
rect 8585 15895 8619 15997
rect 8861 15351 8895 15589
rect 14749 15487 14783 15657
rect 8861 15317 8953 15351
rect 20729 14807 20763 14977
rect 13369 14263 13403 14433
rect 19349 14263 19383 14365
rect 21741 13855 21775 13957
rect 17785 12631 17819 12733
rect 9505 12155 9539 12257
rect 11345 12087 11379 12257
rect 3985 11747 4019 11849
rect 16865 11543 16899 11645
rect 6653 10455 6687 10625
rect 8401 10455 8435 10693
rect 9413 9979 9447 10217
rect 9505 10115 9539 10217
rect 16037 9367 16071 9673
rect 19993 9367 20027 9605
rect 10609 8279 10643 8517
rect 18797 8415 18831 8517
rect 19717 8483 19751 8585
rect 7849 7939 7883 8041
rect 9505 7871 9539 8041
rect 7389 7191 7423 7361
rect 16221 7191 16255 7293
rect 14197 6647 14231 6817
rect 23397 5899 23431 6817
rect 9413 5695 9447 5865
rect 12909 5763 12943 5865
rect 12909 5559 12943 5729
rect 14657 3927 14691 4097
<< viali >>
rect 12357 22117 12391 22151
rect 11713 21981 11747 22015
rect 12357 21913 12391 21947
rect 19257 22117 19291 22151
rect 19257 21913 19291 21947
rect 11713 21845 11747 21879
rect 5917 21641 5951 21675
rect 9137 21641 9171 21675
rect 10057 21641 10091 21675
rect 17325 21641 17359 21675
rect 17693 21641 17727 21675
rect 20913 21641 20947 21675
rect 2421 21505 2455 21539
rect 3341 21505 3375 21539
rect 4721 21505 4755 21539
rect 5549 21505 5583 21539
rect 5733 21505 5767 21539
rect 6929 21573 6963 21607
rect 15025 21573 15059 21607
rect 7481 21505 7515 21539
rect 8585 21505 8619 21539
rect 10517 21505 10551 21539
rect 10701 21505 10735 21539
rect 11621 21505 11655 21539
rect 13185 21505 13219 21539
rect 14197 21505 14231 21539
rect 16129 21505 16163 21539
rect 17141 21505 17175 21539
rect 5457 21437 5491 21471
rect 5917 21437 5951 21471
rect 6101 21437 6135 21471
rect 8401 21437 8435 21471
rect 8953 21437 8987 21471
rect 14841 21437 14875 21471
rect 15945 21437 15979 21471
rect 16957 21437 16991 21471
rect 20177 21505 20211 21539
rect 17509 21437 17543 21471
rect 18337 21437 18371 21471
rect 22201 21573 22235 21607
rect 21833 21505 21867 21539
rect 22845 21505 22879 21539
rect 22661 21437 22695 21471
rect 2145 21369 2179 21403
rect 4445 21369 4479 21403
rect 8309 21369 8343 21403
rect 10425 21369 10459 21403
rect 14105 21369 14139 21403
rect 15853 21369 15887 21403
rect 17325 21369 17359 21403
rect 19165 21369 19199 21403
rect 19993 21369 20027 21403
rect 20913 21369 20947 21403
rect 21557 21369 21591 21403
rect 1777 21301 1811 21335
rect 2237 21301 2271 21335
rect 2789 21301 2823 21335
rect 3157 21301 3191 21335
rect 3249 21301 3283 21335
rect 4077 21301 4111 21335
rect 4537 21301 4571 21335
rect 5089 21301 5123 21335
rect 6285 21301 6319 21335
rect 7297 21301 7331 21335
rect 7389 21301 7423 21335
rect 7941 21301 7975 21335
rect 11069 21301 11103 21335
rect 11437 21301 11471 21335
rect 11529 21301 11563 21335
rect 12081 21301 12115 21335
rect 12633 21301 12667 21335
rect 13001 21301 13035 21335
rect 13093 21301 13127 21335
rect 13645 21301 13679 21335
rect 14013 21301 14047 21335
rect 15485 21301 15519 21335
rect 16497 21301 16531 21335
rect 16865 21301 16899 21335
rect 19625 21301 19659 21335
rect 20085 21301 20119 21335
rect 20637 21301 20671 21335
rect 21189 21301 21223 21335
rect 21649 21301 21683 21335
rect 22569 21301 22603 21335
rect 1777 21097 1811 21131
rect 3525 21097 3559 21131
rect 5457 21097 5491 21131
rect 6101 21097 6135 21131
rect 8125 21097 8159 21131
rect 8953 21097 8987 21131
rect 14473 21097 14507 21131
rect 17325 21097 17359 21131
rect 19809 21097 19843 21131
rect 21281 21097 21315 21131
rect 11590 21029 11624 21063
rect 14565 21029 14599 21063
rect 14749 21029 14783 21063
rect 15568 21029 15602 21063
rect 20177 21029 20211 21063
rect 22293 21029 22327 21063
rect 1593 20961 1627 20995
rect 2412 20961 2446 20995
rect 4344 20961 4378 20995
rect 6193 20961 6227 20995
rect 7012 20961 7046 20995
rect 9956 20961 9990 20995
rect 13360 20961 13394 20995
rect 2145 20893 2179 20927
rect 4077 20893 4111 20927
rect 6285 20893 6319 20927
rect 6745 20893 6779 20927
rect 9045 20893 9079 20927
rect 9229 20893 9263 20927
rect 9689 20893 9723 20927
rect 11345 20893 11379 20927
rect 13093 20893 13127 20927
rect 18420 20961 18454 20995
rect 22201 20961 22235 20995
rect 22661 20961 22695 20995
rect 15301 20893 15335 20927
rect 17417 20893 17451 20927
rect 17601 20893 17635 20927
rect 18153 20893 18187 20927
rect 20269 20893 20303 20927
rect 20361 20893 20395 20927
rect 21373 20893 21407 20927
rect 21465 20893 21499 20927
rect 22385 20893 22419 20927
rect 14565 20825 14599 20859
rect 16957 20825 16991 20859
rect 5733 20757 5767 20791
rect 8585 20757 8619 20791
rect 11069 20757 11103 20791
rect 12725 20757 12759 20791
rect 16681 20757 16715 20791
rect 19533 20757 19567 20791
rect 20913 20757 20947 20791
rect 21833 20757 21867 20791
rect 22845 20757 22879 20791
rect 3157 20553 3191 20587
rect 4813 20553 4847 20587
rect 4997 20553 5031 20587
rect 8217 20553 8251 20587
rect 10241 20553 10275 20587
rect 11897 20553 11931 20587
rect 14105 20553 14139 20587
rect 19441 20553 19475 20587
rect 21189 20553 21223 20587
rect 22017 20553 22051 20587
rect 5733 20417 5767 20451
rect 10517 20417 10551 20451
rect 12725 20417 12759 20451
rect 14381 20417 14415 20451
rect 21741 20417 21775 20451
rect 22661 20417 22695 20451
rect 1777 20349 1811 20383
rect 3433 20349 3467 20383
rect 3689 20349 3723 20383
rect 4997 20349 5031 20383
rect 6285 20349 6319 20383
rect 6837 20349 6871 20383
rect 8861 20349 8895 20383
rect 14637 20349 14671 20383
rect 16037 20349 16071 20383
rect 18061 20349 18095 20383
rect 18328 20349 18362 20383
rect 19717 20349 19751 20383
rect 19984 20349 20018 20383
rect 2044 20281 2078 20315
rect 5549 20281 5583 20315
rect 6101 20281 6135 20315
rect 7104 20281 7138 20315
rect 9128 20281 9162 20315
rect 10784 20281 10818 20315
rect 12992 20281 13026 20315
rect 16304 20281 16338 20315
rect 21649 20281 21683 20315
rect 22477 20281 22511 20315
rect 5089 20213 5123 20247
rect 5457 20213 5491 20247
rect 6469 20213 6503 20247
rect 15761 20213 15795 20247
rect 17417 20213 17451 20247
rect 21097 20213 21131 20247
rect 21557 20213 21591 20247
rect 22385 20213 22419 20247
rect 2973 20009 3007 20043
rect 3433 20009 3467 20043
rect 4077 20009 4111 20043
rect 9873 20009 9907 20043
rect 11075 20009 11109 20043
rect 14105 20009 14139 20043
rect 15669 20009 15703 20043
rect 17877 20009 17911 20043
rect 1860 19941 1894 19975
rect 4445 19941 4479 19975
rect 5273 19941 5307 19975
rect 5632 19941 5666 19975
rect 7472 19941 7506 19975
rect 14749 19941 14783 19975
rect 15761 19941 15795 19975
rect 16764 19941 16798 19975
rect 19073 19941 19107 19975
rect 19432 19941 19466 19975
rect 1593 19873 1627 19907
rect 3157 19873 3191 19907
rect 3249 19873 3283 19907
rect 4537 19873 4571 19907
rect 7205 19873 7239 19907
rect 8861 19873 8895 19907
rect 9689 19873 9723 19907
rect 10425 19873 10459 19907
rect 11345 19873 11379 19907
rect 12992 19873 13026 19907
rect 14565 19873 14599 19907
rect 18521 19873 18555 19907
rect 21456 19873 21490 19907
rect 22661 19873 22695 19907
rect 4629 19805 4663 19839
rect 5273 19805 5307 19839
rect 5365 19805 5399 19839
rect 10609 19805 10643 19839
rect 11115 19805 11149 19839
rect 12725 19805 12759 19839
rect 15945 19805 15979 19839
rect 16497 19805 16531 19839
rect 18613 19805 18647 19839
rect 18705 19805 18739 19839
rect 19073 19805 19107 19839
rect 19165 19805 19199 19839
rect 21189 19805 21223 19839
rect 9045 19737 9079 19771
rect 3157 19669 3191 19703
rect 6745 19669 6779 19703
rect 8585 19669 8619 19703
rect 10241 19669 10275 19703
rect 12449 19669 12483 19703
rect 14933 19669 14967 19703
rect 15301 19669 15335 19703
rect 18153 19669 18187 19703
rect 20545 19669 20579 19703
rect 22569 19669 22603 19703
rect 22845 19669 22879 19703
rect 2605 19465 2639 19499
rect 20085 19465 20119 19499
rect 2145 19329 2179 19363
rect 3157 19329 3191 19363
rect 4169 19329 4203 19363
rect 7896 19329 7930 19363
rect 8079 19329 8113 19363
rect 10241 19329 10275 19363
rect 13001 19329 13035 19363
rect 14013 19329 14047 19363
rect 15117 19329 15151 19363
rect 16129 19329 16163 19363
rect 17141 19329 17175 19363
rect 18524 19329 18558 19363
rect 18751 19329 18785 19363
rect 20637 19329 20671 19363
rect 4629 19261 4663 19295
rect 4896 19261 4930 19295
rect 6285 19261 6319 19295
rect 6837 19261 6871 19295
rect 7573 19261 7607 19295
rect 8309 19261 8343 19295
rect 10701 19261 10735 19295
rect 10968 19261 11002 19295
rect 13829 19261 13863 19295
rect 16957 19261 16991 19295
rect 17509 19261 17543 19295
rect 18069 19261 18103 19295
rect 20453 19261 20487 19295
rect 20913 19261 20947 19295
rect 2053 19193 2087 19227
rect 3985 19193 4019 19227
rect 10149 19193 10183 19227
rect 16865 19193 16899 19227
rect 21180 19193 21214 19227
rect 1593 19125 1627 19159
rect 1961 19125 1995 19159
rect 2973 19125 3007 19159
rect 3065 19125 3099 19159
rect 3617 19125 3651 19159
rect 4077 19125 4111 19159
rect 6009 19125 6043 19159
rect 7021 19125 7055 19159
rect 9413 19125 9447 19159
rect 9689 19125 9723 19159
rect 10057 19125 10091 19159
rect 12081 19125 12115 19159
rect 12449 19125 12483 19159
rect 12817 19125 12851 19159
rect 12909 19125 12943 19159
rect 13461 19125 13495 19159
rect 13921 19125 13955 19159
rect 14473 19125 14507 19159
rect 14841 19125 14875 19159
rect 14933 19125 14967 19159
rect 15485 19125 15519 19159
rect 15853 19125 15887 19159
rect 15945 19125 15979 19159
rect 16497 19125 16531 19159
rect 18527 19125 18561 19159
rect 19901 19125 19935 19159
rect 20545 19125 20579 19159
rect 22293 19125 22327 19159
rect 2973 18921 3007 18955
rect 3433 18921 3467 18955
rect 4077 18921 4111 18955
rect 5549 18921 5583 18955
rect 14013 18921 14047 18955
rect 7104 18853 7138 18887
rect 16028 18853 16062 18887
rect 1593 18785 1627 18819
rect 1860 18785 1894 18819
rect 3249 18785 3283 18819
rect 4445 18785 4479 18819
rect 5641 18785 5675 18819
rect 6193 18785 6227 18819
rect 6837 18785 6871 18819
rect 8861 18785 8895 18819
rect 9689 18785 9723 18819
rect 10425 18785 10459 18819
rect 11805 18785 11839 18819
rect 12900 18785 12934 18819
rect 14657 18785 14691 18819
rect 17601 18785 17635 18819
rect 17960 18785 17994 18819
rect 19533 18785 19567 18819
rect 21741 18785 21775 18819
rect 4537 18717 4571 18751
rect 4721 18717 4755 18751
rect 5825 18717 5859 18751
rect 8953 18717 8987 18751
rect 9137 18717 9171 18751
rect 10012 18717 10046 18751
rect 10152 18717 10186 18751
rect 12633 18717 12667 18751
rect 15301 18717 15335 18751
rect 15761 18717 15795 18751
rect 17693 18717 17727 18751
rect 19625 18717 19659 18751
rect 19717 18717 19751 18751
rect 20361 18717 20395 18751
rect 21833 18717 21867 18751
rect 21925 18717 21959 18751
rect 22569 18717 22603 18751
rect 5181 18649 5215 18683
rect 11529 18649 11563 18683
rect 14841 18649 14875 18683
rect 6377 18581 6411 18615
rect 8217 18581 8251 18615
rect 8493 18581 8527 18615
rect 11989 18581 12023 18615
rect 17141 18581 17175 18615
rect 17417 18581 17451 18615
rect 19073 18581 19107 18615
rect 19165 18581 19199 18615
rect 20177 18581 20211 18615
rect 21373 18581 21407 18615
rect 22385 18581 22419 18615
rect 3065 18377 3099 18411
rect 5273 18377 5307 18411
rect 9137 18377 9171 18411
rect 9413 18377 9447 18411
rect 14289 18377 14323 18411
rect 17509 18377 17543 18411
rect 11897 18309 11931 18343
rect 14565 18309 14599 18343
rect 5825 18241 5859 18275
rect 7297 18241 7331 18275
rect 7620 18241 7654 18275
rect 7803 18241 7837 18275
rect 9873 18241 9907 18275
rect 9965 18241 9999 18275
rect 15025 18241 15059 18275
rect 15209 18241 15243 18275
rect 15992 18241 16026 18275
rect 16175 18241 16209 18275
rect 18061 18241 18095 18275
rect 22477 18241 22511 18275
rect 1685 18173 1719 18207
rect 3341 18173 3375 18207
rect 3608 18173 3642 18207
rect 8033 18173 8067 18207
rect 9781 18173 9815 18207
rect 10517 18173 10551 18207
rect 12909 18173 12943 18207
rect 13176 18173 13210 18207
rect 15669 18173 15703 18207
rect 16405 18173 16439 18207
rect 18521 18173 18555 18207
rect 20177 18173 20211 18207
rect 1952 18105 1986 18139
rect 5733 18105 5767 18139
rect 6285 18105 6319 18139
rect 10784 18105 10818 18139
rect 14933 18105 14967 18139
rect 18788 18105 18822 18139
rect 20422 18105 20456 18139
rect 4721 18037 4755 18071
rect 5641 18037 5675 18071
rect 6837 18037 6871 18071
rect 12449 18037 12483 18071
rect 19901 18037 19935 18071
rect 21557 18037 21591 18071
rect 21925 18037 21959 18071
rect 22293 18037 22327 18071
rect 22385 18037 22419 18071
rect 3157 17833 3191 17867
rect 3617 17833 3651 17867
rect 4261 17833 4295 17867
rect 8125 17833 8159 17867
rect 8861 17833 8895 17867
rect 9689 17833 9723 17867
rect 11437 17833 11471 17867
rect 11805 17833 11839 17867
rect 14381 17833 14415 17867
rect 14841 17833 14875 17867
rect 16681 17833 16715 17867
rect 20269 17833 20303 17867
rect 22293 17833 22327 17867
rect 2044 17765 2078 17799
rect 8769 17765 8803 17799
rect 1777 17697 1811 17731
rect 3433 17697 3467 17731
rect 4077 17697 4111 17731
rect 5264 17697 5298 17731
rect 7012 17697 7046 17731
rect 13268 17765 13302 17799
rect 15546 17765 15580 17799
rect 18420 17765 18454 17799
rect 21158 17765 21192 17799
rect 10048 17697 10082 17731
rect 11897 17697 11931 17731
rect 12449 17697 12483 17731
rect 14657 17697 14691 17731
rect 17325 17697 17359 17731
rect 20177 17697 20211 17731
rect 4997 17629 5031 17663
rect 6745 17629 6779 17663
rect 9045 17629 9079 17663
rect 9689 17629 9723 17663
rect 9781 17629 9815 17663
rect 11989 17629 12023 17663
rect 13001 17629 13035 17663
rect 15301 17629 15335 17663
rect 17417 17629 17451 17663
rect 17601 17629 17635 17663
rect 18153 17629 18187 17663
rect 20453 17629 20487 17663
rect 20913 17629 20947 17663
rect 22569 17629 22603 17663
rect 12633 17561 12667 17595
rect 6377 17493 6411 17527
rect 8401 17493 8435 17527
rect 11161 17493 11195 17527
rect 16957 17493 16991 17527
rect 19533 17493 19567 17527
rect 19809 17493 19843 17527
rect 9413 17289 9447 17323
rect 11069 17289 11103 17323
rect 12449 17289 12483 17323
rect 3709 17221 3743 17255
rect 7021 17221 7055 17255
rect 15485 17221 15519 17255
rect 21097 17221 21131 17255
rect 4905 17153 4939 17187
rect 7665 17153 7699 17187
rect 9597 17153 9631 17187
rect 11805 17153 11839 17187
rect 11897 17153 11931 17187
rect 13001 17153 13035 17187
rect 16037 17153 16071 17187
rect 17049 17153 17083 17187
rect 17325 17153 17359 17187
rect 20177 17153 20211 17187
rect 20269 17153 20303 17187
rect 1777 17085 1811 17119
rect 2237 17085 2271 17119
rect 2329 17085 2363 17119
rect 2596 17085 2630 17119
rect 4261 17085 4295 17119
rect 4353 17085 4387 17119
rect 5172 17085 5206 17119
rect 8033 17085 8067 17119
rect 8289 17085 8323 17119
rect 9689 17085 9723 17119
rect 13737 17085 13771 17119
rect 13829 17085 13863 17119
rect 14096 17085 14130 17119
rect 16865 17085 16899 17119
rect 9956 17017 9990 17051
rect 11713 17017 11747 17051
rect 12817 17017 12851 17051
rect 15945 17017 15979 17051
rect 17509 17085 17543 17119
rect 18061 17085 18095 17119
rect 20085 17085 20119 17119
rect 20729 17085 20763 17119
rect 21373 17085 21407 17119
rect 18306 17017 18340 17051
rect 20913 17017 20947 17051
rect 21640 17017 21674 17051
rect 1961 16949 1995 16983
rect 2237 16949 2271 16983
rect 4077 16949 4111 16983
rect 4537 16949 4571 16983
rect 6285 16949 6319 16983
rect 7389 16949 7423 16983
rect 7481 16949 7515 16983
rect 9597 16949 9631 16983
rect 11345 16949 11379 16983
rect 12909 16949 12943 16983
rect 13553 16949 13587 16983
rect 15209 16949 15243 16983
rect 15853 16949 15887 16983
rect 16497 16949 16531 16983
rect 16957 16949 16991 16983
rect 17325 16949 17359 16983
rect 19441 16949 19475 16983
rect 19717 16949 19751 16983
rect 22753 16949 22787 16983
rect 1777 16745 1811 16779
rect 3525 16745 3559 16779
rect 4445 16745 4479 16779
rect 6193 16745 6227 16779
rect 8493 16745 8527 16779
rect 8585 16745 8619 16779
rect 9873 16745 9907 16779
rect 12173 16745 12207 16779
rect 14381 16745 14415 16779
rect 14473 16745 14507 16779
rect 20269 16745 20303 16779
rect 20913 16745 20947 16779
rect 21281 16745 21315 16779
rect 21925 16745 21959 16779
rect 2412 16677 2446 16711
rect 5080 16677 5114 16711
rect 6469 16677 6503 16711
rect 6837 16677 6871 16711
rect 1593 16609 1627 16643
rect 4261 16609 4295 16643
rect 6653 16609 6687 16643
rect 7380 16609 7414 16643
rect 8585 16609 8619 16643
rect 8769 16609 8803 16643
rect 9137 16609 9171 16643
rect 9505 16609 9539 16643
rect 9689 16609 9723 16643
rect 10564 16609 10598 16643
rect 2145 16541 2179 16575
rect 4813 16541 4847 16575
rect 7113 16541 7147 16575
rect 15568 16677 15602 16711
rect 20361 16677 20395 16711
rect 22385 16677 22419 16711
rect 12624 16609 12658 16643
rect 15301 16609 15335 16643
rect 17224 16609 17258 16643
rect 18429 16609 18463 16643
rect 18685 16609 18719 16643
rect 21373 16609 21407 16643
rect 22293 16609 22327 16643
rect 10241 16541 10275 16575
rect 10704 16541 10738 16575
rect 10977 16541 11011 16575
rect 12173 16541 12207 16575
rect 12357 16541 12391 16575
rect 14565 16541 14599 16575
rect 16957 16541 16991 16575
rect 20453 16541 20487 16575
rect 21465 16541 21499 16575
rect 22477 16541 22511 16575
rect 12081 16473 12115 16507
rect 14013 16473 14047 16507
rect 16681 16473 16715 16507
rect 19809 16473 19843 16507
rect 8953 16405 8987 16439
rect 9137 16405 9171 16439
rect 9321 16405 9355 16439
rect 13737 16405 13771 16439
rect 18337 16405 18371 16439
rect 19901 16405 19935 16439
rect 2881 16201 2915 16235
rect 6469 16201 6503 16235
rect 7389 16201 7423 16235
rect 10793 16201 10827 16235
rect 15209 16201 15243 16235
rect 17601 16201 17635 16235
rect 17785 16201 17819 16235
rect 20545 16201 20579 16235
rect 4445 16133 4479 16167
rect 12449 16133 12483 16167
rect 1501 16065 1535 16099
rect 3801 16065 3835 16099
rect 8033 16065 8067 16099
rect 9000 16065 9034 16099
rect 9183 16065 9217 16099
rect 11437 16065 11471 16099
rect 13001 16065 13035 16099
rect 13829 16065 13863 16099
rect 15485 16065 15519 16099
rect 19717 16133 19751 16167
rect 20269 16065 20303 16099
rect 21097 16065 21131 16099
rect 4261 15997 4295 16031
rect 4813 15997 4847 16031
rect 5080 15997 5114 16031
rect 6653 15997 6687 16031
rect 6837 15997 6871 16031
rect 8585 15997 8619 16031
rect 8677 15997 8711 16031
rect 9413 15997 9447 16031
rect 11161 15997 11195 16031
rect 11805 15997 11839 16031
rect 13737 15997 13771 16031
rect 17325 15997 17359 16031
rect 17417 15997 17451 16031
rect 17785 15997 17819 16031
rect 20085 15997 20119 16031
rect 21373 15997 21407 16031
rect 1768 15929 1802 15963
rect 7849 15929 7883 15963
rect 12909 15929 12943 15963
rect 14096 15929 14130 15963
rect 15730 15929 15764 15963
rect 19533 15929 19567 15963
rect 20177 15929 20211 15963
rect 20913 15929 20947 15963
rect 21640 15929 21674 15963
rect 3157 15861 3191 15895
rect 3525 15861 3559 15895
rect 3617 15861 3651 15895
rect 6193 15861 6227 15895
rect 7021 15861 7055 15895
rect 7757 15861 7791 15895
rect 8585 15861 8619 15895
rect 10517 15861 10551 15895
rect 11253 15861 11287 15895
rect 11989 15861 12023 15895
rect 12817 15861 12851 15895
rect 13553 15861 13587 15895
rect 16865 15861 16899 15895
rect 17141 15861 17175 15895
rect 21005 15861 21039 15895
rect 22753 15861 22787 15895
rect 3157 15657 3191 15691
rect 7113 15657 7147 15691
rect 9229 15657 9263 15691
rect 9689 15657 9723 15691
rect 10149 15657 10183 15691
rect 14749 15657 14783 15691
rect 14933 15657 14967 15691
rect 2044 15589 2078 15623
rect 6000 15589 6034 15623
rect 7634 15589 7668 15623
rect 8861 15589 8895 15623
rect 3433 15521 3467 15555
rect 4077 15521 4111 15555
rect 4997 15521 5031 15555
rect 5733 15521 5767 15555
rect 7389 15521 7423 15555
rect 1777 15453 1811 15487
rect 5089 15453 5123 15487
rect 5181 15453 5215 15487
rect 3617 15385 3651 15419
rect 4629 15385 4663 15419
rect 9045 15521 9079 15555
rect 10057 15521 10091 15555
rect 10968 15521 11002 15555
rect 12633 15521 12667 15555
rect 12992 15521 13026 15555
rect 14381 15521 14415 15555
rect 15546 15589 15580 15623
rect 15117 15521 15151 15555
rect 17224 15521 17258 15555
rect 18880 15521 18914 15555
rect 20085 15521 20119 15555
rect 20453 15521 20487 15555
rect 21005 15521 21039 15555
rect 21261 15521 21295 15555
rect 10241 15453 10275 15487
rect 10701 15453 10735 15487
rect 12725 15453 12759 15487
rect 14749 15453 14783 15487
rect 15301 15453 15335 15487
rect 16957 15453 16991 15487
rect 18613 15453 18647 15487
rect 12449 15385 12483 15419
rect 20269 15385 20303 15419
rect 20637 15385 20671 15419
rect 4261 15317 4295 15351
rect 8769 15317 8803 15351
rect 8953 15317 8987 15351
rect 12081 15317 12115 15351
rect 14105 15317 14139 15351
rect 14565 15317 14599 15351
rect 16681 15317 16715 15351
rect 18337 15317 18371 15351
rect 19993 15317 20027 15351
rect 22385 15317 22419 15351
rect 1593 15113 1627 15147
rect 3341 15113 3375 15147
rect 3617 15113 3651 15147
rect 4629 15113 4663 15147
rect 5641 15113 5675 15147
rect 7849 15113 7883 15147
rect 10241 15113 10275 15147
rect 19625 15113 19659 15147
rect 21925 15113 21959 15147
rect 6837 15045 6871 15079
rect 12081 15045 12115 15079
rect 15485 15045 15519 15079
rect 19901 15045 19935 15079
rect 4169 14977 4203 15011
rect 5181 14977 5215 15011
rect 6193 14977 6227 15011
rect 7297 14977 7331 15011
rect 7481 14977 7515 15011
rect 8401 14977 8435 15011
rect 8861 14977 8895 15011
rect 12456 14977 12490 15011
rect 20453 14977 20487 15011
rect 20729 14977 20763 15011
rect 21465 14977 21499 15011
rect 22477 14977 22511 15011
rect 1409 14909 1443 14943
rect 1961 14909 1995 14943
rect 2228 14909 2262 14943
rect 3985 14909 4019 14943
rect 6101 14909 6135 14943
rect 7205 14909 7239 14943
rect 8309 14909 8343 14943
rect 10701 14909 10735 14943
rect 10968 14909 11002 14943
rect 14105 14909 14139 14943
rect 14372 14909 14406 14943
rect 15761 14909 15795 14943
rect 16313 14909 16347 14943
rect 16580 14909 16614 14943
rect 18245 14909 18279 14943
rect 20361 14909 20395 14943
rect 4997 14841 5031 14875
rect 8217 14841 8251 14875
rect 9128 14841 9162 14875
rect 12716 14841 12750 14875
rect 18512 14841 18546 14875
rect 21281 14909 21315 14943
rect 22385 14841 22419 14875
rect 4077 14773 4111 14807
rect 5089 14773 5123 14807
rect 6009 14773 6043 14807
rect 13829 14773 13863 14807
rect 15945 14773 15979 14807
rect 17693 14773 17727 14807
rect 20269 14773 20303 14807
rect 20729 14773 20763 14807
rect 20913 14773 20947 14807
rect 21373 14773 21407 14807
rect 22293 14773 22327 14807
rect 3617 14569 3651 14603
rect 7113 14569 7147 14603
rect 7389 14569 7423 14603
rect 11069 14569 11103 14603
rect 12909 14569 12943 14603
rect 14289 14569 14323 14603
rect 15761 14569 15795 14603
rect 16129 14569 16163 14603
rect 16957 14569 16991 14603
rect 19533 14569 19567 14603
rect 22569 14569 22603 14603
rect 9956 14501 9990 14535
rect 13829 14501 13863 14535
rect 13921 14501 13955 14535
rect 14749 14501 14783 14535
rect 16497 14501 16531 14535
rect 19901 14501 19935 14535
rect 19993 14501 20027 14535
rect 21456 14501 21490 14535
rect 1501 14433 1535 14467
rect 1768 14433 1802 14467
rect 3341 14433 3375 14467
rect 3433 14433 3467 14467
rect 4344 14433 4378 14467
rect 6000 14433 6034 14467
rect 7757 14433 7791 14467
rect 8769 14433 8803 14467
rect 11796 14433 11830 14467
rect 13001 14433 13035 14467
rect 13369 14433 13403 14467
rect 14657 14433 14691 14467
rect 15669 14433 15703 14467
rect 17325 14433 17359 14467
rect 17877 14433 17911 14467
rect 18144 14433 18178 14467
rect 20729 14433 20763 14467
rect 4077 14365 4111 14399
rect 5733 14365 5767 14399
rect 7849 14365 7883 14399
rect 7941 14365 7975 14399
rect 8861 14365 8895 14399
rect 9045 14365 9079 14399
rect 9689 14365 9723 14399
rect 11529 14365 11563 14399
rect 14105 14365 14139 14399
rect 14933 14365 14967 14399
rect 15853 14365 15887 14399
rect 16589 14365 16623 14399
rect 16681 14365 16715 14399
rect 17417 14365 17451 14399
rect 17509 14365 17543 14399
rect 19349 14365 19383 14399
rect 20085 14365 20119 14399
rect 21189 14365 21223 14399
rect 13461 14297 13495 14331
rect 15301 14297 15335 14331
rect 2881 14229 2915 14263
rect 3157 14229 3191 14263
rect 5457 14229 5491 14263
rect 8401 14229 8435 14263
rect 13185 14229 13219 14263
rect 13369 14229 13403 14263
rect 19257 14229 19291 14263
rect 19349 14229 19383 14263
rect 20545 14229 20579 14263
rect 5089 14025 5123 14059
rect 8677 14025 8711 14059
rect 11989 14025 12023 14059
rect 15577 14025 15611 14059
rect 21925 14025 21959 14059
rect 1685 13957 1719 13991
rect 3433 13957 3467 13991
rect 5365 13957 5399 13991
rect 9781 13957 9815 13991
rect 12449 13957 12483 13991
rect 16405 13957 16439 13991
rect 17509 13957 17543 13991
rect 19441 13957 19475 13991
rect 21649 13957 21683 13991
rect 21741 13957 21775 13991
rect 6009 13889 6043 13923
rect 9229 13889 9263 13923
rect 10425 13889 10459 13923
rect 11437 13889 11471 13923
rect 12909 13889 12943 13923
rect 13093 13889 13127 13923
rect 16037 13889 16071 13923
rect 16129 13889 16163 13923
rect 16957 13889 16991 13923
rect 17693 13889 17727 13923
rect 18061 13889 18095 13923
rect 19809 13889 19843 13923
rect 20315 13889 20349 13923
rect 22477 13889 22511 13923
rect 1501 13821 1535 13855
rect 2053 13821 2087 13855
rect 2320 13821 2354 13855
rect 3709 13821 3743 13855
rect 3976 13821 4010 13855
rect 7021 13821 7055 13855
rect 7288 13821 7322 13855
rect 9137 13821 9171 13855
rect 11805 13821 11839 13855
rect 17325 13821 17359 13855
rect 18328 13821 18362 13855
rect 20545 13821 20579 13855
rect 21741 13821 21775 13855
rect 10149 13753 10183 13787
rect 11161 13753 11195 13787
rect 12817 13753 12851 13787
rect 13737 13753 13771 13787
rect 16773 13753 16807 13787
rect 22293 13753 22327 13787
rect 5733 13685 5767 13719
rect 5825 13685 5859 13719
rect 8401 13685 8435 13719
rect 9045 13685 9079 13719
rect 10241 13685 10275 13719
rect 10793 13685 10827 13719
rect 11253 13685 11287 13719
rect 15209 13685 15243 13719
rect 15945 13685 15979 13719
rect 16865 13685 16899 13719
rect 20275 13685 20309 13719
rect 22385 13685 22419 13719
rect 3065 13481 3099 13515
rect 5917 13481 5951 13515
rect 6377 13481 6411 13515
rect 8769 13481 8803 13515
rect 9781 13481 9815 13515
rect 11989 13481 12023 13515
rect 13461 13481 13495 13515
rect 16681 13481 16715 13515
rect 18797 13481 18831 13515
rect 1952 13413 1986 13447
rect 4804 13413 4838 13447
rect 7380 13413 7414 13447
rect 12326 13413 12360 13447
rect 1685 13345 1719 13379
rect 3433 13345 3467 13379
rect 4077 13345 4111 13379
rect 4537 13345 4571 13379
rect 6193 13345 6227 13379
rect 7113 13345 7147 13379
rect 8953 13345 8987 13379
rect 9045 13345 9079 13379
rect 10149 13345 10183 13379
rect 10241 13345 10275 13379
rect 10876 13345 10910 13379
rect 13820 13345 13854 13379
rect 15557 13345 15591 13379
rect 17224 13345 17258 13379
rect 18613 13345 18647 13379
rect 19421 13345 19455 13379
rect 20913 13345 20947 13379
rect 21189 13345 21223 13379
rect 21373 13345 21407 13379
rect 21640 13345 21674 13379
rect 10425 13277 10459 13311
rect 10609 13277 10643 13311
rect 12081 13277 12115 13311
rect 13553 13277 13587 13311
rect 15301 13277 15335 13311
rect 16957 13277 16991 13311
rect 19165 13277 19199 13311
rect 14933 13209 14967 13243
rect 3617 13141 3651 13175
rect 8493 13141 8527 13175
rect 9229 13141 9263 13175
rect 18337 13141 18371 13175
rect 20545 13141 20579 13175
rect 22753 13141 22787 13175
rect 2789 12937 2823 12971
rect 3249 12937 3283 12971
rect 8677 12937 8711 12971
rect 9689 12937 9723 12971
rect 11713 12937 11747 12971
rect 12173 12937 12207 12971
rect 19901 12937 19935 12971
rect 21741 12937 21775 12971
rect 6469 12869 6503 12903
rect 14381 12869 14415 12903
rect 18061 12869 18095 12903
rect 18889 12869 18923 12903
rect 1409 12801 1443 12835
rect 4169 12801 4203 12835
rect 4721 12801 4755 12835
rect 7021 12801 7055 12835
rect 9321 12801 9355 12835
rect 18613 12801 18647 12835
rect 19441 12801 19475 12835
rect 20269 12801 20303 12835
rect 22385 12801 22419 12835
rect 3065 12733 3099 12767
rect 4988 12733 5022 12767
rect 6653 12733 6687 12767
rect 7288 12733 7322 12767
rect 9873 12733 9907 12767
rect 9990 12733 10024 12767
rect 10333 12733 10367 12767
rect 10600 12733 10634 12767
rect 11989 12733 12023 12767
rect 12449 12733 12483 12767
rect 13001 12733 13035 12767
rect 14657 12733 14691 12767
rect 14924 12733 14958 12767
rect 16313 12733 16347 12767
rect 16580 12733 16614 12767
rect 17785 12733 17819 12767
rect 18429 12733 18463 12767
rect 19257 12733 19291 12767
rect 20085 12733 20119 12767
rect 20525 12733 20559 12767
rect 1676 12665 1710 12699
rect 3985 12665 4019 12699
rect 9137 12665 9171 12699
rect 12633 12665 12667 12699
rect 13268 12665 13302 12699
rect 18521 12665 18555 12699
rect 19349 12665 19383 12699
rect 22109 12665 22143 12699
rect 3617 12597 3651 12631
rect 4077 12597 4111 12631
rect 6101 12597 6135 12631
rect 8401 12597 8435 12631
rect 9045 12597 9079 12631
rect 10149 12597 10183 12631
rect 12817 12597 12851 12631
rect 16037 12597 16071 12631
rect 17693 12597 17727 12631
rect 17785 12597 17819 12631
rect 21649 12597 21683 12631
rect 22201 12597 22235 12631
rect 2053 12393 2087 12427
rect 4261 12393 4295 12427
rect 6009 12393 6043 12427
rect 8861 12393 8895 12427
rect 9229 12393 9263 12427
rect 9873 12393 9907 12427
rect 12725 12393 12759 12427
rect 14933 12393 14967 12427
rect 15669 12393 15703 12427
rect 17417 12393 17451 12427
rect 19165 12393 19199 12427
rect 3157 12325 3191 12359
rect 7288 12325 7322 12359
rect 18052 12325 18086 12359
rect 19901 12325 19935 12359
rect 21272 12325 21306 12359
rect 2145 12257 2179 12291
rect 3065 12257 3099 12291
rect 4077 12257 4111 12291
rect 4896 12257 4930 12291
rect 6469 12257 6503 12291
rect 7021 12257 7055 12291
rect 8677 12257 8711 12291
rect 9413 12257 9447 12291
rect 9505 12257 9539 12291
rect 9689 12257 9723 12291
rect 10425 12257 10459 12291
rect 11161 12257 11195 12291
rect 11345 12257 11379 12291
rect 11437 12257 11471 12291
rect 13544 12257 13578 12291
rect 14749 12257 14783 12291
rect 15485 12257 15519 12291
rect 16037 12257 16071 12291
rect 16304 12257 16338 12291
rect 17785 12257 17819 12291
rect 19809 12257 19843 12291
rect 21005 12257 21039 12291
rect 2329 12189 2363 12223
rect 3249 12189 3283 12223
rect 4629 12189 4663 12223
rect 1685 12121 1719 12155
rect 9505 12121 9539 12155
rect 10977 12121 11011 12155
rect 13277 12189 13311 12223
rect 19993 12189 20027 12223
rect 2697 12053 2731 12087
rect 6653 12053 6687 12087
rect 8401 12053 8435 12087
rect 10241 12053 10275 12087
rect 11345 12053 11379 12087
rect 14657 12053 14691 12087
rect 19441 12053 19475 12087
rect 22385 12053 22419 12087
rect 1501 11849 1535 11883
rect 3893 11849 3927 11883
rect 3985 11849 4019 11883
rect 5825 11849 5859 11883
rect 6377 11849 6411 11883
rect 11621 11849 11655 11883
rect 14197 11849 14231 11883
rect 15853 11849 15887 11883
rect 22477 11849 22511 11883
rect 4169 11781 4203 11815
rect 8493 11781 8527 11815
rect 16957 11781 16991 11815
rect 1961 11713 1995 11747
rect 2145 11713 2179 11747
rect 3985 11713 4019 11747
rect 9137 11713 9171 11747
rect 10241 11713 10275 11747
rect 12817 11713 12851 11747
rect 17417 11713 17451 11747
rect 17601 11713 17635 11747
rect 20177 11713 20211 11747
rect 20640 11713 20674 11747
rect 2513 11645 2547 11679
rect 4353 11645 4387 11679
rect 4445 11645 4479 11679
rect 6193 11645 6227 11679
rect 6837 11645 6871 11679
rect 8861 11645 8895 11679
rect 9689 11645 9723 11679
rect 10508 11645 10542 11679
rect 14473 11645 14507 11679
rect 14740 11645 14774 11679
rect 16497 11645 16531 11679
rect 16865 11645 16899 11679
rect 17325 11645 17359 11679
rect 18245 11645 18279 11679
rect 18512 11645 18546 11679
rect 20913 11645 20947 11679
rect 22293 11645 22327 11679
rect 2780 11577 2814 11611
rect 4712 11577 4746 11611
rect 7104 11577 7138 11611
rect 13084 11577 13118 11611
rect 16313 11577 16347 11611
rect 1869 11509 1903 11543
rect 8217 11509 8251 11543
rect 8953 11509 8987 11543
rect 9873 11509 9907 11543
rect 11897 11509 11931 11543
rect 16681 11509 16715 11543
rect 16865 11509 16899 11543
rect 19625 11509 19659 11543
rect 20643 11509 20677 11543
rect 22017 11509 22051 11543
rect 1593 11305 1627 11339
rect 5457 11305 5491 11339
rect 6101 11305 6135 11339
rect 11345 11305 11379 11339
rect 20913 11305 20947 11339
rect 2228 11237 2262 11271
rect 4322 11237 4356 11271
rect 6193 11237 6227 11271
rect 8953 11237 8987 11271
rect 14565 11237 14599 11271
rect 15844 11237 15878 11271
rect 19156 11237 19190 11271
rect 1409 11169 1443 11203
rect 4077 11169 4111 11203
rect 6929 11169 6963 11203
rect 7196 11169 7230 11203
rect 10232 11169 10266 11203
rect 11621 11169 11655 11203
rect 12449 11169 12483 11203
rect 12541 11169 12575 11203
rect 12808 11169 12842 11203
rect 15577 11169 15611 11203
rect 17233 11169 17267 11203
rect 17489 11169 17523 11203
rect 18889 11169 18923 11203
rect 21629 11169 21663 11203
rect 1961 11101 1995 11135
rect 6377 11101 6411 11135
rect 9045 11101 9079 11135
rect 9229 11101 9263 11135
rect 9965 11101 9999 11135
rect 14657 11101 14691 11135
rect 14749 11101 14783 11135
rect 21373 11101 21407 11135
rect 3341 11033 3375 11067
rect 8585 11033 8619 11067
rect 11805 11033 11839 11067
rect 18613 11033 18647 11067
rect 22753 11033 22787 11067
rect 5733 10965 5767 10999
rect 8309 10965 8343 10999
rect 12265 10965 12299 10999
rect 13921 10965 13955 10999
rect 14197 10965 14231 10999
rect 16957 10965 16991 10999
rect 20269 10965 20303 10999
rect 1501 10761 1535 10795
rect 1777 10761 1811 10795
rect 2145 10761 2179 10795
rect 4537 10761 4571 10795
rect 4813 10761 4847 10795
rect 5917 10761 5951 10795
rect 8217 10761 8251 10795
rect 11161 10761 11195 10795
rect 11621 10761 11655 10795
rect 18061 10761 18095 10795
rect 19073 10761 19107 10795
rect 21189 10761 21223 10795
rect 8401 10693 8435 10727
rect 9505 10693 9539 10727
rect 13829 10693 13863 10727
rect 16589 10693 16623 10727
rect 2789 10625 2823 10659
rect 5365 10625 5399 10659
rect 6653 10625 6687 10659
rect 1593 10557 1627 10591
rect 3157 10557 3191 10591
rect 5181 10557 5215 10591
rect 5273 10557 5307 10591
rect 6101 10557 6135 10591
rect 6193 10557 6227 10591
rect 3424 10489 3458 10523
rect 6837 10557 6871 10591
rect 7104 10557 7138 10591
rect 2513 10421 2547 10455
rect 2605 10421 2639 10455
rect 6377 10421 6411 10455
rect 6653 10421 6687 10455
rect 9137 10625 9171 10659
rect 14749 10625 14783 10659
rect 17509 10625 17543 10659
rect 18613 10625 18647 10659
rect 19812 10625 19846 10659
rect 22201 10625 22235 10659
rect 9689 10557 9723 10591
rect 9781 10557 9815 10591
rect 11437 10557 11471 10591
rect 12449 10557 12483 10591
rect 12716 10557 12750 10591
rect 14565 10557 14599 10591
rect 15209 10557 15243 10591
rect 15465 10557 15499 10591
rect 17325 10557 17359 10591
rect 19257 10557 19291 10591
rect 19349 10557 19383 10591
rect 20085 10557 20119 10591
rect 8953 10489 8987 10523
rect 10048 10489 10082 10523
rect 14657 10489 14691 10523
rect 18521 10489 18555 10523
rect 22109 10489 22143 10523
rect 8401 10421 8435 10455
rect 8493 10421 8527 10455
rect 8861 10421 8895 10455
rect 14197 10421 14231 10455
rect 16957 10421 16991 10455
rect 17417 10421 17451 10455
rect 18429 10421 18463 10455
rect 19815 10421 19849 10455
rect 21649 10421 21683 10455
rect 22017 10421 22051 10455
rect 2605 10217 2639 10251
rect 4077 10217 4111 10251
rect 4445 10217 4479 10251
rect 4537 10217 4571 10251
rect 5457 10217 5491 10251
rect 8493 10217 8527 10251
rect 9229 10217 9263 10251
rect 9413 10217 9447 10251
rect 3341 10149 3375 10183
rect 5549 10149 5583 10183
rect 7380 10149 7414 10183
rect 1869 10081 1903 10115
rect 2421 10081 2455 10115
rect 3433 10081 3467 10115
rect 6469 10081 6503 10115
rect 6561 10081 6595 10115
rect 9045 10081 9079 10115
rect 3617 10013 3651 10047
rect 4721 10013 4755 10047
rect 5733 10013 5767 10047
rect 6745 10013 6779 10047
rect 7113 10013 7147 10047
rect 9505 10217 9539 10251
rect 11069 10217 11103 10251
rect 11805 10217 11839 10251
rect 16681 10217 16715 10251
rect 18429 10217 18463 10251
rect 20545 10217 20579 10251
rect 22569 10217 22603 10251
rect 9934 10149 9968 10183
rect 11713 10149 11747 10183
rect 18705 10149 18739 10183
rect 21180 10149 21214 10183
rect 9505 10081 9539 10115
rect 9689 10081 9723 10115
rect 12633 10081 12667 10115
rect 12992 10081 13026 10115
rect 14381 10081 14415 10115
rect 15117 10081 15151 10115
rect 15301 10081 15335 10115
rect 15557 10081 15591 10115
rect 17049 10081 17083 10115
rect 17316 10081 17350 10115
rect 19165 10081 19199 10115
rect 19432 10081 19466 10115
rect 11897 10013 11931 10047
rect 12725 10013 12759 10047
rect 20913 10013 20947 10047
rect 9413 9945 9447 9979
rect 11345 9945 11379 9979
rect 14105 9945 14139 9979
rect 14565 9945 14599 9979
rect 22293 9945 22327 9979
rect 2053 9877 2087 9911
rect 2973 9877 3007 9911
rect 5089 9877 5123 9911
rect 6101 9877 6135 9911
rect 12449 9877 12483 9911
rect 14933 9877 14967 9911
rect 4537 9673 4571 9707
rect 10793 9673 10827 9707
rect 15853 9673 15887 9707
rect 16037 9673 16071 9707
rect 2789 9605 2823 9639
rect 3341 9605 3375 9639
rect 9137 9605 9171 9639
rect 11345 9605 11379 9639
rect 13461 9605 13495 9639
rect 4261 9537 4295 9571
rect 5181 9537 5215 9571
rect 6193 9537 6227 9571
rect 6377 9537 6411 9571
rect 7757 9537 7791 9571
rect 9413 9537 9447 9571
rect 11897 9537 11931 9571
rect 13093 9537 13127 9571
rect 14013 9537 14047 9571
rect 1409 9469 1443 9503
rect 3157 9469 3191 9503
rect 4905 9469 4939 9503
rect 4997 9469 5031 9503
rect 5641 9469 5675 9503
rect 6101 9469 6135 9503
rect 7205 9469 7239 9503
rect 8024 9469 8058 9503
rect 9669 9469 9703 9503
rect 11713 9469 11747 9503
rect 14473 9469 14507 9503
rect 14740 9469 14774 9503
rect 1654 9401 1688 9435
rect 4169 9401 4203 9435
rect 12817 9401 12851 9435
rect 16129 9605 16163 9639
rect 19993 9605 20027 9639
rect 20177 9605 20211 9639
rect 16773 9537 16807 9571
rect 18524 9537 18558 9571
rect 18797 9537 18831 9571
rect 17141 9469 17175 9503
rect 17877 9469 17911 9503
rect 18061 9469 18095 9503
rect 18384 9469 18418 9503
rect 16497 9401 16531 9435
rect 20729 9537 20763 9571
rect 21373 9537 21407 9571
rect 20545 9469 20579 9503
rect 21640 9469 21674 9503
rect 20637 9401 20671 9435
rect 3709 9333 3743 9367
rect 4077 9333 4111 9367
rect 5733 9333 5767 9367
rect 7389 9333 7423 9367
rect 11805 9333 11839 9367
rect 12449 9333 12483 9367
rect 12909 9333 12943 9367
rect 13829 9333 13863 9367
rect 13921 9333 13955 9367
rect 16037 9333 16071 9367
rect 16589 9333 16623 9367
rect 17325 9333 17359 9367
rect 17693 9333 17727 9367
rect 19901 9333 19935 9367
rect 19993 9333 20027 9367
rect 22753 9333 22787 9367
rect 2973 9129 3007 9163
rect 4721 9129 4755 9163
rect 6193 9129 6227 9163
rect 6745 9129 6779 9163
rect 7113 9129 7147 9163
rect 7757 9129 7791 9163
rect 8125 9129 8159 9163
rect 8769 9129 8803 9163
rect 9689 9129 9723 9163
rect 10057 9129 10091 9163
rect 12633 9129 12667 9163
rect 13185 9129 13219 9163
rect 14933 9129 14967 9163
rect 15301 9129 15335 9163
rect 15669 9129 15703 9163
rect 16497 9129 16531 9163
rect 21925 9129 21959 9163
rect 5089 9061 5123 9095
rect 7205 9061 7239 9095
rect 17224 9061 17258 9095
rect 21281 9061 21315 9095
rect 22385 9061 22419 9095
rect 3433 8993 3467 9027
rect 4169 8993 4203 9027
rect 5181 8993 5215 9027
rect 6101 8993 6135 9027
rect 8217 8993 8251 9027
rect 8961 8993 8995 9027
rect 9070 8993 9104 9027
rect 10149 8993 10183 9027
rect 10701 8993 10735 9027
rect 11520 8993 11554 9027
rect 13001 8993 13035 9027
rect 13553 8993 13587 9027
rect 13820 8993 13854 9027
rect 16313 8993 16347 9027
rect 16957 8993 16991 9027
rect 19053 8993 19087 9027
rect 22293 8993 22327 9027
rect 5273 8925 5307 8959
rect 6377 8925 6411 8959
rect 7389 8925 7423 8959
rect 8401 8925 8435 8959
rect 10241 8925 10275 8959
rect 11253 8925 11287 8959
rect 15761 8925 15795 8959
rect 15853 8925 15887 8959
rect 18797 8925 18831 8959
rect 21373 8925 21407 8959
rect 21465 8925 21499 8959
rect 22477 8925 22511 8959
rect 3617 8857 3651 8891
rect 4353 8789 4387 8823
rect 5733 8789 5767 8823
rect 9229 8789 9263 8823
rect 10885 8789 10919 8823
rect 18337 8789 18371 8823
rect 20177 8789 20211 8823
rect 20913 8789 20947 8823
rect 4353 8585 4387 8619
rect 7021 8585 7055 8619
rect 10333 8585 10367 8619
rect 12081 8585 12115 8619
rect 15485 8585 15519 8619
rect 18889 8585 18923 8619
rect 19717 8585 19751 8619
rect 4721 8517 4755 8551
rect 5733 8517 5767 8551
rect 7389 8517 7423 8551
rect 10609 8517 10643 8551
rect 13829 8517 13863 8551
rect 17693 8517 17727 8551
rect 18797 8517 18831 8551
rect 1961 8449 1995 8483
rect 5365 8449 5399 8483
rect 6285 8449 6319 8483
rect 7941 8449 7975 8483
rect 1777 8381 1811 8415
rect 4169 8381 4203 8415
rect 6837 8381 6871 8415
rect 8401 8381 8435 8415
rect 10149 8381 10183 8415
rect 5181 8313 5215 8347
rect 6193 8313 6227 8347
rect 7849 8313 7883 8347
rect 8668 8313 8702 8347
rect 12449 8449 12483 8483
rect 14105 8449 14139 8483
rect 15853 8449 15887 8483
rect 16316 8449 16350 8483
rect 16589 8449 16623 8483
rect 18429 8449 18463 8483
rect 19349 8449 19383 8483
rect 19441 8449 19475 8483
rect 19717 8449 19751 8483
rect 20224 8449 20258 8483
rect 20364 8449 20398 8483
rect 20637 8449 20671 8483
rect 22477 8449 22511 8483
rect 22661 8449 22695 8483
rect 10701 8381 10735 8415
rect 18153 8381 18187 8415
rect 18797 8381 18831 8415
rect 19901 8381 19935 8415
rect 10968 8313 11002 8347
rect 12694 8313 12728 8347
rect 14372 8313 14406 8347
rect 22385 8313 22419 8347
rect 5089 8245 5123 8279
rect 6101 8245 6135 8279
rect 7757 8245 7791 8279
rect 9781 8245 9815 8279
rect 10609 8245 10643 8279
rect 16319 8245 16353 8279
rect 19257 8245 19291 8279
rect 21741 8245 21775 8279
rect 22017 8245 22051 8279
rect 4629 8041 4663 8075
rect 5089 8041 5123 8075
rect 5549 8041 5583 8075
rect 6009 8041 6043 8075
rect 7849 8041 7883 8075
rect 6101 7973 6135 8007
rect 9505 8041 9539 8075
rect 9689 8041 9723 8075
rect 12541 8041 12575 8075
rect 13277 8041 13311 8075
rect 14197 8041 14231 8075
rect 14841 8041 14875 8075
rect 15767 8041 15801 8075
rect 17141 8041 17175 8075
rect 17969 8041 18003 8075
rect 20453 8041 20487 8075
rect 4905 7905 4939 7939
rect 6837 7905 6871 7939
rect 7481 7905 7515 7939
rect 7849 7905 7883 7939
rect 8208 7905 8242 7939
rect 11428 7973 11462 8007
rect 14289 7973 14323 8007
rect 21548 7973 21582 8007
rect 10057 7905 10091 7939
rect 11161 7905 11195 7939
rect 13185 7905 13219 7939
rect 15025 7905 15059 7939
rect 15301 7905 15335 7939
rect 16037 7905 16071 7939
rect 18061 7905 18095 7939
rect 18613 7905 18647 7939
rect 18936 7905 18970 7939
rect 19349 7905 19383 7939
rect 21281 7905 21315 7939
rect 6285 7837 6319 7871
rect 7941 7837 7975 7871
rect 9505 7837 9539 7871
rect 10149 7837 10183 7871
rect 10241 7837 10275 7871
rect 10701 7837 10735 7871
rect 13369 7837 13403 7871
rect 14381 7837 14415 7871
rect 15764 7837 15798 7871
rect 18245 7837 18279 7871
rect 19119 7837 19153 7871
rect 5641 7769 5675 7803
rect 12817 7769 12851 7803
rect 9321 7701 9355 7735
rect 13829 7701 13863 7735
rect 17601 7701 17635 7735
rect 22661 7701 22695 7735
rect 6377 7497 6411 7531
rect 7205 7497 7239 7531
rect 7573 7497 7607 7531
rect 9965 7497 9999 7531
rect 15669 7497 15703 7531
rect 17693 7497 17727 7531
rect 20177 7497 20211 7531
rect 22569 7497 22603 7531
rect 18429 7429 18463 7463
rect 7389 7361 7423 7395
rect 8125 7361 8159 7395
rect 10241 7361 10275 7395
rect 13001 7361 13035 7395
rect 20729 7361 20763 7395
rect 5641 7293 5675 7327
rect 6193 7293 6227 7327
rect 7021 7293 7055 7327
rect 8585 7293 8619 7327
rect 8852 7293 8886 7327
rect 11897 7293 11931 7327
rect 13645 7293 13679 7327
rect 13737 7293 13771 7327
rect 14289 7293 14323 7327
rect 16129 7293 16163 7327
rect 16221 7293 16255 7327
rect 16313 7293 16347 7327
rect 18245 7293 18279 7327
rect 18797 7293 18831 7327
rect 20453 7293 20487 7327
rect 21189 7293 21223 7327
rect 21456 7293 21490 7327
rect 8033 7225 8067 7259
rect 10486 7225 10520 7259
rect 12909 7225 12943 7259
rect 14556 7225 14590 7259
rect 16580 7225 16614 7259
rect 19064 7225 19098 7259
rect 5825 7157 5859 7191
rect 7389 7157 7423 7191
rect 7941 7157 7975 7191
rect 11621 7157 11655 7191
rect 12449 7157 12483 7191
rect 12817 7157 12851 7191
rect 13461 7157 13495 7191
rect 13921 7157 13955 7191
rect 15945 7157 15979 7191
rect 16221 7157 16255 7191
rect 7481 6953 7515 6987
rect 13737 6953 13771 6987
rect 19165 6953 19199 6987
rect 19809 6953 19843 6987
rect 22293 6953 22327 6987
rect 9045 6885 9079 6919
rect 12725 6885 12759 6919
rect 6469 6817 6503 6851
rect 6837 6817 6871 6851
rect 7941 6817 7975 6851
rect 8033 6817 8067 6851
rect 8953 6817 8987 6851
rect 9956 6817 9990 6851
rect 11713 6817 11747 6851
rect 14197 6817 14231 6851
rect 14381 6817 14415 6851
rect 14565 6817 14599 6851
rect 15568 6817 15602 6851
rect 17213 6817 17247 6851
rect 20177 6817 20211 6851
rect 21180 6817 21214 6851
rect 22569 6817 22603 6851
rect 23397 6817 23431 6851
rect 8217 6749 8251 6783
rect 9229 6749 9263 6783
rect 9689 6749 9723 6783
rect 11805 6749 11839 6783
rect 11897 6749 11931 6783
rect 12817 6749 12851 6783
rect 13001 6749 13035 6783
rect 13829 6749 13863 6783
rect 14013 6749 14047 6783
rect 7573 6681 7607 6715
rect 8585 6681 8619 6715
rect 15301 6749 15335 6783
rect 16957 6749 16991 6783
rect 19257 6749 19291 6783
rect 19349 6749 19383 6783
rect 20269 6749 20303 6783
rect 20361 6749 20395 6783
rect 20913 6749 20947 6783
rect 14749 6681 14783 6715
rect 16681 6681 16715 6715
rect 6653 6613 6687 6647
rect 7021 6613 7055 6647
rect 11069 6613 11103 6647
rect 11345 6613 11379 6647
rect 12357 6613 12391 6647
rect 13369 6613 13403 6647
rect 14197 6613 14231 6647
rect 18337 6613 18371 6647
rect 18797 6613 18831 6647
rect 7849 6409 7883 6443
rect 10149 6409 10183 6443
rect 14289 6409 14323 6443
rect 15945 6409 15979 6443
rect 16957 6409 16991 6443
rect 20913 6409 20947 6443
rect 8401 6341 8435 6375
rect 8769 6273 8803 6307
rect 10885 6273 10919 6307
rect 10977 6273 11011 6307
rect 12909 6273 12943 6307
rect 17601 6273 17635 6307
rect 19073 6273 19107 6307
rect 19533 6273 19567 6307
rect 22109 6273 22143 6307
rect 7665 6205 7699 6239
rect 8217 6205 8251 6239
rect 10793 6205 10827 6239
rect 11621 6205 11655 6239
rect 11805 6205 11839 6239
rect 12449 6205 12483 6239
rect 14565 6205 14599 6239
rect 14821 6205 14855 6239
rect 16405 6205 16439 6239
rect 22569 6205 22603 6239
rect 9014 6137 9048 6171
rect 13176 6137 13210 6171
rect 18981 6137 19015 6171
rect 19778 6137 19812 6171
rect 21925 6137 21959 6171
rect 10425 6069 10459 6103
rect 11437 6069 11471 6103
rect 11989 6069 12023 6103
rect 16589 6069 16623 6103
rect 17325 6069 17359 6103
rect 17417 6069 17451 6103
rect 18061 6069 18095 6103
rect 18521 6069 18555 6103
rect 18889 6069 18923 6103
rect 21557 6069 21591 6103
rect 22017 6069 22051 6103
rect 8125 5865 8159 5899
rect 9413 5865 9447 5899
rect 8953 5797 8987 5831
rect 12909 5865 12943 5899
rect 14381 5865 14415 5899
rect 17509 5865 17543 5899
rect 18245 5865 18279 5899
rect 20177 5865 20211 5899
rect 23397 5865 23431 5899
rect 22569 5797 22603 5831
rect 9956 5729 9990 5763
rect 11612 5729 11646 5763
rect 12909 5729 12943 5763
rect 13001 5729 13035 5763
rect 13268 5729 13302 5763
rect 14657 5729 14691 5763
rect 15577 5729 15611 5763
rect 16396 5729 16430 5763
rect 18153 5729 18187 5763
rect 18797 5729 18831 5763
rect 19064 5729 19098 5763
rect 21649 5729 21683 5763
rect 22293 5729 22327 5763
rect 9045 5661 9079 5695
rect 9229 5661 9263 5695
rect 9413 5661 9447 5695
rect 9689 5661 9723 5695
rect 11345 5661 11379 5695
rect 8585 5593 8619 5627
rect 11069 5593 11103 5627
rect 12725 5593 12759 5627
rect 16129 5661 16163 5695
rect 18337 5661 18371 5695
rect 21741 5661 21775 5695
rect 21833 5661 21867 5695
rect 14841 5593 14875 5627
rect 12909 5525 12943 5559
rect 15761 5525 15795 5559
rect 17785 5525 17819 5559
rect 21281 5525 21315 5559
rect 9597 5321 9631 5355
rect 11345 5321 11379 5355
rect 15117 5321 15151 5355
rect 17693 5321 17727 5355
rect 18061 5321 18095 5355
rect 20361 5321 20395 5355
rect 13829 5253 13863 5287
rect 19257 5253 19291 5287
rect 14565 5185 14599 5219
rect 14657 5185 14691 5219
rect 15669 5185 15703 5219
rect 16313 5185 16347 5219
rect 18521 5185 18555 5219
rect 18613 5185 18647 5219
rect 19809 5185 19843 5219
rect 20821 5185 20855 5219
rect 20913 5185 20947 5219
rect 9413 5117 9447 5151
rect 9965 5117 9999 5151
rect 10232 5117 10266 5151
rect 11805 5117 11839 5151
rect 12449 5117 12483 5151
rect 12716 5117 12750 5151
rect 16580 5117 16614 5151
rect 20729 5117 20763 5151
rect 21373 5117 21407 5151
rect 15485 5049 15519 5083
rect 21618 5049 21652 5083
rect 8953 4981 8987 5015
rect 11989 4981 12023 5015
rect 14105 4981 14139 5015
rect 14473 4981 14507 5015
rect 15577 4981 15611 5015
rect 18429 4981 18463 5015
rect 19625 4981 19659 5015
rect 19717 4981 19751 5015
rect 22753 4981 22787 5015
rect 10149 4777 10183 4811
rect 10609 4777 10643 4811
rect 12725 4777 12759 4811
rect 13001 4777 13035 4811
rect 13369 4777 13403 4811
rect 13461 4777 13495 4811
rect 14381 4777 14415 4811
rect 15485 4777 15519 4811
rect 17509 4777 17543 4811
rect 19717 4777 19751 4811
rect 22753 4777 22787 4811
rect 10517 4709 10551 4743
rect 11612 4709 11646 4743
rect 16120 4709 16154 4743
rect 20913 4709 20947 4743
rect 15301 4641 15335 4675
rect 17877 4641 17911 4675
rect 18889 4641 18923 4675
rect 20085 4641 20119 4675
rect 21640 4641 21674 4675
rect 10793 4573 10827 4607
rect 11345 4573 11379 4607
rect 13553 4573 13587 4607
rect 14473 4573 14507 4607
rect 14657 4573 14691 4607
rect 15853 4573 15887 4607
rect 17969 4573 18003 4607
rect 18061 4573 18095 4607
rect 18981 4573 19015 4607
rect 19073 4573 19107 4607
rect 20177 4573 20211 4607
rect 20269 4573 20303 4607
rect 21373 4573 21407 4607
rect 14013 4505 14047 4539
rect 17233 4437 17267 4471
rect 18521 4437 18555 4471
rect 13737 4233 13771 4267
rect 17141 4233 17175 4267
rect 19717 4233 19751 4267
rect 11897 4097 11931 4131
rect 13277 4097 13311 4131
rect 14289 4097 14323 4131
rect 14657 4097 14691 4131
rect 15301 4097 15335 4131
rect 20269 4097 20303 4131
rect 10793 4029 10827 4063
rect 11713 4029 11747 4063
rect 13185 4029 13219 4063
rect 14197 4029 14231 4063
rect 11805 3961 11839 3995
rect 15117 4029 15151 4063
rect 15761 4029 15795 4063
rect 16028 4029 16062 4063
rect 17417 4029 17451 4063
rect 18061 4029 18095 4063
rect 20729 4029 20763 4063
rect 20913 4029 20947 4063
rect 21373 4029 21407 4063
rect 21640 4029 21674 4063
rect 18328 3961 18362 3995
rect 20177 3961 20211 3995
rect 21097 3961 21131 3995
rect 10977 3893 11011 3927
rect 11345 3893 11379 3927
rect 12725 3893 12759 3927
rect 13093 3893 13127 3927
rect 14105 3893 14139 3927
rect 14657 3893 14691 3927
rect 14749 3893 14783 3927
rect 15209 3893 15243 3927
rect 17601 3893 17635 3927
rect 19441 3893 19475 3927
rect 20085 3893 20119 3927
rect 22753 3893 22787 3927
rect 12817 3689 12851 3723
rect 18889 3689 18923 3723
rect 22293 3689 22327 3723
rect 3249 3621 3283 3655
rect 14657 3621 14691 3655
rect 16120 3621 16154 3655
rect 19432 3621 19466 3655
rect 21180 3621 21214 3655
rect 2513 3553 2547 3587
rect 11989 3553 12023 3587
rect 12633 3553 12667 3587
rect 13553 3553 13587 3587
rect 14565 3553 14599 3587
rect 15301 3553 15335 3587
rect 17776 3553 17810 3587
rect 19165 3553 19199 3587
rect 13645 3485 13679 3519
rect 13829 3485 13863 3519
rect 14749 3485 14783 3519
rect 15853 3485 15887 3519
rect 17509 3485 17543 3519
rect 20913 3485 20947 3519
rect 12173 3417 12207 3451
rect 14197 3417 14231 3451
rect 17233 3417 17267 3451
rect 13185 3349 13219 3383
rect 15485 3349 15519 3383
rect 20545 3349 20579 3383
rect 13093 3145 13127 3179
rect 14013 3145 14047 3179
rect 17417 3145 17451 3179
rect 20269 3145 20303 3179
rect 21925 3145 21959 3179
rect 15025 3077 15059 3111
rect 18521 3077 18555 3111
rect 1961 3009 1995 3043
rect 14657 3009 14691 3043
rect 15577 3009 15611 3043
rect 16037 3009 16071 3043
rect 1777 2941 1811 2975
rect 2513 2941 2547 2975
rect 5089 2941 5123 2975
rect 12909 2941 12943 2975
rect 13461 2941 13495 2975
rect 15393 2941 15427 2975
rect 16304 2941 16338 2975
rect 18337 2941 18371 2975
rect 18889 2941 18923 2975
rect 19156 2941 19190 2975
rect 20545 2941 20579 2975
rect 20812 2941 20846 2975
rect 22201 2941 22235 2975
rect 14381 2873 14415 2907
rect 15485 2873 15519 2907
rect 22477 2873 22511 2907
rect 2697 2805 2731 2839
rect 13645 2805 13679 2839
rect 14473 2805 14507 2839
rect 14013 2601 14047 2635
rect 14749 2601 14783 2635
rect 15853 2601 15887 2635
rect 17877 2601 17911 2635
rect 18705 2601 18739 2635
rect 20729 2601 20763 2635
rect 22569 2601 22603 2635
rect 16764 2533 16798 2567
rect 18797 2533 18831 2567
rect 19616 2533 19650 2567
rect 21456 2533 21490 2567
rect 13829 2465 13863 2499
rect 15945 2465 15979 2499
rect 16497 2465 16531 2499
rect 19349 2465 19383 2499
rect 21189 2465 21223 2499
rect 14841 2397 14875 2431
rect 15025 2397 15059 2431
rect 16037 2397 16071 2431
rect 18981 2397 19015 2431
rect 15485 2329 15519 2363
rect 14381 2261 14415 2295
rect 18337 2261 18371 2295
<< metal1 >>
rect 8570 22856 8576 22908
rect 8628 22896 8634 22908
rect 9490 22896 9496 22908
rect 8628 22868 9496 22896
rect 8628 22856 8634 22868
rect 9490 22856 9496 22868
rect 9548 22856 9554 22908
rect 15378 22856 15384 22908
rect 15436 22896 15442 22908
rect 19426 22896 19432 22908
rect 15436 22868 19432 22896
rect 15436 22856 15442 22868
rect 19426 22856 19432 22868
rect 19484 22856 19490 22908
rect 17678 22584 17684 22636
rect 17736 22624 17742 22636
rect 19334 22624 19340 22636
rect 17736 22596 19340 22624
rect 17736 22584 17742 22596
rect 19334 22584 19340 22596
rect 19392 22584 19398 22636
rect 18322 22312 18328 22364
rect 18380 22352 18386 22364
rect 19794 22352 19800 22364
rect 18380 22324 19800 22352
rect 18380 22312 18386 22324
rect 19794 22312 19800 22324
rect 19852 22312 19858 22364
rect 9214 22108 9220 22160
rect 9272 22148 9278 22160
rect 10962 22148 10968 22160
rect 9272 22120 10968 22148
rect 9272 22108 9278 22120
rect 10962 22108 10968 22120
rect 11020 22108 11026 22160
rect 12345 22151 12403 22157
rect 12345 22117 12357 22151
rect 12391 22148 12403 22151
rect 19245 22151 19303 22157
rect 19245 22148 19257 22151
rect 12391 22120 19257 22148
rect 12391 22117 12403 22120
rect 12345 22111 12403 22117
rect 19245 22117 19257 22120
rect 19291 22117 19303 22151
rect 19245 22111 19303 22117
rect 7926 22040 7932 22092
rect 7984 22080 7990 22092
rect 9398 22080 9404 22092
rect 7984 22052 9404 22080
rect 7984 22040 7990 22052
rect 9398 22040 9404 22052
rect 9456 22040 9462 22092
rect 9674 22040 9680 22092
rect 9732 22080 9738 22092
rect 21634 22080 21640 22092
rect 9732 22052 21640 22080
rect 9732 22040 9738 22052
rect 21634 22040 21640 22052
rect 21692 22040 21698 22092
rect 8754 21972 8760 22024
rect 8812 22012 8818 22024
rect 11701 22015 11759 22021
rect 11701 22012 11713 22015
rect 8812 21984 11713 22012
rect 8812 21972 8818 21984
rect 11701 21981 11713 21984
rect 11747 21981 11759 22015
rect 11701 21975 11759 21981
rect 12710 21972 12716 22024
rect 12768 22012 12774 22024
rect 16942 22012 16948 22024
rect 12768 21984 16948 22012
rect 12768 21972 12774 21984
rect 16942 21972 16948 21984
rect 17000 21972 17006 22024
rect 2038 21904 2044 21956
rect 2096 21944 2102 21956
rect 10042 21944 10048 21956
rect 2096 21916 10048 21944
rect 2096 21904 2102 21916
rect 10042 21904 10048 21916
rect 10100 21944 10106 21956
rect 12345 21947 12403 21953
rect 12345 21944 12357 21947
rect 10100 21916 12357 21944
rect 10100 21904 10106 21916
rect 12345 21913 12357 21916
rect 12391 21913 12403 21947
rect 12345 21907 12403 21913
rect 13446 21904 13452 21956
rect 13504 21944 13510 21956
rect 19150 21944 19156 21956
rect 13504 21916 19156 21944
rect 13504 21904 13510 21916
rect 19150 21904 19156 21916
rect 19208 21904 19214 21956
rect 19245 21947 19303 21953
rect 19245 21913 19257 21947
rect 19291 21944 19303 21947
rect 19610 21944 19616 21956
rect 19291 21916 19616 21944
rect 19291 21913 19303 21916
rect 19245 21907 19303 21913
rect 19610 21904 19616 21916
rect 19668 21904 19674 21956
rect 6638 21836 6644 21888
rect 6696 21876 6702 21888
rect 7742 21876 7748 21888
rect 6696 21848 7748 21876
rect 6696 21836 6702 21848
rect 7742 21836 7748 21848
rect 7800 21836 7806 21888
rect 8202 21836 8208 21888
rect 8260 21876 8266 21888
rect 11606 21876 11612 21888
rect 8260 21848 11612 21876
rect 8260 21836 8266 21848
rect 11606 21836 11612 21848
rect 11664 21836 11670 21888
rect 11701 21879 11759 21885
rect 11701 21845 11713 21879
rect 11747 21876 11759 21879
rect 14182 21876 14188 21888
rect 11747 21848 14188 21876
rect 11747 21845 11759 21848
rect 11701 21839 11759 21845
rect 14182 21836 14188 21848
rect 14240 21836 14246 21888
rect 19794 21836 19800 21888
rect 19852 21876 19858 21888
rect 20622 21876 20628 21888
rect 19852 21848 20628 21876
rect 19852 21836 19858 21848
rect 20622 21836 20628 21848
rect 20680 21836 20686 21888
rect 1104 21786 23276 21808
rect 1104 21734 4680 21786
rect 4732 21734 4744 21786
rect 4796 21734 4808 21786
rect 4860 21734 4872 21786
rect 4924 21734 12078 21786
rect 12130 21734 12142 21786
rect 12194 21734 12206 21786
rect 12258 21734 12270 21786
rect 12322 21734 19475 21786
rect 19527 21734 19539 21786
rect 19591 21734 19603 21786
rect 19655 21734 19667 21786
rect 19719 21734 23276 21786
rect 1104 21712 23276 21734
rect 5905 21675 5963 21681
rect 2700 21644 4752 21672
rect 2409 21539 2467 21545
rect 2409 21505 2421 21539
rect 2455 21536 2467 21539
rect 2700 21536 2728 21644
rect 4724 21604 4752 21644
rect 5905 21641 5917 21675
rect 5951 21672 5963 21675
rect 9125 21675 9183 21681
rect 9125 21672 9137 21675
rect 5951 21644 9137 21672
rect 5951 21641 5963 21644
rect 5905 21635 5963 21641
rect 9125 21641 9137 21644
rect 9171 21641 9183 21675
rect 10042 21672 10048 21684
rect 10003 21644 10048 21672
rect 9125 21635 9183 21641
rect 10042 21632 10048 21644
rect 10100 21632 10106 21684
rect 17313 21675 17371 21681
rect 17313 21672 17325 21675
rect 10152 21644 17325 21672
rect 5626 21604 5632 21616
rect 4724 21576 5632 21604
rect 2455 21508 2728 21536
rect 2455 21505 2467 21508
rect 2409 21499 2467 21505
rect 3050 21496 3056 21548
rect 3108 21536 3114 21548
rect 4724 21545 4752 21576
rect 5626 21564 5632 21576
rect 5684 21564 5690 21616
rect 6917 21607 6975 21613
rect 6917 21573 6929 21607
rect 6963 21604 6975 21607
rect 8386 21604 8392 21616
rect 6963 21576 8392 21604
rect 6963 21573 6975 21576
rect 6917 21567 6975 21573
rect 8386 21564 8392 21576
rect 8444 21564 8450 21616
rect 10152 21604 10180 21644
rect 17313 21641 17325 21644
rect 17359 21641 17371 21675
rect 17313 21635 17371 21641
rect 17586 21632 17592 21684
rect 17644 21672 17650 21684
rect 17681 21675 17739 21681
rect 17681 21672 17693 21675
rect 17644 21644 17693 21672
rect 17644 21632 17650 21644
rect 17681 21641 17693 21644
rect 17727 21641 17739 21675
rect 17681 21635 17739 21641
rect 18966 21632 18972 21684
rect 19024 21672 19030 21684
rect 20901 21675 20959 21681
rect 20901 21672 20913 21675
rect 19024 21644 20913 21672
rect 19024 21632 19030 21644
rect 20901 21641 20913 21644
rect 20947 21641 20959 21675
rect 24026 21672 24032 21684
rect 20901 21635 20959 21641
rect 21100 21644 24032 21672
rect 11330 21604 11336 21616
rect 8496 21576 10180 21604
rect 10520 21576 11336 21604
rect 3329 21539 3387 21545
rect 3329 21536 3341 21539
rect 3108 21508 3341 21536
rect 3108 21496 3114 21508
rect 3329 21505 3341 21508
rect 3375 21505 3387 21539
rect 3329 21499 3387 21505
rect 4709 21539 4767 21545
rect 4709 21505 4721 21539
rect 4755 21505 4767 21539
rect 4709 21499 4767 21505
rect 5258 21496 5264 21548
rect 5316 21536 5322 21548
rect 5537 21539 5595 21545
rect 5537 21536 5549 21539
rect 5316 21508 5549 21536
rect 5316 21496 5322 21508
rect 5537 21505 5549 21508
rect 5583 21505 5595 21539
rect 5537 21499 5595 21505
rect 5721 21539 5779 21545
rect 5721 21505 5733 21539
rect 5767 21536 5779 21539
rect 6638 21536 6644 21548
rect 5767 21508 6644 21536
rect 5767 21505 5779 21508
rect 5721 21499 5779 21505
rect 6638 21496 6644 21508
rect 6696 21496 6702 21548
rect 6730 21496 6736 21548
rect 6788 21536 6794 21548
rect 7469 21539 7527 21545
rect 7469 21536 7481 21539
rect 6788 21508 7481 21536
rect 6788 21496 6794 21508
rect 7469 21505 7481 21508
rect 7515 21505 7527 21539
rect 7469 21499 7527 21505
rect 7650 21496 7656 21548
rect 7708 21536 7714 21548
rect 8496 21536 8524 21576
rect 7708 21508 8524 21536
rect 8573 21539 8631 21545
rect 7708 21496 7714 21508
rect 8573 21505 8585 21539
rect 8619 21536 8631 21539
rect 8662 21536 8668 21548
rect 8619 21508 8668 21536
rect 8619 21505 8631 21508
rect 8573 21499 8631 21505
rect 8662 21496 8668 21508
rect 8720 21496 8726 21548
rect 10520 21545 10548 21576
rect 11330 21564 11336 21576
rect 11388 21564 11394 21616
rect 11422 21564 11428 21616
rect 11480 21604 11486 21616
rect 11882 21604 11888 21616
rect 11480 21576 11888 21604
rect 11480 21564 11486 21576
rect 11882 21564 11888 21576
rect 11940 21564 11946 21616
rect 15013 21607 15071 21613
rect 15013 21573 15025 21607
rect 15059 21604 15071 21607
rect 20530 21604 20536 21616
rect 15059 21576 17080 21604
rect 15059 21573 15071 21576
rect 15013 21567 15071 21573
rect 10505 21539 10563 21545
rect 10505 21505 10517 21539
rect 10551 21505 10563 21539
rect 10505 21499 10563 21505
rect 10689 21539 10747 21545
rect 10689 21505 10701 21539
rect 10735 21536 10747 21539
rect 11514 21536 11520 21548
rect 10735 21508 11520 21536
rect 10735 21505 10747 21508
rect 10689 21499 10747 21505
rect 11514 21496 11520 21508
rect 11572 21496 11578 21548
rect 11606 21496 11612 21548
rect 11664 21536 11670 21548
rect 11664 21508 11709 21536
rect 11664 21496 11670 21508
rect 11974 21496 11980 21548
rect 12032 21536 12038 21548
rect 13173 21539 13231 21545
rect 13173 21536 13185 21539
rect 12032 21508 13185 21536
rect 12032 21496 12038 21508
rect 13173 21505 13185 21508
rect 13219 21505 13231 21539
rect 14182 21536 14188 21548
rect 14143 21508 14188 21536
rect 13173 21499 13231 21505
rect 14182 21496 14188 21508
rect 14240 21496 14246 21548
rect 16117 21539 16175 21545
rect 14844 21508 16068 21536
rect 2866 21428 2872 21480
rect 2924 21468 2930 21480
rect 5445 21471 5503 21477
rect 2924 21440 4568 21468
rect 2924 21428 2930 21440
rect 1578 21360 1584 21412
rect 1636 21400 1642 21412
rect 2133 21403 2191 21409
rect 2133 21400 2145 21403
rect 1636 21372 2145 21400
rect 1636 21360 1642 21372
rect 2133 21369 2145 21372
rect 2179 21369 2191 21403
rect 4433 21403 4491 21409
rect 4433 21400 4445 21403
rect 2133 21363 2191 21369
rect 2792 21372 4445 21400
rect 1394 21292 1400 21344
rect 1452 21332 1458 21344
rect 1765 21335 1823 21341
rect 1765 21332 1777 21335
rect 1452 21304 1777 21332
rect 1452 21292 1458 21304
rect 1765 21301 1777 21304
rect 1811 21301 1823 21335
rect 2222 21332 2228 21344
rect 2183 21304 2228 21332
rect 1765 21295 1823 21301
rect 2222 21292 2228 21304
rect 2280 21292 2286 21344
rect 2792 21341 2820 21372
rect 4433 21369 4445 21372
rect 4479 21369 4491 21403
rect 4540 21400 4568 21440
rect 5445 21437 5457 21471
rect 5491 21468 5503 21471
rect 5905 21471 5963 21477
rect 5905 21468 5917 21471
rect 5491 21440 5917 21468
rect 5491 21437 5503 21440
rect 5445 21431 5503 21437
rect 5905 21437 5917 21440
rect 5951 21437 5963 21471
rect 6086 21468 6092 21480
rect 6047 21440 6092 21468
rect 5905 21431 5963 21437
rect 6086 21428 6092 21440
rect 6144 21428 6150 21480
rect 6270 21428 6276 21480
rect 6328 21468 6334 21480
rect 8386 21468 8392 21480
rect 6328 21440 8110 21468
rect 8347 21440 8392 21468
rect 6328 21428 6334 21440
rect 8082 21400 8110 21440
rect 8386 21428 8392 21440
rect 8444 21428 8450 21480
rect 8938 21468 8944 21480
rect 8899 21440 8944 21468
rect 8938 21428 8944 21440
rect 8996 21428 9002 21480
rect 9030 21428 9036 21480
rect 9088 21468 9094 21480
rect 14642 21468 14648 21480
rect 9088 21440 14648 21468
rect 9088 21428 9094 21440
rect 14642 21428 14648 21440
rect 14700 21428 14706 21480
rect 14844 21477 14872 21508
rect 14829 21471 14887 21477
rect 14829 21437 14841 21471
rect 14875 21437 14887 21471
rect 14829 21431 14887 21437
rect 15102 21428 15108 21480
rect 15160 21468 15166 21480
rect 15933 21471 15991 21477
rect 15933 21468 15945 21471
rect 15160 21440 15945 21468
rect 15160 21428 15166 21440
rect 15933 21437 15945 21440
rect 15979 21437 15991 21471
rect 16040 21468 16068 21508
rect 16117 21505 16129 21539
rect 16163 21536 16175 21539
rect 16206 21536 16212 21548
rect 16163 21508 16212 21536
rect 16163 21505 16175 21508
rect 16117 21499 16175 21505
rect 16206 21496 16212 21508
rect 16264 21496 16270 21548
rect 16758 21468 16764 21480
rect 16040 21440 16764 21468
rect 15933 21431 15991 21437
rect 16758 21428 16764 21440
rect 16816 21428 16822 21480
rect 16850 21428 16856 21480
rect 16908 21468 16914 21480
rect 16945 21471 17003 21477
rect 16945 21468 16957 21471
rect 16908 21440 16957 21468
rect 16908 21428 16914 21440
rect 16945 21437 16957 21440
rect 16991 21437 17003 21471
rect 16945 21431 17003 21437
rect 8297 21403 8355 21409
rect 8297 21400 8309 21403
rect 4540 21372 5948 21400
rect 8082 21372 8309 21400
rect 4433 21363 4491 21369
rect 2777 21335 2835 21341
rect 2777 21301 2789 21335
rect 2823 21301 2835 21335
rect 3142 21332 3148 21344
rect 3103 21304 3148 21332
rect 2777 21295 2835 21301
rect 3142 21292 3148 21304
rect 3200 21292 3206 21344
rect 3234 21292 3240 21344
rect 3292 21332 3298 21344
rect 4065 21335 4123 21341
rect 3292 21304 3337 21332
rect 3292 21292 3298 21304
rect 4065 21301 4077 21335
rect 4111 21332 4123 21335
rect 4338 21332 4344 21344
rect 4111 21304 4344 21332
rect 4111 21301 4123 21304
rect 4065 21295 4123 21301
rect 4338 21292 4344 21304
rect 4396 21292 4402 21344
rect 4522 21332 4528 21344
rect 4483 21304 4528 21332
rect 4522 21292 4528 21304
rect 4580 21292 4586 21344
rect 5077 21335 5135 21341
rect 5077 21301 5089 21335
rect 5123 21332 5135 21335
rect 5534 21332 5540 21344
rect 5123 21304 5540 21332
rect 5123 21301 5135 21304
rect 5077 21295 5135 21301
rect 5534 21292 5540 21304
rect 5592 21292 5598 21344
rect 5920 21332 5948 21372
rect 8297 21369 8309 21372
rect 8343 21369 8355 21403
rect 8297 21363 8355 21369
rect 10413 21403 10471 21409
rect 10413 21369 10425 21403
rect 10459 21400 10471 21403
rect 12526 21400 12532 21412
rect 10459 21372 12532 21400
rect 10459 21369 10471 21372
rect 10413 21363 10471 21369
rect 12526 21360 12532 21372
rect 12584 21360 12590 21412
rect 14093 21403 14151 21409
rect 14093 21400 14105 21403
rect 12636 21372 14105 21400
rect 6273 21335 6331 21341
rect 6273 21332 6285 21335
rect 5920 21304 6285 21332
rect 6273 21301 6285 21304
rect 6319 21301 6331 21335
rect 6273 21295 6331 21301
rect 6914 21292 6920 21344
rect 6972 21332 6978 21344
rect 7285 21335 7343 21341
rect 7285 21332 7297 21335
rect 6972 21304 7297 21332
rect 6972 21292 6978 21304
rect 7285 21301 7297 21304
rect 7331 21301 7343 21335
rect 7285 21295 7343 21301
rect 7374 21292 7380 21344
rect 7432 21332 7438 21344
rect 7929 21335 7987 21341
rect 7432 21304 7477 21332
rect 7432 21292 7438 21304
rect 7929 21301 7941 21335
rect 7975 21332 7987 21335
rect 9766 21332 9772 21344
rect 7975 21304 9772 21332
rect 7975 21301 7987 21304
rect 7929 21295 7987 21301
rect 9766 21292 9772 21304
rect 9824 21292 9830 21344
rect 11057 21335 11115 21341
rect 11057 21301 11069 21335
rect 11103 21332 11115 21335
rect 11238 21332 11244 21344
rect 11103 21304 11244 21332
rect 11103 21301 11115 21304
rect 11057 21295 11115 21301
rect 11238 21292 11244 21304
rect 11296 21292 11302 21344
rect 11422 21332 11428 21344
rect 11383 21304 11428 21332
rect 11422 21292 11428 21304
rect 11480 21292 11486 21344
rect 11517 21335 11575 21341
rect 11517 21301 11529 21335
rect 11563 21332 11575 21335
rect 11606 21332 11612 21344
rect 11563 21304 11612 21332
rect 11563 21301 11575 21304
rect 11517 21295 11575 21301
rect 11606 21292 11612 21304
rect 11664 21292 11670 21344
rect 12066 21332 12072 21344
rect 12027 21304 12072 21332
rect 12066 21292 12072 21304
rect 12124 21292 12130 21344
rect 12636 21341 12664 21372
rect 14093 21369 14105 21372
rect 14139 21369 14151 21403
rect 14093 21363 14151 21369
rect 14458 21360 14464 21412
rect 14516 21400 14522 21412
rect 15841 21403 15899 21409
rect 15841 21400 15853 21403
rect 14516 21372 15853 21400
rect 14516 21360 14522 21372
rect 15841 21369 15853 21372
rect 15887 21369 15899 21403
rect 17052 21400 17080 21576
rect 17144 21576 20536 21604
rect 17144 21545 17172 21576
rect 20530 21564 20536 21576
rect 20588 21564 20594 21616
rect 20622 21564 20628 21616
rect 20680 21604 20686 21616
rect 21100 21604 21128 21644
rect 24026 21632 24032 21644
rect 24084 21632 24090 21684
rect 20680 21576 21128 21604
rect 20680 21564 20686 21576
rect 21634 21564 21640 21616
rect 21692 21604 21698 21616
rect 22189 21607 22247 21613
rect 22189 21604 22201 21607
rect 21692 21576 22201 21604
rect 21692 21564 21698 21576
rect 22189 21573 22201 21576
rect 22235 21573 22247 21607
rect 22189 21567 22247 21573
rect 17129 21539 17187 21545
rect 17129 21505 17141 21539
rect 17175 21505 17187 21539
rect 19334 21536 19340 21548
rect 17129 21499 17187 21505
rect 17236 21508 19340 21536
rect 17236 21400 17264 21508
rect 19334 21496 19340 21508
rect 19392 21496 19398 21548
rect 19886 21496 19892 21548
rect 19944 21536 19950 21548
rect 20165 21539 20223 21545
rect 20165 21536 20177 21539
rect 19944 21508 20177 21536
rect 19944 21496 19950 21508
rect 20165 21505 20177 21508
rect 20211 21505 20223 21539
rect 20165 21499 20223 21505
rect 21821 21539 21879 21545
rect 21821 21505 21833 21539
rect 21867 21536 21879 21539
rect 22002 21536 22008 21548
rect 21867 21508 22008 21536
rect 21867 21505 21879 21508
rect 21821 21499 21879 21505
rect 22002 21496 22008 21508
rect 22060 21496 22066 21548
rect 22833 21539 22891 21545
rect 22833 21505 22845 21539
rect 22879 21536 22891 21539
rect 22922 21536 22928 21548
rect 22879 21508 22928 21536
rect 22879 21505 22891 21508
rect 22833 21499 22891 21505
rect 22922 21496 22928 21508
rect 22980 21496 22986 21548
rect 17402 21428 17408 21480
rect 17460 21468 17466 21480
rect 17497 21471 17555 21477
rect 17497 21468 17509 21471
rect 17460 21440 17509 21468
rect 17460 21428 17466 21440
rect 17497 21437 17509 21440
rect 17543 21437 17555 21471
rect 17497 21431 17555 21437
rect 18230 21428 18236 21480
rect 18288 21468 18294 21480
rect 18325 21471 18383 21477
rect 18325 21468 18337 21471
rect 18288 21440 18337 21468
rect 18288 21428 18294 21440
rect 18325 21437 18337 21440
rect 18371 21437 18383 21471
rect 20346 21468 20352 21480
rect 18325 21431 18383 21437
rect 18432 21440 20352 21468
rect 17052 21372 17264 21400
rect 17313 21403 17371 21409
rect 15841 21363 15899 21369
rect 17313 21369 17325 21403
rect 17359 21400 17371 21403
rect 18432 21400 18460 21440
rect 20346 21428 20352 21440
rect 20404 21428 20410 21480
rect 21266 21428 21272 21480
rect 21324 21468 21330 21480
rect 22649 21471 22707 21477
rect 22649 21468 22661 21471
rect 21324 21440 22661 21468
rect 21324 21428 21330 21440
rect 22649 21437 22661 21440
rect 22695 21437 22707 21471
rect 22649 21431 22707 21437
rect 19150 21400 19156 21412
rect 17359 21372 18460 21400
rect 19111 21372 19156 21400
rect 17359 21369 17371 21372
rect 17313 21363 17371 21369
rect 19150 21360 19156 21372
rect 19208 21360 19214 21412
rect 19981 21403 20039 21409
rect 19981 21400 19993 21403
rect 19260 21372 19993 21400
rect 12621 21335 12679 21341
rect 12621 21301 12633 21335
rect 12667 21301 12679 21335
rect 12986 21332 12992 21344
rect 12947 21304 12992 21332
rect 12621 21295 12679 21301
rect 12986 21292 12992 21304
rect 13044 21292 13050 21344
rect 13078 21292 13084 21344
rect 13136 21332 13142 21344
rect 13633 21335 13691 21341
rect 13136 21304 13181 21332
rect 13136 21292 13142 21304
rect 13633 21301 13645 21335
rect 13679 21332 13691 21335
rect 13814 21332 13820 21344
rect 13679 21304 13820 21332
rect 13679 21301 13691 21304
rect 13633 21295 13691 21301
rect 13814 21292 13820 21304
rect 13872 21292 13878 21344
rect 13998 21332 14004 21344
rect 13959 21304 14004 21332
rect 13998 21292 14004 21304
rect 14056 21292 14062 21344
rect 15470 21332 15476 21344
rect 15431 21304 15476 21332
rect 15470 21292 15476 21304
rect 15528 21292 15534 21344
rect 16482 21332 16488 21344
rect 16443 21304 16488 21332
rect 16482 21292 16488 21304
rect 16540 21292 16546 21344
rect 16853 21335 16911 21341
rect 16853 21301 16865 21335
rect 16899 21332 16911 21335
rect 17770 21332 17776 21344
rect 16899 21304 17776 21332
rect 16899 21301 16911 21304
rect 16853 21295 16911 21301
rect 17770 21292 17776 21304
rect 17828 21292 17834 21344
rect 18046 21292 18052 21344
rect 18104 21332 18110 21344
rect 19260 21332 19288 21372
rect 19981 21369 19993 21372
rect 20027 21369 20039 21403
rect 19981 21363 20039 21369
rect 20901 21403 20959 21409
rect 20901 21369 20913 21403
rect 20947 21400 20959 21403
rect 21545 21403 21603 21409
rect 21545 21400 21557 21403
rect 20947 21372 21557 21400
rect 20947 21369 20959 21372
rect 20901 21363 20959 21369
rect 21545 21369 21557 21372
rect 21591 21369 21603 21403
rect 21545 21363 21603 21369
rect 18104 21304 19288 21332
rect 18104 21292 18110 21304
rect 19426 21292 19432 21344
rect 19484 21332 19490 21344
rect 19613 21335 19671 21341
rect 19613 21332 19625 21335
rect 19484 21304 19625 21332
rect 19484 21292 19490 21304
rect 19613 21301 19625 21304
rect 19659 21332 19671 21335
rect 19794 21332 19800 21344
rect 19659 21304 19800 21332
rect 19659 21301 19671 21304
rect 19613 21295 19671 21301
rect 19794 21292 19800 21304
rect 19852 21292 19858 21344
rect 20070 21332 20076 21344
rect 20031 21304 20076 21332
rect 20070 21292 20076 21304
rect 20128 21292 20134 21344
rect 20622 21332 20628 21344
rect 20583 21304 20628 21332
rect 20622 21292 20628 21304
rect 20680 21292 20686 21344
rect 21174 21332 21180 21344
rect 21135 21304 21180 21332
rect 21174 21292 21180 21304
rect 21232 21292 21238 21344
rect 21637 21335 21695 21341
rect 21637 21301 21649 21335
rect 21683 21332 21695 21335
rect 21726 21332 21732 21344
rect 21683 21304 21732 21332
rect 21683 21301 21695 21304
rect 21637 21295 21695 21301
rect 21726 21292 21732 21304
rect 21784 21292 21790 21344
rect 22557 21335 22615 21341
rect 22557 21301 22569 21335
rect 22603 21332 22615 21335
rect 23198 21332 23204 21344
rect 22603 21304 23204 21332
rect 22603 21301 22615 21304
rect 22557 21295 22615 21301
rect 23198 21292 23204 21304
rect 23256 21292 23262 21344
rect 1104 21242 23276 21264
rect 1104 21190 8379 21242
rect 8431 21190 8443 21242
rect 8495 21190 8507 21242
rect 8559 21190 8571 21242
rect 8623 21190 15776 21242
rect 15828 21190 15840 21242
rect 15892 21190 15904 21242
rect 15956 21190 15968 21242
rect 16020 21190 23276 21242
rect 1104 21168 23276 21190
rect 290 21088 296 21140
rect 348 21128 354 21140
rect 1765 21131 1823 21137
rect 1765 21128 1777 21131
rect 348 21100 1777 21128
rect 348 21088 354 21100
rect 1765 21097 1777 21100
rect 1811 21097 1823 21131
rect 1765 21091 1823 21097
rect 3142 21088 3148 21140
rect 3200 21128 3206 21140
rect 3510 21128 3516 21140
rect 3200 21100 3516 21128
rect 3200 21088 3206 21100
rect 3510 21088 3516 21100
rect 3568 21088 3574 21140
rect 5445 21131 5503 21137
rect 5445 21097 5457 21131
rect 5491 21097 5503 21131
rect 5445 21091 5503 21097
rect 5166 21020 5172 21072
rect 5224 21060 5230 21072
rect 5460 21060 5488 21091
rect 5534 21088 5540 21140
rect 5592 21128 5598 21140
rect 6089 21131 6147 21137
rect 6089 21128 6101 21131
rect 5592 21100 6101 21128
rect 5592 21088 5598 21100
rect 6089 21097 6101 21100
rect 6135 21128 6147 21131
rect 7834 21128 7840 21140
rect 6135 21100 7840 21128
rect 6135 21097 6147 21100
rect 6089 21091 6147 21097
rect 7834 21088 7840 21100
rect 7892 21088 7898 21140
rect 8113 21131 8171 21137
rect 8113 21097 8125 21131
rect 8159 21097 8171 21131
rect 8113 21091 8171 21097
rect 8941 21131 8999 21137
rect 8941 21097 8953 21131
rect 8987 21128 8999 21131
rect 12066 21128 12072 21140
rect 8987 21100 12072 21128
rect 8987 21097 8999 21100
rect 8941 21091 8999 21097
rect 6730 21060 6736 21072
rect 5224 21032 6736 21060
rect 5224 21020 5230 21032
rect 6730 21020 6736 21032
rect 6788 21020 6794 21072
rect 7190 21020 7196 21072
rect 7248 21060 7254 21072
rect 7374 21060 7380 21072
rect 7248 21032 7380 21060
rect 7248 21020 7254 21032
rect 7374 21020 7380 21032
rect 7432 21020 7438 21072
rect 7466 21020 7472 21072
rect 7524 21060 7530 21072
rect 8128 21060 8156 21091
rect 12066 21088 12072 21100
rect 12124 21088 12130 21140
rect 13354 21088 13360 21140
rect 13412 21128 13418 21140
rect 14458 21128 14464 21140
rect 13412 21100 14320 21128
rect 14419 21100 14464 21128
rect 13412 21088 13418 21100
rect 7524 21032 11468 21060
rect 7524 21020 7530 21032
rect 1581 20995 1639 21001
rect 1581 20961 1593 20995
rect 1627 20992 1639 20995
rect 2038 20992 2044 21004
rect 1627 20964 2044 20992
rect 1627 20961 1639 20964
rect 1581 20955 1639 20961
rect 2038 20952 2044 20964
rect 2096 20952 2102 21004
rect 2400 20995 2458 21001
rect 2400 20961 2412 20995
rect 2446 20992 2458 20995
rect 3234 20992 3240 21004
rect 2446 20964 3240 20992
rect 2446 20961 2458 20964
rect 2400 20955 2458 20961
rect 3234 20952 3240 20964
rect 3292 20952 3298 21004
rect 4338 21001 4344 21004
rect 4332 20955 4344 21001
rect 4396 20992 4402 21004
rect 6181 20995 6239 21001
rect 4396 20964 4432 20992
rect 4338 20952 4344 20955
rect 4396 20952 4402 20964
rect 6181 20961 6193 20995
rect 6227 20992 6239 20995
rect 6546 20992 6552 21004
rect 6227 20964 6552 20992
rect 6227 20961 6239 20964
rect 6181 20955 6239 20961
rect 6546 20952 6552 20964
rect 6604 20952 6610 21004
rect 7000 20995 7058 21001
rect 7000 20961 7012 20995
rect 7046 20992 7058 20995
rect 8018 20992 8024 21004
rect 7046 20964 8024 20992
rect 7046 20961 7058 20964
rect 7000 20955 7058 20961
rect 8018 20952 8024 20964
rect 8076 20952 8082 21004
rect 9944 20995 10002 21001
rect 9944 20992 9956 20995
rect 9232 20964 9956 20992
rect 2133 20927 2191 20933
rect 2133 20893 2145 20927
rect 2179 20893 2191 20927
rect 2133 20887 2191 20893
rect 2148 20788 2176 20887
rect 3326 20884 3332 20936
rect 3384 20924 3390 20936
rect 4065 20927 4123 20933
rect 4065 20924 4077 20927
rect 3384 20896 4077 20924
rect 3384 20884 3390 20896
rect 4065 20893 4077 20896
rect 4111 20893 4123 20927
rect 4065 20887 4123 20893
rect 5074 20884 5080 20936
rect 5132 20924 5138 20936
rect 6273 20927 6331 20933
rect 6273 20924 6285 20927
rect 5132 20896 6285 20924
rect 5132 20884 5138 20896
rect 6273 20893 6285 20896
rect 6319 20893 6331 20927
rect 6273 20887 6331 20893
rect 6454 20884 6460 20936
rect 6512 20924 6518 20936
rect 6733 20927 6791 20933
rect 6733 20924 6745 20927
rect 6512 20896 6745 20924
rect 6512 20884 6518 20896
rect 6733 20893 6745 20896
rect 6779 20893 6791 20927
rect 6733 20887 6791 20893
rect 7834 20884 7840 20936
rect 7892 20924 7898 20936
rect 9030 20924 9036 20936
rect 7892 20896 8800 20924
rect 8991 20896 9036 20924
rect 7892 20884 7898 20896
rect 5258 20816 5264 20868
rect 5316 20856 5322 20868
rect 5442 20856 5448 20868
rect 5316 20828 5448 20856
rect 5316 20816 5322 20828
rect 5442 20816 5448 20828
rect 5500 20816 5506 20868
rect 8662 20856 8668 20868
rect 7668 20828 8668 20856
rect 2774 20788 2780 20800
rect 2148 20760 2780 20788
rect 2774 20748 2780 20760
rect 2832 20748 2838 20800
rect 4430 20748 4436 20800
rect 4488 20788 4494 20800
rect 5721 20791 5779 20797
rect 5721 20788 5733 20791
rect 4488 20760 5733 20788
rect 4488 20748 4494 20760
rect 5721 20757 5733 20760
rect 5767 20757 5779 20791
rect 5721 20751 5779 20757
rect 5810 20748 5816 20800
rect 5868 20788 5874 20800
rect 7668 20788 7696 20828
rect 8662 20816 8668 20828
rect 8720 20816 8726 20868
rect 8772 20856 8800 20896
rect 9030 20884 9036 20896
rect 9088 20884 9094 20936
rect 9232 20933 9260 20964
rect 9944 20961 9956 20964
rect 9990 20992 10002 20995
rect 10226 20992 10232 21004
rect 9990 20964 10232 20992
rect 9990 20961 10002 20964
rect 9944 20955 10002 20961
rect 10226 20952 10232 20964
rect 10284 20952 10290 21004
rect 11440 20992 11468 21032
rect 11514 21020 11520 21072
rect 11572 21069 11578 21072
rect 11572 21063 11636 21069
rect 11572 21029 11590 21063
rect 11624 21029 11636 21063
rect 11572 21023 11636 21029
rect 11572 21020 11578 21023
rect 12526 21020 12532 21072
rect 12584 21060 12590 21072
rect 12584 21032 14228 21060
rect 12584 21020 12590 21032
rect 11974 20992 11980 21004
rect 11440 20964 11980 20992
rect 11974 20952 11980 20964
rect 12032 20952 12038 21004
rect 13348 20995 13406 21001
rect 13348 20961 13360 20995
rect 13394 20992 13406 20995
rect 14090 20992 14096 21004
rect 13394 20964 14096 20992
rect 13394 20961 13406 20964
rect 13348 20955 13406 20961
rect 14090 20952 14096 20964
rect 14148 20952 14154 21004
rect 9217 20927 9275 20933
rect 9217 20893 9229 20927
rect 9263 20893 9275 20927
rect 9217 20887 9275 20893
rect 9677 20927 9735 20933
rect 9677 20893 9689 20927
rect 9723 20893 9735 20927
rect 11333 20927 11391 20933
rect 11333 20924 11345 20927
rect 9677 20887 9735 20893
rect 10704 20896 11345 20924
rect 9582 20856 9588 20868
rect 8772 20828 9588 20856
rect 9582 20816 9588 20828
rect 9640 20816 9646 20868
rect 8570 20788 8576 20800
rect 5868 20760 7696 20788
rect 8531 20760 8576 20788
rect 5868 20748 5874 20760
rect 8570 20748 8576 20760
rect 8628 20748 8634 20800
rect 8846 20748 8852 20800
rect 8904 20788 8910 20800
rect 9692 20788 9720 20887
rect 9950 20788 9956 20800
rect 8904 20760 9956 20788
rect 8904 20748 8910 20760
rect 9950 20748 9956 20760
rect 10008 20788 10014 20800
rect 10704 20788 10732 20896
rect 11333 20893 11345 20896
rect 11379 20893 11391 20927
rect 11333 20887 11391 20893
rect 13081 20927 13139 20933
rect 13081 20893 13093 20927
rect 13127 20893 13139 20927
rect 13081 20887 13139 20893
rect 12434 20816 12440 20868
rect 12492 20856 12498 20868
rect 12894 20856 12900 20868
rect 12492 20828 12900 20856
rect 12492 20816 12498 20828
rect 12894 20816 12900 20828
rect 12952 20856 12958 20868
rect 13096 20856 13124 20887
rect 12952 20828 13124 20856
rect 14200 20856 14228 21032
rect 14292 20992 14320 21100
rect 14458 21088 14464 21100
rect 14516 21088 14522 21140
rect 14642 21088 14648 21140
rect 14700 21128 14706 21140
rect 15194 21128 15200 21140
rect 14700 21100 15200 21128
rect 14700 21088 14706 21100
rect 15194 21088 15200 21100
rect 15252 21088 15258 21140
rect 15470 21088 15476 21140
rect 15528 21128 15534 21140
rect 17313 21131 17371 21137
rect 17313 21128 17325 21131
rect 15528 21100 17325 21128
rect 15528 21088 15534 21100
rect 17313 21097 17325 21100
rect 17359 21097 17371 21131
rect 17313 21091 17371 21097
rect 19797 21131 19855 21137
rect 19797 21097 19809 21131
rect 19843 21128 19855 21131
rect 20070 21128 20076 21140
rect 19843 21100 20076 21128
rect 19843 21097 19855 21100
rect 19797 21091 19855 21097
rect 20070 21088 20076 21100
rect 20128 21088 20134 21140
rect 20622 21088 20628 21140
rect 20680 21128 20686 21140
rect 21269 21131 21327 21137
rect 21269 21128 21281 21131
rect 20680 21100 21281 21128
rect 20680 21088 20686 21100
rect 21269 21097 21281 21100
rect 21315 21097 21327 21131
rect 21269 21091 21327 21097
rect 15562 21069 15568 21072
rect 14553 21063 14611 21069
rect 14553 21029 14565 21063
rect 14599 21060 14611 21063
rect 14737 21063 14795 21069
rect 14737 21060 14749 21063
rect 14599 21032 14749 21060
rect 14599 21029 14611 21032
rect 14553 21023 14611 21029
rect 14737 21029 14749 21032
rect 14783 21029 14795 21063
rect 14737 21023 14795 21029
rect 15556 21023 15568 21069
rect 15620 21060 15626 21072
rect 15620 21032 15656 21060
rect 15562 21020 15568 21023
rect 15620 21020 15626 21032
rect 18782 21020 18788 21072
rect 18840 21060 18846 21072
rect 20165 21063 20223 21069
rect 18840 21032 20015 21060
rect 18840 21020 18846 21032
rect 18408 20995 18466 21001
rect 14292 20964 16988 20992
rect 14366 20884 14372 20936
rect 14424 20924 14430 20936
rect 15289 20927 15347 20933
rect 15289 20924 15301 20927
rect 14424 20896 15301 20924
rect 14424 20884 14430 20896
rect 15289 20893 15301 20896
rect 15335 20893 15347 20927
rect 15289 20887 15347 20893
rect 16960 20865 16988 20964
rect 18408 20961 18420 20995
rect 18454 20992 18466 20995
rect 19886 20992 19892 21004
rect 18454 20964 19892 20992
rect 18454 20961 18466 20964
rect 18408 20955 18466 20961
rect 19886 20952 19892 20964
rect 19944 20952 19950 21004
rect 19987 20992 20015 21032
rect 20165 21029 20177 21063
rect 20211 21060 20223 21063
rect 20254 21060 20260 21072
rect 20211 21032 20260 21060
rect 20211 21029 20223 21032
rect 20165 21023 20223 21029
rect 20254 21020 20260 21032
rect 20312 21020 20318 21072
rect 20346 21020 20352 21072
rect 20404 21060 20410 21072
rect 22281 21063 22339 21069
rect 22281 21060 22293 21063
rect 20404 21032 22293 21060
rect 20404 21020 20410 21032
rect 22281 21029 22293 21032
rect 22327 21029 22339 21063
rect 22281 21023 22339 21029
rect 22189 20995 22247 21001
rect 19987 20964 20300 20992
rect 17402 20924 17408 20936
rect 17363 20896 17408 20924
rect 17402 20884 17408 20896
rect 17460 20884 17466 20936
rect 17586 20924 17592 20936
rect 17547 20896 17592 20924
rect 17586 20884 17592 20896
rect 17644 20884 17650 20936
rect 17954 20884 17960 20936
rect 18012 20924 18018 20936
rect 20272 20933 20300 20964
rect 22189 20961 22201 20995
rect 22235 20992 22247 20995
rect 22462 20992 22468 21004
rect 22235 20964 22468 20992
rect 22235 20961 22247 20964
rect 22189 20955 22247 20961
rect 22462 20952 22468 20964
rect 22520 20952 22526 21004
rect 22646 20992 22652 21004
rect 22607 20964 22652 20992
rect 22646 20952 22652 20964
rect 22704 20952 22710 21004
rect 18141 20927 18199 20933
rect 18141 20924 18153 20927
rect 18012 20896 18153 20924
rect 18012 20884 18018 20896
rect 18141 20893 18153 20896
rect 18187 20893 18199 20927
rect 18141 20887 18199 20893
rect 20257 20927 20315 20933
rect 20257 20893 20269 20927
rect 20303 20893 20315 20927
rect 20257 20887 20315 20893
rect 20349 20927 20407 20933
rect 20349 20893 20361 20927
rect 20395 20893 20407 20927
rect 21358 20924 21364 20936
rect 21319 20896 21364 20924
rect 20349 20887 20407 20893
rect 14553 20859 14611 20865
rect 14553 20856 14565 20859
rect 14200 20828 14565 20856
rect 12952 20816 12958 20828
rect 11054 20788 11060 20800
rect 10008 20760 10732 20788
rect 11015 20760 11060 20788
rect 10008 20748 10014 20760
rect 11054 20748 11060 20760
rect 11112 20748 11118 20800
rect 11238 20748 11244 20800
rect 11296 20788 11302 20800
rect 11974 20788 11980 20800
rect 11296 20760 11980 20788
rect 11296 20748 11302 20760
rect 11974 20748 11980 20760
rect 12032 20748 12038 20800
rect 12526 20748 12532 20800
rect 12584 20788 12590 20800
rect 12713 20791 12771 20797
rect 12713 20788 12725 20791
rect 12584 20760 12725 20788
rect 12584 20748 12590 20760
rect 12713 20757 12725 20760
rect 12759 20757 12771 20791
rect 13096 20788 13124 20828
rect 14553 20825 14565 20828
rect 14599 20825 14611 20859
rect 14553 20819 14611 20825
rect 16945 20859 17003 20865
rect 16945 20825 16957 20859
rect 16991 20825 17003 20859
rect 16945 20819 17003 20825
rect 19150 20816 19156 20868
rect 19208 20856 19214 20868
rect 20364 20856 20392 20887
rect 21358 20884 21364 20896
rect 21416 20884 21422 20936
rect 21453 20927 21511 20933
rect 21453 20893 21465 20927
rect 21499 20893 21511 20927
rect 21453 20887 21511 20893
rect 22373 20927 22431 20933
rect 22373 20893 22385 20927
rect 22419 20924 22431 20927
rect 23014 20924 23020 20936
rect 22419 20896 23020 20924
rect 22419 20893 22431 20896
rect 22373 20887 22431 20893
rect 19208 20828 20392 20856
rect 19208 20816 19214 20828
rect 21082 20816 21088 20868
rect 21140 20856 21146 20868
rect 21468 20856 21496 20887
rect 23014 20884 23020 20896
rect 23072 20884 23078 20936
rect 21140 20828 21496 20856
rect 21140 20816 21146 20828
rect 14366 20788 14372 20800
rect 13096 20760 14372 20788
rect 12713 20751 12771 20757
rect 14366 20748 14372 20760
rect 14424 20748 14430 20800
rect 15470 20748 15476 20800
rect 15528 20788 15534 20800
rect 16482 20788 16488 20800
rect 15528 20760 16488 20788
rect 15528 20748 15534 20760
rect 16482 20748 16488 20760
rect 16540 20748 16546 20800
rect 16574 20748 16580 20800
rect 16632 20788 16638 20800
rect 16669 20791 16727 20797
rect 16669 20788 16681 20791
rect 16632 20760 16681 20788
rect 16632 20748 16638 20760
rect 16669 20757 16681 20760
rect 16715 20757 16727 20791
rect 16669 20751 16727 20757
rect 19521 20791 19579 20797
rect 19521 20757 19533 20791
rect 19567 20788 19579 20791
rect 19794 20788 19800 20800
rect 19567 20760 19800 20788
rect 19567 20757 19579 20760
rect 19521 20751 19579 20757
rect 19794 20748 19800 20760
rect 19852 20748 19858 20800
rect 20898 20788 20904 20800
rect 20859 20760 20904 20788
rect 20898 20748 20904 20760
rect 20956 20748 20962 20800
rect 21174 20748 21180 20800
rect 21232 20788 21238 20800
rect 21821 20791 21879 20797
rect 21821 20788 21833 20791
rect 21232 20760 21833 20788
rect 21232 20748 21238 20760
rect 21821 20757 21833 20760
rect 21867 20757 21879 20791
rect 22830 20788 22836 20800
rect 22791 20760 22836 20788
rect 21821 20751 21879 20757
rect 22830 20748 22836 20760
rect 22888 20748 22894 20800
rect 1104 20698 23276 20720
rect 1104 20646 4680 20698
rect 4732 20646 4744 20698
rect 4796 20646 4808 20698
rect 4860 20646 4872 20698
rect 4924 20646 12078 20698
rect 12130 20646 12142 20698
rect 12194 20646 12206 20698
rect 12258 20646 12270 20698
rect 12322 20646 19475 20698
rect 19527 20646 19539 20698
rect 19591 20646 19603 20698
rect 19655 20646 19667 20698
rect 19719 20646 23276 20698
rect 1104 20624 23276 20646
rect 842 20544 848 20596
rect 900 20584 906 20596
rect 3050 20584 3056 20596
rect 900 20556 3056 20584
rect 900 20544 906 20556
rect 3050 20544 3056 20556
rect 3108 20544 3114 20596
rect 3145 20587 3203 20593
rect 3145 20553 3157 20587
rect 3191 20584 3203 20587
rect 3234 20584 3240 20596
rect 3191 20556 3240 20584
rect 3191 20553 3203 20556
rect 3145 20547 3203 20553
rect 3234 20544 3240 20556
rect 3292 20544 3298 20596
rect 4338 20544 4344 20596
rect 4396 20584 4402 20596
rect 4801 20587 4859 20593
rect 4801 20584 4813 20587
rect 4396 20556 4813 20584
rect 4396 20544 4402 20556
rect 4801 20553 4813 20556
rect 4847 20584 4859 20587
rect 4985 20587 5043 20593
rect 4985 20584 4997 20587
rect 4847 20556 4997 20584
rect 4847 20553 4859 20556
rect 4801 20547 4859 20553
rect 4985 20553 4997 20556
rect 5031 20553 5043 20587
rect 4985 20547 5043 20553
rect 5258 20544 5264 20596
rect 5316 20584 5322 20596
rect 5316 20556 8064 20584
rect 5316 20544 5322 20556
rect 5994 20516 6000 20528
rect 4724 20488 6000 20516
rect 1765 20383 1823 20389
rect 1765 20349 1777 20383
rect 1811 20380 1823 20383
rect 2774 20380 2780 20392
rect 1811 20352 2780 20380
rect 1811 20349 1823 20352
rect 1765 20343 1823 20349
rect 2774 20340 2780 20352
rect 2832 20380 2838 20392
rect 3326 20380 3332 20392
rect 2832 20352 3332 20380
rect 2832 20340 2838 20352
rect 3326 20340 3332 20352
rect 3384 20380 3390 20392
rect 3421 20383 3479 20389
rect 3421 20380 3433 20383
rect 3384 20352 3433 20380
rect 3384 20340 3390 20352
rect 3421 20349 3433 20352
rect 3467 20349 3479 20383
rect 3421 20343 3479 20349
rect 3510 20340 3516 20392
rect 3568 20380 3574 20392
rect 3677 20383 3735 20389
rect 3677 20380 3689 20383
rect 3568 20352 3689 20380
rect 3568 20340 3574 20352
rect 3677 20349 3689 20352
rect 3723 20349 3735 20383
rect 3677 20343 3735 20349
rect 3970 20340 3976 20392
rect 4028 20380 4034 20392
rect 4724 20380 4752 20488
rect 5994 20476 6000 20488
rect 6052 20476 6058 20528
rect 5718 20448 5724 20460
rect 5679 20420 5724 20448
rect 5718 20408 5724 20420
rect 5776 20408 5782 20460
rect 8036 20448 8064 20556
rect 8110 20544 8116 20596
rect 8168 20584 8174 20596
rect 8205 20587 8263 20593
rect 8205 20584 8217 20587
rect 8168 20556 8217 20584
rect 8168 20544 8174 20556
rect 8205 20553 8217 20556
rect 8251 20553 8263 20587
rect 8205 20547 8263 20553
rect 8570 20544 8576 20596
rect 8628 20584 8634 20596
rect 10226 20584 10232 20596
rect 8628 20556 10088 20584
rect 10187 20556 10232 20584
rect 8628 20544 8634 20556
rect 10060 20516 10088 20556
rect 10226 20544 10232 20556
rect 10284 20544 10290 20596
rect 10336 20556 11468 20584
rect 10336 20516 10364 20556
rect 10060 20488 10364 20516
rect 11440 20516 11468 20556
rect 11514 20544 11520 20596
rect 11572 20584 11578 20596
rect 11885 20587 11943 20593
rect 11885 20584 11897 20587
rect 11572 20556 11897 20584
rect 11572 20544 11578 20556
rect 11885 20553 11897 20556
rect 11931 20553 11943 20587
rect 14090 20584 14096 20596
rect 11885 20547 11943 20553
rect 11992 20556 13952 20584
rect 14003 20556 14096 20584
rect 11992 20516 12020 20556
rect 11440 20488 12020 20516
rect 12434 20476 12440 20528
rect 12492 20516 12498 20528
rect 13924 20516 13952 20556
rect 14090 20544 14096 20556
rect 14148 20584 14154 20596
rect 15102 20584 15108 20596
rect 14148 20556 15108 20584
rect 14148 20544 14154 20556
rect 15102 20544 15108 20556
rect 15160 20544 15166 20596
rect 19334 20584 19340 20596
rect 15948 20556 19340 20584
rect 12492 20488 12756 20516
rect 13924 20488 14136 20516
rect 12492 20476 12498 20488
rect 8036 20420 8984 20448
rect 4028 20352 4752 20380
rect 4985 20383 5043 20389
rect 4028 20340 4034 20352
rect 4985 20349 4997 20383
rect 5031 20380 5043 20383
rect 6273 20383 6331 20389
rect 6273 20380 6285 20383
rect 5031 20352 6285 20380
rect 5031 20349 5043 20352
rect 4985 20343 5043 20349
rect 6273 20349 6285 20352
rect 6319 20349 6331 20383
rect 6273 20343 6331 20349
rect 6454 20340 6460 20392
rect 6512 20380 6518 20392
rect 6825 20383 6883 20389
rect 6825 20380 6837 20383
rect 6512 20352 6837 20380
rect 6512 20340 6518 20352
rect 6825 20349 6837 20352
rect 6871 20349 6883 20383
rect 8846 20380 8852 20392
rect 8807 20352 8852 20380
rect 6825 20343 6883 20349
rect 8846 20340 8852 20352
rect 8904 20340 8910 20392
rect 8956 20380 8984 20420
rect 9950 20408 9956 20460
rect 10008 20448 10014 20460
rect 10226 20448 10232 20460
rect 10008 20420 10232 20448
rect 10008 20408 10014 20420
rect 10226 20408 10232 20420
rect 10284 20448 10290 20460
rect 12728 20457 12756 20488
rect 10505 20451 10563 20457
rect 10505 20448 10517 20451
rect 10284 20420 10517 20448
rect 10284 20408 10290 20420
rect 10505 20417 10517 20420
rect 10551 20417 10563 20451
rect 10505 20411 10563 20417
rect 12713 20451 12771 20457
rect 12713 20417 12725 20451
rect 12759 20417 12771 20451
rect 12713 20411 12771 20417
rect 10410 20380 10416 20392
rect 8956 20352 10416 20380
rect 10410 20340 10416 20352
rect 10468 20340 10474 20392
rect 12434 20380 12440 20392
rect 10612 20352 12440 20380
rect 2032 20315 2090 20321
rect 2032 20281 2044 20315
rect 2078 20312 2090 20315
rect 2958 20312 2964 20324
rect 2078 20284 2964 20312
rect 2078 20281 2090 20284
rect 2032 20275 2090 20281
rect 2958 20272 2964 20284
rect 3016 20272 3022 20324
rect 4154 20272 4160 20324
rect 4212 20312 4218 20324
rect 7098 20321 7104 20324
rect 5537 20315 5595 20321
rect 5537 20312 5549 20315
rect 4212 20284 5549 20312
rect 4212 20272 4218 20284
rect 5537 20281 5549 20284
rect 5583 20281 5595 20315
rect 5537 20275 5595 20281
rect 6089 20315 6147 20321
rect 6089 20281 6101 20315
rect 6135 20312 6147 20315
rect 7092 20312 7104 20321
rect 6135 20284 6960 20312
rect 7059 20284 7104 20312
rect 6135 20281 6147 20284
rect 6089 20275 6147 20281
rect 2130 20204 2136 20256
rect 2188 20244 2194 20256
rect 3602 20244 3608 20256
rect 2188 20216 3608 20244
rect 2188 20204 2194 20216
rect 3602 20204 3608 20216
rect 3660 20204 3666 20256
rect 4338 20204 4344 20256
rect 4396 20244 4402 20256
rect 5077 20247 5135 20253
rect 5077 20244 5089 20247
rect 4396 20216 5089 20244
rect 4396 20204 4402 20216
rect 5077 20213 5089 20216
rect 5123 20213 5135 20247
rect 5442 20244 5448 20256
rect 5403 20216 5448 20244
rect 5077 20207 5135 20213
rect 5442 20204 5448 20216
rect 5500 20204 5506 20256
rect 5626 20204 5632 20256
rect 5684 20244 5690 20256
rect 6457 20247 6515 20253
rect 6457 20244 6469 20247
rect 5684 20216 6469 20244
rect 5684 20204 5690 20216
rect 6457 20213 6469 20216
rect 6503 20213 6515 20247
rect 6932 20244 6960 20284
rect 7092 20275 7104 20284
rect 7098 20272 7104 20275
rect 7156 20272 7162 20324
rect 9116 20315 9174 20321
rect 9116 20281 9128 20315
rect 9162 20312 9174 20315
rect 9306 20312 9312 20324
rect 9162 20284 9312 20312
rect 9162 20281 9174 20284
rect 9116 20275 9174 20281
rect 9306 20272 9312 20284
rect 9364 20272 9370 20324
rect 9490 20272 9496 20324
rect 9548 20312 9554 20324
rect 10612 20312 10640 20352
rect 12434 20340 12440 20352
rect 12492 20340 12498 20392
rect 13906 20380 13912 20392
rect 12912 20352 13912 20380
rect 9548 20284 10640 20312
rect 10772 20315 10830 20321
rect 9548 20272 9554 20284
rect 10772 20281 10784 20315
rect 10818 20312 10830 20315
rect 11054 20312 11060 20324
rect 10818 20284 11060 20312
rect 10818 20281 10830 20284
rect 10772 20275 10830 20281
rect 11054 20272 11060 20284
rect 11112 20312 11118 20324
rect 11698 20312 11704 20324
rect 11112 20284 11704 20312
rect 11112 20272 11118 20284
rect 11698 20272 11704 20284
rect 11756 20272 11762 20324
rect 11974 20272 11980 20324
rect 12032 20312 12038 20324
rect 12912 20312 12940 20352
rect 13906 20340 13912 20352
rect 13964 20340 13970 20392
rect 12032 20284 12940 20312
rect 12980 20315 13038 20321
rect 12032 20272 12038 20284
rect 12980 20281 12992 20315
rect 13026 20312 13038 20315
rect 13998 20312 14004 20324
rect 13026 20284 14004 20312
rect 13026 20281 13038 20284
rect 12980 20275 13038 20281
rect 13998 20272 14004 20284
rect 14056 20272 14062 20324
rect 14108 20312 14136 20488
rect 14366 20448 14372 20460
rect 14327 20420 14372 20448
rect 14366 20408 14372 20420
rect 14424 20408 14430 20460
rect 14458 20340 14464 20392
rect 14516 20380 14522 20392
rect 14625 20383 14683 20389
rect 14625 20380 14637 20383
rect 14516 20352 14637 20380
rect 14516 20340 14522 20352
rect 14625 20349 14637 20352
rect 14671 20349 14683 20383
rect 14625 20343 14683 20349
rect 14918 20340 14924 20392
rect 14976 20380 14982 20392
rect 15948 20380 15976 20556
rect 19334 20544 19340 20556
rect 19392 20544 19398 20596
rect 19429 20587 19487 20593
rect 19429 20553 19441 20587
rect 19475 20584 19487 20587
rect 19886 20584 19892 20596
rect 19475 20556 19892 20584
rect 19475 20553 19487 20556
rect 19429 20547 19487 20553
rect 19886 20544 19892 20556
rect 19944 20544 19950 20596
rect 20346 20544 20352 20596
rect 20404 20584 20410 20596
rect 21177 20587 21235 20593
rect 21177 20584 21189 20587
rect 20404 20556 21189 20584
rect 20404 20544 20410 20556
rect 21177 20553 21189 20556
rect 21223 20553 21235 20587
rect 21177 20547 21235 20553
rect 21358 20544 21364 20596
rect 21416 20584 21422 20596
rect 22005 20587 22063 20593
rect 22005 20584 22017 20587
rect 21416 20556 22017 20584
rect 21416 20544 21422 20556
rect 22005 20553 22017 20556
rect 22051 20553 22063 20587
rect 22005 20547 22063 20553
rect 20898 20476 20904 20528
rect 20956 20516 20962 20528
rect 23382 20516 23388 20528
rect 20956 20488 23388 20516
rect 20956 20476 20962 20488
rect 23382 20476 23388 20488
rect 23440 20476 23446 20528
rect 20714 20408 20720 20460
rect 20772 20448 20778 20460
rect 21729 20451 21787 20457
rect 21729 20448 21741 20451
rect 20772 20420 21741 20448
rect 20772 20408 20778 20420
rect 21729 20417 21741 20420
rect 21775 20417 21787 20451
rect 21729 20411 21787 20417
rect 22649 20451 22707 20457
rect 22649 20417 22661 20451
rect 22695 20417 22707 20451
rect 22649 20411 22707 20417
rect 14976 20352 15976 20380
rect 16025 20383 16083 20389
rect 14976 20340 14982 20352
rect 16025 20349 16037 20383
rect 16071 20380 16083 20383
rect 16114 20380 16120 20392
rect 16071 20352 16120 20380
rect 16071 20349 16083 20352
rect 16025 20343 16083 20349
rect 16114 20340 16120 20352
rect 16172 20380 16178 20392
rect 17954 20380 17960 20392
rect 16172 20352 17960 20380
rect 16172 20340 16178 20352
rect 17954 20340 17960 20352
rect 18012 20380 18018 20392
rect 18049 20383 18107 20389
rect 18049 20380 18061 20383
rect 18012 20352 18061 20380
rect 18012 20340 18018 20352
rect 18049 20349 18061 20352
rect 18095 20349 18107 20383
rect 18049 20343 18107 20349
rect 18138 20340 18144 20392
rect 18196 20380 18202 20392
rect 18316 20383 18374 20389
rect 18316 20380 18328 20383
rect 18196 20352 18328 20380
rect 18196 20340 18202 20352
rect 18316 20349 18328 20352
rect 18362 20380 18374 20383
rect 19150 20380 19156 20392
rect 18362 20352 19156 20380
rect 18362 20349 18374 20352
rect 18316 20343 18374 20349
rect 19150 20340 19156 20352
rect 19208 20340 19214 20392
rect 19702 20380 19708 20392
rect 19663 20352 19708 20380
rect 19702 20340 19708 20352
rect 19760 20340 19766 20392
rect 19794 20340 19800 20392
rect 19852 20380 19858 20392
rect 19972 20383 20030 20389
rect 19972 20380 19984 20383
rect 19852 20352 19984 20380
rect 19852 20340 19858 20352
rect 19972 20349 19984 20352
rect 20018 20380 20030 20383
rect 22664 20380 22692 20411
rect 20018 20352 22692 20380
rect 20018 20349 20030 20352
rect 19972 20343 20030 20349
rect 16292 20315 16350 20321
rect 14108 20284 15884 20312
rect 9858 20244 9864 20256
rect 6932 20216 9864 20244
rect 6457 20207 6515 20213
rect 9858 20204 9864 20216
rect 9916 20204 9922 20256
rect 11146 20204 11152 20256
rect 11204 20244 11210 20256
rect 11606 20244 11612 20256
rect 11204 20216 11612 20244
rect 11204 20204 11210 20216
rect 11606 20204 11612 20216
rect 11664 20204 11670 20256
rect 15562 20204 15568 20256
rect 15620 20244 15626 20256
rect 15749 20247 15807 20253
rect 15749 20244 15761 20247
rect 15620 20216 15761 20244
rect 15620 20204 15626 20216
rect 15749 20213 15761 20216
rect 15795 20213 15807 20247
rect 15856 20244 15884 20284
rect 16292 20281 16304 20315
rect 16338 20312 16350 20315
rect 16574 20312 16580 20324
rect 16338 20284 16580 20312
rect 16338 20281 16350 20284
rect 16292 20275 16350 20281
rect 16574 20272 16580 20284
rect 16632 20272 16638 20324
rect 19886 20312 19892 20324
rect 16684 20284 19892 20312
rect 16684 20244 16712 20284
rect 19886 20272 19892 20284
rect 19944 20272 19950 20324
rect 20070 20272 20076 20324
rect 20128 20312 20134 20324
rect 21637 20315 21695 20321
rect 21637 20312 21649 20315
rect 20128 20284 21649 20312
rect 20128 20272 20134 20284
rect 21637 20281 21649 20284
rect 21683 20281 21695 20315
rect 21637 20275 21695 20281
rect 21910 20272 21916 20324
rect 21968 20312 21974 20324
rect 22465 20315 22523 20321
rect 22465 20312 22477 20315
rect 21968 20284 22477 20312
rect 21968 20272 21974 20284
rect 22465 20281 22477 20284
rect 22511 20281 22523 20315
rect 22465 20275 22523 20281
rect 15856 20216 16712 20244
rect 15749 20207 15807 20213
rect 16758 20204 16764 20256
rect 16816 20244 16822 20256
rect 17405 20247 17463 20253
rect 17405 20244 17417 20247
rect 16816 20216 17417 20244
rect 16816 20204 16822 20216
rect 17405 20213 17417 20216
rect 17451 20244 17463 20247
rect 20714 20244 20720 20256
rect 17451 20216 20720 20244
rect 17451 20213 17463 20216
rect 17405 20207 17463 20213
rect 20714 20204 20720 20216
rect 20772 20204 20778 20256
rect 21082 20244 21088 20256
rect 21043 20216 21088 20244
rect 21082 20204 21088 20216
rect 21140 20204 21146 20256
rect 21542 20244 21548 20256
rect 21503 20216 21548 20244
rect 21542 20204 21548 20216
rect 21600 20204 21606 20256
rect 22370 20244 22376 20256
rect 22331 20216 22376 20244
rect 22370 20204 22376 20216
rect 22428 20204 22434 20256
rect 1104 20154 23276 20176
rect 1104 20102 8379 20154
rect 8431 20102 8443 20154
rect 8495 20102 8507 20154
rect 8559 20102 8571 20154
rect 8623 20102 15776 20154
rect 15828 20102 15840 20154
rect 15892 20102 15904 20154
rect 15956 20102 15968 20154
rect 16020 20102 23276 20154
rect 1104 20080 23276 20102
rect 2958 20040 2964 20052
rect 2871 20012 2964 20040
rect 2958 20000 2964 20012
rect 3016 20000 3022 20052
rect 3050 20000 3056 20052
rect 3108 20040 3114 20052
rect 3421 20043 3479 20049
rect 3421 20040 3433 20043
rect 3108 20012 3433 20040
rect 3108 20000 3114 20012
rect 3421 20009 3433 20012
rect 3467 20009 3479 20043
rect 3421 20003 3479 20009
rect 4065 20043 4123 20049
rect 4065 20009 4077 20043
rect 4111 20040 4123 20043
rect 4522 20040 4528 20052
rect 4111 20012 4528 20040
rect 4111 20009 4123 20012
rect 4065 20003 4123 20009
rect 4522 20000 4528 20012
rect 4580 20000 4586 20052
rect 6454 20040 6460 20052
rect 5276 20012 6460 20040
rect 1854 19981 1860 19984
rect 1848 19972 1860 19981
rect 1815 19944 1860 19972
rect 1848 19935 1860 19944
rect 1854 19932 1860 19935
rect 1912 19932 1918 19984
rect 2976 19972 3004 20000
rect 4433 19975 4491 19981
rect 4433 19972 4445 19975
rect 2976 19944 4445 19972
rect 4433 19941 4445 19944
rect 4479 19941 4491 19975
rect 4433 19935 4491 19941
rect 4614 19932 4620 19984
rect 4672 19972 4678 19984
rect 5276 19981 5304 20012
rect 6454 20000 6460 20012
rect 6512 20000 6518 20052
rect 8662 20040 8668 20052
rect 6564 20012 8668 20040
rect 5261 19975 5319 19981
rect 5261 19972 5273 19975
rect 4672 19944 5273 19972
rect 4672 19932 4678 19944
rect 5261 19941 5273 19944
rect 5307 19941 5319 19975
rect 5261 19935 5319 19941
rect 5620 19975 5678 19981
rect 5620 19941 5632 19975
rect 5666 19972 5678 19975
rect 5810 19972 5816 19984
rect 5666 19944 5816 19972
rect 5666 19941 5678 19944
rect 5620 19935 5678 19941
rect 5810 19932 5816 19944
rect 5868 19932 5874 19984
rect 1581 19907 1639 19913
rect 1581 19873 1593 19907
rect 1627 19904 1639 19907
rect 1670 19904 1676 19916
rect 1627 19876 1676 19904
rect 1627 19873 1639 19876
rect 1581 19867 1639 19873
rect 1670 19864 1676 19876
rect 1728 19864 1734 19916
rect 3145 19907 3203 19913
rect 3145 19873 3157 19907
rect 3191 19904 3203 19907
rect 3237 19907 3295 19913
rect 3237 19904 3249 19907
rect 3191 19876 3249 19904
rect 3191 19873 3203 19876
rect 3145 19867 3203 19873
rect 3237 19873 3249 19876
rect 3283 19873 3295 19907
rect 3237 19867 3295 19873
rect 3418 19864 3424 19916
rect 3476 19904 3482 19916
rect 4246 19904 4252 19916
rect 3476 19876 4252 19904
rect 3476 19864 3482 19876
rect 4246 19864 4252 19876
rect 4304 19864 4310 19916
rect 4525 19907 4583 19913
rect 4525 19873 4537 19907
rect 4571 19904 4583 19907
rect 4798 19904 4804 19916
rect 4571 19876 4804 19904
rect 4571 19873 4583 19876
rect 4525 19867 4583 19873
rect 4798 19864 4804 19876
rect 4856 19864 4862 19916
rect 6362 19904 6368 19916
rect 5184 19876 6368 19904
rect 3878 19796 3884 19848
rect 3936 19836 3942 19848
rect 4617 19839 4675 19845
rect 4617 19836 4629 19839
rect 3936 19808 4629 19836
rect 3936 19796 3942 19808
rect 4617 19805 4629 19808
rect 4663 19805 4675 19839
rect 4617 19799 4675 19805
rect 4062 19728 4068 19780
rect 4120 19768 4126 19780
rect 5184 19768 5212 19876
rect 6362 19864 6368 19876
rect 6420 19864 6426 19916
rect 5261 19839 5319 19845
rect 5261 19805 5273 19839
rect 5307 19836 5319 19839
rect 5353 19839 5411 19845
rect 5353 19836 5365 19839
rect 5307 19808 5365 19836
rect 5307 19805 5319 19808
rect 5261 19799 5319 19805
rect 5353 19805 5365 19808
rect 5399 19805 5411 19839
rect 5353 19799 5411 19805
rect 4120 19740 5212 19768
rect 4120 19728 4126 19740
rect 3145 19703 3203 19709
rect 3145 19669 3157 19703
rect 3191 19700 3203 19703
rect 6564 19700 6592 20012
rect 8662 20000 8668 20012
rect 8720 20000 8726 20052
rect 9674 20000 9680 20052
rect 9732 20040 9738 20052
rect 9858 20040 9864 20052
rect 9732 20012 9864 20040
rect 9732 20000 9738 20012
rect 9858 20000 9864 20012
rect 9916 20000 9922 20052
rect 10594 20000 10600 20052
rect 10652 20040 10658 20052
rect 11063 20043 11121 20049
rect 11063 20040 11075 20043
rect 10652 20012 11075 20040
rect 10652 20000 10658 20012
rect 11063 20009 11075 20012
rect 11109 20009 11121 20043
rect 11063 20003 11121 20009
rect 13998 20000 14004 20052
rect 14056 20040 14062 20052
rect 14093 20043 14151 20049
rect 14093 20040 14105 20043
rect 14056 20012 14105 20040
rect 14056 20000 14062 20012
rect 14093 20009 14105 20012
rect 14139 20040 14151 20043
rect 15657 20043 15715 20049
rect 15657 20040 15669 20043
rect 14139 20012 15669 20040
rect 14139 20009 14151 20012
rect 14093 20003 14151 20009
rect 15657 20009 15669 20012
rect 15703 20009 15715 20043
rect 15657 20003 15715 20009
rect 17865 20043 17923 20049
rect 17865 20009 17877 20043
rect 17911 20040 17923 20043
rect 18138 20040 18144 20052
rect 17911 20012 18144 20040
rect 17911 20009 17923 20012
rect 17865 20003 17923 20009
rect 18138 20000 18144 20012
rect 18196 20000 18202 20052
rect 18230 20000 18236 20052
rect 18288 20040 18294 20052
rect 20806 20040 20812 20052
rect 18288 20012 20812 20040
rect 18288 20000 18294 20012
rect 20806 20000 20812 20012
rect 20864 20000 20870 20052
rect 21450 20000 21456 20052
rect 21508 20000 21514 20052
rect 7466 19981 7472 19984
rect 7460 19935 7472 19981
rect 7524 19972 7530 19984
rect 7524 19944 7560 19972
rect 7466 19932 7472 19935
rect 7524 19932 7530 19944
rect 7742 19932 7748 19984
rect 7800 19972 7806 19984
rect 12710 19972 12716 19984
rect 7800 19944 8892 19972
rect 7800 19932 7806 19944
rect 7006 19864 7012 19916
rect 7064 19904 7070 19916
rect 7193 19907 7251 19913
rect 7193 19904 7205 19907
rect 7064 19876 7205 19904
rect 7064 19864 7070 19876
rect 7193 19873 7205 19876
rect 7239 19873 7251 19907
rect 7193 19867 7251 19873
rect 7834 19864 7840 19916
rect 7892 19904 7898 19916
rect 8864 19913 8892 19944
rect 9508 19944 10456 19972
rect 8849 19907 8907 19913
rect 7892 19876 8248 19904
rect 7892 19864 7898 19876
rect 8220 19768 8248 19876
rect 8849 19873 8861 19907
rect 8895 19873 8907 19907
rect 8849 19867 8907 19873
rect 9214 19864 9220 19916
rect 9272 19904 9278 19916
rect 9508 19904 9536 19944
rect 9272 19876 9536 19904
rect 9272 19864 9278 19876
rect 9674 19864 9680 19916
rect 9732 19904 9738 19916
rect 10428 19913 10456 19944
rect 12636 19944 12716 19972
rect 10413 19907 10471 19913
rect 9732 19876 9777 19904
rect 9732 19864 9738 19876
rect 10413 19873 10425 19907
rect 10459 19873 10471 19907
rect 10413 19867 10471 19873
rect 11333 19907 11391 19913
rect 11333 19873 11345 19907
rect 11379 19904 11391 19907
rect 12636 19904 12664 19944
rect 12710 19932 12716 19944
rect 12768 19932 12774 19984
rect 12894 19932 12900 19984
rect 12952 19932 12958 19984
rect 13170 19932 13176 19984
rect 13228 19972 13234 19984
rect 14642 19972 14648 19984
rect 13228 19944 14648 19972
rect 13228 19932 13234 19944
rect 14642 19932 14648 19944
rect 14700 19932 14706 19984
rect 14737 19975 14795 19981
rect 14737 19941 14749 19975
rect 14783 19972 14795 19975
rect 15562 19972 15568 19984
rect 14783 19944 15568 19972
rect 14783 19941 14795 19944
rect 14737 19935 14795 19941
rect 15562 19932 15568 19944
rect 15620 19932 15626 19984
rect 16758 19981 16764 19984
rect 15749 19975 15807 19981
rect 15749 19941 15761 19975
rect 15795 19941 15807 19975
rect 16752 19972 16764 19981
rect 16719 19944 16764 19972
rect 15749 19935 15807 19941
rect 16752 19935 16764 19944
rect 12912 19904 12940 19932
rect 11379 19876 12664 19904
rect 12728 19876 12940 19904
rect 12980 19907 13038 19913
rect 11379 19873 11391 19876
rect 11333 19867 11391 19873
rect 10597 19839 10655 19845
rect 10597 19805 10609 19839
rect 10643 19805 10655 19839
rect 10597 19799 10655 19805
rect 11103 19839 11161 19845
rect 11103 19805 11115 19839
rect 11149 19836 11161 19839
rect 11422 19836 11428 19848
rect 11149 19808 11428 19836
rect 11149 19805 11161 19808
rect 11103 19799 11161 19805
rect 9033 19771 9091 19777
rect 9033 19768 9045 19771
rect 8220 19740 9045 19768
rect 9033 19737 9045 19740
rect 9079 19737 9091 19771
rect 9033 19731 9091 19737
rect 10410 19728 10416 19780
rect 10468 19768 10474 19780
rect 10612 19768 10640 19799
rect 11422 19796 11428 19808
rect 11480 19796 11486 19848
rect 12728 19845 12756 19876
rect 12980 19873 12992 19907
rect 13026 19904 13038 19907
rect 14553 19907 14611 19913
rect 13026 19876 14320 19904
rect 13026 19873 13038 19876
rect 12980 19867 13038 19873
rect 14016 19848 14044 19876
rect 12713 19839 12771 19845
rect 12713 19805 12725 19839
rect 12759 19805 12771 19839
rect 12713 19799 12771 19805
rect 13998 19796 14004 19848
rect 14056 19796 14062 19848
rect 14292 19836 14320 19876
rect 14553 19873 14565 19907
rect 14599 19904 14611 19907
rect 15010 19904 15016 19916
rect 14599 19876 15016 19904
rect 14599 19873 14611 19876
rect 14553 19867 14611 19873
rect 15010 19864 15016 19876
rect 15068 19864 15074 19916
rect 15764 19836 15792 19935
rect 16758 19932 16764 19935
rect 16816 19932 16822 19984
rect 17954 19932 17960 19984
rect 18012 19972 18018 19984
rect 18598 19972 18604 19984
rect 18012 19944 18604 19972
rect 18012 19932 18018 19944
rect 18598 19932 18604 19944
rect 18656 19972 18662 19984
rect 19061 19975 19119 19981
rect 19061 19972 19073 19975
rect 18656 19944 19073 19972
rect 18656 19932 18662 19944
rect 19061 19941 19073 19944
rect 19107 19941 19119 19975
rect 19061 19935 19119 19941
rect 19420 19975 19478 19981
rect 19420 19941 19432 19975
rect 19466 19972 19478 19975
rect 21082 19972 21088 19984
rect 19466 19944 21088 19972
rect 19466 19941 19478 19944
rect 19420 19935 19478 19941
rect 21082 19932 21088 19944
rect 21140 19932 21146 19984
rect 21468 19972 21496 20000
rect 21192 19944 21496 19972
rect 16022 19864 16028 19916
rect 16080 19904 16086 19916
rect 18509 19907 18567 19913
rect 18509 19904 18521 19907
rect 16080 19876 18521 19904
rect 16080 19864 16086 19876
rect 18509 19873 18521 19876
rect 18555 19873 18567 19907
rect 21192 19904 21220 19944
rect 21450 19913 21456 19916
rect 21444 19904 21456 19913
rect 18509 19867 18567 19873
rect 18892 19876 21220 19904
rect 21411 19876 21456 19904
rect 14292 19808 15792 19836
rect 15933 19839 15991 19845
rect 15933 19805 15945 19839
rect 15979 19805 15991 19839
rect 15933 19799 15991 19805
rect 10468 19740 10640 19768
rect 15948 19768 15976 19799
rect 16114 19796 16120 19848
rect 16172 19836 16178 19848
rect 16485 19839 16543 19845
rect 16485 19836 16497 19839
rect 16172 19808 16497 19836
rect 16172 19796 16178 19808
rect 16485 19805 16497 19808
rect 16531 19805 16543 19839
rect 16485 19799 16543 19805
rect 18230 19796 18236 19848
rect 18288 19836 18294 19848
rect 18601 19839 18659 19845
rect 18601 19836 18613 19839
rect 18288 19808 18613 19836
rect 18288 19796 18294 19808
rect 18601 19805 18613 19808
rect 18647 19805 18659 19839
rect 18601 19799 18659 19805
rect 18690 19796 18696 19848
rect 18748 19836 18754 19848
rect 18748 19808 18793 19836
rect 18748 19796 18754 19808
rect 16206 19768 16212 19780
rect 15948 19740 16212 19768
rect 10468 19728 10474 19740
rect 16206 19728 16212 19740
rect 16264 19728 16270 19780
rect 17494 19728 17500 19780
rect 17552 19768 17558 19780
rect 18892 19768 18920 19876
rect 21444 19867 21456 19876
rect 21450 19864 21456 19867
rect 21508 19864 21514 19916
rect 21818 19864 21824 19916
rect 21876 19904 21882 19916
rect 22649 19907 22707 19913
rect 22649 19904 22661 19907
rect 21876 19876 22661 19904
rect 21876 19864 21882 19876
rect 22649 19873 22661 19876
rect 22695 19873 22707 19907
rect 22649 19867 22707 19873
rect 19061 19839 19119 19845
rect 19061 19805 19073 19839
rect 19107 19836 19119 19839
rect 19153 19839 19211 19845
rect 19153 19836 19165 19839
rect 19107 19808 19165 19836
rect 19107 19805 19119 19808
rect 19061 19799 19119 19805
rect 19153 19805 19165 19808
rect 19199 19805 19211 19839
rect 19153 19799 19211 19805
rect 17552 19740 18920 19768
rect 17552 19728 17558 19740
rect 3191 19672 6592 19700
rect 6733 19703 6791 19709
rect 3191 19669 3203 19672
rect 3145 19663 3203 19669
rect 6733 19669 6745 19703
rect 6779 19700 6791 19703
rect 7098 19700 7104 19712
rect 6779 19672 7104 19700
rect 6779 19669 6791 19672
rect 6733 19663 6791 19669
rect 7098 19660 7104 19672
rect 7156 19700 7162 19712
rect 8110 19700 8116 19712
rect 7156 19672 8116 19700
rect 7156 19660 7162 19672
rect 8110 19660 8116 19672
rect 8168 19660 8174 19712
rect 8294 19660 8300 19712
rect 8352 19700 8358 19712
rect 8573 19703 8631 19709
rect 8573 19700 8585 19703
rect 8352 19672 8585 19700
rect 8352 19660 8358 19672
rect 8573 19669 8585 19672
rect 8619 19700 8631 19703
rect 8754 19700 8760 19712
rect 8619 19672 8760 19700
rect 8619 19669 8631 19672
rect 8573 19663 8631 19669
rect 8754 19660 8760 19672
rect 8812 19660 8818 19712
rect 10226 19700 10232 19712
rect 10187 19672 10232 19700
rect 10226 19660 10232 19672
rect 10284 19660 10290 19712
rect 11054 19660 11060 19712
rect 11112 19700 11118 19712
rect 12437 19703 12495 19709
rect 12437 19700 12449 19703
rect 11112 19672 12449 19700
rect 11112 19660 11118 19672
rect 12437 19669 12449 19672
rect 12483 19669 12495 19703
rect 12437 19663 12495 19669
rect 14458 19660 14464 19712
rect 14516 19700 14522 19712
rect 14921 19703 14979 19709
rect 14921 19700 14933 19703
rect 14516 19672 14933 19700
rect 14516 19660 14522 19672
rect 14921 19669 14933 19672
rect 14967 19669 14979 19703
rect 14921 19663 14979 19669
rect 15289 19703 15347 19709
rect 15289 19669 15301 19703
rect 15335 19700 15347 19703
rect 17402 19700 17408 19712
rect 15335 19672 17408 19700
rect 15335 19669 15347 19672
rect 15289 19663 15347 19669
rect 17402 19660 17408 19672
rect 17460 19660 17466 19712
rect 17770 19660 17776 19712
rect 17828 19700 17834 19712
rect 18141 19703 18199 19709
rect 18141 19700 18153 19703
rect 17828 19672 18153 19700
rect 17828 19660 17834 19672
rect 18141 19669 18153 19672
rect 18187 19669 18199 19703
rect 18141 19663 18199 19669
rect 18414 19660 18420 19712
rect 18472 19700 18478 19712
rect 18874 19700 18880 19712
rect 18472 19672 18880 19700
rect 18472 19660 18478 19672
rect 18874 19660 18880 19672
rect 18932 19660 18938 19712
rect 19168 19700 19196 19799
rect 20530 19796 20536 19848
rect 20588 19796 20594 19848
rect 20990 19796 20996 19848
rect 21048 19836 21054 19848
rect 21177 19839 21235 19845
rect 21177 19836 21189 19839
rect 21048 19808 21189 19836
rect 21048 19796 21054 19808
rect 21177 19805 21189 19808
rect 21223 19805 21235 19839
rect 21177 19799 21235 19805
rect 19794 19700 19800 19712
rect 19168 19672 19800 19700
rect 19794 19660 19800 19672
rect 19852 19660 19858 19712
rect 20548 19709 20576 19796
rect 20533 19703 20591 19709
rect 20533 19669 20545 19703
rect 20579 19669 20591 19703
rect 22554 19700 22560 19712
rect 22515 19672 22560 19700
rect 20533 19663 20591 19669
rect 22554 19660 22560 19672
rect 22612 19660 22618 19712
rect 22830 19700 22836 19712
rect 22791 19672 22836 19700
rect 22830 19660 22836 19672
rect 22888 19660 22894 19712
rect 1104 19610 23276 19632
rect 1104 19558 4680 19610
rect 4732 19558 4744 19610
rect 4796 19558 4808 19610
rect 4860 19558 4872 19610
rect 4924 19558 12078 19610
rect 12130 19558 12142 19610
rect 12194 19558 12206 19610
rect 12258 19558 12270 19610
rect 12322 19558 19475 19610
rect 19527 19558 19539 19610
rect 19591 19558 19603 19610
rect 19655 19558 19667 19610
rect 19719 19558 23276 19610
rect 1104 19536 23276 19558
rect 2593 19499 2651 19505
rect 2593 19465 2605 19499
rect 2639 19496 2651 19499
rect 4154 19496 4160 19508
rect 2639 19468 4160 19496
rect 2639 19465 2651 19468
rect 2593 19459 2651 19465
rect 4154 19456 4160 19468
rect 4212 19456 4218 19508
rect 4982 19456 4988 19508
rect 5040 19496 5046 19508
rect 13170 19496 13176 19508
rect 5040 19468 5948 19496
rect 5040 19456 5046 19468
rect 1486 19388 1492 19440
rect 1544 19428 1550 19440
rect 3050 19428 3056 19440
rect 1544 19400 3056 19428
rect 1544 19388 1550 19400
rect 3050 19388 3056 19400
rect 3108 19388 3114 19440
rect 3878 19428 3884 19440
rect 3160 19400 3884 19428
rect 3160 19372 3188 19400
rect 3878 19388 3884 19400
rect 3936 19428 3942 19440
rect 4614 19428 4620 19440
rect 3936 19400 4620 19428
rect 3936 19388 3942 19400
rect 2133 19363 2191 19369
rect 2133 19329 2145 19363
rect 2179 19360 2191 19363
rect 3142 19360 3148 19372
rect 2179 19332 3148 19360
rect 2179 19329 2191 19332
rect 2133 19323 2191 19329
rect 3142 19320 3148 19332
rect 3200 19320 3206 19372
rect 3326 19320 3332 19372
rect 3384 19360 3390 19372
rect 4172 19369 4200 19400
rect 4614 19388 4620 19400
rect 4672 19388 4678 19440
rect 4157 19363 4215 19369
rect 3384 19332 4108 19360
rect 3384 19320 3390 19332
rect 2222 19252 2228 19304
rect 2280 19292 2286 19304
rect 4080 19292 4108 19332
rect 4157 19329 4169 19363
rect 4203 19329 4215 19363
rect 4157 19323 4215 19329
rect 4522 19320 4528 19372
rect 4580 19320 4586 19372
rect 4540 19292 4568 19320
rect 4617 19295 4675 19301
rect 4617 19292 4629 19295
rect 2280 19264 3648 19292
rect 4080 19264 4629 19292
rect 2280 19252 2286 19264
rect 2041 19227 2099 19233
rect 2041 19193 2053 19227
rect 2087 19224 2099 19227
rect 3142 19224 3148 19236
rect 2087 19196 3148 19224
rect 2087 19193 2099 19196
rect 2041 19187 2099 19193
rect 3142 19184 3148 19196
rect 3200 19184 3206 19236
rect 1578 19156 1584 19168
rect 1539 19128 1584 19156
rect 1578 19116 1584 19128
rect 1636 19116 1642 19168
rect 1946 19156 1952 19168
rect 1907 19128 1952 19156
rect 1946 19116 1952 19128
rect 2004 19116 2010 19168
rect 2866 19116 2872 19168
rect 2924 19156 2930 19168
rect 2961 19159 3019 19165
rect 2961 19156 2973 19159
rect 2924 19128 2973 19156
rect 2924 19116 2930 19128
rect 2961 19125 2973 19128
rect 3007 19125 3019 19159
rect 2961 19119 3019 19125
rect 3053 19159 3111 19165
rect 3053 19125 3065 19159
rect 3099 19156 3111 19159
rect 3510 19156 3516 19168
rect 3099 19128 3516 19156
rect 3099 19125 3111 19128
rect 3053 19119 3111 19125
rect 3510 19116 3516 19128
rect 3568 19116 3574 19168
rect 3620 19165 3648 19264
rect 4617 19261 4629 19264
rect 4663 19261 4675 19295
rect 4617 19255 4675 19261
rect 4884 19295 4942 19301
rect 4884 19261 4896 19295
rect 4930 19292 4942 19295
rect 5166 19292 5172 19304
rect 4930 19264 5172 19292
rect 4930 19261 4942 19264
rect 4884 19255 4942 19261
rect 5166 19252 5172 19264
rect 5224 19252 5230 19304
rect 3878 19184 3884 19236
rect 3936 19224 3942 19236
rect 3973 19227 4031 19233
rect 3973 19224 3985 19227
rect 3936 19196 3985 19224
rect 3936 19184 3942 19196
rect 3973 19193 3985 19196
rect 4019 19193 4031 19227
rect 5920 19224 5948 19468
rect 6840 19468 13176 19496
rect 6270 19292 6276 19304
rect 6231 19264 6276 19292
rect 6270 19252 6276 19264
rect 6328 19252 6334 19304
rect 6840 19301 6868 19468
rect 13170 19456 13176 19468
rect 13228 19456 13234 19508
rect 14090 19496 14096 19508
rect 13372 19468 14096 19496
rect 9122 19388 9128 19440
rect 9180 19388 9186 19440
rect 9398 19388 9404 19440
rect 9456 19428 9462 19440
rect 9456 19400 10272 19428
rect 9456 19388 9462 19400
rect 7742 19320 7748 19372
rect 7800 19360 7806 19372
rect 7926 19369 7932 19372
rect 7884 19363 7932 19369
rect 7884 19360 7896 19363
rect 7800 19332 7896 19360
rect 7800 19320 7806 19332
rect 7884 19329 7896 19332
rect 7930 19329 7932 19363
rect 7884 19323 7932 19329
rect 7926 19320 7932 19323
rect 7984 19320 7990 19372
rect 8067 19363 8125 19369
rect 8067 19329 8079 19363
rect 8113 19360 8125 19363
rect 9131 19360 9159 19388
rect 10244 19369 10272 19400
rect 11790 19388 11796 19440
rect 11848 19428 11854 19440
rect 13372 19428 13400 19468
rect 14090 19456 14096 19468
rect 14148 19456 14154 19508
rect 14182 19456 14188 19508
rect 14240 19496 14246 19508
rect 14240 19468 15792 19496
rect 14240 19456 14246 19468
rect 11848 19400 13400 19428
rect 11848 19388 11854 19400
rect 13722 19388 13728 19440
rect 13780 19428 13786 19440
rect 14550 19428 14556 19440
rect 13780 19400 14556 19428
rect 13780 19388 13786 19400
rect 14550 19388 14556 19400
rect 14608 19388 14614 19440
rect 15654 19428 15660 19440
rect 14936 19400 15660 19428
rect 10229 19363 10287 19369
rect 8113 19332 9159 19360
rect 9232 19332 9812 19360
rect 8113 19329 8125 19332
rect 8067 19323 8125 19329
rect 6825 19295 6883 19301
rect 6825 19261 6837 19295
rect 6871 19261 6883 19295
rect 6825 19255 6883 19261
rect 7561 19295 7619 19301
rect 7561 19261 7573 19295
rect 7607 19261 7619 19295
rect 7561 19255 7619 19261
rect 5920 19196 7052 19224
rect 3973 19187 4031 19193
rect 3605 19159 3663 19165
rect 3605 19125 3617 19159
rect 3651 19125 3663 19159
rect 4062 19156 4068 19168
rect 4023 19128 4068 19156
rect 3605 19119 3663 19125
rect 4062 19116 4068 19128
rect 4120 19116 4126 19168
rect 5810 19116 5816 19168
rect 5868 19156 5874 19168
rect 7024 19165 7052 19196
rect 5997 19159 6055 19165
rect 5997 19156 6009 19159
rect 5868 19128 6009 19156
rect 5868 19116 5874 19128
rect 5997 19125 6009 19128
rect 6043 19125 6055 19159
rect 5997 19119 6055 19125
rect 7009 19159 7067 19165
rect 7009 19125 7021 19159
rect 7055 19125 7067 19159
rect 7009 19119 7067 19125
rect 7098 19116 7104 19168
rect 7156 19156 7162 19168
rect 7576 19156 7604 19255
rect 7650 19252 7656 19304
rect 7708 19292 7714 19304
rect 8202 19292 8208 19304
rect 7708 19264 8208 19292
rect 7708 19252 7714 19264
rect 8202 19252 8208 19264
rect 8260 19252 8266 19304
rect 8297 19295 8355 19301
rect 8297 19261 8309 19295
rect 8343 19292 8355 19295
rect 9122 19292 9128 19304
rect 8343 19264 9128 19292
rect 8343 19261 8355 19264
rect 8297 19255 8355 19261
rect 9122 19252 9128 19264
rect 9180 19252 9186 19304
rect 9030 19184 9036 19236
rect 9088 19224 9094 19236
rect 9232 19224 9260 19332
rect 9674 19292 9680 19304
rect 9088 19196 9260 19224
rect 9324 19264 9680 19292
rect 9088 19184 9094 19196
rect 9324 19156 9352 19264
rect 9674 19252 9680 19264
rect 9732 19252 9738 19304
rect 7156 19128 9352 19156
rect 9401 19159 9459 19165
rect 7156 19116 7162 19128
rect 9401 19125 9413 19159
rect 9447 19156 9459 19159
rect 9582 19156 9588 19168
rect 9447 19128 9588 19156
rect 9447 19125 9459 19128
rect 9401 19119 9459 19125
rect 9582 19116 9588 19128
rect 9640 19116 9646 19168
rect 9677 19159 9735 19165
rect 9677 19125 9689 19159
rect 9723 19156 9735 19159
rect 9784 19156 9812 19332
rect 10229 19329 10241 19363
rect 10275 19329 10287 19363
rect 10229 19323 10287 19329
rect 11698 19320 11704 19372
rect 11756 19360 11762 19372
rect 12989 19363 13047 19369
rect 12989 19360 13001 19363
rect 11756 19332 13001 19360
rect 11756 19320 11762 19332
rect 12989 19329 13001 19332
rect 13035 19329 13047 19363
rect 14001 19363 14059 19369
rect 14001 19360 14013 19363
rect 12989 19323 13047 19329
rect 13096 19332 14013 19360
rect 10318 19252 10324 19304
rect 10376 19292 10382 19304
rect 10502 19292 10508 19304
rect 10376 19264 10508 19292
rect 10376 19252 10382 19264
rect 10502 19252 10508 19264
rect 10560 19292 10566 19304
rect 10689 19295 10747 19301
rect 10689 19292 10701 19295
rect 10560 19264 10701 19292
rect 10560 19252 10566 19264
rect 10689 19261 10701 19264
rect 10735 19261 10747 19295
rect 10689 19255 10747 19261
rect 10956 19295 11014 19301
rect 10956 19261 10968 19295
rect 11002 19292 11014 19295
rect 12526 19292 12532 19304
rect 11002 19264 12532 19292
rect 11002 19261 11014 19264
rect 10956 19255 11014 19261
rect 12526 19252 12532 19264
rect 12584 19292 12590 19304
rect 13096 19292 13124 19332
rect 14001 19329 14013 19332
rect 14047 19329 14059 19363
rect 14936 19360 14964 19400
rect 15654 19388 15660 19400
rect 15712 19388 15718 19440
rect 15764 19428 15792 19468
rect 16574 19456 16580 19508
rect 16632 19496 16638 19508
rect 20070 19496 20076 19508
rect 16632 19468 19472 19496
rect 20031 19468 20076 19496
rect 16632 19456 16638 19468
rect 17494 19428 17500 19440
rect 15764 19400 17500 19428
rect 17494 19388 17500 19400
rect 17552 19388 17558 19440
rect 19444 19428 19472 19468
rect 20070 19456 20076 19468
rect 20128 19456 20134 19508
rect 21634 19456 21640 19508
rect 21692 19496 21698 19508
rect 22094 19496 22100 19508
rect 21692 19468 22100 19496
rect 21692 19456 21698 19468
rect 22094 19456 22100 19468
rect 22152 19456 22158 19508
rect 19444 19400 20668 19428
rect 14001 19323 14059 19329
rect 14384 19332 14964 19360
rect 15105 19363 15163 19369
rect 12584 19264 13124 19292
rect 13817 19295 13875 19301
rect 12584 19252 12590 19264
rect 13817 19261 13829 19295
rect 13863 19292 13875 19295
rect 14384 19292 14412 19332
rect 15105 19329 15117 19363
rect 15151 19360 15163 19363
rect 15194 19360 15200 19372
rect 15151 19332 15200 19360
rect 15151 19329 15163 19332
rect 15105 19323 15163 19329
rect 15194 19320 15200 19332
rect 15252 19360 15258 19372
rect 16117 19363 16175 19369
rect 16117 19360 16129 19363
rect 15252 19332 16129 19360
rect 15252 19320 15258 19332
rect 16117 19329 16129 19332
rect 16163 19360 16175 19363
rect 16206 19360 16212 19372
rect 16163 19332 16212 19360
rect 16163 19329 16175 19332
rect 16117 19323 16175 19329
rect 16206 19320 16212 19332
rect 16264 19320 16270 19372
rect 17129 19363 17187 19369
rect 17129 19329 17141 19363
rect 17175 19360 17187 19363
rect 17586 19360 17592 19372
rect 17175 19332 17592 19360
rect 17175 19329 17187 19332
rect 17129 19323 17187 19329
rect 17586 19320 17592 19332
rect 17644 19320 17650 19372
rect 18506 19320 18512 19372
rect 18564 19360 18570 19372
rect 18782 19369 18788 19372
rect 18739 19363 18788 19369
rect 18564 19332 18609 19360
rect 18564 19320 18570 19332
rect 18739 19329 18751 19363
rect 18785 19329 18788 19363
rect 18739 19323 18788 19329
rect 18782 19320 18788 19323
rect 18840 19320 18846 19372
rect 19794 19320 19800 19372
rect 19852 19360 19858 19372
rect 20640 19369 20668 19400
rect 20625 19363 20683 19369
rect 19852 19332 20576 19360
rect 19852 19320 19858 19332
rect 16945 19295 17003 19301
rect 16945 19292 16957 19295
rect 13863 19264 14412 19292
rect 14476 19264 16957 19292
rect 13863 19261 13875 19264
rect 13817 19255 13875 19261
rect 10137 19227 10195 19233
rect 10137 19193 10149 19227
rect 10183 19224 10195 19227
rect 11054 19224 11060 19236
rect 10183 19196 11060 19224
rect 10183 19193 10195 19196
rect 10137 19187 10195 19193
rect 11054 19184 11060 19196
rect 11112 19184 11118 19236
rect 11330 19184 11336 19236
rect 11388 19224 11394 19236
rect 11388 19196 12480 19224
rect 11388 19184 11394 19196
rect 9723 19128 9812 19156
rect 9723 19125 9735 19128
rect 9677 19119 9735 19125
rect 9858 19116 9864 19168
rect 9916 19156 9922 19168
rect 10045 19159 10103 19165
rect 10045 19156 10057 19159
rect 9916 19128 10057 19156
rect 9916 19116 9922 19128
rect 10045 19125 10057 19128
rect 10091 19156 10103 19159
rect 11698 19156 11704 19168
rect 10091 19128 11704 19156
rect 10091 19125 10103 19128
rect 10045 19119 10103 19125
rect 11698 19116 11704 19128
rect 11756 19116 11762 19168
rect 11974 19116 11980 19168
rect 12032 19156 12038 19168
rect 12452 19165 12480 19196
rect 12069 19159 12127 19165
rect 12069 19156 12081 19159
rect 12032 19128 12081 19156
rect 12032 19116 12038 19128
rect 12069 19125 12081 19128
rect 12115 19125 12127 19159
rect 12069 19119 12127 19125
rect 12437 19159 12495 19165
rect 12437 19125 12449 19159
rect 12483 19125 12495 19159
rect 12437 19119 12495 19125
rect 12710 19116 12716 19168
rect 12768 19156 12774 19168
rect 12805 19159 12863 19165
rect 12805 19156 12817 19159
rect 12768 19128 12817 19156
rect 12768 19116 12774 19128
rect 12805 19125 12817 19128
rect 12851 19125 12863 19159
rect 12805 19119 12863 19125
rect 12897 19159 12955 19165
rect 12897 19125 12909 19159
rect 12943 19156 12955 19159
rect 12986 19156 12992 19168
rect 12943 19128 12992 19156
rect 12943 19125 12955 19128
rect 12897 19119 12955 19125
rect 12986 19116 12992 19128
rect 13044 19116 13050 19168
rect 13078 19116 13084 19168
rect 13136 19156 13142 19168
rect 13449 19159 13507 19165
rect 13449 19156 13461 19159
rect 13136 19128 13461 19156
rect 13136 19116 13142 19128
rect 13449 19125 13461 19128
rect 13495 19125 13507 19159
rect 13449 19119 13507 19125
rect 13538 19116 13544 19168
rect 13596 19156 13602 19168
rect 14476 19165 14504 19264
rect 16945 19261 16957 19264
rect 16991 19261 17003 19295
rect 16945 19255 17003 19261
rect 17497 19295 17555 19301
rect 17497 19261 17509 19295
rect 17543 19292 17555 19295
rect 17954 19292 17960 19304
rect 17543 19264 17960 19292
rect 17543 19261 17555 19264
rect 17497 19255 17555 19261
rect 17954 19252 17960 19264
rect 18012 19252 18018 19304
rect 18057 19295 18115 19301
rect 18057 19261 18069 19295
rect 18103 19261 18115 19295
rect 20441 19295 20499 19301
rect 20441 19292 20453 19295
rect 18057 19255 18115 19261
rect 19720 19264 20453 19292
rect 16853 19227 16911 19233
rect 16853 19224 16865 19227
rect 15488 19196 16865 19224
rect 13909 19159 13967 19165
rect 13909 19156 13921 19159
rect 13596 19128 13921 19156
rect 13596 19116 13602 19128
rect 13909 19125 13921 19128
rect 13955 19125 13967 19159
rect 13909 19119 13967 19125
rect 14461 19159 14519 19165
rect 14461 19125 14473 19159
rect 14507 19125 14519 19159
rect 14826 19156 14832 19168
rect 14787 19128 14832 19156
rect 14461 19119 14519 19125
rect 14826 19116 14832 19128
rect 14884 19116 14890 19168
rect 14921 19159 14979 19165
rect 14921 19125 14933 19159
rect 14967 19156 14979 19159
rect 15286 19156 15292 19168
rect 14967 19128 15292 19156
rect 14967 19125 14979 19128
rect 14921 19119 14979 19125
rect 15286 19116 15292 19128
rect 15344 19116 15350 19168
rect 15488 19165 15516 19196
rect 16853 19193 16865 19196
rect 16899 19193 16911 19227
rect 18072 19224 18100 19255
rect 18072 19196 18184 19224
rect 16853 19187 16911 19193
rect 18156 19168 18184 19196
rect 15473 19159 15531 19165
rect 15473 19125 15485 19159
rect 15519 19125 15531 19159
rect 15473 19119 15531 19125
rect 15562 19116 15568 19168
rect 15620 19156 15626 19168
rect 15841 19159 15899 19165
rect 15841 19156 15853 19159
rect 15620 19128 15853 19156
rect 15620 19116 15626 19128
rect 15841 19125 15853 19128
rect 15887 19125 15899 19159
rect 15841 19119 15899 19125
rect 15933 19159 15991 19165
rect 15933 19125 15945 19159
rect 15979 19156 15991 19159
rect 16114 19156 16120 19168
rect 15979 19128 16120 19156
rect 15979 19125 15991 19128
rect 15933 19119 15991 19125
rect 16114 19116 16120 19128
rect 16172 19116 16178 19168
rect 16206 19116 16212 19168
rect 16264 19156 16270 19168
rect 16485 19159 16543 19165
rect 16485 19156 16497 19159
rect 16264 19128 16497 19156
rect 16264 19116 16270 19128
rect 16485 19125 16497 19128
rect 16531 19125 16543 19159
rect 16485 19119 16543 19125
rect 18138 19116 18144 19168
rect 18196 19116 18202 19168
rect 18515 19159 18573 19165
rect 18515 19125 18527 19159
rect 18561 19156 18573 19159
rect 18782 19156 18788 19168
rect 18561 19128 18788 19156
rect 18561 19125 18573 19128
rect 18515 19119 18573 19125
rect 18782 19116 18788 19128
rect 18840 19116 18846 19168
rect 19058 19116 19064 19168
rect 19116 19156 19122 19168
rect 19720 19156 19748 19264
rect 20441 19261 20453 19264
rect 20487 19261 20499 19295
rect 20441 19255 20499 19261
rect 20548 19224 20576 19332
rect 20625 19329 20637 19363
rect 20671 19329 20683 19363
rect 20625 19323 20683 19329
rect 20901 19295 20959 19301
rect 20901 19261 20913 19295
rect 20947 19261 20959 19295
rect 20901 19255 20959 19261
rect 20916 19224 20944 19255
rect 20548 19196 20944 19224
rect 20916 19168 20944 19196
rect 21168 19227 21226 19233
rect 21168 19193 21180 19227
rect 21214 19224 21226 19227
rect 21634 19224 21640 19236
rect 21214 19196 21640 19224
rect 21214 19193 21226 19196
rect 21168 19187 21226 19193
rect 21634 19184 21640 19196
rect 21692 19184 21698 19236
rect 19116 19128 19748 19156
rect 19889 19159 19947 19165
rect 19116 19116 19122 19128
rect 19889 19125 19901 19159
rect 19935 19156 19947 19159
rect 20070 19156 20076 19168
rect 19935 19128 20076 19156
rect 19935 19125 19947 19128
rect 19889 19119 19947 19125
rect 20070 19116 20076 19128
rect 20128 19116 20134 19168
rect 20346 19116 20352 19168
rect 20404 19156 20410 19168
rect 20533 19159 20591 19165
rect 20533 19156 20545 19159
rect 20404 19128 20545 19156
rect 20404 19116 20410 19128
rect 20533 19125 20545 19128
rect 20579 19125 20591 19159
rect 20533 19119 20591 19125
rect 20898 19116 20904 19168
rect 20956 19116 20962 19168
rect 22186 19116 22192 19168
rect 22244 19156 22250 19168
rect 22281 19159 22339 19165
rect 22281 19156 22293 19159
rect 22244 19128 22293 19156
rect 22244 19116 22250 19128
rect 22281 19125 22293 19128
rect 22327 19125 22339 19159
rect 22281 19119 22339 19125
rect 1104 19066 23276 19088
rect 1104 19014 8379 19066
rect 8431 19014 8443 19066
rect 8495 19014 8507 19066
rect 8559 19014 8571 19066
rect 8623 19014 15776 19066
rect 15828 19014 15840 19066
rect 15892 19014 15904 19066
rect 15956 19014 15968 19066
rect 16020 19014 23276 19066
rect 1104 18992 23276 19014
rect 2774 18912 2780 18964
rect 2832 18952 2838 18964
rect 2961 18955 3019 18961
rect 2961 18952 2973 18955
rect 2832 18924 2973 18952
rect 2832 18912 2838 18924
rect 2961 18921 2973 18924
rect 3007 18921 3019 18955
rect 2961 18915 3019 18921
rect 3050 18912 3056 18964
rect 3108 18952 3114 18964
rect 3421 18955 3479 18961
rect 3421 18952 3433 18955
rect 3108 18924 3433 18952
rect 3108 18912 3114 18924
rect 3421 18921 3433 18924
rect 3467 18921 3479 18955
rect 3421 18915 3479 18921
rect 3510 18912 3516 18964
rect 3568 18952 3574 18964
rect 3694 18952 3700 18964
rect 3568 18924 3700 18952
rect 3568 18912 3574 18924
rect 3694 18912 3700 18924
rect 3752 18912 3758 18964
rect 4065 18955 4123 18961
rect 4065 18921 4077 18955
rect 4111 18952 4123 18955
rect 5442 18952 5448 18964
rect 4111 18924 5448 18952
rect 4111 18921 4123 18924
rect 4065 18915 4123 18921
rect 5442 18912 5448 18924
rect 5500 18912 5506 18964
rect 5537 18955 5595 18961
rect 5537 18921 5549 18955
rect 5583 18952 5595 18955
rect 5626 18952 5632 18964
rect 5583 18924 5632 18952
rect 5583 18921 5595 18924
rect 5537 18915 5595 18921
rect 5626 18912 5632 18924
rect 5684 18912 5690 18964
rect 13998 18952 14004 18964
rect 6196 18924 13860 18952
rect 13959 18924 14004 18952
rect 1946 18844 1952 18896
rect 2004 18844 2010 18896
rect 5258 18884 5264 18896
rect 3252 18856 5264 18884
rect 1581 18819 1639 18825
rect 1581 18785 1593 18819
rect 1627 18816 1639 18819
rect 1670 18816 1676 18828
rect 1627 18788 1676 18816
rect 1627 18785 1639 18788
rect 1581 18779 1639 18785
rect 1670 18776 1676 18788
rect 1728 18776 1734 18828
rect 1848 18819 1906 18825
rect 1848 18785 1860 18819
rect 1894 18816 1906 18819
rect 1964 18816 1992 18844
rect 3050 18816 3056 18828
rect 1894 18788 3056 18816
rect 1894 18785 1906 18788
rect 1848 18779 1906 18785
rect 3050 18776 3056 18788
rect 3108 18776 3114 18828
rect 3252 18825 3280 18856
rect 5258 18844 5264 18856
rect 5316 18844 5322 18896
rect 3237 18819 3295 18825
rect 3237 18785 3249 18819
rect 3283 18785 3295 18819
rect 3237 18779 3295 18785
rect 3510 18776 3516 18828
rect 3568 18816 3574 18828
rect 4433 18819 4491 18825
rect 4433 18816 4445 18819
rect 3568 18788 4445 18816
rect 3568 18776 3574 18788
rect 4433 18785 4445 18788
rect 4479 18785 4491 18819
rect 4433 18779 4491 18785
rect 5629 18819 5687 18825
rect 5629 18785 5641 18819
rect 5675 18816 5687 18819
rect 6086 18816 6092 18828
rect 5675 18788 6092 18816
rect 5675 18785 5687 18788
rect 5629 18779 5687 18785
rect 6086 18776 6092 18788
rect 6144 18776 6150 18828
rect 6196 18825 6224 18924
rect 7092 18887 7150 18893
rect 7092 18853 7104 18887
rect 7138 18884 7150 18887
rect 7650 18884 7656 18896
rect 7138 18856 7656 18884
rect 7138 18853 7150 18856
rect 7092 18847 7150 18853
rect 7650 18844 7656 18856
rect 7708 18844 7714 18896
rect 8018 18844 8024 18896
rect 8076 18884 8082 18896
rect 8076 18856 9628 18884
rect 8076 18844 8082 18856
rect 6181 18819 6239 18825
rect 6181 18785 6193 18819
rect 6227 18785 6239 18819
rect 6181 18779 6239 18785
rect 6454 18776 6460 18828
rect 6512 18816 6518 18828
rect 6825 18819 6883 18825
rect 6825 18816 6837 18819
rect 6512 18788 6837 18816
rect 6512 18776 6518 18788
rect 6825 18785 6837 18788
rect 6871 18785 6883 18819
rect 7374 18816 7380 18828
rect 6825 18779 6883 18785
rect 6932 18788 7380 18816
rect 3418 18708 3424 18760
rect 3476 18748 3482 18760
rect 4525 18751 4583 18757
rect 4525 18748 4537 18751
rect 3476 18720 4537 18748
rect 3476 18708 3482 18720
rect 4525 18717 4537 18720
rect 4571 18717 4583 18751
rect 4525 18711 4583 18717
rect 4614 18708 4620 18760
rect 4672 18748 4678 18760
rect 4709 18751 4767 18757
rect 4709 18748 4721 18751
rect 4672 18720 4721 18748
rect 4672 18708 4678 18720
rect 4709 18717 4721 18720
rect 4755 18748 4767 18751
rect 5810 18748 5816 18760
rect 4755 18720 5816 18748
rect 4755 18717 4767 18720
rect 4709 18711 4767 18717
rect 5810 18708 5816 18720
rect 5868 18748 5874 18760
rect 6932 18748 6960 18788
rect 7374 18776 7380 18788
rect 7432 18776 7438 18828
rect 7466 18776 7472 18828
rect 7524 18816 7530 18828
rect 8849 18819 8907 18825
rect 8849 18816 8861 18819
rect 7524 18788 8861 18816
rect 7524 18776 7530 18788
rect 8849 18785 8861 18788
rect 8895 18785 8907 18819
rect 8849 18779 8907 18785
rect 5868 18720 6960 18748
rect 5868 18708 5874 18720
rect 7926 18708 7932 18760
rect 7984 18748 7990 18760
rect 8941 18751 8999 18757
rect 8941 18748 8953 18751
rect 7984 18720 8953 18748
rect 7984 18708 7990 18720
rect 8941 18717 8953 18720
rect 8987 18717 8999 18751
rect 8941 18711 8999 18717
rect 9125 18751 9183 18757
rect 9125 18717 9137 18751
rect 9171 18748 9183 18751
rect 9490 18748 9496 18760
rect 9171 18720 9496 18748
rect 9171 18717 9183 18720
rect 9125 18711 9183 18717
rect 9490 18708 9496 18720
rect 9548 18708 9554 18760
rect 5169 18683 5227 18689
rect 5169 18649 5181 18683
rect 5215 18680 5227 18683
rect 8754 18680 8760 18692
rect 5215 18652 6868 18680
rect 5215 18649 5227 18652
rect 5169 18643 5227 18649
rect 6362 18612 6368 18624
rect 6323 18584 6368 18612
rect 6362 18572 6368 18584
rect 6420 18572 6426 18624
rect 6840 18612 6868 18652
rect 8128 18652 8760 18680
rect 8128 18612 8156 18652
rect 8754 18640 8760 18652
rect 8812 18640 8818 18692
rect 6840 18584 8156 18612
rect 8202 18572 8208 18624
rect 8260 18612 8266 18624
rect 8478 18612 8484 18624
rect 8260 18584 8305 18612
rect 8439 18584 8484 18612
rect 8260 18572 8266 18584
rect 8478 18572 8484 18584
rect 8536 18572 8542 18624
rect 9600 18612 9628 18856
rect 11698 18844 11704 18896
rect 11756 18884 11762 18896
rect 13538 18884 13544 18896
rect 11756 18856 13544 18884
rect 11756 18844 11762 18856
rect 13538 18844 13544 18856
rect 13596 18844 13602 18896
rect 13832 18884 13860 18924
rect 13998 18912 14004 18924
rect 14056 18912 14062 18964
rect 14366 18912 14372 18964
rect 14424 18952 14430 18964
rect 16114 18952 16120 18964
rect 14424 18924 16120 18952
rect 14424 18912 14430 18924
rect 16114 18912 16120 18924
rect 16172 18912 16178 18964
rect 18138 18912 18144 18964
rect 18196 18952 18202 18964
rect 19978 18952 19984 18964
rect 18196 18924 19984 18952
rect 18196 18912 18202 18924
rect 19978 18912 19984 18924
rect 20036 18912 20042 18964
rect 20162 18912 20168 18964
rect 20220 18952 20226 18964
rect 21174 18952 21180 18964
rect 20220 18924 21180 18952
rect 20220 18912 20226 18924
rect 21174 18912 21180 18924
rect 21232 18912 21238 18964
rect 21726 18912 21732 18964
rect 21784 18912 21790 18964
rect 14274 18884 14280 18896
rect 13832 18856 14280 18884
rect 14274 18844 14280 18856
rect 14332 18844 14338 18896
rect 15562 18884 15568 18896
rect 14384 18856 15568 18884
rect 9674 18776 9680 18828
rect 9732 18816 9738 18828
rect 10318 18816 10324 18828
rect 9732 18788 10324 18816
rect 9732 18776 9738 18788
rect 10318 18776 10324 18788
rect 10376 18776 10382 18828
rect 10413 18819 10471 18825
rect 10413 18785 10425 18819
rect 10459 18816 10471 18819
rect 11054 18816 11060 18828
rect 10459 18788 11060 18816
rect 10459 18785 10471 18788
rect 10413 18779 10471 18785
rect 11054 18776 11060 18788
rect 11112 18776 11118 18828
rect 11146 18776 11152 18828
rect 11204 18816 11210 18828
rect 11793 18819 11851 18825
rect 11793 18816 11805 18819
rect 11204 18788 11805 18816
rect 11204 18776 11210 18788
rect 11793 18785 11805 18788
rect 11839 18785 11851 18819
rect 12710 18816 12716 18828
rect 11793 18779 11851 18785
rect 12544 18788 12716 18816
rect 10042 18757 10048 18760
rect 10000 18751 10048 18757
rect 10000 18717 10012 18751
rect 10046 18717 10048 18751
rect 10000 18711 10048 18717
rect 10042 18708 10048 18711
rect 10100 18708 10106 18760
rect 10134 18708 10140 18760
rect 10192 18748 10198 18760
rect 12544 18748 12572 18788
rect 12710 18776 12716 18788
rect 12768 18776 12774 18828
rect 12888 18819 12946 18825
rect 12888 18785 12900 18819
rect 12934 18816 12946 18819
rect 14384 18816 14412 18856
rect 15562 18844 15568 18856
rect 15620 18844 15626 18896
rect 16016 18887 16074 18893
rect 16016 18853 16028 18887
rect 16062 18884 16074 18887
rect 20530 18884 20536 18896
rect 16062 18856 20536 18884
rect 16062 18853 16074 18856
rect 16016 18847 16074 18853
rect 20530 18844 20536 18856
rect 20588 18844 20594 18896
rect 21744 18884 21772 18912
rect 20640 18856 21772 18884
rect 12934 18788 14412 18816
rect 14645 18819 14703 18825
rect 12934 18785 12946 18788
rect 12888 18779 12946 18785
rect 14645 18785 14657 18819
rect 14691 18816 14703 18819
rect 15102 18816 15108 18828
rect 14691 18788 15108 18816
rect 14691 18785 14703 18788
rect 14645 18779 14703 18785
rect 15102 18776 15108 18788
rect 15160 18776 15166 18828
rect 16482 18816 16488 18828
rect 15212 18788 16488 18816
rect 10192 18720 12572 18748
rect 12621 18751 12679 18757
rect 10192 18708 10198 18720
rect 12621 18717 12633 18751
rect 12667 18717 12679 18751
rect 12621 18711 12679 18717
rect 11517 18683 11575 18689
rect 11517 18649 11529 18683
rect 11563 18680 11575 18683
rect 11698 18680 11704 18692
rect 11563 18652 11704 18680
rect 11563 18649 11575 18652
rect 11517 18643 11575 18649
rect 11532 18612 11560 18643
rect 11698 18640 11704 18652
rect 11756 18680 11762 18692
rect 12066 18680 12072 18692
rect 11756 18652 12072 18680
rect 11756 18640 11762 18652
rect 12066 18640 12072 18652
rect 12124 18640 12130 18692
rect 9600 18584 11560 18612
rect 11790 18572 11796 18624
rect 11848 18612 11854 18624
rect 11977 18615 12035 18621
rect 11977 18612 11989 18615
rect 11848 18584 11989 18612
rect 11848 18572 11854 18584
rect 11977 18581 11989 18584
rect 12023 18581 12035 18615
rect 12636 18612 12664 18711
rect 14829 18683 14887 18689
rect 14829 18649 14841 18683
rect 14875 18680 14887 18683
rect 15212 18680 15240 18788
rect 16482 18776 16488 18788
rect 16540 18776 16546 18828
rect 16574 18776 16580 18828
rect 16632 18816 16638 18828
rect 16850 18816 16856 18828
rect 16632 18788 16856 18816
rect 16632 18776 16638 18788
rect 16850 18776 16856 18788
rect 16908 18776 16914 18828
rect 17494 18776 17500 18828
rect 17552 18816 17558 18828
rect 17954 18825 17960 18828
rect 17589 18819 17647 18825
rect 17589 18816 17601 18819
rect 17552 18788 17601 18816
rect 17552 18776 17558 18788
rect 17589 18785 17601 18788
rect 17635 18785 17647 18819
rect 17948 18816 17960 18825
rect 17915 18788 17960 18816
rect 17589 18779 17647 18785
rect 17948 18779 17960 18788
rect 17954 18776 17960 18779
rect 18012 18776 18018 18828
rect 18322 18776 18328 18828
rect 18380 18816 18386 18828
rect 18506 18816 18512 18828
rect 18380 18788 18512 18816
rect 18380 18776 18386 18788
rect 18506 18776 18512 18788
rect 18564 18776 18570 18828
rect 19521 18819 19579 18825
rect 19521 18785 19533 18819
rect 19567 18816 19579 18819
rect 19794 18816 19800 18828
rect 19567 18788 19800 18816
rect 19567 18785 19579 18788
rect 19521 18779 19579 18785
rect 19794 18776 19800 18788
rect 19852 18776 19858 18828
rect 19886 18776 19892 18828
rect 19944 18816 19950 18828
rect 20640 18816 20668 18856
rect 19944 18788 20668 18816
rect 19944 18776 19950 18788
rect 21174 18776 21180 18828
rect 21232 18816 21238 18828
rect 21729 18819 21787 18825
rect 21729 18816 21741 18819
rect 21232 18788 21741 18816
rect 21232 18776 21238 18788
rect 21729 18785 21741 18788
rect 21775 18785 21787 18819
rect 21729 18779 21787 18785
rect 15289 18751 15347 18757
rect 15289 18717 15301 18751
rect 15335 18717 15347 18751
rect 15746 18748 15752 18760
rect 15707 18720 15752 18748
rect 15289 18711 15347 18717
rect 14875 18652 15240 18680
rect 14875 18649 14887 18652
rect 14829 18643 14887 18649
rect 12894 18612 12900 18624
rect 12636 18584 12900 18612
rect 11977 18575 12035 18581
rect 12894 18572 12900 18584
rect 12952 18572 12958 18624
rect 15304 18612 15332 18711
rect 15746 18708 15752 18720
rect 15804 18708 15810 18760
rect 17681 18751 17739 18757
rect 17681 18748 17693 18751
rect 17420 18720 17693 18748
rect 17420 18624 17448 18720
rect 17681 18717 17693 18720
rect 17727 18717 17739 18751
rect 17681 18711 17739 18717
rect 19242 18708 19248 18760
rect 19300 18748 19306 18760
rect 19613 18751 19671 18757
rect 19613 18748 19625 18751
rect 19300 18720 19625 18748
rect 19300 18708 19306 18720
rect 19613 18717 19625 18720
rect 19659 18717 19671 18751
rect 19613 18711 19671 18717
rect 19705 18751 19763 18757
rect 19705 18717 19717 18751
rect 19751 18717 19763 18751
rect 19705 18711 19763 18717
rect 20349 18751 20407 18757
rect 20349 18717 20361 18751
rect 20395 18717 20407 18751
rect 20349 18711 20407 18717
rect 18690 18640 18696 18692
rect 18748 18680 18754 18692
rect 19720 18680 19748 18711
rect 18748 18652 19748 18680
rect 18748 18640 18754 18652
rect 17034 18612 17040 18624
rect 15304 18584 17040 18612
rect 17034 18572 17040 18584
rect 17092 18572 17098 18624
rect 17126 18572 17132 18624
rect 17184 18612 17190 18624
rect 17402 18612 17408 18624
rect 17184 18584 17229 18612
rect 17363 18584 17408 18612
rect 17184 18572 17190 18584
rect 17402 18572 17408 18584
rect 17460 18572 17466 18624
rect 18598 18572 18604 18624
rect 18656 18612 18662 18624
rect 19061 18615 19119 18621
rect 19061 18612 19073 18615
rect 18656 18584 19073 18612
rect 18656 18572 18662 18584
rect 19061 18581 19073 18584
rect 19107 18581 19119 18615
rect 19061 18575 19119 18581
rect 19150 18572 19156 18624
rect 19208 18612 19214 18624
rect 20162 18612 20168 18624
rect 19208 18584 19253 18612
rect 20123 18584 20168 18612
rect 19208 18572 19214 18584
rect 20162 18572 20168 18584
rect 20220 18612 20226 18624
rect 20364 18612 20392 18711
rect 20806 18708 20812 18760
rect 20864 18748 20870 18760
rect 21821 18751 21879 18757
rect 21821 18748 21833 18751
rect 20864 18720 21833 18748
rect 20864 18708 20870 18720
rect 21821 18717 21833 18720
rect 21867 18717 21879 18751
rect 21821 18711 21879 18717
rect 21913 18751 21971 18757
rect 21913 18717 21925 18751
rect 21959 18748 21971 18751
rect 22002 18748 22008 18760
rect 21959 18720 22008 18748
rect 21959 18717 21971 18720
rect 21913 18711 21971 18717
rect 20990 18640 20996 18692
rect 21048 18680 21054 18692
rect 21928 18680 21956 18711
rect 22002 18708 22008 18720
rect 22060 18708 22066 18760
rect 22557 18751 22615 18757
rect 22557 18717 22569 18751
rect 22603 18717 22615 18751
rect 22557 18711 22615 18717
rect 21048 18652 21956 18680
rect 21048 18640 21054 18652
rect 21358 18612 21364 18624
rect 20220 18584 20392 18612
rect 21319 18584 21364 18612
rect 20220 18572 20226 18584
rect 21358 18572 21364 18584
rect 21416 18572 21422 18624
rect 22094 18572 22100 18624
rect 22152 18612 22158 18624
rect 22373 18615 22431 18621
rect 22373 18612 22385 18615
rect 22152 18584 22385 18612
rect 22152 18572 22158 18584
rect 22373 18581 22385 18584
rect 22419 18612 22431 18615
rect 22572 18612 22600 18711
rect 22419 18584 22600 18612
rect 22419 18581 22431 18584
rect 22373 18575 22431 18581
rect 1104 18522 23276 18544
rect 1104 18470 4680 18522
rect 4732 18470 4744 18522
rect 4796 18470 4808 18522
rect 4860 18470 4872 18522
rect 4924 18470 12078 18522
rect 12130 18470 12142 18522
rect 12194 18470 12206 18522
rect 12258 18470 12270 18522
rect 12322 18470 19475 18522
rect 19527 18470 19539 18522
rect 19591 18470 19603 18522
rect 19655 18470 19667 18522
rect 19719 18470 23276 18522
rect 1104 18448 23276 18470
rect 3050 18408 3056 18420
rect 3011 18380 3056 18408
rect 3050 18368 3056 18380
rect 3108 18368 3114 18420
rect 5261 18411 5319 18417
rect 5261 18377 5273 18411
rect 5307 18408 5319 18411
rect 8846 18408 8852 18420
rect 5307 18380 8852 18408
rect 5307 18377 5319 18380
rect 5261 18371 5319 18377
rect 8846 18368 8852 18380
rect 8904 18368 8910 18420
rect 9122 18408 9128 18420
rect 9083 18380 9128 18408
rect 9122 18368 9128 18380
rect 9180 18368 9186 18420
rect 9401 18411 9459 18417
rect 9401 18377 9413 18411
rect 9447 18408 9459 18411
rect 11514 18408 11520 18420
rect 9447 18380 11520 18408
rect 9447 18377 9459 18380
rect 9401 18371 9459 18377
rect 11514 18368 11520 18380
rect 11572 18368 11578 18420
rect 14277 18411 14335 18417
rect 14277 18377 14289 18411
rect 14323 18408 14335 18411
rect 15562 18408 15568 18420
rect 14323 18380 15568 18408
rect 14323 18377 14335 18380
rect 14277 18371 14335 18377
rect 15562 18368 15568 18380
rect 15620 18368 15626 18420
rect 17497 18411 17555 18417
rect 15672 18380 17448 18408
rect 4982 18300 4988 18352
rect 5040 18340 5046 18352
rect 6546 18340 6552 18352
rect 5040 18312 6552 18340
rect 5040 18300 5046 18312
rect 6546 18300 6552 18312
rect 6604 18300 6610 18352
rect 5810 18272 5816 18284
rect 5771 18244 5816 18272
rect 5810 18232 5816 18244
rect 5868 18232 5874 18284
rect 7098 18232 7104 18284
rect 7156 18272 7162 18284
rect 7650 18281 7656 18284
rect 7285 18275 7343 18281
rect 7285 18272 7297 18275
rect 7156 18244 7297 18272
rect 7156 18232 7162 18244
rect 7285 18241 7297 18244
rect 7331 18241 7343 18275
rect 7285 18235 7343 18241
rect 7608 18275 7656 18281
rect 7608 18241 7620 18275
rect 7654 18241 7656 18275
rect 7608 18235 7656 18241
rect 7650 18232 7656 18235
rect 7708 18232 7714 18284
rect 7791 18275 7849 18281
rect 7791 18241 7803 18275
rect 7837 18272 7849 18275
rect 9140 18272 9168 18368
rect 11885 18343 11943 18349
rect 11885 18309 11897 18343
rect 11931 18340 11943 18343
rect 12894 18340 12900 18352
rect 11931 18312 12900 18340
rect 11931 18309 11943 18312
rect 11885 18303 11943 18309
rect 12894 18300 12900 18312
rect 12952 18300 12958 18352
rect 14553 18343 14611 18349
rect 14553 18309 14565 18343
rect 14599 18340 14611 18343
rect 15672 18340 15700 18380
rect 14599 18312 15700 18340
rect 17420 18340 17448 18380
rect 17497 18377 17509 18411
rect 17543 18408 17555 18411
rect 18782 18408 18788 18420
rect 17543 18380 18788 18408
rect 17543 18377 17555 18380
rect 17497 18371 17555 18377
rect 18782 18368 18788 18380
rect 18840 18368 18846 18420
rect 18874 18368 18880 18420
rect 18932 18408 18938 18420
rect 19242 18408 19248 18420
rect 18932 18380 19248 18408
rect 18932 18368 18938 18380
rect 19242 18368 19248 18380
rect 19300 18368 19306 18420
rect 20346 18408 20352 18420
rect 19536 18380 20352 18408
rect 19536 18352 19564 18380
rect 20346 18368 20352 18380
rect 20404 18368 20410 18420
rect 17420 18312 18558 18340
rect 14599 18309 14611 18312
rect 14553 18303 14611 18309
rect 9861 18275 9919 18281
rect 9861 18272 9873 18275
rect 7837 18244 9076 18272
rect 9140 18244 9873 18272
rect 7837 18241 7849 18244
rect 7791 18235 7849 18241
rect 1673 18207 1731 18213
rect 1673 18173 1685 18207
rect 1719 18204 1731 18207
rect 1762 18204 1768 18216
rect 1719 18176 1768 18204
rect 1719 18173 1731 18176
rect 1673 18167 1731 18173
rect 1762 18164 1768 18176
rect 1820 18164 1826 18216
rect 3326 18204 3332 18216
rect 3287 18176 3332 18204
rect 3326 18164 3332 18176
rect 3384 18164 3390 18216
rect 3596 18207 3654 18213
rect 3596 18173 3608 18207
rect 3642 18204 3654 18207
rect 4062 18204 4068 18216
rect 3642 18176 4068 18204
rect 3642 18173 3654 18176
rect 3596 18167 3654 18173
rect 4062 18164 4068 18176
rect 4120 18164 4126 18216
rect 4522 18164 4528 18216
rect 4580 18204 4586 18216
rect 6914 18204 6920 18216
rect 4580 18176 6920 18204
rect 4580 18164 4586 18176
rect 6914 18164 6920 18176
rect 6972 18164 6978 18216
rect 8018 18204 8024 18216
rect 7979 18176 8024 18204
rect 8018 18164 8024 18176
rect 8076 18164 8082 18216
rect 8110 18164 8116 18216
rect 8168 18204 8174 18216
rect 9048 18204 9076 18244
rect 9861 18241 9873 18244
rect 9907 18241 9919 18275
rect 9861 18235 9919 18241
rect 9953 18275 10011 18281
rect 9953 18241 9965 18275
rect 9999 18241 10011 18275
rect 9953 18235 10011 18241
rect 9674 18204 9680 18216
rect 8168 18176 8708 18204
rect 9048 18176 9680 18204
rect 8168 18164 8174 18176
rect 1940 18139 1998 18145
rect 1940 18105 1952 18139
rect 1986 18136 1998 18139
rect 3142 18136 3148 18148
rect 1986 18108 3148 18136
rect 1986 18105 1998 18108
rect 1940 18099 1998 18105
rect 3142 18096 3148 18108
rect 3200 18096 3206 18148
rect 5166 18096 5172 18148
rect 5224 18136 5230 18148
rect 5718 18136 5724 18148
rect 5224 18108 5724 18136
rect 5224 18096 5230 18108
rect 5718 18096 5724 18108
rect 5776 18096 5782 18148
rect 6273 18139 6331 18145
rect 6273 18105 6285 18139
rect 6319 18136 6331 18139
rect 8680 18136 8708 18176
rect 9674 18164 9680 18176
rect 9732 18164 9738 18216
rect 9766 18164 9772 18216
rect 9824 18204 9830 18216
rect 9824 18176 9869 18204
rect 9824 18164 9830 18176
rect 9968 18136 9996 18235
rect 14918 18232 14924 18284
rect 14976 18272 14982 18284
rect 15013 18275 15071 18281
rect 15013 18272 15025 18275
rect 14976 18244 15025 18272
rect 14976 18232 14982 18244
rect 15013 18241 15025 18244
rect 15059 18241 15071 18275
rect 15194 18272 15200 18284
rect 15155 18244 15200 18272
rect 15013 18235 15071 18241
rect 15194 18232 15200 18244
rect 15252 18232 15258 18284
rect 16022 18281 16028 18284
rect 15980 18275 16028 18281
rect 15980 18272 15992 18275
rect 15304 18244 15992 18272
rect 10502 18204 10508 18216
rect 10463 18176 10508 18204
rect 10502 18164 10508 18176
rect 10560 18164 10566 18216
rect 10704 18176 12020 18204
rect 6319 18108 7420 18136
rect 8680 18108 9996 18136
rect 6319 18105 6331 18108
rect 6273 18099 6331 18105
rect 3878 18028 3884 18080
rect 3936 18068 3942 18080
rect 4709 18071 4767 18077
rect 4709 18068 4721 18071
rect 3936 18040 4721 18068
rect 3936 18028 3942 18040
rect 4709 18037 4721 18040
rect 4755 18037 4767 18071
rect 5626 18068 5632 18080
rect 5587 18040 5632 18068
rect 4709 18031 4767 18037
rect 5626 18028 5632 18040
rect 5684 18028 5690 18080
rect 6825 18071 6883 18077
rect 6825 18037 6837 18071
rect 6871 18068 6883 18071
rect 7098 18068 7104 18080
rect 6871 18040 7104 18068
rect 6871 18037 6883 18040
rect 6825 18031 6883 18037
rect 7098 18028 7104 18040
rect 7156 18028 7162 18080
rect 7392 18068 7420 18108
rect 10042 18096 10048 18148
rect 10100 18136 10106 18148
rect 10704 18136 10732 18176
rect 10100 18108 10732 18136
rect 10772 18139 10830 18145
rect 10100 18096 10106 18108
rect 10772 18105 10784 18139
rect 10818 18136 10830 18139
rect 11238 18136 11244 18148
rect 10818 18108 11244 18136
rect 10818 18105 10830 18108
rect 10772 18099 10830 18105
rect 11238 18096 11244 18108
rect 11296 18096 11302 18148
rect 11992 18136 12020 18176
rect 12802 18164 12808 18216
rect 12860 18204 12866 18216
rect 12897 18207 12955 18213
rect 12897 18204 12909 18207
rect 12860 18176 12909 18204
rect 12860 18164 12866 18176
rect 12897 18173 12909 18176
rect 12943 18173 12955 18207
rect 12897 18167 12955 18173
rect 13164 18207 13222 18213
rect 13164 18173 13176 18207
rect 13210 18204 13222 18207
rect 14366 18204 14372 18216
rect 13210 18176 14372 18204
rect 13210 18173 13222 18176
rect 13164 18167 13222 18173
rect 14366 18164 14372 18176
rect 14424 18164 14430 18216
rect 15304 18204 15332 18244
rect 15980 18241 15992 18244
rect 16026 18241 16028 18275
rect 15980 18235 16028 18241
rect 16022 18232 16028 18235
rect 16080 18272 16086 18284
rect 16163 18275 16221 18281
rect 16080 18244 16128 18272
rect 16080 18232 16086 18244
rect 16163 18241 16175 18275
rect 16209 18272 16221 18275
rect 17862 18272 17868 18284
rect 16209 18244 17868 18272
rect 16209 18241 16221 18244
rect 16163 18235 16221 18241
rect 17862 18232 17868 18244
rect 17920 18232 17926 18284
rect 18046 18272 18052 18284
rect 18007 18244 18052 18272
rect 18046 18232 18052 18244
rect 18104 18232 18110 18284
rect 18530 18272 18558 18312
rect 19518 18300 19524 18352
rect 19576 18300 19582 18352
rect 18530 18244 18644 18272
rect 14476 18176 15332 18204
rect 15657 18207 15715 18213
rect 14476 18136 14504 18176
rect 15657 18173 15669 18207
rect 15703 18173 15715 18207
rect 15657 18167 15715 18173
rect 16393 18207 16451 18213
rect 16393 18173 16405 18207
rect 16439 18204 16451 18207
rect 16482 18204 16488 18216
rect 16439 18176 16488 18204
rect 16439 18173 16451 18176
rect 16393 18167 16451 18173
rect 11992 18108 14504 18136
rect 14921 18139 14979 18145
rect 14921 18105 14933 18139
rect 14967 18136 14979 18139
rect 15562 18136 15568 18148
rect 14967 18108 15568 18136
rect 14967 18105 14979 18108
rect 14921 18099 14979 18105
rect 15562 18096 15568 18108
rect 15620 18096 15626 18148
rect 11882 18068 11888 18080
rect 7392 18040 11888 18068
rect 11882 18028 11888 18040
rect 11940 18028 11946 18080
rect 12434 18028 12440 18080
rect 12492 18068 12498 18080
rect 12492 18040 12537 18068
rect 12492 18028 12498 18040
rect 12802 18028 12808 18080
rect 12860 18068 12866 18080
rect 15672 18068 15700 18167
rect 16482 18164 16488 18176
rect 16540 18204 16546 18216
rect 18506 18204 18512 18216
rect 16540 18176 17080 18204
rect 18419 18176 18512 18204
rect 16540 18164 16546 18176
rect 12860 18040 15700 18068
rect 17052 18068 17080 18176
rect 18506 18164 18512 18176
rect 18564 18164 18570 18216
rect 18616 18204 18644 18244
rect 21910 18232 21916 18284
rect 21968 18272 21974 18284
rect 22465 18275 22523 18281
rect 22465 18272 22477 18275
rect 21968 18244 22477 18272
rect 21968 18232 21974 18244
rect 22465 18241 22477 18244
rect 22511 18241 22523 18275
rect 22465 18235 22523 18241
rect 20070 18204 20076 18216
rect 18616 18176 20076 18204
rect 20070 18164 20076 18176
rect 20128 18164 20134 18216
rect 20165 18207 20223 18213
rect 20165 18173 20177 18207
rect 20211 18204 20223 18207
rect 20898 18204 20904 18216
rect 20211 18176 20904 18204
rect 20211 18173 20223 18176
rect 20165 18167 20223 18173
rect 20898 18164 20904 18176
rect 20956 18164 20962 18216
rect 17402 18096 17408 18148
rect 17460 18136 17466 18148
rect 18046 18136 18052 18148
rect 17460 18108 18052 18136
rect 17460 18096 17466 18108
rect 18046 18096 18052 18108
rect 18104 18136 18110 18148
rect 18524 18136 18552 18164
rect 18104 18108 18552 18136
rect 18776 18139 18834 18145
rect 18104 18096 18110 18108
rect 18776 18105 18788 18139
rect 18822 18136 18834 18139
rect 19150 18136 19156 18148
rect 18822 18108 19156 18136
rect 18822 18105 18834 18108
rect 18776 18099 18834 18105
rect 19150 18096 19156 18108
rect 19208 18096 19214 18148
rect 20346 18136 20352 18148
rect 19904 18108 20352 18136
rect 19242 18068 19248 18080
rect 17052 18040 19248 18068
rect 12860 18028 12866 18040
rect 19242 18028 19248 18040
rect 19300 18028 19306 18080
rect 19904 18077 19932 18108
rect 20346 18096 20352 18108
rect 20404 18145 20410 18148
rect 20404 18139 20468 18145
rect 20404 18105 20422 18139
rect 20456 18105 20468 18139
rect 20404 18099 20468 18105
rect 20404 18096 20410 18099
rect 19889 18071 19947 18077
rect 19889 18037 19901 18071
rect 19935 18037 19947 18071
rect 19889 18031 19947 18037
rect 21545 18071 21603 18077
rect 21545 18037 21557 18071
rect 21591 18068 21603 18071
rect 21634 18068 21640 18080
rect 21591 18040 21640 18068
rect 21591 18037 21603 18040
rect 21545 18031 21603 18037
rect 21634 18028 21640 18040
rect 21692 18028 21698 18080
rect 21913 18071 21971 18077
rect 21913 18037 21925 18071
rect 21959 18068 21971 18071
rect 22002 18068 22008 18080
rect 21959 18040 22008 18068
rect 21959 18037 21971 18040
rect 21913 18031 21971 18037
rect 22002 18028 22008 18040
rect 22060 18028 22066 18080
rect 22278 18068 22284 18080
rect 22239 18040 22284 18068
rect 22278 18028 22284 18040
rect 22336 18028 22342 18080
rect 22370 18028 22376 18080
rect 22428 18068 22434 18080
rect 22428 18040 22473 18068
rect 22428 18028 22434 18040
rect 1104 17978 23276 18000
rect 1104 17926 8379 17978
rect 8431 17926 8443 17978
rect 8495 17926 8507 17978
rect 8559 17926 8571 17978
rect 8623 17926 15776 17978
rect 15828 17926 15840 17978
rect 15892 17926 15904 17978
rect 15956 17926 15968 17978
rect 16020 17926 23276 17978
rect 1104 17904 23276 17926
rect 3142 17864 3148 17876
rect 3103 17836 3148 17864
rect 3142 17824 3148 17836
rect 3200 17824 3206 17876
rect 3602 17864 3608 17876
rect 3563 17836 3608 17864
rect 3602 17824 3608 17836
rect 3660 17824 3666 17876
rect 4246 17864 4252 17876
rect 4207 17836 4252 17864
rect 4246 17824 4252 17836
rect 4304 17824 4310 17876
rect 5258 17824 5264 17876
rect 5316 17864 5322 17876
rect 7466 17864 7472 17876
rect 5316 17836 7472 17864
rect 5316 17824 5322 17836
rect 7466 17824 7472 17836
rect 7524 17824 7530 17876
rect 7558 17824 7564 17876
rect 7616 17864 7622 17876
rect 8113 17867 8171 17873
rect 8113 17864 8125 17867
rect 7616 17836 8125 17864
rect 7616 17824 7622 17836
rect 8113 17833 8125 17836
rect 8159 17833 8171 17867
rect 8846 17864 8852 17876
rect 8807 17836 8852 17864
rect 8113 17827 8171 17833
rect 8846 17824 8852 17836
rect 8904 17824 8910 17876
rect 9677 17867 9735 17873
rect 9677 17833 9689 17867
rect 9723 17864 9735 17867
rect 10502 17864 10508 17876
rect 9723 17836 10508 17864
rect 9723 17833 9735 17836
rect 9677 17827 9735 17833
rect 10502 17824 10508 17836
rect 10560 17824 10566 17876
rect 10594 17824 10600 17876
rect 10652 17864 10658 17876
rect 11422 17864 11428 17876
rect 10652 17836 11284 17864
rect 11383 17836 11428 17864
rect 10652 17824 10658 17836
rect 2032 17799 2090 17805
rect 2032 17765 2044 17799
rect 2078 17796 2090 17799
rect 3878 17796 3884 17808
rect 2078 17768 3884 17796
rect 2078 17765 2090 17768
rect 2032 17759 2090 17765
rect 3878 17756 3884 17768
rect 3936 17756 3942 17808
rect 8754 17796 8760 17808
rect 8715 17768 8760 17796
rect 8754 17756 8760 17768
rect 8812 17756 8818 17808
rect 9858 17796 9864 17808
rect 8864 17768 9864 17796
rect 1765 17731 1823 17737
rect 1765 17697 1777 17731
rect 1811 17728 1823 17731
rect 1854 17728 1860 17740
rect 1811 17700 1860 17728
rect 1811 17697 1823 17700
rect 1765 17691 1823 17697
rect 1854 17688 1860 17700
rect 1912 17688 1918 17740
rect 3421 17731 3479 17737
rect 3421 17697 3433 17731
rect 3467 17728 3479 17731
rect 3786 17728 3792 17740
rect 3467 17700 3792 17728
rect 3467 17697 3479 17700
rect 3421 17691 3479 17697
rect 3786 17688 3792 17700
rect 3844 17688 3850 17740
rect 4065 17731 4123 17737
rect 4065 17697 4077 17731
rect 4111 17728 4123 17731
rect 4890 17728 4896 17740
rect 4111 17700 4896 17728
rect 4111 17697 4123 17700
rect 4065 17691 4123 17697
rect 4890 17688 4896 17700
rect 4948 17688 4954 17740
rect 5252 17731 5310 17737
rect 5252 17697 5264 17731
rect 5298 17728 5310 17731
rect 7000 17731 7058 17737
rect 5298 17700 6592 17728
rect 5298 17697 5310 17700
rect 5252 17691 5310 17697
rect 3326 17620 3332 17672
rect 3384 17660 3390 17672
rect 4985 17663 5043 17669
rect 4985 17660 4997 17663
rect 3384 17632 4997 17660
rect 3384 17620 3390 17632
rect 4985 17629 4997 17632
rect 5031 17629 5043 17663
rect 4985 17623 5043 17629
rect 1762 17484 1768 17536
rect 1820 17524 1826 17536
rect 5258 17524 5264 17536
rect 1820 17496 5264 17524
rect 1820 17484 1826 17496
rect 5258 17484 5264 17496
rect 5316 17484 5322 17536
rect 5718 17484 5724 17536
rect 5776 17524 5782 17536
rect 6365 17527 6423 17533
rect 6365 17524 6377 17527
rect 5776 17496 6377 17524
rect 5776 17484 5782 17496
rect 6365 17493 6377 17496
rect 6411 17493 6423 17527
rect 6564 17524 6592 17700
rect 7000 17697 7012 17731
rect 7046 17728 7058 17731
rect 8110 17728 8116 17740
rect 7046 17700 8116 17728
rect 7046 17697 7058 17700
rect 7000 17691 7058 17697
rect 8110 17688 8116 17700
rect 8168 17688 8174 17740
rect 6638 17620 6644 17672
rect 6696 17660 6702 17672
rect 6733 17663 6791 17669
rect 6733 17660 6745 17663
rect 6696 17632 6745 17660
rect 6696 17620 6702 17632
rect 6733 17629 6745 17632
rect 6779 17629 6791 17663
rect 6733 17623 6791 17629
rect 7742 17620 7748 17672
rect 7800 17660 7806 17672
rect 8864 17660 8892 17768
rect 9858 17756 9864 17768
rect 9916 17756 9922 17808
rect 11146 17796 11152 17808
rect 9968 17768 11152 17796
rect 9122 17688 9128 17740
rect 9180 17728 9186 17740
rect 9968 17728 9996 17768
rect 11146 17756 11152 17768
rect 11204 17756 11210 17808
rect 11256 17796 11284 17836
rect 11422 17824 11428 17836
rect 11480 17824 11486 17876
rect 11793 17867 11851 17873
rect 11793 17833 11805 17867
rect 11839 17864 11851 17867
rect 12434 17864 12440 17876
rect 11839 17836 12440 17864
rect 11839 17833 11851 17836
rect 11793 17827 11851 17833
rect 12434 17824 12440 17836
rect 12492 17824 12498 17876
rect 14182 17864 14188 17876
rect 13188 17836 14188 17864
rect 13188 17796 13216 17836
rect 14182 17824 14188 17836
rect 14240 17824 14246 17876
rect 14366 17864 14372 17876
rect 14327 17836 14372 17864
rect 14366 17824 14372 17836
rect 14424 17824 14430 17876
rect 14829 17867 14887 17873
rect 14829 17833 14841 17867
rect 14875 17864 14887 17867
rect 15378 17864 15384 17876
rect 14875 17836 15384 17864
rect 14875 17833 14887 17836
rect 14829 17827 14887 17833
rect 15378 17824 15384 17836
rect 15436 17824 15442 17876
rect 16669 17867 16727 17873
rect 16669 17833 16681 17867
rect 16715 17833 16727 17867
rect 16669 17827 16727 17833
rect 11256 17768 13216 17796
rect 13256 17799 13314 17805
rect 13256 17765 13268 17799
rect 13302 17796 13314 17799
rect 13302 17768 14872 17796
rect 13302 17765 13314 17768
rect 13256 17759 13314 17765
rect 14844 17740 14872 17768
rect 14918 17756 14924 17808
rect 14976 17796 14982 17808
rect 15194 17796 15200 17808
rect 14976 17768 15200 17796
rect 14976 17756 14982 17768
rect 15194 17756 15200 17768
rect 15252 17756 15258 17808
rect 15286 17756 15292 17808
rect 15344 17796 15350 17808
rect 15534 17799 15592 17805
rect 15534 17796 15546 17799
rect 15344 17768 15546 17796
rect 15344 17756 15350 17768
rect 15534 17765 15546 17768
rect 15580 17765 15592 17799
rect 15534 17759 15592 17765
rect 9180 17700 9996 17728
rect 10036 17731 10094 17737
rect 9180 17688 9186 17700
rect 10036 17697 10048 17731
rect 10082 17728 10094 17731
rect 11054 17728 11060 17740
rect 10082 17700 11060 17728
rect 10082 17697 10094 17700
rect 10036 17691 10094 17697
rect 11054 17688 11060 17700
rect 11112 17688 11118 17740
rect 11885 17731 11943 17737
rect 11885 17697 11897 17731
rect 11931 17728 11943 17731
rect 12437 17731 12495 17737
rect 11931 17700 12204 17728
rect 11931 17697 11943 17700
rect 11885 17691 11943 17697
rect 7800 17632 8892 17660
rect 7800 17620 7806 17632
rect 8938 17620 8944 17672
rect 8996 17660 9002 17672
rect 9033 17663 9091 17669
rect 9033 17660 9045 17663
rect 8996 17632 9045 17660
rect 8996 17620 9002 17632
rect 9033 17629 9045 17632
rect 9079 17660 9091 17663
rect 9306 17660 9312 17672
rect 9079 17632 9312 17660
rect 9079 17629 9091 17632
rect 9033 17623 9091 17629
rect 9306 17620 9312 17632
rect 9364 17620 9370 17672
rect 9490 17620 9496 17672
rect 9548 17660 9554 17672
rect 9677 17663 9735 17669
rect 9677 17660 9689 17663
rect 9548 17632 9689 17660
rect 9548 17620 9554 17632
rect 9677 17629 9689 17632
rect 9723 17660 9735 17663
rect 9769 17663 9827 17669
rect 9769 17660 9781 17663
rect 9723 17632 9781 17660
rect 9723 17629 9735 17632
rect 9677 17623 9735 17629
rect 9769 17629 9781 17632
rect 9815 17629 9827 17663
rect 11974 17660 11980 17672
rect 9769 17623 9827 17629
rect 10796 17632 11980 17660
rect 8220 17564 9812 17592
rect 8220 17524 8248 17564
rect 8386 17524 8392 17536
rect 6564 17496 8248 17524
rect 8347 17496 8392 17524
rect 6365 17487 6423 17493
rect 8386 17484 8392 17496
rect 8444 17484 8450 17536
rect 9784 17524 9812 17564
rect 10796 17524 10824 17632
rect 11974 17620 11980 17632
rect 12032 17620 12038 17672
rect 12176 17660 12204 17700
rect 12437 17697 12449 17731
rect 12483 17728 12495 17731
rect 12526 17728 12532 17740
rect 12483 17700 12532 17728
rect 12483 17697 12495 17700
rect 12437 17691 12495 17697
rect 12526 17688 12532 17700
rect 12584 17688 12590 17740
rect 13078 17728 13084 17740
rect 12912 17700 13084 17728
rect 12912 17660 12940 17700
rect 13078 17688 13084 17700
rect 13136 17688 13142 17740
rect 13814 17688 13820 17740
rect 13872 17728 13878 17740
rect 14642 17728 14648 17740
rect 13872 17700 14044 17728
rect 14603 17700 14648 17728
rect 13872 17688 13878 17700
rect 12176 17632 12940 17660
rect 12989 17663 13047 17669
rect 12989 17629 13001 17663
rect 13035 17629 13047 17663
rect 14016 17660 14044 17700
rect 14642 17688 14648 17700
rect 14700 17688 14706 17740
rect 14826 17688 14832 17740
rect 14884 17728 14890 17740
rect 16684 17728 16712 17827
rect 17034 17824 17040 17876
rect 17092 17864 17098 17876
rect 19334 17864 19340 17876
rect 17092 17836 19340 17864
rect 17092 17824 17098 17836
rect 19334 17824 19340 17836
rect 19392 17824 19398 17876
rect 20254 17864 20260 17876
rect 20215 17836 20260 17864
rect 20254 17824 20260 17836
rect 20312 17824 20318 17876
rect 21450 17824 21456 17876
rect 21508 17864 21514 17876
rect 22281 17867 22339 17873
rect 22281 17864 22293 17867
rect 21508 17836 22293 17864
rect 21508 17824 21514 17836
rect 22281 17833 22293 17836
rect 22327 17833 22339 17867
rect 22281 17827 22339 17833
rect 16758 17756 16764 17808
rect 16816 17796 16822 17808
rect 18408 17799 18466 17805
rect 16816 17768 18368 17796
rect 16816 17756 16822 17768
rect 14884 17700 16712 17728
rect 14884 17688 14890 17700
rect 16850 17688 16856 17740
rect 16908 17728 16914 17740
rect 17034 17728 17040 17740
rect 16908 17700 17040 17728
rect 16908 17688 16914 17700
rect 17034 17688 17040 17700
rect 17092 17688 17098 17740
rect 17310 17728 17316 17740
rect 17271 17700 17316 17728
rect 17310 17688 17316 17700
rect 17368 17688 17374 17740
rect 18340 17728 18368 17768
rect 18408 17765 18420 17799
rect 18454 17796 18466 17799
rect 18598 17796 18604 17808
rect 18454 17768 18604 17796
rect 18454 17765 18466 17768
rect 18408 17759 18466 17765
rect 18598 17756 18604 17768
rect 18656 17756 18662 17808
rect 18782 17756 18788 17808
rect 18840 17796 18846 17808
rect 19058 17796 19064 17808
rect 18840 17768 19064 17796
rect 18840 17756 18846 17768
rect 19058 17756 19064 17768
rect 19116 17756 19122 17808
rect 20990 17796 20996 17808
rect 20088 17768 20996 17796
rect 20088 17728 20116 17768
rect 20990 17756 20996 17768
rect 21048 17756 21054 17808
rect 21082 17756 21088 17808
rect 21140 17805 21146 17808
rect 21140 17799 21204 17805
rect 21140 17765 21158 17799
rect 21192 17796 21204 17799
rect 22186 17796 22192 17808
rect 21192 17768 22192 17796
rect 21192 17765 21204 17768
rect 21140 17759 21204 17765
rect 21140 17756 21146 17759
rect 22186 17756 22192 17768
rect 22244 17756 22250 17808
rect 18340 17700 20116 17728
rect 20165 17731 20223 17737
rect 20165 17697 20177 17731
rect 20211 17697 20223 17731
rect 20165 17691 20223 17697
rect 14016 17632 14596 17660
rect 12989 17623 13047 17629
rect 12526 17552 12532 17604
rect 12584 17592 12590 17604
rect 12621 17595 12679 17601
rect 12621 17592 12633 17595
rect 12584 17564 12633 17592
rect 12584 17552 12590 17564
rect 12621 17561 12633 17564
rect 12667 17561 12679 17595
rect 12621 17555 12679 17561
rect 12710 17552 12716 17604
rect 12768 17592 12774 17604
rect 12894 17592 12900 17604
rect 12768 17564 12900 17592
rect 12768 17552 12774 17564
rect 12894 17552 12900 17564
rect 12952 17592 12958 17604
rect 13004 17592 13032 17623
rect 12952 17564 13032 17592
rect 14568 17592 14596 17632
rect 15102 17620 15108 17672
rect 15160 17660 15166 17672
rect 15289 17663 15347 17669
rect 15289 17660 15301 17663
rect 15160 17632 15301 17660
rect 15160 17620 15166 17632
rect 15289 17629 15301 17632
rect 15335 17629 15347 17663
rect 15289 17623 15347 17629
rect 16390 17620 16396 17672
rect 16448 17660 16454 17672
rect 17405 17663 17463 17669
rect 17405 17660 17417 17663
rect 16448 17632 17417 17660
rect 16448 17620 16454 17632
rect 17405 17629 17417 17632
rect 17451 17629 17463 17663
rect 17586 17660 17592 17672
rect 17547 17632 17592 17660
rect 17405 17623 17463 17629
rect 17586 17620 17592 17632
rect 17644 17620 17650 17672
rect 18046 17620 18052 17672
rect 18104 17660 18110 17672
rect 18141 17663 18199 17669
rect 18141 17660 18153 17663
rect 18104 17632 18153 17660
rect 18104 17620 18110 17632
rect 18141 17629 18153 17632
rect 18187 17629 18199 17663
rect 18141 17623 18199 17629
rect 19242 17620 19248 17672
rect 19300 17660 19306 17672
rect 20180 17660 20208 17691
rect 19300 17632 20208 17660
rect 20441 17663 20499 17669
rect 19300 17620 19306 17632
rect 20441 17629 20453 17663
rect 20487 17660 20499 17663
rect 20530 17660 20536 17672
rect 20487 17632 20536 17660
rect 20487 17629 20499 17632
rect 20441 17623 20499 17629
rect 20530 17620 20536 17632
rect 20588 17620 20594 17672
rect 20898 17660 20904 17672
rect 20859 17632 20904 17660
rect 20898 17620 20904 17632
rect 20956 17620 20962 17672
rect 22557 17663 22615 17669
rect 22557 17629 22569 17663
rect 22603 17660 22615 17663
rect 22830 17660 22836 17672
rect 22603 17632 22836 17660
rect 22603 17629 22615 17632
rect 22557 17623 22615 17629
rect 22830 17620 22836 17632
rect 22888 17620 22894 17672
rect 14568 17564 15240 17592
rect 12952 17552 12958 17564
rect 9784 17496 10824 17524
rect 11149 17527 11207 17533
rect 11149 17493 11161 17527
rect 11195 17524 11207 17527
rect 11238 17524 11244 17536
rect 11195 17496 11244 17524
rect 11195 17493 11207 17496
rect 11149 17487 11207 17493
rect 11238 17484 11244 17496
rect 11296 17484 11302 17536
rect 13004 17524 13032 17564
rect 13722 17524 13728 17536
rect 13004 17496 13728 17524
rect 13722 17484 13728 17496
rect 13780 17484 13786 17536
rect 15212 17524 15240 17564
rect 16224 17564 17540 17592
rect 16224 17524 16252 17564
rect 15212 17496 16252 17524
rect 16945 17527 17003 17533
rect 16945 17493 16957 17527
rect 16991 17524 17003 17527
rect 17402 17524 17408 17536
rect 16991 17496 17408 17524
rect 16991 17493 17003 17496
rect 16945 17487 17003 17493
rect 17402 17484 17408 17496
rect 17460 17484 17466 17536
rect 17512 17524 17540 17564
rect 19076 17564 20300 17592
rect 19076 17524 19104 17564
rect 17512 17496 19104 17524
rect 19150 17484 19156 17536
rect 19208 17524 19214 17536
rect 19521 17527 19579 17533
rect 19521 17524 19533 17527
rect 19208 17496 19533 17524
rect 19208 17484 19214 17496
rect 19521 17493 19533 17496
rect 19567 17493 19579 17527
rect 19521 17487 19579 17493
rect 19797 17527 19855 17533
rect 19797 17493 19809 17527
rect 19843 17524 19855 17527
rect 20162 17524 20168 17536
rect 19843 17496 20168 17524
rect 19843 17493 19855 17496
rect 19797 17487 19855 17493
rect 20162 17484 20168 17496
rect 20220 17484 20226 17536
rect 20272 17524 20300 17564
rect 22738 17524 22744 17536
rect 20272 17496 22744 17524
rect 22738 17484 22744 17496
rect 22796 17484 22802 17536
rect 1104 17434 23276 17456
rect 1104 17382 4680 17434
rect 4732 17382 4744 17434
rect 4796 17382 4808 17434
rect 4860 17382 4872 17434
rect 4924 17382 12078 17434
rect 12130 17382 12142 17434
rect 12194 17382 12206 17434
rect 12258 17382 12270 17434
rect 12322 17382 19475 17434
rect 19527 17382 19539 17434
rect 19591 17382 19603 17434
rect 19655 17382 19667 17434
rect 19719 17382 23276 17434
rect 1104 17360 23276 17382
rect 8386 17320 8392 17332
rect 1780 17292 8392 17320
rect 1780 17125 1808 17292
rect 8386 17280 8392 17292
rect 8444 17280 8450 17332
rect 9398 17320 9404 17332
rect 9359 17292 9404 17320
rect 9398 17280 9404 17292
rect 9456 17280 9462 17332
rect 9858 17280 9864 17332
rect 9916 17320 9922 17332
rect 11054 17320 11060 17332
rect 9916 17292 10732 17320
rect 11015 17292 11060 17320
rect 9916 17280 9922 17292
rect 3697 17255 3755 17261
rect 3697 17221 3709 17255
rect 3743 17252 3755 17255
rect 4062 17252 4068 17264
rect 3743 17224 4068 17252
rect 3743 17221 3755 17224
rect 3697 17215 3755 17221
rect 4062 17212 4068 17224
rect 4120 17212 4126 17264
rect 4246 17212 4252 17264
rect 4304 17252 4310 17264
rect 7009 17255 7067 17261
rect 4304 17224 4936 17252
rect 4304 17212 4310 17224
rect 4908 17193 4936 17224
rect 7009 17221 7021 17255
rect 7055 17252 7067 17255
rect 7742 17252 7748 17264
rect 7055 17224 7748 17252
rect 7055 17221 7067 17224
rect 7009 17215 7067 17221
rect 7742 17212 7748 17224
rect 7800 17212 7806 17264
rect 4893 17187 4951 17193
rect 4893 17153 4905 17187
rect 4939 17153 4951 17187
rect 4893 17147 4951 17153
rect 5902 17144 5908 17196
rect 5960 17184 5966 17196
rect 7190 17184 7196 17196
rect 5960 17156 7196 17184
rect 5960 17144 5966 17156
rect 7190 17144 7196 17156
rect 7248 17144 7254 17196
rect 7653 17187 7711 17193
rect 7653 17153 7665 17187
rect 7699 17184 7711 17187
rect 9585 17187 9643 17193
rect 7699 17156 8156 17184
rect 7699 17153 7711 17156
rect 7653 17147 7711 17153
rect 1765 17119 1823 17125
rect 1765 17085 1777 17119
rect 1811 17085 1823 17119
rect 1765 17079 1823 17085
rect 1854 17076 1860 17128
rect 1912 17116 1918 17128
rect 2225 17119 2283 17125
rect 2225 17116 2237 17119
rect 1912 17088 2237 17116
rect 1912 17076 1918 17088
rect 2225 17085 2237 17088
rect 2271 17116 2283 17119
rect 2317 17119 2375 17125
rect 2317 17116 2329 17119
rect 2271 17088 2329 17116
rect 2271 17085 2283 17088
rect 2225 17079 2283 17085
rect 2317 17085 2329 17088
rect 2363 17085 2375 17119
rect 2317 17079 2375 17085
rect 2584 17119 2642 17125
rect 2584 17085 2596 17119
rect 2630 17116 2642 17119
rect 3510 17116 3516 17128
rect 2630 17088 3516 17116
rect 2630 17085 2642 17088
rect 2584 17079 2642 17085
rect 3510 17076 3516 17088
rect 3568 17076 3574 17128
rect 4154 17076 4160 17128
rect 4212 17116 4218 17128
rect 4249 17119 4307 17125
rect 4249 17116 4261 17119
rect 4212 17088 4261 17116
rect 4212 17076 4218 17088
rect 4249 17085 4261 17088
rect 4295 17085 4307 17119
rect 4249 17079 4307 17085
rect 4341 17119 4399 17125
rect 4341 17085 4353 17119
rect 4387 17116 4399 17119
rect 4982 17116 4988 17128
rect 4387 17088 4988 17116
rect 4387 17085 4399 17088
rect 4341 17079 4399 17085
rect 4982 17076 4988 17088
rect 5040 17076 5046 17128
rect 5166 17125 5172 17128
rect 5160 17079 5172 17125
rect 5224 17116 5230 17128
rect 5224 17088 5260 17116
rect 5166 17076 5172 17079
rect 5224 17076 5230 17088
rect 7006 17076 7012 17128
rect 7064 17116 7070 17128
rect 8021 17119 8079 17125
rect 8021 17116 8033 17119
rect 7064 17088 8033 17116
rect 7064 17076 7070 17088
rect 8021 17085 8033 17088
rect 8067 17085 8079 17119
rect 8128 17116 8156 17156
rect 9585 17153 9597 17187
rect 9631 17184 9643 17187
rect 10704 17184 10732 17292
rect 11054 17280 11060 17292
rect 11112 17280 11118 17332
rect 11146 17280 11152 17332
rect 11204 17320 11210 17332
rect 12437 17323 12495 17329
rect 12437 17320 12449 17323
rect 11204 17292 12449 17320
rect 11204 17280 11210 17292
rect 12437 17289 12449 17292
rect 12483 17320 12495 17323
rect 12483 17292 12848 17320
rect 12483 17289 12495 17292
rect 12437 17283 12495 17289
rect 11072 17252 11100 17280
rect 12820 17252 12848 17292
rect 12894 17280 12900 17332
rect 12952 17320 12958 17332
rect 22094 17320 22100 17332
rect 12952 17292 22100 17320
rect 12952 17280 12958 17292
rect 22094 17280 22100 17292
rect 22152 17280 22158 17332
rect 13814 17252 13820 17264
rect 11072 17224 12296 17252
rect 12820 17224 13820 17252
rect 11793 17187 11851 17193
rect 11793 17184 11805 17187
rect 9631 17156 9812 17184
rect 10704 17156 11805 17184
rect 9631 17153 9643 17156
rect 9585 17147 9643 17153
rect 8294 17125 8300 17128
rect 8277 17119 8300 17125
rect 8277 17116 8289 17119
rect 8128 17088 8289 17116
rect 8021 17079 8079 17085
rect 8277 17085 8289 17088
rect 8352 17116 8358 17128
rect 9490 17116 9496 17128
rect 8352 17088 8425 17116
rect 9048 17088 9496 17116
rect 8277 17079 8300 17085
rect 7926 17048 7932 17060
rect 1964 17020 5488 17048
rect 1964 16989 1992 17020
rect 1949 16983 2007 16989
rect 1949 16949 1961 16983
rect 1995 16949 2007 16983
rect 1949 16943 2007 16949
rect 2130 16940 2136 16992
rect 2188 16980 2194 16992
rect 2225 16983 2283 16989
rect 2225 16980 2237 16983
rect 2188 16952 2237 16980
rect 2188 16940 2194 16952
rect 2225 16949 2237 16952
rect 2271 16980 2283 16983
rect 3326 16980 3332 16992
rect 2271 16952 3332 16980
rect 2271 16949 2283 16952
rect 2225 16943 2283 16949
rect 3326 16940 3332 16952
rect 3384 16980 3390 16992
rect 4065 16983 4123 16989
rect 4065 16980 4077 16983
rect 3384 16952 4077 16980
rect 3384 16940 3390 16952
rect 4065 16949 4077 16952
rect 4111 16949 4123 16983
rect 4522 16980 4528 16992
rect 4483 16952 4528 16980
rect 4065 16943 4123 16949
rect 4522 16940 4528 16952
rect 4580 16940 4586 16992
rect 5460 16980 5488 17020
rect 5828 17020 7932 17048
rect 5828 16980 5856 17020
rect 7926 17008 7932 17020
rect 7984 17008 7990 17060
rect 8036 17048 8064 17079
rect 8294 17076 8300 17079
rect 8352 17076 8358 17088
rect 9048 17048 9076 17088
rect 9490 17076 9496 17088
rect 9548 17116 9554 17128
rect 9677 17119 9735 17125
rect 9677 17116 9689 17119
rect 9548 17088 9689 17116
rect 9548 17076 9554 17088
rect 9677 17085 9689 17088
rect 9723 17085 9735 17119
rect 9784 17116 9812 17156
rect 11793 17153 11805 17156
rect 11839 17153 11851 17187
rect 11793 17147 11851 17153
rect 11885 17187 11943 17193
rect 11885 17153 11897 17187
rect 11931 17153 11943 17187
rect 12268 17184 12296 17224
rect 13814 17212 13820 17224
rect 13872 17212 13878 17264
rect 15010 17212 15016 17264
rect 15068 17252 15074 17264
rect 15473 17255 15531 17261
rect 15473 17252 15485 17255
rect 15068 17224 15485 17252
rect 15068 17212 15074 17224
rect 15473 17221 15485 17224
rect 15519 17221 15531 17255
rect 15473 17215 15531 17221
rect 19058 17212 19064 17264
rect 19116 17252 19122 17264
rect 21085 17255 21143 17261
rect 21085 17252 21097 17255
rect 19116 17224 21097 17252
rect 19116 17212 19122 17224
rect 21085 17221 21097 17224
rect 21131 17221 21143 17255
rect 21085 17215 21143 17221
rect 12989 17187 13047 17193
rect 12989 17184 13001 17187
rect 12268 17156 13001 17184
rect 11885 17147 11943 17153
rect 12989 17153 13001 17156
rect 13035 17153 13047 17187
rect 12989 17147 13047 17153
rect 11900 17116 11928 17147
rect 14826 17144 14832 17196
rect 14884 17184 14890 17196
rect 16025 17187 16083 17193
rect 16025 17184 16037 17187
rect 14884 17156 16037 17184
rect 14884 17144 14890 17156
rect 16025 17153 16037 17156
rect 16071 17153 16083 17187
rect 16025 17147 16083 17153
rect 16298 17144 16304 17196
rect 16356 17184 16362 17196
rect 16758 17184 16764 17196
rect 16356 17156 16764 17184
rect 16356 17144 16362 17156
rect 16758 17144 16764 17156
rect 16816 17184 16822 17196
rect 17037 17187 17095 17193
rect 17037 17184 17049 17187
rect 16816 17156 17049 17184
rect 16816 17144 16822 17156
rect 17037 17153 17049 17156
rect 17083 17153 17095 17187
rect 17037 17147 17095 17153
rect 17313 17187 17371 17193
rect 17313 17153 17325 17187
rect 17359 17184 17371 17187
rect 17359 17156 18175 17184
rect 17359 17153 17371 17156
rect 17313 17147 17371 17153
rect 9784 17088 11928 17116
rect 9677 17079 9735 17085
rect 11974 17076 11980 17128
rect 12032 17116 12038 17128
rect 12434 17116 12440 17128
rect 12032 17088 12440 17116
rect 12032 17076 12038 17088
rect 12434 17076 12440 17088
rect 12492 17076 12498 17128
rect 13262 17076 13268 17128
rect 13320 17116 13326 17128
rect 13725 17119 13783 17125
rect 13725 17116 13737 17119
rect 13320 17088 13737 17116
rect 13320 17076 13326 17088
rect 13725 17085 13737 17088
rect 13771 17085 13783 17119
rect 13725 17079 13783 17085
rect 13817 17119 13875 17125
rect 13817 17085 13829 17119
rect 13863 17085 13875 17119
rect 13817 17079 13875 17085
rect 14084 17119 14142 17125
rect 14084 17085 14096 17119
rect 14130 17116 14142 17119
rect 16666 17116 16672 17128
rect 14130 17088 16672 17116
rect 14130 17085 14142 17088
rect 14084 17079 14142 17085
rect 9950 17057 9956 17060
rect 8036 17020 9076 17048
rect 9944 17011 9956 17057
rect 10008 17048 10014 17060
rect 11698 17048 11704 17060
rect 10008 17020 10044 17048
rect 11659 17020 11704 17048
rect 9950 17008 9956 17011
rect 10008 17008 10014 17020
rect 11698 17008 11704 17020
rect 11756 17008 11762 17060
rect 12805 17051 12863 17057
rect 12805 17017 12817 17051
rect 12851 17048 12863 17051
rect 13354 17048 13360 17060
rect 12851 17020 13360 17048
rect 12851 17017 12863 17020
rect 12805 17011 12863 17017
rect 13354 17008 13360 17020
rect 13412 17008 13418 17060
rect 13832 17048 13860 17079
rect 16666 17076 16672 17088
rect 16724 17116 16730 17128
rect 16853 17119 16911 17125
rect 16853 17116 16865 17119
rect 16724 17088 16865 17116
rect 16724 17076 16730 17088
rect 16853 17085 16865 17088
rect 16899 17085 16911 17119
rect 16853 17079 16911 17085
rect 17218 17076 17224 17128
rect 17276 17116 17282 17128
rect 17497 17119 17555 17125
rect 17497 17116 17509 17119
rect 17276 17088 17509 17116
rect 17276 17076 17282 17088
rect 17497 17085 17509 17088
rect 17543 17085 17555 17119
rect 18046 17116 18052 17128
rect 18007 17088 18052 17116
rect 17497 17079 17555 17085
rect 18046 17076 18052 17088
rect 18104 17076 18110 17128
rect 18147 17116 18175 17156
rect 19334 17144 19340 17196
rect 19392 17184 19398 17196
rect 20162 17184 20168 17196
rect 19392 17156 20024 17184
rect 20123 17156 20168 17184
rect 19392 17144 19398 17156
rect 19886 17116 19892 17128
rect 18147 17088 19892 17116
rect 19886 17076 19892 17088
rect 19944 17076 19950 17128
rect 19996 17116 20024 17156
rect 20162 17144 20168 17156
rect 20220 17144 20226 17196
rect 20254 17144 20260 17196
rect 20312 17184 20318 17196
rect 20312 17156 20357 17184
rect 20312 17144 20318 17156
rect 20898 17144 20904 17196
rect 20956 17184 20962 17196
rect 20956 17156 21404 17184
rect 20956 17144 20962 17156
rect 20073 17119 20131 17125
rect 20073 17116 20085 17119
rect 19996 17088 20085 17116
rect 20073 17085 20085 17088
rect 20119 17085 20131 17119
rect 20714 17116 20720 17128
rect 20675 17088 20720 17116
rect 20073 17079 20131 17085
rect 20714 17076 20720 17088
rect 20772 17076 20778 17128
rect 21174 17116 21180 17128
rect 20824 17088 21180 17116
rect 13740 17020 13860 17048
rect 13740 16992 13768 17020
rect 13998 17008 14004 17060
rect 14056 17048 14062 17060
rect 15933 17051 15991 17057
rect 15933 17048 15945 17051
rect 14056 17020 15945 17048
rect 14056 17008 14062 17020
rect 15933 17017 15945 17020
rect 15979 17017 15991 17051
rect 15933 17011 15991 17017
rect 18138 17008 18144 17060
rect 18196 17048 18202 17060
rect 18294 17051 18352 17057
rect 18294 17048 18306 17051
rect 18196 17020 18306 17048
rect 18196 17008 18202 17020
rect 18294 17017 18306 17020
rect 18340 17017 18352 17051
rect 18294 17011 18352 17017
rect 18432 17020 19748 17048
rect 6270 16980 6276 16992
rect 5460 16952 5856 16980
rect 6231 16952 6276 16980
rect 6270 16940 6276 16952
rect 6328 16940 6334 16992
rect 7098 16940 7104 16992
rect 7156 16980 7162 16992
rect 7377 16983 7435 16989
rect 7377 16980 7389 16983
rect 7156 16952 7389 16980
rect 7156 16940 7162 16952
rect 7377 16949 7389 16952
rect 7423 16949 7435 16983
rect 7377 16943 7435 16949
rect 7466 16940 7472 16992
rect 7524 16980 7530 16992
rect 7524 16952 7569 16980
rect 7524 16940 7530 16952
rect 8110 16940 8116 16992
rect 8168 16980 8174 16992
rect 9585 16983 9643 16989
rect 9585 16980 9597 16983
rect 8168 16952 9597 16980
rect 8168 16940 8174 16952
rect 9585 16949 9597 16952
rect 9631 16949 9643 16983
rect 11330 16980 11336 16992
rect 11291 16952 11336 16980
rect 9585 16943 9643 16949
rect 11330 16940 11336 16952
rect 11388 16940 11394 16992
rect 12342 16940 12348 16992
rect 12400 16980 12406 16992
rect 12710 16980 12716 16992
rect 12400 16952 12716 16980
rect 12400 16940 12406 16952
rect 12710 16940 12716 16952
rect 12768 16940 12774 16992
rect 12894 16940 12900 16992
rect 12952 16980 12958 16992
rect 13541 16983 13599 16989
rect 12952 16952 12997 16980
rect 12952 16940 12958 16952
rect 13541 16949 13553 16983
rect 13587 16980 13599 16983
rect 13722 16980 13728 16992
rect 13587 16952 13728 16980
rect 13587 16949 13599 16952
rect 13541 16943 13599 16949
rect 13722 16940 13728 16952
rect 13780 16980 13786 16992
rect 15102 16980 15108 16992
rect 13780 16952 15108 16980
rect 13780 16940 13786 16952
rect 15102 16940 15108 16952
rect 15160 16940 15166 16992
rect 15197 16983 15255 16989
rect 15197 16949 15209 16983
rect 15243 16980 15255 16983
rect 15286 16980 15292 16992
rect 15243 16952 15292 16980
rect 15243 16949 15255 16952
rect 15197 16943 15255 16949
rect 15286 16940 15292 16952
rect 15344 16940 15350 16992
rect 15841 16983 15899 16989
rect 15841 16949 15853 16983
rect 15887 16980 15899 16983
rect 16298 16980 16304 16992
rect 15887 16952 16304 16980
rect 15887 16949 15899 16952
rect 15841 16943 15899 16949
rect 16298 16940 16304 16952
rect 16356 16940 16362 16992
rect 16482 16980 16488 16992
rect 16443 16952 16488 16980
rect 16482 16940 16488 16952
rect 16540 16940 16546 16992
rect 16942 16980 16948 16992
rect 16903 16952 16948 16980
rect 16942 16940 16948 16952
rect 17000 16940 17006 16992
rect 17034 16940 17040 16992
rect 17092 16980 17098 16992
rect 17313 16983 17371 16989
rect 17313 16980 17325 16983
rect 17092 16952 17325 16980
rect 17092 16940 17098 16952
rect 17313 16949 17325 16952
rect 17359 16949 17371 16983
rect 17313 16943 17371 16949
rect 17862 16940 17868 16992
rect 17920 16980 17926 16992
rect 18432 16980 18460 17020
rect 17920 16952 18460 16980
rect 17920 16940 17926 16952
rect 18506 16940 18512 16992
rect 18564 16980 18570 16992
rect 19058 16980 19064 16992
rect 18564 16952 19064 16980
rect 18564 16940 18570 16952
rect 19058 16940 19064 16952
rect 19116 16940 19122 16992
rect 19242 16940 19248 16992
rect 19300 16980 19306 16992
rect 19720 16989 19748 17020
rect 19429 16983 19487 16989
rect 19429 16980 19441 16983
rect 19300 16952 19441 16980
rect 19300 16940 19306 16952
rect 19429 16949 19441 16952
rect 19475 16949 19487 16983
rect 19429 16943 19487 16949
rect 19705 16983 19763 16989
rect 19705 16949 19717 16983
rect 19751 16949 19763 16983
rect 19705 16943 19763 16949
rect 19886 16940 19892 16992
rect 19944 16980 19950 16992
rect 20824 16980 20852 17088
rect 21174 17076 21180 17088
rect 21232 17076 21238 17128
rect 21376 17125 21404 17156
rect 21361 17119 21419 17125
rect 21361 17085 21373 17119
rect 21407 17116 21419 17119
rect 22186 17116 22192 17128
rect 21407 17088 22192 17116
rect 21407 17085 21419 17088
rect 21361 17079 21419 17085
rect 22186 17076 22192 17088
rect 22244 17076 22250 17128
rect 21634 17057 21640 17060
rect 20901 17051 20959 17057
rect 20901 17017 20913 17051
rect 20947 17048 20959 17051
rect 20947 17020 21588 17048
rect 20947 17017 20959 17020
rect 20901 17011 20959 17017
rect 19944 16952 20852 16980
rect 19944 16940 19950 16952
rect 21174 16940 21180 16992
rect 21232 16980 21238 16992
rect 21450 16980 21456 16992
rect 21232 16952 21456 16980
rect 21232 16940 21238 16952
rect 21450 16940 21456 16952
rect 21508 16940 21514 16992
rect 21560 16980 21588 17020
rect 21628 17011 21640 17057
rect 21692 17048 21698 17060
rect 22554 17048 22560 17060
rect 21692 17020 22560 17048
rect 21634 17008 21640 17011
rect 21692 17008 21698 17020
rect 22554 17008 22560 17020
rect 22612 17008 22618 17060
rect 21726 16980 21732 16992
rect 21560 16952 21732 16980
rect 21726 16940 21732 16952
rect 21784 16980 21790 16992
rect 22741 16983 22799 16989
rect 22741 16980 22753 16983
rect 21784 16952 22753 16980
rect 21784 16940 21790 16952
rect 22741 16949 22753 16952
rect 22787 16949 22799 16983
rect 22741 16943 22799 16949
rect 1104 16890 23276 16912
rect 1104 16838 8379 16890
rect 8431 16838 8443 16890
rect 8495 16838 8507 16890
rect 8559 16838 8571 16890
rect 8623 16838 15776 16890
rect 15828 16838 15840 16890
rect 15892 16838 15904 16890
rect 15956 16838 15968 16890
rect 16020 16838 23276 16890
rect 1104 16816 23276 16838
rect 1762 16776 1768 16788
rect 1723 16748 1768 16776
rect 1762 16736 1768 16748
rect 1820 16736 1826 16788
rect 3510 16776 3516 16788
rect 3471 16748 3516 16776
rect 3510 16736 3516 16748
rect 3568 16736 3574 16788
rect 4433 16779 4491 16785
rect 4433 16745 4445 16779
rect 4479 16776 4491 16779
rect 5902 16776 5908 16788
rect 4479 16748 5908 16776
rect 4479 16745 4491 16748
rect 4433 16739 4491 16745
rect 5902 16736 5908 16748
rect 5960 16736 5966 16788
rect 6086 16736 6092 16788
rect 6144 16776 6150 16788
rect 6181 16779 6239 16785
rect 6181 16776 6193 16779
rect 6144 16748 6193 16776
rect 6144 16736 6150 16748
rect 6181 16745 6193 16748
rect 6227 16745 6239 16779
rect 7282 16776 7288 16788
rect 6181 16739 6239 16745
rect 6472 16748 7288 16776
rect 2400 16711 2458 16717
rect 2400 16677 2412 16711
rect 2446 16708 2458 16711
rect 3418 16708 3424 16720
rect 2446 16680 3424 16708
rect 2446 16677 2458 16680
rect 2400 16671 2458 16677
rect 3418 16668 3424 16680
rect 3476 16668 3482 16720
rect 4338 16708 4344 16720
rect 3896 16680 4344 16708
rect 1581 16643 1639 16649
rect 1581 16609 1593 16643
rect 1627 16640 1639 16643
rect 3896 16640 3924 16680
rect 4338 16668 4344 16680
rect 4396 16668 4402 16720
rect 5068 16711 5126 16717
rect 5068 16677 5080 16711
rect 5114 16708 5126 16711
rect 5626 16708 5632 16720
rect 5114 16680 5632 16708
rect 5114 16677 5126 16680
rect 5068 16671 5126 16677
rect 5626 16668 5632 16680
rect 5684 16708 5690 16720
rect 6270 16708 6276 16720
rect 5684 16680 6276 16708
rect 5684 16668 5690 16680
rect 6270 16668 6276 16680
rect 6328 16668 6334 16720
rect 6472 16717 6500 16748
rect 7282 16736 7288 16748
rect 7340 16736 7346 16788
rect 8202 16736 8208 16788
rect 8260 16776 8266 16788
rect 8481 16779 8539 16785
rect 8481 16776 8493 16779
rect 8260 16748 8493 16776
rect 8260 16736 8266 16748
rect 8481 16745 8493 16748
rect 8527 16745 8539 16779
rect 8481 16739 8539 16745
rect 8573 16779 8631 16785
rect 8573 16745 8585 16779
rect 8619 16776 8631 16779
rect 9861 16779 9919 16785
rect 9861 16776 9873 16779
rect 8619 16748 9873 16776
rect 8619 16745 8631 16748
rect 8573 16739 8631 16745
rect 9861 16745 9873 16748
rect 9907 16745 9919 16779
rect 9861 16739 9919 16745
rect 12161 16779 12219 16785
rect 12161 16745 12173 16779
rect 12207 16776 12219 16779
rect 14369 16779 14427 16785
rect 14369 16776 14381 16779
rect 12207 16748 14381 16776
rect 12207 16745 12219 16748
rect 12161 16739 12219 16745
rect 14369 16745 14381 16748
rect 14415 16745 14427 16779
rect 14369 16739 14427 16745
rect 14461 16779 14519 16785
rect 14461 16745 14473 16779
rect 14507 16776 14519 16779
rect 14918 16776 14924 16788
rect 14507 16748 14924 16776
rect 14507 16745 14519 16748
rect 14461 16739 14519 16745
rect 14918 16736 14924 16748
rect 14976 16736 14982 16788
rect 16482 16736 16488 16788
rect 16540 16776 16546 16788
rect 20257 16779 20315 16785
rect 20257 16776 20269 16779
rect 16540 16748 20269 16776
rect 16540 16736 16546 16748
rect 20257 16745 20269 16748
rect 20303 16745 20315 16779
rect 20898 16776 20904 16788
rect 20859 16748 20904 16776
rect 20257 16739 20315 16745
rect 20898 16736 20904 16748
rect 20956 16736 20962 16788
rect 20990 16736 20996 16788
rect 21048 16776 21054 16788
rect 21269 16779 21327 16785
rect 21269 16776 21281 16779
rect 21048 16748 21281 16776
rect 21048 16736 21054 16748
rect 21269 16745 21281 16748
rect 21315 16776 21327 16779
rect 21913 16779 21971 16785
rect 21913 16776 21925 16779
rect 21315 16748 21925 16776
rect 21315 16745 21327 16748
rect 21269 16739 21327 16745
rect 21913 16745 21925 16748
rect 21959 16745 21971 16779
rect 21913 16739 21971 16745
rect 6457 16711 6515 16717
rect 6457 16677 6469 16711
rect 6503 16677 6515 16711
rect 6457 16671 6515 16677
rect 6825 16711 6883 16717
rect 6825 16677 6837 16711
rect 6871 16708 6883 16711
rect 6871 16680 9720 16708
rect 6871 16677 6883 16680
rect 6825 16671 6883 16677
rect 1627 16612 3924 16640
rect 4249 16643 4307 16649
rect 1627 16609 1639 16612
rect 1581 16603 1639 16609
rect 4249 16609 4261 16643
rect 4295 16640 4307 16643
rect 4430 16640 4436 16652
rect 4295 16612 4436 16640
rect 4295 16609 4307 16612
rect 4249 16603 4307 16609
rect 4430 16600 4436 16612
rect 4488 16600 4494 16652
rect 6641 16643 6699 16649
rect 6641 16609 6653 16643
rect 6687 16640 6699 16643
rect 7006 16640 7012 16652
rect 6687 16612 7012 16640
rect 6687 16609 6699 16612
rect 6641 16603 6699 16609
rect 7006 16600 7012 16612
rect 7064 16600 7070 16652
rect 7368 16643 7426 16649
rect 7368 16609 7380 16643
rect 7414 16640 7426 16643
rect 7926 16640 7932 16652
rect 7414 16612 7932 16640
rect 7414 16609 7426 16612
rect 7368 16603 7426 16609
rect 7926 16600 7932 16612
rect 7984 16600 7990 16652
rect 8202 16600 8208 16652
rect 8260 16640 8266 16652
rect 8573 16643 8631 16649
rect 8573 16640 8585 16643
rect 8260 16612 8585 16640
rect 8260 16600 8266 16612
rect 8573 16609 8585 16612
rect 8619 16609 8631 16643
rect 8754 16640 8760 16652
rect 8715 16612 8760 16640
rect 8573 16603 8631 16609
rect 8754 16600 8760 16612
rect 8812 16600 8818 16652
rect 9125 16643 9183 16649
rect 9125 16609 9137 16643
rect 9171 16640 9183 16643
rect 9490 16640 9496 16652
rect 9171 16612 9352 16640
rect 9451 16612 9496 16640
rect 9171 16609 9183 16612
rect 9125 16603 9183 16609
rect 1486 16532 1492 16584
rect 1544 16572 1550 16584
rect 2130 16572 2136 16584
rect 1544 16544 2136 16572
rect 1544 16532 1550 16544
rect 2130 16532 2136 16544
rect 2188 16532 2194 16584
rect 4798 16572 4804 16584
rect 4759 16544 4804 16572
rect 4798 16532 4804 16544
rect 4856 16532 4862 16584
rect 6914 16532 6920 16584
rect 6972 16572 6978 16584
rect 7101 16575 7159 16581
rect 7101 16572 7113 16575
rect 6972 16544 7113 16572
rect 6972 16532 6978 16544
rect 7101 16541 7113 16544
rect 7147 16541 7159 16575
rect 9324 16572 9352 16612
rect 9490 16600 9496 16612
rect 9548 16600 9554 16652
rect 9692 16649 9720 16680
rect 10042 16668 10048 16720
rect 10100 16708 10106 16720
rect 14182 16708 14188 16720
rect 10100 16680 10364 16708
rect 10100 16668 10106 16680
rect 10336 16652 10364 16680
rect 12544 16680 14188 16708
rect 9677 16643 9735 16649
rect 9677 16609 9689 16643
rect 9723 16609 9735 16643
rect 10134 16640 10140 16652
rect 9677 16603 9735 16609
rect 9784 16612 10140 16640
rect 9784 16572 9812 16612
rect 10134 16600 10140 16612
rect 10192 16600 10198 16652
rect 10318 16600 10324 16652
rect 10376 16640 10382 16652
rect 10552 16643 10610 16649
rect 10552 16640 10564 16643
rect 10376 16612 10564 16640
rect 10376 16600 10382 16612
rect 10552 16609 10564 16612
rect 10598 16609 10610 16643
rect 10552 16603 10610 16609
rect 10796 16612 11192 16640
rect 9324 16544 9812 16572
rect 10229 16575 10287 16581
rect 7101 16535 7159 16541
rect 10229 16541 10241 16575
rect 10275 16572 10287 16575
rect 10410 16572 10416 16584
rect 10275 16544 10416 16572
rect 10275 16541 10287 16544
rect 10229 16535 10287 16541
rect 10410 16532 10416 16544
rect 10468 16532 10474 16584
rect 10686 16532 10692 16584
rect 10744 16572 10750 16584
rect 10796 16572 10824 16612
rect 10962 16572 10968 16584
rect 10744 16544 10824 16572
rect 10923 16544 10968 16572
rect 10744 16532 10750 16544
rect 10962 16532 10968 16544
rect 11020 16532 11026 16584
rect 11164 16572 11192 16612
rect 11238 16600 11244 16652
rect 11296 16640 11302 16652
rect 12544 16640 12572 16680
rect 14182 16668 14188 16680
rect 14240 16668 14246 16720
rect 15556 16711 15614 16717
rect 15556 16677 15568 16711
rect 15602 16708 15614 16711
rect 16022 16708 16028 16720
rect 15602 16680 16028 16708
rect 15602 16677 15614 16680
rect 15556 16671 15614 16677
rect 16022 16668 16028 16680
rect 16080 16708 16086 16720
rect 16942 16708 16948 16720
rect 16080 16680 16948 16708
rect 16080 16668 16086 16680
rect 16942 16668 16948 16680
rect 17000 16668 17006 16720
rect 17052 16680 17908 16708
rect 11296 16612 12572 16640
rect 12612 16643 12670 16649
rect 11296 16600 11302 16612
rect 12612 16609 12624 16643
rect 12658 16640 12670 16643
rect 12986 16640 12992 16652
rect 12658 16612 12992 16640
rect 12658 16609 12670 16612
rect 12612 16603 12670 16609
rect 12986 16600 12992 16612
rect 13044 16640 13050 16652
rect 14826 16640 14832 16652
rect 13044 16612 14832 16640
rect 13044 16600 13050 16612
rect 14826 16600 14832 16612
rect 14884 16600 14890 16652
rect 15102 16600 15108 16652
rect 15160 16640 15166 16652
rect 15289 16643 15347 16649
rect 15289 16640 15301 16643
rect 15160 16612 15301 16640
rect 15160 16600 15166 16612
rect 15289 16609 15301 16612
rect 15335 16609 15347 16643
rect 15289 16603 15347 16609
rect 15396 16612 16335 16640
rect 12161 16575 12219 16581
rect 12161 16572 12173 16575
rect 11164 16544 12173 16572
rect 12161 16541 12173 16544
rect 12207 16541 12219 16575
rect 12342 16572 12348 16584
rect 12303 16544 12348 16572
rect 12161 16535 12219 16541
rect 12342 16532 12348 16544
rect 12400 16532 12406 16584
rect 14553 16575 14611 16581
rect 14553 16541 14565 16575
rect 14599 16541 14611 16575
rect 14553 16535 14611 16541
rect 12069 16507 12127 16513
rect 8036 16476 9444 16504
rect 4522 16396 4528 16448
rect 4580 16436 4586 16448
rect 8036 16436 8064 16476
rect 4580 16408 8064 16436
rect 8941 16439 8999 16445
rect 4580 16396 4586 16408
rect 8941 16405 8953 16439
rect 8987 16436 8999 16439
rect 9125 16439 9183 16445
rect 9125 16436 9137 16439
rect 8987 16408 9137 16436
rect 8987 16405 8999 16408
rect 8941 16399 8999 16405
rect 9125 16405 9137 16408
rect 9171 16405 9183 16439
rect 9125 16399 9183 16405
rect 9214 16396 9220 16448
rect 9272 16436 9278 16448
rect 9309 16439 9367 16445
rect 9309 16436 9321 16439
rect 9272 16408 9321 16436
rect 9272 16396 9278 16408
rect 9309 16405 9321 16408
rect 9355 16405 9367 16439
rect 9416 16436 9444 16476
rect 12069 16473 12081 16507
rect 12115 16504 12127 16507
rect 12250 16504 12256 16516
rect 12115 16476 12256 16504
rect 12115 16473 12127 16476
rect 12069 16467 12127 16473
rect 12250 16464 12256 16476
rect 12308 16464 12314 16516
rect 13998 16504 14004 16516
rect 13280 16476 13860 16504
rect 13959 16476 14004 16504
rect 11882 16436 11888 16448
rect 9416 16408 11888 16436
rect 9309 16399 9367 16405
rect 11882 16396 11888 16408
rect 11940 16396 11946 16448
rect 12710 16396 12716 16448
rect 12768 16436 12774 16448
rect 13280 16436 13308 16476
rect 13722 16436 13728 16448
rect 12768 16408 13308 16436
rect 13683 16408 13728 16436
rect 12768 16396 12774 16408
rect 13722 16396 13728 16408
rect 13780 16396 13786 16448
rect 13832 16436 13860 16476
rect 13998 16464 14004 16476
rect 14056 16464 14062 16516
rect 14182 16464 14188 16516
rect 14240 16504 14246 16516
rect 14568 16504 14596 16535
rect 14734 16532 14740 16584
rect 14792 16572 14798 16584
rect 15396 16572 15424 16612
rect 14792 16544 15424 16572
rect 16307 16572 16335 16612
rect 16482 16600 16488 16652
rect 16540 16640 16546 16652
rect 16758 16640 16764 16652
rect 16540 16612 16764 16640
rect 16540 16600 16546 16612
rect 16758 16600 16764 16612
rect 16816 16600 16822 16652
rect 17052 16640 17080 16680
rect 17218 16649 17224 16652
rect 17212 16640 17224 16649
rect 16960 16612 17080 16640
rect 17179 16612 17224 16640
rect 16960 16584 16988 16612
rect 17212 16603 17224 16612
rect 17218 16600 17224 16603
rect 17276 16600 17282 16652
rect 17880 16640 17908 16680
rect 18138 16668 18144 16720
rect 18196 16708 18202 16720
rect 18196 16680 19840 16708
rect 18196 16668 18202 16680
rect 18046 16640 18052 16652
rect 17880 16612 18052 16640
rect 18046 16600 18052 16612
rect 18104 16640 18110 16652
rect 18417 16643 18475 16649
rect 18417 16640 18429 16643
rect 18104 16612 18429 16640
rect 18104 16600 18110 16612
rect 18417 16609 18429 16612
rect 18463 16609 18475 16643
rect 18673 16643 18731 16649
rect 18673 16640 18685 16643
rect 18417 16603 18475 16609
rect 18515 16612 18685 16640
rect 16942 16572 16948 16584
rect 16307 16544 16804 16572
rect 16903 16544 16948 16572
rect 14792 16532 14798 16544
rect 16776 16516 16804 16544
rect 16942 16532 16948 16544
rect 17000 16532 17006 16584
rect 18515 16572 18543 16612
rect 18673 16609 18685 16612
rect 18719 16609 18731 16643
rect 18673 16603 18731 16609
rect 18966 16600 18972 16652
rect 19024 16640 19030 16652
rect 19024 16612 19748 16640
rect 19024 16600 19030 16612
rect 18340 16544 18543 16572
rect 16666 16504 16672 16516
rect 14240 16476 14596 16504
rect 16627 16476 16672 16504
rect 14240 16464 14246 16476
rect 16666 16464 16672 16476
rect 16724 16464 16730 16516
rect 16758 16464 16764 16516
rect 16816 16464 16822 16516
rect 17862 16436 17868 16448
rect 13832 16408 17868 16436
rect 17862 16396 17868 16408
rect 17920 16396 17926 16448
rect 18138 16396 18144 16448
rect 18196 16436 18202 16448
rect 18340 16445 18368 16544
rect 18325 16439 18383 16445
rect 18325 16436 18337 16439
rect 18196 16408 18337 16436
rect 18196 16396 18202 16408
rect 18325 16405 18337 16408
rect 18371 16405 18383 16439
rect 19720 16436 19748 16612
rect 19812 16513 19840 16680
rect 20070 16668 20076 16720
rect 20128 16708 20134 16720
rect 20349 16711 20407 16717
rect 20349 16708 20361 16711
rect 20128 16680 20361 16708
rect 20128 16668 20134 16680
rect 20349 16677 20361 16680
rect 20395 16677 20407 16711
rect 20349 16671 20407 16677
rect 22094 16668 22100 16720
rect 22152 16708 22158 16720
rect 22373 16711 22431 16717
rect 22373 16708 22385 16711
rect 22152 16680 22385 16708
rect 22152 16668 22158 16680
rect 22373 16677 22385 16680
rect 22419 16677 22431 16711
rect 22373 16671 22431 16677
rect 21358 16640 21364 16652
rect 21319 16612 21364 16640
rect 21358 16600 21364 16612
rect 21416 16600 21422 16652
rect 22281 16643 22339 16649
rect 22281 16609 22293 16643
rect 22327 16640 22339 16643
rect 23106 16640 23112 16652
rect 22327 16612 23112 16640
rect 22327 16609 22339 16612
rect 22281 16603 22339 16609
rect 23106 16600 23112 16612
rect 23164 16600 23170 16652
rect 20162 16532 20168 16584
rect 20220 16572 20226 16584
rect 20441 16575 20499 16581
rect 20441 16572 20453 16575
rect 20220 16544 20453 16572
rect 20220 16532 20226 16544
rect 20441 16541 20453 16544
rect 20487 16541 20499 16575
rect 21450 16572 21456 16584
rect 21411 16544 21456 16572
rect 20441 16535 20499 16541
rect 21450 16532 21456 16544
rect 21508 16532 21514 16584
rect 22465 16575 22523 16581
rect 22465 16541 22477 16575
rect 22511 16541 22523 16575
rect 22465 16535 22523 16541
rect 19797 16507 19855 16513
rect 19797 16473 19809 16507
rect 19843 16473 19855 16507
rect 19797 16467 19855 16473
rect 20254 16464 20260 16516
rect 20312 16504 20318 16516
rect 22480 16504 22508 16535
rect 20312 16476 22508 16504
rect 20312 16464 20318 16476
rect 19889 16439 19947 16445
rect 19889 16436 19901 16439
rect 19720 16408 19901 16436
rect 18325 16399 18383 16405
rect 19889 16405 19901 16408
rect 19935 16405 19947 16439
rect 19889 16399 19947 16405
rect 1104 16346 23276 16368
rect 1104 16294 4680 16346
rect 4732 16294 4744 16346
rect 4796 16294 4808 16346
rect 4860 16294 4872 16346
rect 4924 16294 12078 16346
rect 12130 16294 12142 16346
rect 12194 16294 12206 16346
rect 12258 16294 12270 16346
rect 12322 16294 19475 16346
rect 19527 16294 19539 16346
rect 19591 16294 19603 16346
rect 19655 16294 19667 16346
rect 19719 16294 23276 16346
rect 1104 16272 23276 16294
rect 2774 16192 2780 16244
rect 2832 16232 2838 16244
rect 2869 16235 2927 16241
rect 2869 16232 2881 16235
rect 2832 16204 2881 16232
rect 2832 16192 2838 16204
rect 2869 16201 2881 16204
rect 2915 16232 2927 16235
rect 3694 16232 3700 16244
rect 2915 16204 3700 16232
rect 2915 16201 2927 16204
rect 2869 16195 2927 16201
rect 3694 16192 3700 16204
rect 3752 16192 3758 16244
rect 4154 16192 4160 16244
rect 4212 16232 4218 16244
rect 6457 16235 6515 16241
rect 6457 16232 6469 16235
rect 4212 16204 6469 16232
rect 4212 16192 4218 16204
rect 6457 16201 6469 16204
rect 6503 16201 6515 16235
rect 6457 16195 6515 16201
rect 7377 16235 7435 16241
rect 7377 16201 7389 16235
rect 7423 16232 7435 16235
rect 7466 16232 7472 16244
rect 7423 16204 7472 16232
rect 7423 16201 7435 16204
rect 7377 16195 7435 16201
rect 7466 16192 7472 16204
rect 7524 16192 7530 16244
rect 9214 16192 9220 16244
rect 9272 16232 9278 16244
rect 10781 16235 10839 16241
rect 10781 16232 10793 16235
rect 9272 16204 10793 16232
rect 9272 16192 9278 16204
rect 10781 16201 10793 16204
rect 10827 16201 10839 16235
rect 12986 16232 12992 16244
rect 10781 16195 10839 16201
rect 10888 16204 12992 16232
rect 4430 16164 4436 16176
rect 4391 16136 4436 16164
rect 4430 16124 4436 16136
rect 4488 16124 4494 16176
rect 7650 16124 7656 16176
rect 7708 16164 7714 16176
rect 8110 16164 8116 16176
rect 7708 16136 8116 16164
rect 7708 16124 7714 16136
rect 8110 16124 8116 16136
rect 8168 16124 8174 16176
rect 10226 16124 10232 16176
rect 10284 16164 10290 16176
rect 10888 16164 10916 16204
rect 12986 16192 12992 16204
rect 13044 16192 13050 16244
rect 15194 16232 15200 16244
rect 13832 16204 15056 16232
rect 15155 16204 15200 16232
rect 10284 16136 10916 16164
rect 12437 16167 12495 16173
rect 10284 16124 10290 16136
rect 12437 16133 12449 16167
rect 12483 16164 12495 16167
rect 12894 16164 12900 16176
rect 12483 16136 12900 16164
rect 12483 16133 12495 16136
rect 12437 16127 12495 16133
rect 12894 16124 12900 16136
rect 12952 16124 12958 16176
rect 13832 16164 13860 16204
rect 13464 16136 13860 16164
rect 15028 16164 15056 16204
rect 15194 16192 15200 16204
rect 15252 16192 15258 16244
rect 17589 16235 17647 16241
rect 15488 16204 16804 16232
rect 15488 16164 15516 16204
rect 15028 16136 15516 16164
rect 1486 16096 1492 16108
rect 1447 16068 1492 16096
rect 1486 16056 1492 16068
rect 1544 16056 1550 16108
rect 3789 16099 3847 16105
rect 3789 16065 3801 16099
rect 3835 16096 3847 16099
rect 4338 16096 4344 16108
rect 3835 16068 4344 16096
rect 3835 16065 3847 16068
rect 3789 16059 3847 16065
rect 4338 16056 4344 16068
rect 4396 16056 4402 16108
rect 6656 16068 7788 16096
rect 4249 16031 4307 16037
rect 4249 15997 4261 16031
rect 4295 15997 4307 16031
rect 4798 16028 4804 16040
rect 4759 16000 4804 16028
rect 4249 15991 4307 15997
rect 1756 15963 1814 15969
rect 1756 15929 1768 15963
rect 1802 15960 1814 15963
rect 4264 15960 4292 15991
rect 4798 15988 4804 16000
rect 4856 15988 4862 16040
rect 5068 16031 5126 16037
rect 5068 15997 5080 16031
rect 5114 16028 5126 16031
rect 6086 16028 6092 16040
rect 5114 16000 6092 16028
rect 5114 15997 5126 16000
rect 5068 15991 5126 15997
rect 6086 15988 6092 16000
rect 6144 15988 6150 16040
rect 6656 16037 6684 16068
rect 6641 16031 6699 16037
rect 6641 15997 6653 16031
rect 6687 15997 6699 16031
rect 6641 15991 6699 15997
rect 6825 16031 6883 16037
rect 6825 15997 6837 16031
rect 6871 16028 6883 16031
rect 7650 16028 7656 16040
rect 6871 16000 7656 16028
rect 6871 15997 6883 16000
rect 6825 15991 6883 15997
rect 7650 15988 7656 16000
rect 7708 15988 7714 16040
rect 7760 16028 7788 16068
rect 7926 16056 7932 16108
rect 7984 16096 7990 16108
rect 8021 16099 8079 16105
rect 8021 16096 8033 16099
rect 7984 16068 8033 16096
rect 7984 16056 7990 16068
rect 8021 16065 8033 16068
rect 8067 16096 8079 16099
rect 8846 16096 8852 16108
rect 8067 16068 8852 16096
rect 8067 16065 8079 16068
rect 8021 16059 8079 16065
rect 8846 16056 8852 16068
rect 8904 16056 8910 16108
rect 8938 16056 8944 16108
rect 8996 16105 9002 16108
rect 8996 16099 9046 16105
rect 8996 16065 9000 16099
rect 9034 16065 9046 16099
rect 8996 16059 9046 16065
rect 9171 16099 9229 16105
rect 9171 16065 9183 16099
rect 9217 16096 9229 16099
rect 11238 16096 11244 16108
rect 9217 16068 11244 16096
rect 9217 16065 9229 16068
rect 9171 16059 9229 16065
rect 8996 16056 9002 16059
rect 11238 16056 11244 16068
rect 11296 16056 11302 16108
rect 11422 16096 11428 16108
rect 11383 16068 11428 16096
rect 11422 16056 11428 16068
rect 11480 16056 11486 16108
rect 11698 16056 11704 16108
rect 11756 16096 11762 16108
rect 12989 16099 13047 16105
rect 12989 16096 13001 16099
rect 11756 16068 13001 16096
rect 11756 16056 11762 16068
rect 12989 16065 13001 16068
rect 13035 16065 13047 16099
rect 12989 16059 13047 16065
rect 8573 16031 8631 16037
rect 7760 16000 8340 16028
rect 5350 15960 5356 15972
rect 1802 15932 4200 15960
rect 4264 15932 5356 15960
rect 1802 15929 1814 15932
rect 1756 15923 1814 15929
rect 3142 15892 3148 15904
rect 3103 15864 3148 15892
rect 3142 15852 3148 15864
rect 3200 15852 3206 15904
rect 3510 15892 3516 15904
rect 3471 15864 3516 15892
rect 3510 15852 3516 15864
rect 3568 15852 3574 15904
rect 3605 15895 3663 15901
rect 3605 15861 3617 15895
rect 3651 15892 3663 15895
rect 3694 15892 3700 15904
rect 3651 15864 3700 15892
rect 3651 15861 3663 15864
rect 3605 15855 3663 15861
rect 3694 15852 3700 15864
rect 3752 15852 3758 15904
rect 4172 15892 4200 15932
rect 5350 15920 5356 15932
rect 5408 15920 5414 15972
rect 7837 15963 7895 15969
rect 7837 15960 7849 15963
rect 7024 15932 7849 15960
rect 5534 15892 5540 15904
rect 4172 15864 5540 15892
rect 5534 15852 5540 15864
rect 5592 15892 5598 15904
rect 7024 15901 7052 15932
rect 7837 15929 7849 15932
rect 7883 15929 7895 15963
rect 8312 15960 8340 16000
rect 8573 15997 8585 16031
rect 8619 16028 8631 16031
rect 8665 16031 8723 16037
rect 8665 16028 8677 16031
rect 8619 16000 8677 16028
rect 8619 15997 8631 16000
rect 8573 15991 8631 15997
rect 8665 15997 8677 16000
rect 8711 15997 8723 16031
rect 9306 16028 9312 16040
rect 8665 15991 8723 15997
rect 8772 16000 9312 16028
rect 8772 15960 8800 16000
rect 9306 15988 9312 16000
rect 9364 15988 9370 16040
rect 9401 16031 9459 16037
rect 9401 15997 9413 16031
rect 9447 16028 9459 16031
rect 9674 16028 9680 16040
rect 9447 16000 9680 16028
rect 9447 15997 9459 16000
rect 9401 15991 9459 15997
rect 9674 15988 9680 16000
rect 9732 15988 9738 16040
rect 10134 15988 10140 16040
rect 10192 16028 10198 16040
rect 11149 16031 11207 16037
rect 11149 16028 11161 16031
rect 10192 16000 11161 16028
rect 10192 15988 10198 16000
rect 11149 15997 11161 16000
rect 11195 15997 11207 16031
rect 11149 15991 11207 15997
rect 11514 15988 11520 16040
rect 11572 16028 11578 16040
rect 11793 16031 11851 16037
rect 11793 16028 11805 16031
rect 11572 16000 11805 16028
rect 11572 15988 11578 16000
rect 11793 15997 11805 16000
rect 11839 15997 11851 16031
rect 11793 15991 11851 15997
rect 11882 15988 11888 16040
rect 11940 16028 11946 16040
rect 13464 16028 13492 16136
rect 13814 16096 13820 16108
rect 13775 16068 13820 16096
rect 13814 16056 13820 16068
rect 13872 16056 13878 16108
rect 15102 16056 15108 16108
rect 15160 16096 15166 16108
rect 15473 16099 15531 16105
rect 15473 16096 15485 16099
rect 15160 16068 15485 16096
rect 15160 16056 15166 16068
rect 15473 16065 15485 16068
rect 15519 16065 15531 16099
rect 16776 16096 16804 16204
rect 17589 16201 17601 16235
rect 17635 16232 17647 16235
rect 17678 16232 17684 16244
rect 17635 16204 17684 16232
rect 17635 16201 17647 16204
rect 17589 16195 17647 16201
rect 17678 16192 17684 16204
rect 17736 16192 17742 16244
rect 17773 16235 17831 16241
rect 17773 16201 17785 16235
rect 17819 16232 17831 16235
rect 20162 16232 20168 16244
rect 17819 16204 20168 16232
rect 17819 16201 17831 16204
rect 17773 16195 17831 16201
rect 20162 16192 20168 16204
rect 20220 16192 20226 16244
rect 20533 16235 20591 16241
rect 20533 16201 20545 16235
rect 20579 16232 20591 16235
rect 22370 16232 22376 16244
rect 20579 16204 22376 16232
rect 20579 16201 20591 16204
rect 20533 16195 20591 16201
rect 22370 16192 22376 16204
rect 22428 16192 22434 16244
rect 17034 16124 17040 16176
rect 17092 16164 17098 16176
rect 19705 16167 19763 16173
rect 19705 16164 19717 16167
rect 17092 16136 19717 16164
rect 17092 16124 17098 16136
rect 19705 16133 19717 16136
rect 19751 16164 19763 16167
rect 21358 16164 21364 16176
rect 19751 16136 21364 16164
rect 19751 16133 19763 16136
rect 19705 16127 19763 16133
rect 21358 16124 21364 16136
rect 21416 16124 21422 16176
rect 20254 16096 20260 16108
rect 16776 16068 20260 16096
rect 15473 16059 15531 16065
rect 20254 16056 20260 16068
rect 20312 16056 20318 16108
rect 20806 16056 20812 16108
rect 20864 16096 20870 16108
rect 21085 16099 21143 16105
rect 21085 16096 21097 16099
rect 20864 16068 21097 16096
rect 20864 16056 20870 16068
rect 21085 16065 21097 16068
rect 21131 16065 21143 16099
rect 21085 16059 21143 16065
rect 11940 16000 13492 16028
rect 13725 16031 13783 16037
rect 11940 15988 11946 16000
rect 13725 15997 13737 16031
rect 13771 16028 13783 16031
rect 14918 16028 14924 16040
rect 13771 16000 14924 16028
rect 13771 15997 13783 16000
rect 13725 15991 13783 15997
rect 14918 15988 14924 16000
rect 14976 16028 14982 16040
rect 17313 16031 17371 16037
rect 17313 16028 17325 16031
rect 14976 16000 17325 16028
rect 14976 15988 14982 16000
rect 17313 15997 17325 16000
rect 17359 15997 17371 16031
rect 17313 15991 17371 15997
rect 17405 16031 17463 16037
rect 17405 15997 17417 16031
rect 17451 16028 17463 16031
rect 17586 16028 17592 16040
rect 17451 16000 17592 16028
rect 17451 15997 17463 16000
rect 17405 15991 17463 15997
rect 17586 15988 17592 16000
rect 17644 15988 17650 16040
rect 17678 15988 17684 16040
rect 17736 16028 17742 16040
rect 17773 16031 17831 16037
rect 17773 16028 17785 16031
rect 17736 16000 17785 16028
rect 17736 15988 17742 16000
rect 17773 15997 17785 16000
rect 17819 15997 17831 16031
rect 17773 15991 17831 15997
rect 17862 15988 17868 16040
rect 17920 16028 17926 16040
rect 20073 16031 20131 16037
rect 20073 16028 20085 16031
rect 17920 16000 20085 16028
rect 17920 15988 17926 16000
rect 20073 15997 20085 16000
rect 20119 15997 20131 16031
rect 21358 16028 21364 16040
rect 21319 16000 21364 16028
rect 20073 15991 20131 15997
rect 21358 15988 21364 16000
rect 21416 16028 21422 16040
rect 22186 16028 22192 16040
rect 21416 16000 22192 16028
rect 21416 15988 21422 16000
rect 22186 15988 22192 16000
rect 22244 15988 22250 16040
rect 10962 15960 10968 15972
rect 8312 15932 8800 15960
rect 10520 15932 10968 15960
rect 7837 15923 7895 15929
rect 6181 15895 6239 15901
rect 6181 15892 6193 15895
rect 5592 15864 6193 15892
rect 5592 15852 5598 15864
rect 6181 15861 6193 15864
rect 6227 15861 6239 15895
rect 6181 15855 6239 15861
rect 7009 15895 7067 15901
rect 7009 15861 7021 15895
rect 7055 15861 7067 15895
rect 7742 15892 7748 15904
rect 7703 15864 7748 15892
rect 7009 15855 7067 15861
rect 7742 15852 7748 15864
rect 7800 15852 7806 15904
rect 8573 15895 8631 15901
rect 8573 15861 8585 15895
rect 8619 15892 8631 15895
rect 10410 15892 10416 15904
rect 8619 15864 10416 15892
rect 8619 15861 8631 15864
rect 8573 15855 8631 15861
rect 10410 15852 10416 15864
rect 10468 15852 10474 15904
rect 10520 15901 10548 15932
rect 10962 15920 10968 15932
rect 11020 15960 11026 15972
rect 12897 15963 12955 15969
rect 12897 15960 12909 15963
rect 11020 15932 12909 15960
rect 11020 15920 11026 15932
rect 12897 15929 12909 15932
rect 12943 15929 12955 15963
rect 12897 15923 12955 15929
rect 14084 15963 14142 15969
rect 14084 15929 14096 15963
rect 14130 15960 14142 15963
rect 15378 15960 15384 15972
rect 14130 15932 15384 15960
rect 14130 15929 14142 15932
rect 14084 15923 14142 15929
rect 15378 15920 15384 15932
rect 15436 15920 15442 15972
rect 15654 15920 15660 15972
rect 15712 15969 15718 15972
rect 15712 15963 15776 15969
rect 15712 15929 15730 15963
rect 15764 15929 15776 15963
rect 15712 15923 15776 15929
rect 15712 15920 15718 15923
rect 15838 15920 15844 15972
rect 15896 15960 15902 15972
rect 19521 15963 19579 15969
rect 19521 15960 19533 15963
rect 15896 15932 19533 15960
rect 15896 15920 15902 15932
rect 19521 15929 19533 15932
rect 19567 15960 19579 15963
rect 20165 15963 20223 15969
rect 20165 15960 20177 15963
rect 19567 15932 20177 15960
rect 19567 15929 19579 15932
rect 19521 15923 19579 15929
rect 20165 15929 20177 15932
rect 20211 15929 20223 15963
rect 20898 15960 20904 15972
rect 20859 15932 20904 15960
rect 20165 15923 20223 15929
rect 20898 15920 20904 15932
rect 20956 15920 20962 15972
rect 21628 15963 21686 15969
rect 21628 15929 21640 15963
rect 21674 15960 21686 15963
rect 21726 15960 21732 15972
rect 21674 15932 21732 15960
rect 21674 15929 21686 15932
rect 21628 15923 21686 15929
rect 21726 15920 21732 15932
rect 21784 15920 21790 15972
rect 10505 15895 10563 15901
rect 10505 15861 10517 15895
rect 10551 15861 10563 15895
rect 11238 15892 11244 15904
rect 11199 15864 11244 15892
rect 10505 15855 10563 15861
rect 11238 15852 11244 15864
rect 11296 15852 11302 15904
rect 11790 15852 11796 15904
rect 11848 15892 11854 15904
rect 11977 15895 12035 15901
rect 11977 15892 11989 15895
rect 11848 15864 11989 15892
rect 11848 15852 11854 15864
rect 11977 15861 11989 15864
rect 12023 15861 12035 15895
rect 11977 15855 12035 15861
rect 12342 15852 12348 15904
rect 12400 15892 12406 15904
rect 12710 15892 12716 15904
rect 12400 15864 12716 15892
rect 12400 15852 12406 15864
rect 12710 15852 12716 15864
rect 12768 15852 12774 15904
rect 12802 15852 12808 15904
rect 12860 15892 12866 15904
rect 12860 15864 12905 15892
rect 12860 15852 12866 15864
rect 13262 15852 13268 15904
rect 13320 15892 13326 15904
rect 13541 15895 13599 15901
rect 13541 15892 13553 15895
rect 13320 15864 13553 15892
rect 13320 15852 13326 15864
rect 13541 15861 13553 15864
rect 13587 15861 13599 15895
rect 13541 15855 13599 15861
rect 13906 15852 13912 15904
rect 13964 15892 13970 15904
rect 16298 15892 16304 15904
rect 13964 15864 16304 15892
rect 13964 15852 13970 15864
rect 16298 15852 16304 15864
rect 16356 15852 16362 15904
rect 16666 15852 16672 15904
rect 16724 15892 16730 15904
rect 16853 15895 16911 15901
rect 16853 15892 16865 15895
rect 16724 15864 16865 15892
rect 16724 15852 16730 15864
rect 16853 15861 16865 15864
rect 16899 15861 16911 15895
rect 16853 15855 16911 15861
rect 17129 15895 17187 15901
rect 17129 15861 17141 15895
rect 17175 15892 17187 15895
rect 17494 15892 17500 15904
rect 17175 15864 17500 15892
rect 17175 15861 17187 15864
rect 17129 15855 17187 15861
rect 17494 15852 17500 15864
rect 17552 15892 17558 15904
rect 20530 15892 20536 15904
rect 17552 15864 20536 15892
rect 17552 15852 17558 15864
rect 20530 15852 20536 15864
rect 20588 15852 20594 15904
rect 20990 15892 20996 15904
rect 20951 15864 20996 15892
rect 20990 15852 20996 15864
rect 21048 15852 21054 15904
rect 22738 15892 22744 15904
rect 22699 15864 22744 15892
rect 22738 15852 22744 15864
rect 22796 15852 22802 15904
rect 1104 15802 23276 15824
rect 1104 15750 8379 15802
rect 8431 15750 8443 15802
rect 8495 15750 8507 15802
rect 8559 15750 8571 15802
rect 8623 15750 15776 15802
rect 15828 15750 15840 15802
rect 15892 15750 15904 15802
rect 15956 15750 15968 15802
rect 16020 15750 23276 15802
rect 1104 15728 23276 15750
rect 2866 15648 2872 15700
rect 2924 15688 2930 15700
rect 3145 15691 3203 15697
rect 3145 15688 3157 15691
rect 2924 15660 3157 15688
rect 2924 15648 2930 15660
rect 3145 15657 3157 15660
rect 3191 15657 3203 15691
rect 3145 15651 3203 15657
rect 7006 15648 7012 15700
rect 7064 15688 7070 15700
rect 7101 15691 7159 15697
rect 7101 15688 7113 15691
rect 7064 15660 7113 15688
rect 7064 15648 7070 15660
rect 7101 15657 7113 15660
rect 7147 15657 7159 15691
rect 7101 15651 7159 15657
rect 2032 15623 2090 15629
rect 2032 15589 2044 15623
rect 2078 15620 2090 15623
rect 2774 15620 2780 15632
rect 2078 15592 2780 15620
rect 2078 15589 2090 15592
rect 2032 15583 2090 15589
rect 2774 15580 2780 15592
rect 2832 15580 2838 15632
rect 4338 15580 4344 15632
rect 4396 15620 4402 15632
rect 4396 15592 4752 15620
rect 4396 15580 4402 15592
rect 3421 15555 3479 15561
rect 3421 15521 3433 15555
rect 3467 15552 3479 15555
rect 3970 15552 3976 15564
rect 3467 15524 3976 15552
rect 3467 15521 3479 15524
rect 3421 15515 3479 15521
rect 3970 15512 3976 15524
rect 4028 15512 4034 15564
rect 4065 15555 4123 15561
rect 4065 15521 4077 15555
rect 4111 15552 4123 15555
rect 4111 15524 4660 15552
rect 4111 15521 4123 15524
rect 4065 15515 4123 15521
rect 1762 15484 1768 15496
rect 1723 15456 1768 15484
rect 1762 15444 1768 15456
rect 1820 15444 1826 15496
rect 4522 15484 4528 15496
rect 3528 15456 4528 15484
rect 1670 15308 1676 15360
rect 1728 15348 1734 15360
rect 3528 15348 3556 15456
rect 4522 15444 4528 15456
rect 4580 15444 4586 15496
rect 3605 15419 3663 15425
rect 3605 15385 3617 15419
rect 3651 15416 3663 15419
rect 4338 15416 4344 15428
rect 3651 15388 4344 15416
rect 3651 15385 3663 15388
rect 3605 15379 3663 15385
rect 4338 15376 4344 15388
rect 4396 15376 4402 15428
rect 4632 15425 4660 15524
rect 4617 15419 4675 15425
rect 4617 15385 4629 15419
rect 4663 15385 4675 15419
rect 4724 15416 4752 15592
rect 4798 15580 4804 15632
rect 4856 15620 4862 15632
rect 5988 15623 6046 15629
rect 4856 15592 5672 15620
rect 4856 15580 4862 15592
rect 4985 15555 5043 15561
rect 4985 15521 4997 15555
rect 5031 15552 5043 15555
rect 5534 15552 5540 15564
rect 5031 15524 5540 15552
rect 5031 15521 5043 15524
rect 4985 15515 5043 15521
rect 5534 15512 5540 15524
rect 5592 15512 5598 15564
rect 5644 15552 5672 15592
rect 5988 15589 6000 15623
rect 6034 15620 6046 15623
rect 6178 15620 6184 15632
rect 6034 15592 6184 15620
rect 6034 15589 6046 15592
rect 5988 15583 6046 15589
rect 6178 15580 6184 15592
rect 6236 15580 6242 15632
rect 6546 15580 6552 15632
rect 6604 15620 6610 15632
rect 6730 15620 6736 15632
rect 6604 15592 6736 15620
rect 6604 15580 6610 15592
rect 6730 15580 6736 15592
rect 6788 15580 6794 15632
rect 7116 15620 7144 15651
rect 7742 15648 7748 15700
rect 7800 15688 7806 15700
rect 9217 15691 9275 15697
rect 9217 15688 9229 15691
rect 7800 15660 9229 15688
rect 7800 15648 7806 15660
rect 9217 15657 9229 15660
rect 9263 15657 9275 15691
rect 9217 15651 9275 15657
rect 9306 15648 9312 15700
rect 9364 15688 9370 15700
rect 9490 15688 9496 15700
rect 9364 15660 9496 15688
rect 9364 15648 9370 15660
rect 9490 15648 9496 15660
rect 9548 15648 9554 15700
rect 9677 15691 9735 15697
rect 9677 15657 9689 15691
rect 9723 15688 9735 15691
rect 9858 15688 9864 15700
rect 9723 15660 9864 15688
rect 9723 15657 9735 15660
rect 9677 15651 9735 15657
rect 9858 15648 9864 15660
rect 9916 15648 9922 15700
rect 10137 15691 10195 15697
rect 10137 15657 10149 15691
rect 10183 15688 10195 15691
rect 11330 15688 11336 15700
rect 10183 15660 11336 15688
rect 10183 15657 10195 15660
rect 10137 15651 10195 15657
rect 11330 15648 11336 15660
rect 11388 15648 11394 15700
rect 14737 15691 14795 15697
rect 14737 15688 14749 15691
rect 11440 15660 14749 15688
rect 7622 15623 7680 15629
rect 7622 15620 7634 15623
rect 7116 15592 7634 15620
rect 7622 15589 7634 15592
rect 7668 15589 7680 15623
rect 8849 15623 8907 15629
rect 8849 15620 8861 15623
rect 7622 15583 7680 15589
rect 7760 15592 8861 15620
rect 5721 15555 5779 15561
rect 5721 15552 5733 15555
rect 5644 15524 5733 15552
rect 5721 15521 5733 15524
rect 5767 15552 5779 15555
rect 6914 15552 6920 15564
rect 5767 15524 6920 15552
rect 5767 15521 5779 15524
rect 5721 15515 5779 15521
rect 6914 15512 6920 15524
rect 6972 15552 6978 15564
rect 7377 15555 7435 15561
rect 7377 15552 7389 15555
rect 6972 15524 7389 15552
rect 6972 15512 6978 15524
rect 7377 15521 7389 15524
rect 7423 15552 7435 15555
rect 7760 15552 7788 15592
rect 8849 15589 8861 15592
rect 8895 15589 8907 15623
rect 8849 15583 8907 15589
rect 8938 15580 8944 15632
rect 8996 15620 9002 15632
rect 10226 15620 10232 15632
rect 8996 15592 10232 15620
rect 8996 15580 9002 15592
rect 10226 15580 10232 15592
rect 10284 15580 10290 15632
rect 11440 15620 11468 15660
rect 14737 15657 14749 15660
rect 14783 15657 14795 15691
rect 14918 15688 14924 15700
rect 14879 15660 14924 15688
rect 14737 15651 14795 15657
rect 14918 15648 14924 15660
rect 14976 15648 14982 15700
rect 15194 15648 15200 15700
rect 15252 15688 15258 15700
rect 15252 15660 15577 15688
rect 15252 15648 15258 15660
rect 10336 15592 11468 15620
rect 7423 15524 7788 15552
rect 7423 15521 7435 15524
rect 7377 15515 7435 15521
rect 8110 15512 8116 15564
rect 8168 15552 8174 15564
rect 8168 15524 8432 15552
rect 8168 15512 8174 15524
rect 5074 15484 5080 15496
rect 5035 15456 5080 15484
rect 5074 15444 5080 15456
rect 5132 15444 5138 15496
rect 5169 15487 5227 15493
rect 5169 15453 5181 15487
rect 5215 15453 5227 15487
rect 8404 15484 8432 15524
rect 8478 15512 8484 15564
rect 8536 15552 8542 15564
rect 9033 15555 9091 15561
rect 9033 15552 9045 15555
rect 8536 15524 9045 15552
rect 8536 15512 8542 15524
rect 9033 15521 9045 15524
rect 9079 15521 9091 15555
rect 10042 15552 10048 15564
rect 10003 15524 10048 15552
rect 9033 15515 9091 15521
rect 10042 15512 10048 15524
rect 10100 15512 10106 15564
rect 10229 15487 10287 15493
rect 10229 15484 10241 15487
rect 8404 15456 10241 15484
rect 5169 15447 5227 15453
rect 10229 15453 10241 15456
rect 10275 15453 10287 15487
rect 10229 15447 10287 15453
rect 5184 15416 5212 15447
rect 4724 15388 5212 15416
rect 4617 15379 4675 15385
rect 6730 15376 6736 15428
rect 6788 15416 6794 15428
rect 10336 15416 10364 15592
rect 11790 15580 11796 15632
rect 11848 15620 11854 15632
rect 13906 15620 13912 15632
rect 11848 15592 13912 15620
rect 11848 15580 11854 15592
rect 13906 15580 13912 15592
rect 13964 15580 13970 15632
rect 15549 15629 15577 15660
rect 16298 15648 16304 15700
rect 16356 15688 16362 15700
rect 20990 15688 20996 15700
rect 16356 15660 20996 15688
rect 16356 15648 16362 15660
rect 20990 15648 20996 15660
rect 21048 15648 21054 15700
rect 15534 15623 15592 15629
rect 15534 15589 15546 15623
rect 15580 15589 15592 15623
rect 15534 15583 15592 15589
rect 15746 15580 15752 15632
rect 15804 15620 15810 15632
rect 19334 15620 19340 15632
rect 15804 15592 19340 15620
rect 15804 15580 15810 15592
rect 19334 15580 19340 15592
rect 19392 15580 19398 15632
rect 19426 15580 19432 15632
rect 19484 15620 19490 15632
rect 20714 15620 20720 15632
rect 19484 15592 20720 15620
rect 19484 15580 19490 15592
rect 20714 15580 20720 15592
rect 20772 15580 20778 15632
rect 21358 15620 21364 15632
rect 21008 15592 21364 15620
rect 10956 15555 11014 15561
rect 10956 15521 10968 15555
rect 11002 15552 11014 15555
rect 12621 15555 12679 15561
rect 11002 15524 12572 15552
rect 11002 15521 11014 15524
rect 10956 15515 11014 15521
rect 10594 15444 10600 15496
rect 10652 15484 10658 15496
rect 10689 15487 10747 15493
rect 10689 15484 10701 15487
rect 10652 15456 10701 15484
rect 10652 15444 10658 15456
rect 10689 15453 10701 15456
rect 10735 15453 10747 15487
rect 10689 15447 10747 15453
rect 10612 15416 10640 15444
rect 12342 15416 12348 15428
rect 6788 15388 6960 15416
rect 6788 15376 6794 15388
rect 1728 15320 3556 15348
rect 4249 15351 4307 15357
rect 1728 15308 1734 15320
rect 4249 15317 4261 15351
rect 4295 15348 4307 15351
rect 6822 15348 6828 15360
rect 4295 15320 6828 15348
rect 4295 15317 4307 15320
rect 4249 15311 4307 15317
rect 6822 15308 6828 15320
rect 6880 15308 6886 15360
rect 6932 15348 6960 15388
rect 8312 15388 10364 15416
rect 10428 15388 10640 15416
rect 11624 15388 12348 15416
rect 8312 15348 8340 15388
rect 6932 15320 8340 15348
rect 8757 15351 8815 15357
rect 8757 15317 8769 15351
rect 8803 15348 8815 15351
rect 8846 15348 8852 15360
rect 8803 15320 8852 15348
rect 8803 15317 8815 15320
rect 8757 15311 8815 15317
rect 8846 15308 8852 15320
rect 8904 15308 8910 15360
rect 8941 15351 8999 15357
rect 8941 15317 8953 15351
rect 8987 15348 8999 15351
rect 9674 15348 9680 15360
rect 8987 15320 9680 15348
rect 8987 15317 8999 15320
rect 8941 15311 8999 15317
rect 9674 15308 9680 15320
rect 9732 15348 9738 15360
rect 10428 15348 10456 15388
rect 9732 15320 10456 15348
rect 9732 15308 9738 15320
rect 10502 15308 10508 15360
rect 10560 15348 10566 15360
rect 11624 15348 11652 15388
rect 12342 15376 12348 15388
rect 12400 15416 12406 15428
rect 12437 15419 12495 15425
rect 12437 15416 12449 15419
rect 12400 15388 12449 15416
rect 12400 15376 12406 15388
rect 12437 15385 12449 15388
rect 12483 15385 12495 15419
rect 12437 15379 12495 15385
rect 10560 15320 11652 15348
rect 10560 15308 10566 15320
rect 11974 15308 11980 15360
rect 12032 15348 12038 15360
rect 12069 15351 12127 15357
rect 12069 15348 12081 15351
rect 12032 15320 12081 15348
rect 12032 15308 12038 15320
rect 12069 15317 12081 15320
rect 12115 15317 12127 15351
rect 12544 15348 12572 15524
rect 12621 15521 12633 15555
rect 12667 15552 12679 15555
rect 12802 15552 12808 15564
rect 12667 15524 12808 15552
rect 12667 15521 12679 15524
rect 12621 15515 12679 15521
rect 12802 15512 12808 15524
rect 12860 15512 12866 15564
rect 12980 15555 13038 15561
rect 12980 15521 12992 15555
rect 13026 15552 13038 15555
rect 13814 15552 13820 15564
rect 13026 15524 13820 15552
rect 13026 15521 13038 15524
rect 12980 15515 13038 15521
rect 13814 15512 13820 15524
rect 13872 15512 13878 15564
rect 14090 15512 14096 15564
rect 14148 15552 14154 15564
rect 14369 15555 14427 15561
rect 14369 15552 14381 15555
rect 14148 15524 14381 15552
rect 14148 15512 14154 15524
rect 14369 15521 14381 15524
rect 14415 15521 14427 15555
rect 14369 15515 14427 15521
rect 14918 15512 14924 15564
rect 14976 15552 14982 15564
rect 15105 15555 15163 15561
rect 15105 15552 15117 15555
rect 14976 15524 15117 15552
rect 14976 15512 14982 15524
rect 15105 15521 15117 15524
rect 15151 15521 15163 15555
rect 17034 15552 17040 15564
rect 15105 15515 15163 15521
rect 15212 15524 17040 15552
rect 12710 15484 12716 15496
rect 12671 15456 12716 15484
rect 12710 15444 12716 15456
rect 12768 15444 12774 15496
rect 13722 15444 13728 15496
rect 13780 15484 13786 15496
rect 13906 15484 13912 15496
rect 13780 15456 13912 15484
rect 13780 15444 13786 15456
rect 13906 15444 13912 15456
rect 13964 15444 13970 15496
rect 14737 15487 14795 15493
rect 14737 15453 14749 15487
rect 14783 15484 14795 15487
rect 15212 15484 15240 15524
rect 17034 15512 17040 15524
rect 17092 15512 17098 15564
rect 17212 15555 17270 15561
rect 17212 15521 17224 15555
rect 17258 15552 17270 15555
rect 17494 15552 17500 15564
rect 17258 15524 17500 15552
rect 17258 15521 17270 15524
rect 17212 15515 17270 15521
rect 17494 15512 17500 15524
rect 17552 15512 17558 15564
rect 17954 15512 17960 15564
rect 18012 15552 18018 15564
rect 18322 15552 18328 15564
rect 18012 15524 18328 15552
rect 18012 15512 18018 15524
rect 18322 15512 18328 15524
rect 18380 15512 18386 15564
rect 18868 15555 18926 15561
rect 18868 15521 18880 15555
rect 18914 15552 18926 15555
rect 19444 15552 19472 15580
rect 18914 15524 19472 15552
rect 20073 15555 20131 15561
rect 18914 15521 18926 15524
rect 18868 15515 18926 15521
rect 20073 15521 20085 15555
rect 20119 15552 20131 15555
rect 20254 15552 20260 15564
rect 20119 15524 20260 15552
rect 20119 15521 20131 15524
rect 20073 15515 20131 15521
rect 20254 15512 20260 15524
rect 20312 15512 20318 15564
rect 21008 15561 21036 15592
rect 21358 15580 21364 15592
rect 21416 15580 21422 15632
rect 20441 15555 20499 15561
rect 20441 15521 20453 15555
rect 20487 15521 20499 15555
rect 20441 15515 20499 15521
rect 20993 15555 21051 15561
rect 20993 15521 21005 15555
rect 21039 15521 21051 15555
rect 21249 15555 21307 15561
rect 21249 15552 21261 15555
rect 20993 15515 21051 15521
rect 21100 15524 21261 15552
rect 14783 15456 15240 15484
rect 15289 15487 15347 15493
rect 14783 15453 14795 15456
rect 14737 15447 14795 15453
rect 15289 15453 15301 15487
rect 15335 15453 15347 15487
rect 16942 15484 16948 15496
rect 16903 15456 16948 15484
rect 15289 15447 15347 15453
rect 13740 15348 13768 15444
rect 13998 15376 14004 15428
rect 14056 15416 14062 15428
rect 15194 15416 15200 15428
rect 14056 15388 15200 15416
rect 14056 15376 14062 15388
rect 15194 15376 15200 15388
rect 15252 15416 15258 15428
rect 15304 15416 15332 15447
rect 16942 15444 16948 15456
rect 17000 15444 17006 15496
rect 18046 15444 18052 15496
rect 18104 15484 18110 15496
rect 18601 15487 18659 15493
rect 18601 15484 18613 15487
rect 18104 15456 18613 15484
rect 18104 15444 18110 15456
rect 18601 15453 18613 15456
rect 18647 15453 18659 15487
rect 18601 15447 18659 15453
rect 19978 15444 19984 15496
rect 20036 15484 20042 15496
rect 20456 15484 20484 15515
rect 21100 15484 21128 15524
rect 21249 15521 21261 15524
rect 21295 15552 21307 15555
rect 22738 15552 22744 15564
rect 21295 15524 22744 15552
rect 21295 15521 21307 15524
rect 21249 15515 21307 15521
rect 22738 15512 22744 15524
rect 22796 15512 22802 15564
rect 20036 15456 20484 15484
rect 21008 15456 21128 15484
rect 20036 15444 20042 15456
rect 15252 15388 15332 15416
rect 20257 15419 20315 15425
rect 15252 15376 15258 15388
rect 20257 15385 20269 15419
rect 20303 15416 20315 15419
rect 20438 15416 20444 15428
rect 20303 15388 20444 15416
rect 20303 15385 20315 15388
rect 20257 15379 20315 15385
rect 20438 15376 20444 15388
rect 20496 15376 20502 15428
rect 20622 15416 20628 15428
rect 20583 15388 20628 15416
rect 20622 15376 20628 15388
rect 20680 15376 20686 15428
rect 12544 15320 13768 15348
rect 14093 15351 14151 15357
rect 12069 15311 12127 15317
rect 14093 15317 14105 15351
rect 14139 15348 14151 15351
rect 14182 15348 14188 15360
rect 14139 15320 14188 15348
rect 14139 15317 14151 15320
rect 14093 15311 14151 15317
rect 14182 15308 14188 15320
rect 14240 15308 14246 15360
rect 14550 15348 14556 15360
rect 14511 15320 14556 15348
rect 14550 15308 14556 15320
rect 14608 15308 14614 15360
rect 15654 15308 15660 15360
rect 15712 15348 15718 15360
rect 16669 15351 16727 15357
rect 16669 15348 16681 15351
rect 15712 15320 16681 15348
rect 15712 15308 15718 15320
rect 16669 15317 16681 15320
rect 16715 15317 16727 15351
rect 16669 15311 16727 15317
rect 16942 15308 16948 15360
rect 17000 15348 17006 15360
rect 17218 15348 17224 15360
rect 17000 15320 17224 15348
rect 17000 15308 17006 15320
rect 17218 15308 17224 15320
rect 17276 15348 17282 15360
rect 18325 15351 18383 15357
rect 18325 15348 18337 15351
rect 17276 15320 18337 15348
rect 17276 15308 17282 15320
rect 18325 15317 18337 15320
rect 18371 15317 18383 15351
rect 18325 15311 18383 15317
rect 19886 15308 19892 15360
rect 19944 15348 19950 15360
rect 19981 15351 20039 15357
rect 19981 15348 19993 15351
rect 19944 15320 19993 15348
rect 19944 15308 19950 15320
rect 19981 15317 19993 15320
rect 20027 15317 20039 15351
rect 19981 15311 20039 15317
rect 20070 15308 20076 15360
rect 20128 15348 20134 15360
rect 21008 15348 21036 15456
rect 22370 15348 22376 15360
rect 20128 15320 21036 15348
rect 22331 15320 22376 15348
rect 20128 15308 20134 15320
rect 22370 15308 22376 15320
rect 22428 15308 22434 15360
rect 1104 15258 23276 15280
rect 1104 15206 4680 15258
rect 4732 15206 4744 15258
rect 4796 15206 4808 15258
rect 4860 15206 4872 15258
rect 4924 15206 12078 15258
rect 12130 15206 12142 15258
rect 12194 15206 12206 15258
rect 12258 15206 12270 15258
rect 12322 15206 19475 15258
rect 19527 15206 19539 15258
rect 19591 15206 19603 15258
rect 19655 15206 19667 15258
rect 19719 15206 23276 15258
rect 1104 15184 23276 15206
rect 1581 15147 1639 15153
rect 1581 15113 1593 15147
rect 1627 15144 1639 15147
rect 3329 15147 3387 15153
rect 1627 15116 3280 15144
rect 1627 15113 1639 15116
rect 1581 15107 1639 15113
rect 3252 15076 3280 15116
rect 3329 15113 3341 15147
rect 3375 15144 3387 15147
rect 3418 15144 3424 15156
rect 3375 15116 3424 15144
rect 3375 15113 3387 15116
rect 3329 15107 3387 15113
rect 3418 15104 3424 15116
rect 3476 15104 3482 15156
rect 3510 15104 3516 15156
rect 3568 15144 3574 15156
rect 3605 15147 3663 15153
rect 3605 15144 3617 15147
rect 3568 15116 3617 15144
rect 3568 15104 3574 15116
rect 3605 15113 3617 15116
rect 3651 15113 3663 15147
rect 3605 15107 3663 15113
rect 4617 15147 4675 15153
rect 4617 15113 4629 15147
rect 4663 15144 4675 15147
rect 5074 15144 5080 15156
rect 4663 15116 5080 15144
rect 4663 15113 4675 15116
rect 4617 15107 4675 15113
rect 5074 15104 5080 15116
rect 5132 15104 5138 15156
rect 5534 15104 5540 15156
rect 5592 15144 5598 15156
rect 5629 15147 5687 15153
rect 5629 15144 5641 15147
rect 5592 15116 5641 15144
rect 5592 15104 5598 15116
rect 5629 15113 5641 15116
rect 5675 15113 5687 15147
rect 5629 15107 5687 15113
rect 7650 15104 7656 15156
rect 7708 15144 7714 15156
rect 7837 15147 7895 15153
rect 7837 15144 7849 15147
rect 7708 15116 7849 15144
rect 7708 15104 7714 15116
rect 7837 15113 7849 15116
rect 7883 15113 7895 15147
rect 7837 15107 7895 15113
rect 7926 15104 7932 15156
rect 7984 15144 7990 15156
rect 7984 15116 8892 15144
rect 7984 15104 7990 15116
rect 5442 15076 5448 15088
rect 3252 15048 5448 15076
rect 5442 15036 5448 15048
rect 5500 15036 5506 15088
rect 5718 15036 5724 15088
rect 5776 15076 5782 15088
rect 6825 15079 6883 15085
rect 5776 15048 6316 15076
rect 5776 15036 5782 15048
rect 3878 14968 3884 15020
rect 3936 15008 3942 15020
rect 4157 15011 4215 15017
rect 4157 15008 4169 15011
rect 3936 14980 4169 15008
rect 3936 14968 3942 14980
rect 4157 14977 4169 14980
rect 4203 15008 4215 15011
rect 4430 15008 4436 15020
rect 4203 14980 4436 15008
rect 4203 14977 4215 14980
rect 4157 14971 4215 14977
rect 4430 14968 4436 14980
rect 4488 15008 4494 15020
rect 5169 15011 5227 15017
rect 5169 15008 5181 15011
rect 4488 14980 5181 15008
rect 4488 14968 4494 14980
rect 5169 14977 5181 14980
rect 5215 15008 5227 15011
rect 6181 15011 6239 15017
rect 6181 15008 6193 15011
rect 5215 14980 6193 15008
rect 5215 14977 5227 14980
rect 5169 14971 5227 14977
rect 6181 14977 6193 14980
rect 6227 14977 6239 15011
rect 6288 15008 6316 15048
rect 6825 15045 6837 15079
rect 6871 15076 6883 15079
rect 8754 15076 8760 15088
rect 6871 15048 8760 15076
rect 6871 15045 6883 15048
rect 6825 15039 6883 15045
rect 8754 15036 8760 15048
rect 8812 15036 8818 15088
rect 7285 15011 7343 15017
rect 7285 15008 7297 15011
rect 6288 14980 7297 15008
rect 6181 14971 6239 14977
rect 7285 14977 7297 14980
rect 7331 14977 7343 15011
rect 7285 14971 7343 14977
rect 7469 15011 7527 15017
rect 7469 14977 7481 15011
rect 7515 15008 7527 15011
rect 7834 15008 7840 15020
rect 7515 14980 7840 15008
rect 7515 14977 7527 14980
rect 7469 14971 7527 14977
rect 7834 14968 7840 14980
rect 7892 15008 7898 15020
rect 8018 15008 8024 15020
rect 7892 14980 8024 15008
rect 7892 14968 7898 14980
rect 8018 14968 8024 14980
rect 8076 14968 8082 15020
rect 8202 14968 8208 15020
rect 8260 15008 8266 15020
rect 8864 15017 8892 15116
rect 9950 15104 9956 15156
rect 10008 15144 10014 15156
rect 10229 15147 10287 15153
rect 10229 15144 10241 15147
rect 10008 15116 10241 15144
rect 10008 15104 10014 15116
rect 10229 15113 10241 15116
rect 10275 15113 10287 15147
rect 11882 15144 11888 15156
rect 10229 15107 10287 15113
rect 10336 15116 11888 15144
rect 8389 15011 8447 15017
rect 8389 15008 8401 15011
rect 8260 14980 8401 15008
rect 8260 14968 8266 14980
rect 8389 14977 8401 14980
rect 8435 14977 8447 15011
rect 8389 14971 8447 14977
rect 8849 15011 8907 15017
rect 8849 14977 8861 15011
rect 8895 14977 8907 15011
rect 8849 14971 8907 14977
rect 1394 14940 1400 14952
rect 1355 14912 1400 14940
rect 1394 14900 1400 14912
rect 1452 14900 1458 14952
rect 1762 14900 1768 14952
rect 1820 14940 1826 14952
rect 1949 14943 2007 14949
rect 1949 14940 1961 14943
rect 1820 14912 1961 14940
rect 1820 14900 1826 14912
rect 1949 14909 1961 14912
rect 1995 14909 2007 14943
rect 1949 14903 2007 14909
rect 2216 14943 2274 14949
rect 2216 14909 2228 14943
rect 2262 14940 2274 14943
rect 2774 14940 2780 14952
rect 2262 14912 2780 14940
rect 2262 14909 2274 14912
rect 2216 14903 2274 14909
rect 1964 14872 1992 14903
rect 2774 14900 2780 14912
rect 2832 14900 2838 14952
rect 3970 14940 3976 14952
rect 3931 14912 3976 14940
rect 3970 14900 3976 14912
rect 4028 14900 4034 14952
rect 4908 14912 5672 14940
rect 2498 14872 2504 14884
rect 1964 14844 2504 14872
rect 2498 14832 2504 14844
rect 2556 14832 2562 14884
rect 2682 14832 2688 14884
rect 2740 14872 2746 14884
rect 4908 14872 4936 14912
rect 2740 14844 4936 14872
rect 4985 14875 5043 14881
rect 2740 14832 2746 14844
rect 4985 14841 4997 14875
rect 5031 14872 5043 14875
rect 5166 14872 5172 14884
rect 5031 14844 5172 14872
rect 5031 14841 5043 14844
rect 4985 14835 5043 14841
rect 5166 14832 5172 14844
rect 5224 14832 5230 14884
rect 5644 14872 5672 14912
rect 5994 14900 6000 14952
rect 6052 14940 6058 14952
rect 6089 14943 6147 14949
rect 6089 14940 6101 14943
rect 6052 14912 6101 14940
rect 6052 14900 6058 14912
rect 6089 14909 6101 14912
rect 6135 14909 6147 14943
rect 6089 14903 6147 14909
rect 6822 14900 6828 14952
rect 6880 14940 6886 14952
rect 7193 14943 7251 14949
rect 7193 14940 7205 14943
rect 6880 14912 7205 14940
rect 6880 14900 6886 14912
rect 7193 14909 7205 14912
rect 7239 14909 7251 14943
rect 8294 14940 8300 14952
rect 8207 14912 8300 14940
rect 7193 14903 7251 14909
rect 8294 14900 8300 14912
rect 8352 14940 8358 14952
rect 8478 14940 8484 14952
rect 8352 14912 8484 14940
rect 8352 14900 8358 14912
rect 8478 14900 8484 14912
rect 8536 14900 8542 14952
rect 8662 14900 8668 14952
rect 8720 14940 8726 14952
rect 10336 14940 10364 15116
rect 11882 15104 11888 15116
rect 11940 15104 11946 15156
rect 12710 15144 12716 15156
rect 12459 15116 12716 15144
rect 12069 15079 12127 15085
rect 12069 15045 12081 15079
rect 12115 15076 12127 15079
rect 12115 15048 12388 15076
rect 12115 15045 12127 15048
rect 12069 15039 12127 15045
rect 8720 14912 10364 14940
rect 8720 14900 8726 14912
rect 10594 14900 10600 14952
rect 10652 14940 10658 14952
rect 10689 14943 10747 14949
rect 10689 14940 10701 14943
rect 10652 14912 10701 14940
rect 10652 14900 10658 14912
rect 10689 14909 10701 14912
rect 10735 14909 10747 14943
rect 10689 14903 10747 14909
rect 10956 14943 11014 14949
rect 10956 14909 10968 14943
rect 11002 14940 11014 14943
rect 11974 14940 11980 14952
rect 11002 14912 11980 14940
rect 11002 14909 11014 14912
rect 10956 14903 11014 14909
rect 11974 14900 11980 14912
rect 12032 14900 12038 14952
rect 12360 14940 12388 15048
rect 12459 15017 12487 15116
rect 12710 15104 12716 15116
rect 12768 15104 12774 15156
rect 12802 15104 12808 15156
rect 12860 15144 12866 15156
rect 18506 15144 18512 15156
rect 12860 15116 18512 15144
rect 12860 15104 12866 15116
rect 18506 15104 18512 15116
rect 18564 15104 18570 15156
rect 19334 15104 19340 15156
rect 19392 15144 19398 15156
rect 19613 15147 19671 15153
rect 19613 15144 19625 15147
rect 19392 15116 19625 15144
rect 19392 15104 19398 15116
rect 19613 15113 19625 15116
rect 19659 15113 19671 15147
rect 21913 15147 21971 15153
rect 21913 15144 21925 15147
rect 19613 15107 19671 15113
rect 19720 15116 21925 15144
rect 13538 15036 13544 15088
rect 13596 15076 13602 15088
rect 13722 15076 13728 15088
rect 13596 15048 13728 15076
rect 13596 15036 13602 15048
rect 13722 15036 13728 15048
rect 13780 15036 13786 15088
rect 15378 15036 15384 15088
rect 15436 15076 15442 15088
rect 15473 15079 15531 15085
rect 15473 15076 15485 15079
rect 15436 15048 15485 15076
rect 15436 15036 15442 15048
rect 15473 15045 15485 15048
rect 15519 15076 15531 15079
rect 16298 15076 16304 15088
rect 15519 15048 16304 15076
rect 15519 15045 15531 15048
rect 15473 15039 15531 15045
rect 16298 15036 16304 15048
rect 16356 15036 16362 15088
rect 12444 15011 12502 15017
rect 12444 14977 12456 15011
rect 12490 15008 12502 15011
rect 12490 14980 12572 15008
rect 12490 14977 12502 14980
rect 12444 14971 12502 14977
rect 12544 14940 12572 14980
rect 15194 14968 15200 15020
rect 15252 15008 15258 15020
rect 16206 15008 16212 15020
rect 15252 14980 16212 15008
rect 15252 14968 15258 14980
rect 16206 14968 16212 14980
rect 16264 14968 16270 15020
rect 17862 14968 17868 15020
rect 17920 14968 17926 15020
rect 19426 14968 19432 15020
rect 19484 15008 19490 15020
rect 19720 15008 19748 15116
rect 21913 15113 21925 15116
rect 21959 15113 21971 15147
rect 21913 15107 21971 15113
rect 19889 15079 19947 15085
rect 19889 15045 19901 15079
rect 19935 15076 19947 15079
rect 19935 15048 20668 15076
rect 19935 15045 19947 15048
rect 19889 15039 19947 15045
rect 19484 14980 19748 15008
rect 20441 15011 20499 15017
rect 19484 14968 19490 14980
rect 20441 14977 20453 15011
rect 20487 14977 20499 15011
rect 20441 14971 20499 14977
rect 12986 14940 12992 14952
rect 12360 14912 12487 14940
rect 12544 14912 12992 14940
rect 8205 14875 8263 14881
rect 5644 14844 7604 14872
rect 4062 14804 4068 14816
rect 4023 14776 4068 14804
rect 4062 14764 4068 14776
rect 4120 14764 4126 14816
rect 5074 14764 5080 14816
rect 5132 14804 5138 14816
rect 5997 14807 6055 14813
rect 5132 14776 5177 14804
rect 5132 14764 5138 14776
rect 5997 14773 6009 14807
rect 6043 14804 6055 14807
rect 6178 14804 6184 14816
rect 6043 14776 6184 14804
rect 6043 14773 6055 14776
rect 5997 14767 6055 14773
rect 6178 14764 6184 14776
rect 6236 14764 6242 14816
rect 7576 14804 7604 14844
rect 8205 14841 8217 14875
rect 8251 14872 8263 14875
rect 8754 14872 8760 14884
rect 8251 14844 8760 14872
rect 8251 14841 8263 14844
rect 8205 14835 8263 14841
rect 8754 14832 8760 14844
rect 8812 14832 8818 14884
rect 9122 14881 9128 14884
rect 9116 14872 9128 14881
rect 9083 14844 9128 14872
rect 9116 14835 9128 14844
rect 9122 14832 9128 14835
rect 9180 14832 9186 14884
rect 12342 14872 12348 14884
rect 9232 14844 12348 14872
rect 9232 14804 9260 14844
rect 12342 14832 12348 14844
rect 12400 14832 12406 14884
rect 12459 14872 12487 14912
rect 12986 14900 12992 14912
rect 13044 14940 13050 14952
rect 13998 14940 14004 14952
rect 13044 14912 14004 14940
rect 13044 14900 13050 14912
rect 13998 14900 14004 14912
rect 14056 14940 14062 14952
rect 14093 14943 14151 14949
rect 14093 14940 14105 14943
rect 14056 14912 14105 14940
rect 14056 14900 14062 14912
rect 14093 14909 14105 14912
rect 14139 14909 14151 14943
rect 14093 14903 14151 14909
rect 14182 14900 14188 14952
rect 14240 14940 14246 14952
rect 14360 14943 14418 14949
rect 14360 14940 14372 14943
rect 14240 14912 14372 14940
rect 14240 14900 14246 14912
rect 14360 14909 14372 14912
rect 14406 14940 14418 14943
rect 15378 14940 15384 14952
rect 14406 14912 15384 14940
rect 14406 14909 14418 14912
rect 14360 14903 14418 14909
rect 15378 14900 15384 14912
rect 15436 14900 15442 14952
rect 15746 14900 15752 14952
rect 15804 14940 15810 14952
rect 15804 14912 15849 14940
rect 15804 14900 15810 14912
rect 15930 14900 15936 14952
rect 15988 14940 15994 14952
rect 16301 14943 16359 14949
rect 16301 14940 16313 14943
rect 15988 14912 16313 14940
rect 15988 14900 15994 14912
rect 16301 14909 16313 14912
rect 16347 14909 16359 14943
rect 16301 14903 16359 14909
rect 16568 14943 16626 14949
rect 16568 14909 16580 14943
rect 16614 14940 16626 14943
rect 17880 14940 17908 14968
rect 16614 14912 17908 14940
rect 16614 14909 16626 14912
rect 16568 14903 16626 14909
rect 18046 14900 18052 14952
rect 18104 14940 18110 14952
rect 18233 14943 18291 14949
rect 18233 14940 18245 14943
rect 18104 14912 18245 14940
rect 18104 14900 18110 14912
rect 18233 14909 18245 14912
rect 18279 14909 18291 14943
rect 20349 14943 20407 14949
rect 20349 14940 20361 14943
rect 18233 14903 18291 14909
rect 18331 14912 20361 14940
rect 12704 14875 12762 14881
rect 12704 14872 12716 14875
rect 12459 14844 12716 14872
rect 12704 14841 12716 14844
rect 12750 14872 12762 14875
rect 13538 14872 13544 14884
rect 12750 14844 13544 14872
rect 12750 14841 12762 14844
rect 12704 14835 12762 14841
rect 13538 14832 13544 14844
rect 13596 14832 13602 14884
rect 13906 14832 13912 14884
rect 13964 14872 13970 14884
rect 13964 14844 14872 14872
rect 13964 14832 13970 14844
rect 7576 14776 9260 14804
rect 10134 14764 10140 14816
rect 10192 14804 10198 14816
rect 13446 14804 13452 14816
rect 10192 14776 13452 14804
rect 10192 14764 10198 14776
rect 13446 14764 13452 14776
rect 13504 14764 13510 14816
rect 13814 14804 13820 14816
rect 13775 14776 13820 14804
rect 13814 14764 13820 14776
rect 13872 14764 13878 14816
rect 14182 14764 14188 14816
rect 14240 14804 14246 14816
rect 14734 14804 14740 14816
rect 14240 14776 14740 14804
rect 14240 14764 14246 14776
rect 14734 14764 14740 14776
rect 14792 14764 14798 14816
rect 14844 14804 14872 14844
rect 15286 14832 15292 14884
rect 15344 14872 15350 14884
rect 16666 14872 16672 14884
rect 15344 14844 16672 14872
rect 15344 14832 15350 14844
rect 16666 14832 16672 14844
rect 16724 14832 16730 14884
rect 17218 14832 17224 14884
rect 17276 14872 17282 14884
rect 17276 14844 17816 14872
rect 17276 14832 17282 14844
rect 15654 14804 15660 14816
rect 14844 14776 15660 14804
rect 15654 14764 15660 14776
rect 15712 14764 15718 14816
rect 15933 14807 15991 14813
rect 15933 14773 15945 14807
rect 15979 14804 15991 14807
rect 16574 14804 16580 14816
rect 15979 14776 16580 14804
rect 15979 14773 15991 14776
rect 15933 14767 15991 14773
rect 16574 14764 16580 14776
rect 16632 14764 16638 14816
rect 16758 14764 16764 14816
rect 16816 14804 16822 14816
rect 17494 14804 17500 14816
rect 16816 14776 17500 14804
rect 16816 14764 16822 14776
rect 17494 14764 17500 14776
rect 17552 14804 17558 14816
rect 17681 14807 17739 14813
rect 17681 14804 17693 14807
rect 17552 14776 17693 14804
rect 17552 14764 17558 14776
rect 17681 14773 17693 14776
rect 17727 14773 17739 14807
rect 17788 14804 17816 14844
rect 17862 14832 17868 14884
rect 17920 14872 17926 14884
rect 18331 14872 18359 14912
rect 20349 14909 20361 14912
rect 20395 14909 20407 14943
rect 20349 14903 20407 14909
rect 17920 14844 18359 14872
rect 18500 14875 18558 14881
rect 17920 14832 17926 14844
rect 18500 14841 18512 14875
rect 18546 14872 18558 14875
rect 19058 14872 19064 14884
rect 18546 14844 19064 14872
rect 18546 14841 18558 14844
rect 18500 14835 18558 14841
rect 19058 14832 19064 14844
rect 19116 14832 19122 14884
rect 19886 14832 19892 14884
rect 19944 14872 19950 14884
rect 20456 14872 20484 14971
rect 20640 14940 20668 15048
rect 20717 15011 20775 15017
rect 20717 14977 20729 15011
rect 20763 15008 20775 15011
rect 21453 15011 21511 15017
rect 21453 15008 21465 15011
rect 20763 14980 21465 15008
rect 20763 14977 20775 14980
rect 20717 14971 20775 14977
rect 21453 14977 21465 14980
rect 21499 15008 21511 15011
rect 22465 15011 22523 15017
rect 22465 15008 22477 15011
rect 21499 14980 22477 15008
rect 21499 14977 21511 14980
rect 21453 14971 21511 14977
rect 22465 14977 22477 14980
rect 22511 14977 22523 15011
rect 22465 14971 22523 14977
rect 21269 14943 21327 14949
rect 21269 14940 21281 14943
rect 20640 14912 21281 14940
rect 21269 14909 21281 14912
rect 21315 14909 21327 14943
rect 21269 14903 21327 14909
rect 19944 14844 20484 14872
rect 19944 14832 19950 14844
rect 21726 14832 21732 14884
rect 21784 14872 21790 14884
rect 22373 14875 22431 14881
rect 22373 14872 22385 14875
rect 21784 14844 22385 14872
rect 21784 14832 21790 14844
rect 22373 14841 22385 14844
rect 22419 14841 22431 14875
rect 22373 14835 22431 14841
rect 20257 14807 20315 14813
rect 20257 14804 20269 14807
rect 17788 14776 20269 14804
rect 17681 14767 17739 14773
rect 20257 14773 20269 14776
rect 20303 14773 20315 14807
rect 20257 14767 20315 14773
rect 20438 14764 20444 14816
rect 20496 14804 20502 14816
rect 20717 14807 20775 14813
rect 20717 14804 20729 14807
rect 20496 14776 20729 14804
rect 20496 14764 20502 14776
rect 20717 14773 20729 14776
rect 20763 14773 20775 14807
rect 20898 14804 20904 14816
rect 20859 14776 20904 14804
rect 20717 14767 20775 14773
rect 20898 14764 20904 14776
rect 20956 14764 20962 14816
rect 21358 14804 21364 14816
rect 21319 14776 21364 14804
rect 21358 14764 21364 14776
rect 21416 14764 21422 14816
rect 22278 14804 22284 14816
rect 22239 14776 22284 14804
rect 22278 14764 22284 14776
rect 22336 14764 22342 14816
rect 1104 14714 23276 14736
rect 1104 14662 8379 14714
rect 8431 14662 8443 14714
rect 8495 14662 8507 14714
rect 8559 14662 8571 14714
rect 8623 14662 15776 14714
rect 15828 14662 15840 14714
rect 15892 14662 15904 14714
rect 15956 14662 15968 14714
rect 16020 14662 23276 14714
rect 1104 14640 23276 14662
rect 1762 14560 1768 14612
rect 1820 14560 1826 14612
rect 3605 14603 3663 14609
rect 3605 14569 3617 14603
rect 3651 14569 3663 14603
rect 3605 14563 3663 14569
rect 1780 14532 1808 14560
rect 1504 14504 1808 14532
rect 1504 14473 1532 14504
rect 3142 14492 3148 14544
rect 3200 14532 3206 14544
rect 3620 14532 3648 14563
rect 4982 14560 4988 14612
rect 5040 14600 5046 14612
rect 5040 14572 5856 14600
rect 5040 14560 5046 14572
rect 5718 14532 5724 14544
rect 3200 14504 3464 14532
rect 3620 14504 5724 14532
rect 3200 14492 3206 14504
rect 1489 14467 1547 14473
rect 1489 14433 1501 14467
rect 1535 14433 1547 14467
rect 1489 14427 1547 14433
rect 1756 14467 1814 14473
rect 1756 14433 1768 14467
rect 1802 14464 1814 14467
rect 2038 14464 2044 14476
rect 1802 14436 2044 14464
rect 1802 14433 1814 14436
rect 1756 14427 1814 14433
rect 2038 14424 2044 14436
rect 2096 14424 2102 14476
rect 3436 14473 3464 14504
rect 5718 14492 5724 14504
rect 5776 14492 5782 14544
rect 5828 14532 5856 14572
rect 6178 14560 6184 14612
rect 6236 14600 6242 14612
rect 7101 14603 7159 14609
rect 7101 14600 7113 14603
rect 6236 14572 7113 14600
rect 6236 14560 6242 14572
rect 7101 14569 7113 14572
rect 7147 14569 7159 14603
rect 7101 14563 7159 14569
rect 7377 14603 7435 14609
rect 7377 14569 7389 14603
rect 7423 14600 7435 14603
rect 8202 14600 8208 14612
rect 7423 14572 8208 14600
rect 7423 14569 7435 14572
rect 7377 14563 7435 14569
rect 8202 14560 8208 14572
rect 8260 14560 8266 14612
rect 9122 14560 9128 14612
rect 9180 14600 9186 14612
rect 11054 14600 11060 14612
rect 9180 14572 11060 14600
rect 9180 14560 9186 14572
rect 11054 14560 11060 14572
rect 11112 14560 11118 14612
rect 11330 14560 11336 14612
rect 11388 14600 11394 14612
rect 12526 14600 12532 14612
rect 11388 14572 12532 14600
rect 11388 14560 11394 14572
rect 12526 14560 12532 14572
rect 12584 14560 12590 14612
rect 12897 14603 12955 14609
rect 12897 14569 12909 14603
rect 12943 14600 12955 14603
rect 14182 14600 14188 14612
rect 12943 14572 14188 14600
rect 12943 14569 12955 14572
rect 12897 14563 12955 14569
rect 8662 14532 8668 14544
rect 5828 14504 8668 14532
rect 8662 14492 8668 14504
rect 8720 14492 8726 14544
rect 9944 14535 10002 14541
rect 9944 14501 9956 14535
rect 9990 14532 10002 14535
rect 12912 14532 12940 14563
rect 14182 14560 14188 14572
rect 14240 14560 14246 14612
rect 14277 14603 14335 14609
rect 14277 14569 14289 14603
rect 14323 14600 14335 14603
rect 15749 14603 15807 14609
rect 15749 14600 15761 14603
rect 14323 14572 15761 14600
rect 14323 14569 14335 14572
rect 14277 14563 14335 14569
rect 15749 14569 15761 14572
rect 15795 14569 15807 14603
rect 16114 14600 16120 14612
rect 16075 14572 16120 14600
rect 15749 14563 15807 14569
rect 16114 14560 16120 14572
rect 16172 14560 16178 14612
rect 16945 14603 17003 14609
rect 16945 14569 16957 14603
rect 16991 14600 17003 14603
rect 17310 14600 17316 14612
rect 16991 14572 17316 14600
rect 16991 14569 17003 14572
rect 16945 14563 17003 14569
rect 17310 14560 17316 14572
rect 17368 14560 17374 14612
rect 18506 14560 18512 14612
rect 18564 14600 18570 14612
rect 19426 14600 19432 14612
rect 18564 14572 19432 14600
rect 18564 14560 18570 14572
rect 19426 14560 19432 14572
rect 19484 14560 19490 14612
rect 19521 14603 19579 14609
rect 19521 14569 19533 14603
rect 19567 14600 19579 14603
rect 21358 14600 21364 14612
rect 19567 14572 21364 14600
rect 19567 14569 19579 14572
rect 19521 14563 19579 14569
rect 21358 14560 21364 14572
rect 21416 14560 21422 14612
rect 21634 14560 21640 14612
rect 21692 14600 21698 14612
rect 22557 14603 22615 14609
rect 22557 14600 22569 14603
rect 21692 14572 22569 14600
rect 21692 14560 21698 14572
rect 22557 14569 22569 14572
rect 22603 14569 22615 14603
rect 22557 14563 22615 14569
rect 9990 14504 12940 14532
rect 9990 14501 10002 14504
rect 9944 14495 10002 14501
rect 13078 14492 13084 14544
rect 13136 14532 13142 14544
rect 13817 14535 13875 14541
rect 13817 14532 13829 14535
rect 13136 14504 13829 14532
rect 13136 14492 13142 14504
rect 13817 14501 13829 14504
rect 13863 14501 13875 14535
rect 13817 14495 13875 14501
rect 13909 14535 13967 14541
rect 13909 14501 13921 14535
rect 13955 14532 13967 14535
rect 13998 14532 14004 14544
rect 13955 14504 14004 14532
rect 13955 14501 13967 14504
rect 13909 14495 13967 14501
rect 13998 14492 14004 14504
rect 14056 14492 14062 14544
rect 14737 14535 14795 14541
rect 14737 14532 14749 14535
rect 14099 14504 14749 14532
rect 3329 14467 3387 14473
rect 3329 14433 3341 14467
rect 3375 14433 3387 14467
rect 3329 14427 3387 14433
rect 3421 14467 3479 14473
rect 3421 14433 3433 14467
rect 3467 14433 3479 14467
rect 4154 14464 4160 14476
rect 3421 14427 3479 14433
rect 3988 14436 4160 14464
rect 3344 14396 3372 14427
rect 3988 14396 4016 14436
rect 4154 14424 4160 14436
rect 4212 14424 4218 14476
rect 4332 14467 4390 14473
rect 4332 14433 4344 14467
rect 4378 14464 4390 14467
rect 5074 14464 5080 14476
rect 4378 14436 5080 14464
rect 4378 14433 4390 14436
rect 4332 14427 4390 14433
rect 5074 14424 5080 14436
rect 5132 14424 5138 14476
rect 5994 14473 6000 14476
rect 5988 14464 6000 14473
rect 5955 14436 6000 14464
rect 5988 14427 6000 14436
rect 5994 14424 6000 14427
rect 6052 14424 6058 14476
rect 7742 14464 7748 14476
rect 7703 14436 7748 14464
rect 7742 14424 7748 14436
rect 7800 14424 7806 14476
rect 8018 14424 8024 14476
rect 8076 14424 8082 14476
rect 8754 14464 8760 14476
rect 8715 14436 8760 14464
rect 8754 14424 8760 14436
rect 8812 14424 8818 14476
rect 11330 14464 11336 14476
rect 8956 14436 11336 14464
rect 3344 14368 4016 14396
rect 4065 14399 4123 14405
rect 4065 14365 4077 14399
rect 4111 14365 4123 14399
rect 5350 14396 5356 14408
rect 4065 14359 4123 14365
rect 5092 14368 5356 14396
rect 2498 14288 2504 14340
rect 2556 14328 2562 14340
rect 2556 14300 3004 14328
rect 2556 14288 2562 14300
rect 2130 14220 2136 14272
rect 2188 14260 2194 14272
rect 2869 14263 2927 14269
rect 2869 14260 2881 14263
rect 2188 14232 2881 14260
rect 2188 14220 2194 14232
rect 2869 14229 2881 14232
rect 2915 14229 2927 14263
rect 2976 14260 3004 14300
rect 3145 14263 3203 14269
rect 3145 14260 3157 14263
rect 2976 14232 3157 14260
rect 2869 14223 2927 14229
rect 3145 14229 3157 14232
rect 3191 14260 3203 14263
rect 3602 14260 3608 14272
rect 3191 14232 3608 14260
rect 3191 14229 3203 14232
rect 3145 14223 3203 14229
rect 3602 14220 3608 14232
rect 3660 14260 3666 14272
rect 4080 14260 4108 14359
rect 4246 14260 4252 14272
rect 3660 14232 4252 14260
rect 3660 14220 3666 14232
rect 4246 14220 4252 14232
rect 4304 14260 4310 14272
rect 5092 14260 5120 14368
rect 5350 14356 5356 14368
rect 5408 14396 5414 14408
rect 5721 14399 5779 14405
rect 5721 14396 5733 14399
rect 5408 14368 5733 14396
rect 5408 14356 5414 14368
rect 5721 14365 5733 14368
rect 5767 14365 5779 14399
rect 5721 14359 5779 14365
rect 7837 14399 7895 14405
rect 7837 14365 7849 14399
rect 7883 14365 7895 14399
rect 7837 14359 7895 14365
rect 7929 14399 7987 14405
rect 7929 14365 7941 14399
rect 7975 14396 7987 14399
rect 8036 14396 8064 14424
rect 7975 14368 8064 14396
rect 7975 14365 7987 14368
rect 7929 14359 7987 14365
rect 5258 14288 5264 14340
rect 5316 14328 5322 14340
rect 5316 14300 5580 14328
rect 5316 14288 5322 14300
rect 4304 14232 5120 14260
rect 4304 14220 4310 14232
rect 5166 14220 5172 14272
rect 5224 14260 5230 14272
rect 5442 14260 5448 14272
rect 5224 14232 5448 14260
rect 5224 14220 5230 14232
rect 5442 14220 5448 14232
rect 5500 14220 5506 14272
rect 5552 14260 5580 14300
rect 7852 14260 7880 14359
rect 8662 14356 8668 14408
rect 8720 14396 8726 14408
rect 8849 14399 8907 14405
rect 8849 14396 8861 14399
rect 8720 14368 8861 14396
rect 8720 14356 8726 14368
rect 8849 14365 8861 14368
rect 8895 14365 8907 14399
rect 8849 14359 8907 14365
rect 8018 14288 8024 14340
rect 8076 14328 8082 14340
rect 8956 14328 8984 14436
rect 11330 14424 11336 14436
rect 11388 14424 11394 14476
rect 11784 14467 11842 14473
rect 11784 14433 11796 14467
rect 11830 14464 11842 14467
rect 12526 14464 12532 14476
rect 11830 14436 12532 14464
rect 11830 14433 11842 14436
rect 11784 14427 11842 14433
rect 12526 14424 12532 14436
rect 12584 14424 12590 14476
rect 12989 14467 13047 14473
rect 12989 14433 13001 14467
rect 13035 14464 13047 14467
rect 13170 14464 13176 14476
rect 13035 14436 13176 14464
rect 13035 14433 13047 14436
rect 12989 14427 13047 14433
rect 13170 14424 13176 14436
rect 13228 14424 13234 14476
rect 13357 14467 13415 14473
rect 13357 14433 13369 14467
rect 13403 14464 13415 14467
rect 14099 14464 14127 14504
rect 14737 14501 14749 14504
rect 14783 14501 14795 14535
rect 14737 14495 14795 14501
rect 14826 14492 14832 14544
rect 14884 14532 14890 14544
rect 16485 14535 16543 14541
rect 16485 14532 16497 14535
rect 14884 14504 16497 14532
rect 14884 14492 14890 14504
rect 16485 14501 16497 14504
rect 16531 14501 16543 14535
rect 16485 14495 16543 14501
rect 17126 14492 17132 14544
rect 17184 14532 17190 14544
rect 18046 14532 18052 14544
rect 17184 14504 17520 14532
rect 17184 14492 17190 14504
rect 13403 14436 14127 14464
rect 14645 14467 14703 14473
rect 13403 14433 13415 14436
rect 13357 14427 13415 14433
rect 14645 14433 14657 14467
rect 14691 14433 14703 14467
rect 14645 14427 14703 14433
rect 9033 14399 9091 14405
rect 9033 14365 9045 14399
rect 9079 14396 9091 14399
rect 9079 14368 9628 14396
rect 9079 14365 9091 14368
rect 9033 14359 9091 14365
rect 8076 14300 8984 14328
rect 8076 14288 8082 14300
rect 5552 14232 7880 14260
rect 8389 14263 8447 14269
rect 8389 14229 8401 14263
rect 8435 14260 8447 14263
rect 8846 14260 8852 14272
rect 8435 14232 8852 14260
rect 8435 14229 8447 14232
rect 8389 14223 8447 14229
rect 8846 14220 8852 14232
rect 8904 14220 8910 14272
rect 9600 14260 9628 14368
rect 9674 14356 9680 14408
rect 9732 14396 9738 14408
rect 11517 14399 11575 14405
rect 9732 14368 9777 14396
rect 9732 14356 9738 14368
rect 11517 14365 11529 14399
rect 11563 14365 11575 14399
rect 11517 14359 11575 14365
rect 10962 14288 10968 14340
rect 11020 14328 11026 14340
rect 11330 14328 11336 14340
rect 11020 14300 11336 14328
rect 11020 14288 11026 14300
rect 11330 14288 11336 14300
rect 11388 14328 11394 14340
rect 11532 14328 11560 14359
rect 12710 14356 12716 14408
rect 12768 14396 12774 14408
rect 14090 14396 14096 14408
rect 12768 14368 13575 14396
rect 14051 14368 14096 14396
rect 12768 14356 12774 14368
rect 11388 14300 11560 14328
rect 11388 14288 11394 14300
rect 12802 14288 12808 14340
rect 12860 14328 12866 14340
rect 13446 14328 13452 14340
rect 12860 14300 13299 14328
rect 13407 14300 13452 14328
rect 12860 14288 12866 14300
rect 10410 14260 10416 14272
rect 9600 14232 10416 14260
rect 10410 14220 10416 14232
rect 10468 14220 10474 14272
rect 11514 14220 11520 14272
rect 11572 14260 11578 14272
rect 13173 14263 13231 14269
rect 13173 14260 13185 14263
rect 11572 14232 13185 14260
rect 11572 14220 11578 14232
rect 13173 14229 13185 14232
rect 13219 14229 13231 14263
rect 13271 14260 13299 14300
rect 13446 14288 13452 14300
rect 13504 14288 13510 14340
rect 13547 14328 13575 14368
rect 14090 14356 14096 14368
rect 14148 14356 14154 14408
rect 14660 14328 14688 14427
rect 15010 14424 15016 14476
rect 15068 14464 15074 14476
rect 15657 14467 15715 14473
rect 15657 14464 15669 14467
rect 15068 14436 15669 14464
rect 15068 14424 15074 14436
rect 15657 14433 15669 14436
rect 15703 14433 15715 14467
rect 15657 14427 15715 14433
rect 16298 14424 16304 14476
rect 16356 14464 16362 14476
rect 17313 14467 17371 14473
rect 17313 14464 17325 14467
rect 16356 14436 17325 14464
rect 16356 14424 16362 14436
rect 17313 14433 17325 14436
rect 17359 14433 17371 14467
rect 17313 14427 17371 14433
rect 14921 14399 14979 14405
rect 14921 14365 14933 14399
rect 14967 14365 14979 14399
rect 15841 14399 15899 14405
rect 15841 14396 15853 14399
rect 14921 14359 14979 14365
rect 15028 14368 15853 14396
rect 13547 14300 14688 14328
rect 14826 14288 14832 14340
rect 14884 14328 14890 14340
rect 14936 14328 14964 14359
rect 14884 14300 14964 14328
rect 14884 14288 14890 14300
rect 13357 14263 13415 14269
rect 13357 14260 13369 14263
rect 13271 14232 13369 14260
rect 13173 14223 13231 14229
rect 13357 14229 13369 14232
rect 13403 14229 13415 14263
rect 13357 14223 13415 14229
rect 14182 14220 14188 14272
rect 14240 14260 14246 14272
rect 15028 14260 15056 14368
rect 15841 14365 15853 14368
rect 15887 14365 15899 14399
rect 16574 14396 16580 14408
rect 16535 14368 16580 14396
rect 15841 14359 15899 14365
rect 16574 14356 16580 14368
rect 16632 14356 16638 14408
rect 16666 14356 16672 14408
rect 16724 14396 16730 14408
rect 17492 14405 17520 14504
rect 17880 14504 18052 14532
rect 17880 14473 17908 14504
rect 18046 14492 18052 14504
rect 18104 14532 18110 14544
rect 18874 14532 18880 14544
rect 18104 14504 18880 14532
rect 18104 14492 18110 14504
rect 18874 14492 18880 14504
rect 18932 14492 18938 14544
rect 19889 14535 19947 14541
rect 19889 14532 19901 14535
rect 19812 14504 19901 14532
rect 17865 14467 17923 14473
rect 17865 14433 17877 14467
rect 17911 14433 17923 14467
rect 17865 14427 17923 14433
rect 18132 14467 18190 14473
rect 18132 14433 18144 14467
rect 18178 14464 18190 14467
rect 19242 14464 19248 14476
rect 18178 14436 19248 14464
rect 18178 14433 18190 14436
rect 18132 14427 18190 14433
rect 19242 14424 19248 14436
rect 19300 14424 19306 14476
rect 19426 14424 19432 14476
rect 19484 14464 19490 14476
rect 19812 14464 19840 14504
rect 19889 14501 19901 14504
rect 19935 14501 19947 14535
rect 19889 14495 19947 14501
rect 19981 14535 20039 14541
rect 19981 14501 19993 14535
rect 20027 14532 20039 14535
rect 20070 14532 20076 14544
rect 20027 14504 20076 14532
rect 20027 14501 20039 14504
rect 19981 14495 20039 14501
rect 20070 14492 20076 14504
rect 20128 14492 20134 14544
rect 21444 14535 21502 14541
rect 21444 14501 21456 14535
rect 21490 14532 21502 14535
rect 22370 14532 22376 14544
rect 21490 14504 22376 14532
rect 21490 14501 21502 14504
rect 21444 14495 21502 14501
rect 20714 14464 20720 14476
rect 19484 14436 19840 14464
rect 20675 14436 20720 14464
rect 19484 14424 19490 14436
rect 20714 14424 20720 14436
rect 20772 14424 20778 14476
rect 17405 14399 17463 14405
rect 16724 14368 16769 14396
rect 16724 14356 16730 14368
rect 17405 14365 17417 14399
rect 17451 14365 17463 14399
rect 17492 14399 17555 14405
rect 17492 14368 17509 14399
rect 17405 14359 17463 14365
rect 17497 14365 17509 14368
rect 17543 14365 17555 14399
rect 17497 14359 17555 14365
rect 15102 14288 15108 14340
rect 15160 14328 15166 14340
rect 15289 14331 15347 14337
rect 15289 14328 15301 14331
rect 15160 14300 15301 14328
rect 15160 14288 15166 14300
rect 15289 14297 15301 14300
rect 15335 14297 15347 14331
rect 15289 14291 15347 14297
rect 15378 14288 15384 14340
rect 15436 14328 15442 14340
rect 17420 14328 17448 14359
rect 18874 14356 18880 14408
rect 18932 14396 18938 14408
rect 19337 14399 19395 14405
rect 19337 14396 19349 14399
rect 18932 14368 19349 14396
rect 18932 14356 18938 14368
rect 19337 14365 19349 14368
rect 19383 14365 19395 14399
rect 19337 14359 19395 14365
rect 19886 14356 19892 14408
rect 19944 14396 19950 14408
rect 20073 14399 20131 14405
rect 20073 14396 20085 14399
rect 19944 14368 20085 14396
rect 19944 14356 19950 14368
rect 20073 14365 20085 14368
rect 20119 14365 20131 14399
rect 21177 14399 21235 14405
rect 21177 14396 21189 14399
rect 20073 14359 20131 14365
rect 21100 14368 21189 14396
rect 20990 14328 20996 14340
rect 15436 14300 17448 14328
rect 18791 14300 20996 14328
rect 15436 14288 15442 14300
rect 14240 14232 15056 14260
rect 14240 14220 14246 14232
rect 15654 14220 15660 14272
rect 15712 14260 15718 14272
rect 16114 14260 16120 14272
rect 15712 14232 16120 14260
rect 15712 14220 15718 14232
rect 16114 14220 16120 14232
rect 16172 14220 16178 14272
rect 17310 14220 17316 14272
rect 17368 14260 17374 14272
rect 18791 14260 18819 14300
rect 20990 14288 20996 14300
rect 21048 14288 21054 14340
rect 17368 14232 18819 14260
rect 17368 14220 17374 14232
rect 19058 14220 19064 14272
rect 19116 14260 19122 14272
rect 19245 14263 19303 14269
rect 19245 14260 19257 14263
rect 19116 14232 19257 14260
rect 19116 14220 19122 14232
rect 19245 14229 19257 14232
rect 19291 14229 19303 14263
rect 19245 14223 19303 14229
rect 19337 14263 19395 14269
rect 19337 14229 19349 14263
rect 19383 14260 19395 14263
rect 20533 14263 20591 14269
rect 20533 14260 20545 14263
rect 19383 14232 20545 14260
rect 19383 14229 19395 14232
rect 19337 14223 19395 14229
rect 20533 14229 20545 14232
rect 20579 14260 20591 14263
rect 21100 14260 21128 14368
rect 21177 14365 21189 14368
rect 21223 14365 21235 14399
rect 21177 14359 21235 14365
rect 21358 14260 21364 14272
rect 20579 14232 21364 14260
rect 20579 14229 20591 14232
rect 20533 14223 20591 14229
rect 21358 14220 21364 14232
rect 21416 14220 21422 14272
rect 22094 14220 22100 14272
rect 22152 14260 22158 14272
rect 22204 14260 22232 14504
rect 22370 14492 22376 14504
rect 22428 14492 22434 14544
rect 22152 14232 22232 14260
rect 22152 14220 22158 14232
rect 1104 14170 23276 14192
rect 1104 14118 4680 14170
rect 4732 14118 4744 14170
rect 4796 14118 4808 14170
rect 4860 14118 4872 14170
rect 4924 14118 12078 14170
rect 12130 14118 12142 14170
rect 12194 14118 12206 14170
rect 12258 14118 12270 14170
rect 12322 14118 19475 14170
rect 19527 14118 19539 14170
rect 19591 14118 19603 14170
rect 19655 14118 19667 14170
rect 19719 14118 23276 14170
rect 1104 14096 23276 14118
rect 5074 14056 5080 14068
rect 1504 14028 4936 14056
rect 5035 14028 5080 14056
rect 1504 13861 1532 14028
rect 1670 13988 1676 14000
rect 1631 13960 1676 13988
rect 1670 13948 1676 13960
rect 1728 13948 1734 14000
rect 3421 13991 3479 13997
rect 3421 13957 3433 13991
rect 3467 13957 3479 13991
rect 3421 13951 3479 13957
rect 3436 13920 3464 13951
rect 4908 13920 4936 14028
rect 5074 14016 5080 14028
rect 5132 14016 5138 14068
rect 8662 14056 8668 14068
rect 5460 14028 7972 14056
rect 8623 14028 8668 14056
rect 5166 13948 5172 14000
rect 5224 13988 5230 14000
rect 5353 13991 5411 13997
rect 5353 13988 5365 13991
rect 5224 13960 5365 13988
rect 5224 13948 5230 13960
rect 5353 13957 5365 13960
rect 5399 13957 5411 13991
rect 5353 13951 5411 13957
rect 5460 13920 5488 14028
rect 6178 13948 6184 14000
rect 6236 13988 6242 14000
rect 6454 13988 6460 14000
rect 6236 13960 6460 13988
rect 6236 13948 6242 13960
rect 6454 13948 6460 13960
rect 6512 13948 6518 14000
rect 7944 13988 7972 14028
rect 8662 14016 8668 14028
rect 8720 14016 8726 14068
rect 11698 14056 11704 14068
rect 8772 14028 11704 14056
rect 8772 13988 8800 14028
rect 11698 14016 11704 14028
rect 11756 14016 11762 14068
rect 11977 14059 12035 14065
rect 11977 14025 11989 14059
rect 12023 14056 12035 14059
rect 12710 14056 12716 14068
rect 12023 14028 12716 14056
rect 12023 14025 12035 14028
rect 11977 14019 12035 14025
rect 12710 14016 12716 14028
rect 12768 14016 12774 14068
rect 15010 14056 15016 14068
rect 12820 14028 15016 14056
rect 9306 13988 9312 14000
rect 7944 13960 8800 13988
rect 9219 13960 9312 13988
rect 3436 13892 3832 13920
rect 4908 13892 5488 13920
rect 5997 13923 6055 13929
rect 1489 13855 1547 13861
rect 1489 13821 1501 13855
rect 1535 13821 1547 13855
rect 1489 13815 1547 13821
rect 2041 13855 2099 13861
rect 2041 13821 2053 13855
rect 2087 13821 2099 13855
rect 2041 13815 2099 13821
rect 2308 13855 2366 13861
rect 2308 13821 2320 13855
rect 2354 13852 2366 13855
rect 3050 13852 3056 13864
rect 2354 13824 3056 13852
rect 2354 13821 2366 13824
rect 2308 13815 2366 13821
rect 1670 13744 1676 13796
rect 1728 13784 1734 13796
rect 2056 13784 2084 13815
rect 3050 13812 3056 13824
rect 3108 13812 3114 13864
rect 3602 13812 3608 13864
rect 3660 13852 3666 13864
rect 3697 13855 3755 13861
rect 3697 13852 3709 13855
rect 3660 13824 3709 13852
rect 3660 13812 3666 13824
rect 3697 13821 3709 13824
rect 3743 13821 3755 13855
rect 3804 13852 3832 13892
rect 5997 13889 6009 13923
rect 6043 13920 6055 13923
rect 6362 13920 6368 13932
rect 6043 13892 6368 13920
rect 6043 13889 6055 13892
rect 5997 13883 6055 13889
rect 6362 13880 6368 13892
rect 6420 13880 6426 13932
rect 9232 13929 9260 13960
rect 9306 13948 9312 13960
rect 9364 13988 9370 14000
rect 9769 13991 9827 13997
rect 9364 13960 9700 13988
rect 9364 13948 9370 13960
rect 9217 13923 9275 13929
rect 9217 13889 9229 13923
rect 9263 13889 9275 13923
rect 9672 13920 9700 13960
rect 9769 13957 9781 13991
rect 9815 13988 9827 13991
rect 11790 13988 11796 14000
rect 9815 13960 11796 13988
rect 9815 13957 9827 13960
rect 9769 13951 9827 13957
rect 11790 13948 11796 13960
rect 11848 13948 11854 14000
rect 12437 13991 12495 13997
rect 12437 13988 12449 13991
rect 11900 13960 12449 13988
rect 10410 13920 10416 13932
rect 9672 13892 10272 13920
rect 10371 13892 10416 13920
rect 9217 13883 9275 13889
rect 3970 13861 3976 13864
rect 3964 13852 3976 13861
rect 3804 13824 3976 13852
rect 3697 13815 3755 13821
rect 3964 13815 3976 13824
rect 3970 13812 3976 13815
rect 4028 13812 4034 13864
rect 5350 13812 5356 13864
rect 5408 13852 5414 13864
rect 7009 13855 7067 13861
rect 7009 13852 7021 13855
rect 5408 13824 7021 13852
rect 5408 13812 5414 13824
rect 7009 13821 7021 13824
rect 7055 13821 7067 13855
rect 7009 13815 7067 13821
rect 7276 13855 7334 13861
rect 7276 13821 7288 13855
rect 7322 13852 7334 13855
rect 7558 13852 7564 13864
rect 7322 13824 7564 13852
rect 7322 13821 7334 13824
rect 7276 13815 7334 13821
rect 7558 13812 7564 13824
rect 7616 13812 7622 13864
rect 8662 13812 8668 13864
rect 8720 13852 8726 13864
rect 9125 13855 9183 13861
rect 9125 13852 9137 13855
rect 8720 13824 9137 13852
rect 8720 13812 8726 13824
rect 9125 13821 9137 13824
rect 9171 13821 9183 13855
rect 10244 13852 10272 13892
rect 10410 13880 10416 13892
rect 10468 13880 10474 13932
rect 10594 13880 10600 13932
rect 10652 13920 10658 13932
rect 11425 13923 11483 13929
rect 11425 13920 11437 13923
rect 10652 13892 11437 13920
rect 10652 13880 10658 13892
rect 11425 13889 11437 13892
rect 11471 13920 11483 13923
rect 11514 13920 11520 13932
rect 11471 13892 11520 13920
rect 11471 13889 11483 13892
rect 11425 13883 11483 13889
rect 11514 13880 11520 13892
rect 11572 13880 11578 13932
rect 11900 13920 11928 13960
rect 12437 13957 12449 13960
rect 12483 13957 12495 13991
rect 12437 13951 12495 13957
rect 11808 13892 11928 13920
rect 10612 13852 10640 13880
rect 10244 13824 10640 13852
rect 9125 13815 9183 13821
rect 11238 13812 11244 13864
rect 11296 13852 11302 13864
rect 11808 13861 11836 13892
rect 12158 13880 12164 13932
rect 12216 13920 12222 13932
rect 12820 13920 12848 14028
rect 15010 14016 15016 14028
rect 15068 14016 15074 14068
rect 15565 14059 15623 14065
rect 15565 14025 15577 14059
rect 15611 14056 15623 14059
rect 16574 14056 16580 14068
rect 15611 14028 16580 14056
rect 15611 14025 15623 14028
rect 15565 14019 15623 14025
rect 16574 14016 16580 14028
rect 16632 14016 16638 14068
rect 19334 14056 19340 14068
rect 16684 14028 19340 14056
rect 13446 13988 13452 14000
rect 12912 13960 13452 13988
rect 12912 13929 12940 13960
rect 13446 13948 13452 13960
rect 13504 13948 13510 14000
rect 13538 13948 13544 14000
rect 13596 13988 13602 14000
rect 16206 13988 16212 14000
rect 13596 13960 16212 13988
rect 13596 13948 13602 13960
rect 16206 13948 16212 13960
rect 16264 13948 16270 14000
rect 16390 13988 16396 14000
rect 16351 13960 16396 13988
rect 16390 13948 16396 13960
rect 16448 13948 16454 14000
rect 16684 13988 16712 14028
rect 19334 14016 19340 14028
rect 19392 14016 19398 14068
rect 21913 14059 21971 14065
rect 21913 14025 21925 14059
rect 21959 14056 21971 14059
rect 22278 14056 22284 14068
rect 21959 14028 22284 14056
rect 21959 14025 21971 14028
rect 21913 14019 21971 14025
rect 22278 14016 22284 14028
rect 22336 14016 22342 14068
rect 16500 13960 16712 13988
rect 17497 13991 17555 13997
rect 12216 13892 12848 13920
rect 12897 13923 12955 13929
rect 12216 13880 12222 13892
rect 12897 13889 12909 13923
rect 12943 13889 12955 13923
rect 12897 13883 12955 13889
rect 13081 13923 13139 13929
rect 13081 13889 13093 13923
rect 13127 13920 13139 13923
rect 14090 13920 14096 13932
rect 13127 13892 14096 13920
rect 13127 13889 13139 13892
rect 13081 13883 13139 13889
rect 14090 13880 14096 13892
rect 14148 13920 14154 13932
rect 14550 13920 14556 13932
rect 14148 13892 14556 13920
rect 14148 13880 14154 13892
rect 14550 13880 14556 13892
rect 14608 13880 14614 13932
rect 15102 13880 15108 13932
rect 15160 13920 15166 13932
rect 16025 13923 16083 13929
rect 16025 13920 16037 13923
rect 15160 13892 16037 13920
rect 15160 13880 15166 13892
rect 16025 13889 16037 13892
rect 16071 13889 16083 13923
rect 16025 13883 16083 13889
rect 16114 13880 16120 13932
rect 16172 13920 16178 13932
rect 16500 13920 16528 13960
rect 17497 13957 17509 13991
rect 17543 13988 17555 13991
rect 17954 13988 17960 14000
rect 17543 13960 17960 13988
rect 17543 13957 17555 13960
rect 17497 13951 17555 13957
rect 17954 13948 17960 13960
rect 18012 13948 18018 14000
rect 19242 13948 19248 14000
rect 19300 13988 19306 14000
rect 19429 13991 19487 13997
rect 19429 13988 19441 13991
rect 19300 13960 19441 13988
rect 19300 13948 19306 13960
rect 19429 13957 19441 13960
rect 19475 13957 19487 13991
rect 19429 13951 19487 13957
rect 21637 13991 21695 13997
rect 21637 13957 21649 13991
rect 21683 13988 21695 13991
rect 21729 13991 21787 13997
rect 21729 13988 21741 13991
rect 21683 13960 21741 13988
rect 21683 13957 21695 13960
rect 21637 13951 21695 13957
rect 21729 13957 21741 13960
rect 21775 13957 21787 13991
rect 21729 13951 21787 13957
rect 16945 13923 17003 13929
rect 16945 13920 16957 13923
rect 16172 13892 16217 13920
rect 16307 13892 16528 13920
rect 16583 13892 16957 13920
rect 16172 13880 16178 13892
rect 11793 13855 11851 13861
rect 11793 13852 11805 13855
rect 11296 13824 11805 13852
rect 11296 13812 11302 13824
rect 11793 13821 11805 13824
rect 11839 13821 11851 13855
rect 11793 13815 11851 13821
rect 11882 13812 11888 13864
rect 11940 13852 11946 13864
rect 12710 13852 12716 13864
rect 11940 13824 12716 13852
rect 11940 13812 11946 13824
rect 12710 13812 12716 13824
rect 12768 13812 12774 13864
rect 14182 13812 14188 13864
rect 14240 13852 14246 13864
rect 16307 13852 16335 13892
rect 14240 13824 16335 13852
rect 14240 13812 14246 13824
rect 16482 13812 16488 13864
rect 16540 13852 16546 13864
rect 16583 13852 16611 13892
rect 16945 13889 16957 13892
rect 16991 13920 17003 13923
rect 17126 13920 17132 13932
rect 16991 13892 17132 13920
rect 16991 13889 17003 13892
rect 16945 13883 17003 13889
rect 17126 13880 17132 13892
rect 17184 13880 17190 13932
rect 17681 13923 17739 13929
rect 17681 13920 17693 13923
rect 17236 13892 17693 13920
rect 16540 13824 16611 13852
rect 16540 13812 16546 13824
rect 16666 13812 16672 13864
rect 16724 13852 16730 13864
rect 17236 13852 17264 13892
rect 17681 13889 17693 13892
rect 17727 13889 17739 13923
rect 18046 13920 18052 13932
rect 18007 13892 18052 13920
rect 17681 13883 17739 13889
rect 18046 13880 18052 13892
rect 18104 13880 18110 13932
rect 19797 13923 19855 13929
rect 19797 13889 19809 13923
rect 19843 13920 19855 13923
rect 20162 13920 20168 13932
rect 19843 13892 20168 13920
rect 19843 13889 19855 13892
rect 19797 13883 19855 13889
rect 20162 13880 20168 13892
rect 20220 13880 20226 13932
rect 20303 13923 20361 13929
rect 20303 13889 20315 13923
rect 20349 13920 20361 13923
rect 20714 13920 20720 13932
rect 20349 13892 20720 13920
rect 20349 13889 20361 13892
rect 20303 13883 20361 13889
rect 20714 13880 20720 13892
rect 20772 13880 20778 13932
rect 22462 13920 22468 13932
rect 22423 13892 22468 13920
rect 22462 13880 22468 13892
rect 22520 13880 22526 13932
rect 16724 13824 17264 13852
rect 17313 13855 17371 13861
rect 16724 13812 16730 13824
rect 17313 13821 17325 13855
rect 17359 13852 17371 13855
rect 17770 13852 17776 13864
rect 17359 13824 17776 13852
rect 17359 13821 17371 13824
rect 17313 13815 17371 13821
rect 17770 13812 17776 13824
rect 17828 13812 17834 13864
rect 18322 13861 18328 13864
rect 18316 13852 18328 13861
rect 18283 13824 18328 13852
rect 18316 13815 18328 13824
rect 18322 13812 18328 13815
rect 18380 13812 18386 13864
rect 20438 13812 20444 13864
rect 20496 13852 20502 13864
rect 20533 13855 20591 13861
rect 20533 13852 20545 13855
rect 20496 13824 20545 13852
rect 20496 13812 20502 13824
rect 20533 13821 20545 13824
rect 20579 13821 20591 13855
rect 20533 13815 20591 13821
rect 21266 13812 21272 13864
rect 21324 13852 21330 13864
rect 21729 13855 21787 13861
rect 21729 13852 21741 13855
rect 21324 13824 21741 13852
rect 21324 13812 21330 13824
rect 21729 13821 21741 13824
rect 21775 13821 21787 13855
rect 21729 13815 21787 13821
rect 2498 13784 2504 13796
rect 1728 13756 2504 13784
rect 1728 13744 1734 13756
rect 2498 13744 2504 13756
rect 2556 13744 2562 13796
rect 4154 13744 4160 13796
rect 4212 13784 4218 13796
rect 10042 13784 10048 13796
rect 4212 13756 10048 13784
rect 4212 13744 4218 13756
rect 10042 13744 10048 13756
rect 10100 13744 10106 13796
rect 10137 13787 10195 13793
rect 10137 13753 10149 13787
rect 10183 13784 10195 13787
rect 11146 13784 11152 13796
rect 10183 13756 10824 13784
rect 11107 13756 11152 13784
rect 10183 13753 10195 13756
rect 10137 13747 10195 13753
rect 5718 13716 5724 13728
rect 5679 13688 5724 13716
rect 5718 13676 5724 13688
rect 5776 13676 5782 13728
rect 5810 13676 5816 13728
rect 5868 13716 5874 13728
rect 5868 13688 5913 13716
rect 5868 13676 5874 13688
rect 7190 13676 7196 13728
rect 7248 13716 7254 13728
rect 7558 13716 7564 13728
rect 7248 13688 7564 13716
rect 7248 13676 7254 13688
rect 7558 13676 7564 13688
rect 7616 13676 7622 13728
rect 8389 13719 8447 13725
rect 8389 13685 8401 13719
rect 8435 13716 8447 13719
rect 8662 13716 8668 13728
rect 8435 13688 8668 13716
rect 8435 13685 8447 13688
rect 8389 13679 8447 13685
rect 8662 13676 8668 13688
rect 8720 13676 8726 13728
rect 9030 13716 9036 13728
rect 8991 13688 9036 13716
rect 9030 13676 9036 13688
rect 9088 13676 9094 13728
rect 10226 13716 10232 13728
rect 10187 13688 10232 13716
rect 10226 13676 10232 13688
rect 10284 13676 10290 13728
rect 10796 13725 10824 13756
rect 11146 13744 11152 13756
rect 11204 13744 11210 13796
rect 12805 13787 12863 13793
rect 12805 13784 12817 13787
rect 12636 13756 12817 13784
rect 10781 13719 10839 13725
rect 10781 13685 10793 13719
rect 10827 13685 10839 13719
rect 11238 13716 11244 13728
rect 11199 13688 11244 13716
rect 10781 13679 10839 13685
rect 11238 13676 11244 13688
rect 11296 13676 11302 13728
rect 11514 13676 11520 13728
rect 11572 13716 11578 13728
rect 12636 13716 12664 13756
rect 12805 13753 12817 13756
rect 12851 13753 12863 13787
rect 13722 13784 13728 13796
rect 13683 13756 13728 13784
rect 12805 13747 12863 13753
rect 13722 13744 13728 13756
rect 13780 13744 13786 13796
rect 13814 13744 13820 13796
rect 13872 13784 13878 13796
rect 16761 13787 16819 13793
rect 16761 13784 16773 13787
rect 13872 13756 16773 13784
rect 13872 13744 13878 13756
rect 16761 13753 16773 13756
rect 16807 13753 16819 13787
rect 16761 13747 16819 13753
rect 17126 13744 17132 13796
rect 17184 13784 17190 13796
rect 19610 13784 19616 13796
rect 17184 13756 19616 13784
rect 17184 13744 17190 13756
rect 19610 13744 19616 13756
rect 19668 13744 19674 13796
rect 22281 13787 22339 13793
rect 22281 13784 22293 13787
rect 21284 13756 22293 13784
rect 21284 13728 21312 13756
rect 22281 13753 22293 13756
rect 22327 13753 22339 13787
rect 22281 13747 22339 13753
rect 11572 13688 12664 13716
rect 11572 13676 11578 13688
rect 12710 13676 12716 13728
rect 12768 13716 12774 13728
rect 13078 13716 13084 13728
rect 12768 13688 13084 13716
rect 12768 13676 12774 13688
rect 13078 13676 13084 13688
rect 13136 13676 13142 13728
rect 14274 13676 14280 13728
rect 14332 13716 14338 13728
rect 15197 13719 15255 13725
rect 15197 13716 15209 13719
rect 14332 13688 15209 13716
rect 14332 13676 14338 13688
rect 15197 13685 15209 13688
rect 15243 13716 15255 13719
rect 15654 13716 15660 13728
rect 15243 13688 15660 13716
rect 15243 13685 15255 13688
rect 15197 13679 15255 13685
rect 15654 13676 15660 13688
rect 15712 13676 15718 13728
rect 15933 13719 15991 13725
rect 15933 13685 15945 13719
rect 15979 13716 15991 13719
rect 16114 13716 16120 13728
rect 15979 13688 16120 13716
rect 15979 13685 15991 13688
rect 15933 13679 15991 13685
rect 16114 13676 16120 13688
rect 16172 13676 16178 13728
rect 16206 13676 16212 13728
rect 16264 13716 16270 13728
rect 16853 13719 16911 13725
rect 16853 13716 16865 13719
rect 16264 13688 16865 13716
rect 16264 13676 16270 13688
rect 16853 13685 16865 13688
rect 16899 13685 16911 13719
rect 16853 13679 16911 13685
rect 19334 13676 19340 13728
rect 19392 13716 19398 13728
rect 20070 13716 20076 13728
rect 19392 13688 20076 13716
rect 19392 13676 19398 13688
rect 20070 13676 20076 13688
rect 20128 13676 20134 13728
rect 20263 13719 20321 13725
rect 20263 13685 20275 13719
rect 20309 13716 20321 13719
rect 20622 13716 20628 13728
rect 20309 13688 20628 13716
rect 20309 13685 20321 13688
rect 20263 13679 20321 13685
rect 20622 13676 20628 13688
rect 20680 13676 20686 13728
rect 21266 13676 21272 13728
rect 21324 13676 21330 13728
rect 22370 13716 22376 13728
rect 22331 13688 22376 13716
rect 22370 13676 22376 13688
rect 22428 13676 22434 13728
rect 1104 13626 23276 13648
rect 1104 13574 8379 13626
rect 8431 13574 8443 13626
rect 8495 13574 8507 13626
rect 8559 13574 8571 13626
rect 8623 13574 15776 13626
rect 15828 13574 15840 13626
rect 15892 13574 15904 13626
rect 15956 13574 15968 13626
rect 16020 13574 23276 13626
rect 1104 13552 23276 13574
rect 3050 13512 3056 13524
rect 2963 13484 3056 13512
rect 3050 13472 3056 13484
rect 3108 13512 3114 13524
rect 4062 13512 4068 13524
rect 3108 13484 4068 13512
rect 3108 13472 3114 13484
rect 4062 13472 4068 13484
rect 4120 13472 4126 13524
rect 5905 13515 5963 13521
rect 5905 13481 5917 13515
rect 5951 13512 5963 13515
rect 5994 13512 6000 13524
rect 5951 13484 6000 13512
rect 5951 13481 5963 13484
rect 5905 13475 5963 13481
rect 5994 13472 6000 13484
rect 6052 13472 6058 13524
rect 6365 13515 6423 13521
rect 6365 13481 6377 13515
rect 6411 13512 6423 13515
rect 7742 13512 7748 13524
rect 6411 13484 7748 13512
rect 6411 13481 6423 13484
rect 6365 13475 6423 13481
rect 7742 13472 7748 13484
rect 7800 13472 7806 13524
rect 8757 13515 8815 13521
rect 8757 13481 8769 13515
rect 8803 13512 8815 13515
rect 9490 13512 9496 13524
rect 8803 13484 9496 13512
rect 8803 13481 8815 13484
rect 8757 13475 8815 13481
rect 9490 13472 9496 13484
rect 9548 13472 9554 13524
rect 9769 13515 9827 13521
rect 9769 13481 9781 13515
rect 9815 13512 9827 13515
rect 10226 13512 10232 13524
rect 9815 13484 10232 13512
rect 9815 13481 9827 13484
rect 9769 13475 9827 13481
rect 10226 13472 10232 13484
rect 10284 13472 10290 13524
rect 10502 13512 10508 13524
rect 10336 13484 10508 13512
rect 1940 13447 1998 13453
rect 1940 13413 1952 13447
rect 1986 13444 1998 13447
rect 2130 13444 2136 13456
rect 1986 13416 2136 13444
rect 1986 13413 1998 13416
rect 1940 13407 1998 13413
rect 2130 13404 2136 13416
rect 2188 13404 2194 13456
rect 4792 13447 4850 13453
rect 4792 13413 4804 13447
rect 4838 13444 4850 13447
rect 5442 13444 5448 13456
rect 4838 13416 5448 13444
rect 4838 13413 4850 13416
rect 4792 13407 4850 13413
rect 5442 13404 5448 13416
rect 5500 13404 5506 13456
rect 7368 13447 7426 13453
rect 7368 13413 7380 13447
rect 7414 13444 7426 13447
rect 8662 13444 8668 13456
rect 7414 13416 8668 13444
rect 7414 13413 7426 13416
rect 7368 13407 7426 13413
rect 8662 13404 8668 13416
rect 8720 13404 8726 13456
rect 9950 13444 9956 13456
rect 8772 13416 9956 13444
rect 1670 13376 1676 13388
rect 1631 13348 1676 13376
rect 1670 13336 1676 13348
rect 1728 13336 1734 13388
rect 3418 13376 3424 13388
rect 3379 13348 3424 13376
rect 3418 13336 3424 13348
rect 3476 13336 3482 13388
rect 4065 13379 4123 13385
rect 4065 13345 4077 13379
rect 4111 13376 4123 13379
rect 4154 13376 4160 13388
rect 4111 13348 4160 13376
rect 4111 13345 4123 13348
rect 4065 13339 4123 13345
rect 4154 13336 4160 13348
rect 4212 13336 4218 13388
rect 4246 13336 4252 13388
rect 4304 13376 4310 13388
rect 4525 13379 4583 13385
rect 4525 13376 4537 13379
rect 4304 13348 4537 13376
rect 4304 13336 4310 13348
rect 4525 13345 4537 13348
rect 4571 13345 4583 13379
rect 4525 13339 4583 13345
rect 5074 13336 5080 13388
rect 5132 13376 5138 13388
rect 6181 13379 6239 13385
rect 6181 13376 6193 13379
rect 5132 13348 6193 13376
rect 5132 13336 5138 13348
rect 6181 13345 6193 13348
rect 6227 13345 6239 13379
rect 6181 13339 6239 13345
rect 7006 13336 7012 13388
rect 7064 13376 7070 13388
rect 7101 13379 7159 13385
rect 7101 13376 7113 13379
rect 7064 13348 7113 13376
rect 7064 13336 7070 13348
rect 7101 13345 7113 13348
rect 7147 13376 7159 13379
rect 7926 13376 7932 13388
rect 7147 13348 7932 13376
rect 7147 13345 7159 13348
rect 7101 13339 7159 13345
rect 7926 13336 7932 13348
rect 7984 13336 7990 13388
rect 8772 13308 8800 13416
rect 9950 13404 9956 13416
rect 10008 13404 10014 13456
rect 10336 13444 10364 13484
rect 10502 13472 10508 13484
rect 10560 13472 10566 13524
rect 11146 13472 11152 13524
rect 11204 13512 11210 13524
rect 11977 13515 12035 13521
rect 11977 13512 11989 13515
rect 11204 13484 11989 13512
rect 11204 13472 11210 13484
rect 11977 13481 11989 13484
rect 12023 13481 12035 13515
rect 11977 13475 12035 13481
rect 10594 13444 10600 13456
rect 10244 13416 10364 13444
rect 10428 13416 10600 13444
rect 8941 13379 8999 13385
rect 8941 13345 8953 13379
rect 8987 13345 8999 13379
rect 8941 13339 8999 13345
rect 9033 13379 9091 13385
rect 9033 13345 9045 13379
rect 9079 13376 9091 13379
rect 9214 13376 9220 13388
rect 9079 13348 9220 13376
rect 9079 13345 9091 13348
rect 9033 13339 9091 13345
rect 8128 13280 8800 13308
rect 8956 13308 8984 13339
rect 9214 13336 9220 13348
rect 9272 13336 9278 13388
rect 10134 13376 10140 13388
rect 10095 13348 10140 13376
rect 10134 13336 10140 13348
rect 10192 13336 10198 13388
rect 10244 13385 10272 13416
rect 10229 13379 10287 13385
rect 10229 13345 10241 13379
rect 10275 13345 10287 13379
rect 10229 13339 10287 13345
rect 9674 13308 9680 13320
rect 8956 13280 9680 13308
rect 3605 13175 3663 13181
rect 3605 13141 3617 13175
rect 3651 13172 3663 13175
rect 5258 13172 5264 13184
rect 3651 13144 5264 13172
rect 3651 13141 3663 13144
rect 3605 13135 3663 13141
rect 5258 13132 5264 13144
rect 5316 13132 5322 13184
rect 5442 13132 5448 13184
rect 5500 13172 5506 13184
rect 8128 13172 8156 13280
rect 9674 13268 9680 13280
rect 9732 13268 9738 13320
rect 10428 13317 10456 13416
rect 10594 13404 10600 13416
rect 10652 13404 10658 13456
rect 10962 13404 10968 13456
rect 11020 13444 11026 13456
rect 11992 13444 12020 13475
rect 12526 13472 12532 13524
rect 12584 13512 12590 13524
rect 13449 13515 13507 13521
rect 13449 13512 13461 13515
rect 12584 13484 13461 13512
rect 12584 13472 12590 13484
rect 13449 13481 13461 13484
rect 13495 13481 13507 13515
rect 13449 13475 13507 13481
rect 14090 13472 14096 13524
rect 14148 13512 14154 13524
rect 14642 13512 14648 13524
rect 14148 13484 14648 13512
rect 14148 13472 14154 13484
rect 14642 13472 14648 13484
rect 14700 13472 14706 13524
rect 14826 13472 14832 13524
rect 14884 13512 14890 13524
rect 16669 13515 16727 13521
rect 14884 13484 16620 13512
rect 14884 13472 14890 13484
rect 16592 13456 16620 13484
rect 16669 13481 16681 13515
rect 16715 13512 16727 13515
rect 16758 13512 16764 13524
rect 16715 13484 16764 13512
rect 16715 13481 16727 13484
rect 16669 13475 16727 13481
rect 16758 13472 16764 13484
rect 16816 13512 16822 13524
rect 18506 13512 18512 13524
rect 16816 13484 18512 13512
rect 16816 13472 16822 13484
rect 18506 13472 18512 13484
rect 18564 13472 18570 13524
rect 18785 13515 18843 13521
rect 18785 13481 18797 13515
rect 18831 13512 18843 13515
rect 19794 13512 19800 13524
rect 18831 13484 19800 13512
rect 18831 13481 18843 13484
rect 18785 13475 18843 13481
rect 19794 13472 19800 13484
rect 19852 13472 19858 13524
rect 12314 13447 12372 13453
rect 12314 13444 12326 13447
rect 11020 13416 11928 13444
rect 11992 13416 12326 13444
rect 11020 13404 11026 13416
rect 10864 13379 10922 13385
rect 10864 13345 10876 13379
rect 10910 13376 10922 13379
rect 11238 13376 11244 13388
rect 10910 13348 11244 13376
rect 10910 13345 10922 13348
rect 10864 13339 10922 13345
rect 11238 13336 11244 13348
rect 11296 13336 11302 13388
rect 11900 13376 11928 13416
rect 12314 13413 12326 13416
rect 12360 13413 12372 13447
rect 16482 13444 16488 13456
rect 12314 13407 12372 13413
rect 13740 13416 16488 13444
rect 13740 13376 13768 13416
rect 16482 13404 16488 13416
rect 16540 13404 16546 13456
rect 16574 13404 16580 13456
rect 16632 13404 16638 13456
rect 22370 13444 22376 13456
rect 17963 13416 22376 13444
rect 11900 13348 13768 13376
rect 13808 13379 13866 13385
rect 13808 13345 13820 13379
rect 13854 13376 13866 13379
rect 13854 13348 14596 13376
rect 13854 13345 13866 13348
rect 13808 13339 13866 13345
rect 10413 13311 10471 13317
rect 10413 13277 10425 13311
rect 10459 13277 10471 13311
rect 10413 13271 10471 13277
rect 10597 13311 10655 13317
rect 10597 13277 10609 13311
rect 10643 13277 10655 13311
rect 12066 13308 12072 13320
rect 12027 13280 12072 13308
rect 10597 13271 10655 13277
rect 9030 13240 9036 13252
rect 8496 13212 9036 13240
rect 8496 13184 8524 13212
rect 9030 13200 9036 13212
rect 9088 13200 9094 13252
rect 10226 13200 10232 13252
rect 10284 13240 10290 13252
rect 10612 13240 10640 13271
rect 12066 13268 12072 13280
rect 12124 13268 12130 13320
rect 13538 13308 13544 13320
rect 13499 13280 13544 13308
rect 13538 13268 13544 13280
rect 13596 13268 13602 13320
rect 14568 13252 14596 13348
rect 15378 13336 15384 13388
rect 15436 13376 15442 13388
rect 17218 13385 17224 13388
rect 15545 13379 15603 13385
rect 15545 13376 15557 13379
rect 15436 13348 15557 13376
rect 15436 13336 15442 13348
rect 15545 13345 15557 13348
rect 15591 13345 15603 13379
rect 17212 13376 17224 13385
rect 17179 13348 17224 13376
rect 15545 13339 15603 13345
rect 17212 13339 17224 13348
rect 17218 13336 17224 13339
rect 17276 13336 17282 13388
rect 15286 13308 15292 13320
rect 15247 13280 15292 13308
rect 15286 13268 15292 13280
rect 15344 13268 15350 13320
rect 16298 13268 16304 13320
rect 16356 13308 16362 13320
rect 16945 13311 17003 13317
rect 16945 13308 16957 13311
rect 16356 13280 16957 13308
rect 16356 13268 16362 13280
rect 16945 13277 16957 13280
rect 16991 13277 17003 13311
rect 16945 13271 17003 13277
rect 10284 13212 10640 13240
rect 10284 13200 10290 13212
rect 14550 13200 14556 13252
rect 14608 13240 14614 13252
rect 14608 13212 14872 13240
rect 14608 13200 14614 13212
rect 8478 13172 8484 13184
rect 5500 13144 8156 13172
rect 8439 13144 8484 13172
rect 5500 13132 5506 13144
rect 8478 13132 8484 13144
rect 8536 13132 8542 13184
rect 9214 13172 9220 13184
rect 9175 13144 9220 13172
rect 9214 13132 9220 13144
rect 9272 13132 9278 13184
rect 9950 13132 9956 13184
rect 10008 13172 10014 13184
rect 12434 13172 12440 13184
rect 10008 13144 12440 13172
rect 10008 13132 10014 13144
rect 12434 13132 12440 13144
rect 12492 13132 12498 13184
rect 14844 13172 14872 13212
rect 14918 13200 14924 13252
rect 14976 13240 14982 13252
rect 14976 13212 15021 13240
rect 14976 13200 14982 13212
rect 17963 13172 17991 13416
rect 22370 13404 22376 13416
rect 22428 13404 22434 13456
rect 18601 13379 18659 13385
rect 18601 13345 18613 13379
rect 18647 13376 18659 13379
rect 18966 13376 18972 13388
rect 18647 13348 18972 13376
rect 18647 13345 18659 13348
rect 18601 13339 18659 13345
rect 18966 13336 18972 13348
rect 19024 13336 19030 13388
rect 19409 13379 19467 13385
rect 19409 13376 19421 13379
rect 19076 13348 19421 13376
rect 18046 13268 18052 13320
rect 18104 13268 18110 13320
rect 18782 13268 18788 13320
rect 18840 13308 18846 13320
rect 19076 13308 19104 13348
rect 19409 13345 19421 13348
rect 19455 13376 19467 13379
rect 20898 13376 20904 13388
rect 19455 13348 20760 13376
rect 20859 13348 20904 13376
rect 19455 13345 19467 13348
rect 19409 13339 19467 13345
rect 18840 13280 19104 13308
rect 19153 13311 19211 13317
rect 18840 13268 18846 13280
rect 19153 13277 19165 13311
rect 19199 13277 19211 13311
rect 19153 13271 19211 13277
rect 18064 13240 18092 13268
rect 19168 13240 19196 13271
rect 18064 13212 19196 13240
rect 14844 13144 17991 13172
rect 18046 13132 18052 13184
rect 18104 13172 18110 13184
rect 18325 13175 18383 13181
rect 18325 13172 18337 13175
rect 18104 13144 18337 13172
rect 18104 13132 18110 13144
rect 18325 13141 18337 13144
rect 18371 13141 18383 13175
rect 18325 13135 18383 13141
rect 18506 13132 18512 13184
rect 18564 13172 18570 13184
rect 19334 13172 19340 13184
rect 18564 13144 19340 13172
rect 18564 13132 18570 13144
rect 19334 13132 19340 13144
rect 19392 13132 19398 13184
rect 19794 13132 19800 13184
rect 19852 13172 19858 13184
rect 20530 13172 20536 13184
rect 19852 13144 20536 13172
rect 19852 13132 19858 13144
rect 20530 13132 20536 13144
rect 20588 13132 20594 13184
rect 20732 13172 20760 13348
rect 20898 13336 20904 13348
rect 20956 13376 20962 13388
rect 21177 13379 21235 13385
rect 21177 13376 21189 13379
rect 20956 13348 21189 13376
rect 20956 13336 20962 13348
rect 21177 13345 21189 13348
rect 21223 13345 21235 13379
rect 21358 13376 21364 13388
rect 21319 13348 21364 13376
rect 21177 13339 21235 13345
rect 21358 13336 21364 13348
rect 21416 13336 21422 13388
rect 21634 13385 21640 13388
rect 21628 13376 21640 13385
rect 21595 13348 21640 13376
rect 21628 13339 21640 13348
rect 21634 13336 21640 13339
rect 21692 13336 21698 13388
rect 22741 13175 22799 13181
rect 22741 13172 22753 13175
rect 20732 13144 22753 13172
rect 22741 13141 22753 13144
rect 22787 13141 22799 13175
rect 22741 13135 22799 13141
rect 1104 13082 23276 13104
rect 1104 13030 4680 13082
rect 4732 13030 4744 13082
rect 4796 13030 4808 13082
rect 4860 13030 4872 13082
rect 4924 13030 12078 13082
rect 12130 13030 12142 13082
rect 12194 13030 12206 13082
rect 12258 13030 12270 13082
rect 12322 13030 19475 13082
rect 19527 13030 19539 13082
rect 19591 13030 19603 13082
rect 19655 13030 19667 13082
rect 19719 13030 23276 13082
rect 1104 13008 23276 13030
rect 1670 12968 1676 12980
rect 1412 12940 1676 12968
rect 1412 12841 1440 12940
rect 1670 12928 1676 12940
rect 1728 12928 1734 12980
rect 2038 12928 2044 12980
rect 2096 12968 2102 12980
rect 2777 12971 2835 12977
rect 2777 12968 2789 12971
rect 2096 12940 2789 12968
rect 2096 12928 2102 12940
rect 2777 12937 2789 12940
rect 2823 12937 2835 12971
rect 2777 12931 2835 12937
rect 3237 12971 3295 12977
rect 3237 12937 3249 12971
rect 3283 12968 3295 12971
rect 3786 12968 3792 12980
rect 3283 12940 3792 12968
rect 3283 12937 3295 12940
rect 3237 12931 3295 12937
rect 3786 12928 3792 12940
rect 3844 12928 3850 12980
rect 7650 12928 7656 12980
rect 7708 12968 7714 12980
rect 8665 12971 8723 12977
rect 7708 12940 7972 12968
rect 7708 12928 7714 12940
rect 6457 12903 6515 12909
rect 6457 12869 6469 12903
rect 6503 12869 6515 12903
rect 7944 12900 7972 12940
rect 8665 12937 8677 12971
rect 8711 12968 8723 12971
rect 8754 12968 8760 12980
rect 8711 12940 8760 12968
rect 8711 12937 8723 12940
rect 8665 12931 8723 12937
rect 8754 12928 8760 12940
rect 8812 12928 8818 12980
rect 9674 12968 9680 12980
rect 9635 12940 9680 12968
rect 9674 12928 9680 12940
rect 9732 12928 9738 12980
rect 11054 12968 11060 12980
rect 10336 12940 11060 12968
rect 10336 12900 10364 12940
rect 11054 12928 11060 12940
rect 11112 12928 11118 12980
rect 11238 12928 11244 12980
rect 11296 12968 11302 12980
rect 11701 12971 11759 12977
rect 11701 12968 11713 12971
rect 11296 12940 11713 12968
rect 11296 12928 11302 12940
rect 11701 12937 11713 12940
rect 11747 12937 11759 12971
rect 11701 12931 11759 12937
rect 12161 12971 12219 12977
rect 12161 12937 12173 12971
rect 12207 12968 12219 12971
rect 12710 12968 12716 12980
rect 12207 12940 12716 12968
rect 12207 12937 12219 12940
rect 12161 12931 12219 12937
rect 12710 12928 12716 12940
rect 12768 12928 12774 12980
rect 19794 12968 19800 12980
rect 13004 12940 19800 12968
rect 7944 12872 9720 12900
rect 6457 12863 6515 12869
rect 1397 12835 1455 12841
rect 1397 12801 1409 12835
rect 1443 12801 1455 12835
rect 1397 12795 1455 12801
rect 3878 12792 3884 12844
rect 3936 12832 3942 12844
rect 4157 12835 4215 12841
rect 4157 12832 4169 12835
rect 3936 12804 4169 12832
rect 3936 12792 3942 12804
rect 4157 12801 4169 12804
rect 4203 12801 4215 12835
rect 4157 12795 4215 12801
rect 4246 12792 4252 12844
rect 4304 12832 4310 12844
rect 4709 12835 4767 12841
rect 4709 12832 4721 12835
rect 4304 12804 4721 12832
rect 4304 12792 4310 12804
rect 4709 12801 4721 12804
rect 4755 12801 4767 12835
rect 6472 12832 6500 12863
rect 7006 12832 7012 12844
rect 6472 12804 7012 12832
rect 4709 12795 4767 12801
rect 7006 12792 7012 12804
rect 7064 12792 7070 12844
rect 9306 12832 9312 12844
rect 9267 12804 9312 12832
rect 9306 12792 9312 12804
rect 9364 12792 9370 12844
rect 9692 12832 9720 12872
rect 10015 12872 10364 12900
rect 10015 12832 10043 12872
rect 11330 12860 11336 12912
rect 11388 12900 11394 12912
rect 13004 12900 13032 12940
rect 19794 12928 19800 12940
rect 19852 12928 19858 12980
rect 19889 12971 19947 12977
rect 19889 12937 19901 12971
rect 19935 12968 19947 12971
rect 20162 12968 20168 12980
rect 19935 12940 20168 12968
rect 19935 12937 19947 12940
rect 19889 12931 19947 12937
rect 20162 12928 20168 12940
rect 20220 12928 20226 12980
rect 20990 12968 20996 12980
rect 20278 12940 20996 12968
rect 11388 12872 13032 12900
rect 14369 12903 14427 12909
rect 11388 12860 11394 12872
rect 14369 12869 14381 12903
rect 14415 12900 14427 12903
rect 14550 12900 14556 12912
rect 14415 12872 14556 12900
rect 14415 12869 14427 12872
rect 14369 12863 14427 12869
rect 14550 12860 14556 12872
rect 14608 12860 14614 12912
rect 17310 12860 17316 12912
rect 17368 12900 17374 12912
rect 18049 12903 18107 12909
rect 18049 12900 18061 12903
rect 17368 12872 18061 12900
rect 17368 12860 17374 12872
rect 18049 12869 18061 12872
rect 18095 12869 18107 12903
rect 18049 12863 18107 12869
rect 18322 12860 18328 12912
rect 18380 12900 18386 12912
rect 18877 12903 18935 12909
rect 18877 12900 18889 12903
rect 18380 12872 18889 12900
rect 18380 12860 18386 12872
rect 18877 12869 18889 12872
rect 18923 12869 18935 12903
rect 18877 12863 18935 12869
rect 9692 12804 10043 12832
rect 10134 12792 10140 12844
rect 10192 12832 10198 12844
rect 12618 12832 12624 12844
rect 10192 12804 10456 12832
rect 10192 12792 10198 12804
rect 3053 12767 3111 12773
rect 3053 12733 3065 12767
rect 3099 12764 3111 12767
rect 3326 12764 3332 12776
rect 3099 12736 3332 12764
rect 3099 12733 3111 12736
rect 3053 12727 3111 12733
rect 3326 12724 3332 12736
rect 3384 12724 3390 12776
rect 4976 12767 5034 12773
rect 3896 12736 4384 12764
rect 1664 12699 1722 12705
rect 1664 12665 1676 12699
rect 1710 12696 1722 12699
rect 3896 12696 3924 12736
rect 1710 12668 3924 12696
rect 3973 12699 4031 12705
rect 1710 12665 1722 12668
rect 1664 12659 1722 12665
rect 3973 12665 3985 12699
rect 4019 12696 4031 12699
rect 4246 12696 4252 12708
rect 4019 12668 4252 12696
rect 4019 12665 4031 12668
rect 3973 12659 4031 12665
rect 4246 12656 4252 12668
rect 4304 12656 4310 12708
rect 3602 12628 3608 12640
rect 3563 12600 3608 12628
rect 3602 12588 3608 12600
rect 3660 12588 3666 12640
rect 4062 12628 4068 12640
rect 4023 12600 4068 12628
rect 4062 12588 4068 12600
rect 4120 12588 4126 12640
rect 4356 12628 4384 12736
rect 4976 12733 4988 12767
rect 5022 12764 5034 12767
rect 5810 12764 5816 12776
rect 5022 12736 5816 12764
rect 5022 12733 5034 12736
rect 4976 12727 5034 12733
rect 5810 12724 5816 12736
rect 5868 12724 5874 12776
rect 5902 12724 5908 12776
rect 5960 12764 5966 12776
rect 6641 12767 6699 12773
rect 6641 12764 6653 12767
rect 5960 12736 6653 12764
rect 5960 12724 5966 12736
rect 6641 12733 6653 12736
rect 6687 12733 6699 12767
rect 6641 12727 6699 12733
rect 7276 12767 7334 12773
rect 7276 12733 7288 12767
rect 7322 12764 7334 12767
rect 8478 12764 8484 12776
rect 7322 12736 8484 12764
rect 7322 12733 7334 12736
rect 7276 12727 7334 12733
rect 8478 12724 8484 12736
rect 8536 12724 8542 12776
rect 10033 12773 10039 12776
rect 9861 12767 9919 12773
rect 9861 12733 9873 12767
rect 9907 12733 9919 12767
rect 9861 12727 9919 12733
rect 9978 12767 10039 12773
rect 9978 12733 9990 12767
rect 10024 12733 10039 12767
rect 9978 12727 10039 12733
rect 4430 12656 4436 12708
rect 4488 12696 4494 12708
rect 5442 12696 5448 12708
rect 4488 12668 5448 12696
rect 4488 12656 4494 12668
rect 5442 12656 5448 12668
rect 5500 12656 5506 12708
rect 9125 12699 9183 12705
rect 9125 12696 9137 12699
rect 8404 12668 9137 12696
rect 5718 12628 5724 12640
rect 4356 12600 5724 12628
rect 5718 12588 5724 12600
rect 5776 12628 5782 12640
rect 6089 12631 6147 12637
rect 6089 12628 6101 12631
rect 5776 12600 6101 12628
rect 5776 12588 5782 12600
rect 6089 12597 6101 12600
rect 6135 12597 6147 12631
rect 6089 12591 6147 12597
rect 8202 12588 8208 12640
rect 8260 12628 8266 12640
rect 8404 12637 8432 12668
rect 9125 12665 9137 12668
rect 9171 12665 9183 12699
rect 9876 12696 9904 12727
rect 10033 12724 10039 12727
rect 10091 12724 10097 12776
rect 10226 12724 10232 12776
rect 10284 12764 10290 12776
rect 10321 12767 10379 12773
rect 10321 12764 10333 12767
rect 10284 12736 10333 12764
rect 10284 12724 10290 12736
rect 10321 12733 10333 12736
rect 10367 12733 10379 12767
rect 10428 12764 10456 12804
rect 12452 12804 12624 12832
rect 10588 12767 10646 12773
rect 10588 12764 10600 12767
rect 10428 12736 10600 12764
rect 10321 12727 10379 12733
rect 10588 12733 10600 12736
rect 10634 12764 10646 12767
rect 11146 12764 11152 12776
rect 10634 12736 11152 12764
rect 10634 12733 10646 12736
rect 10588 12727 10646 12733
rect 11146 12724 11152 12736
rect 11204 12724 11210 12776
rect 11790 12724 11796 12776
rect 11848 12764 11854 12776
rect 12452 12773 12480 12804
rect 12618 12792 12624 12804
rect 12676 12792 12682 12844
rect 17494 12832 17500 12844
rect 17319 12804 17500 12832
rect 11977 12767 12035 12773
rect 11977 12764 11989 12767
rect 11848 12736 11989 12764
rect 11848 12724 11854 12736
rect 11977 12733 11989 12736
rect 12023 12733 12035 12767
rect 11977 12727 12035 12733
rect 12437 12767 12495 12773
rect 12437 12733 12449 12767
rect 12483 12733 12495 12767
rect 12986 12764 12992 12776
rect 12947 12736 12992 12764
rect 12437 12727 12495 12733
rect 12986 12724 12992 12736
rect 13044 12764 13050 12776
rect 13538 12764 13544 12776
rect 13044 12736 13544 12764
rect 13044 12724 13050 12736
rect 13538 12724 13544 12736
rect 13596 12764 13602 12776
rect 14550 12764 14556 12776
rect 13596 12736 14556 12764
rect 13596 12724 13602 12736
rect 14550 12724 14556 12736
rect 14608 12764 14614 12776
rect 14918 12773 14924 12776
rect 14645 12767 14703 12773
rect 14645 12764 14657 12767
rect 14608 12736 14657 12764
rect 14608 12724 14614 12736
rect 14645 12733 14657 12736
rect 14691 12733 14703 12767
rect 14912 12764 14924 12773
rect 14879 12736 14924 12764
rect 14645 12727 14703 12733
rect 14912 12727 14924 12736
rect 14918 12724 14924 12727
rect 14976 12724 14982 12776
rect 15286 12724 15292 12776
rect 15344 12764 15350 12776
rect 16298 12764 16304 12776
rect 15344 12736 16304 12764
rect 15344 12724 15350 12736
rect 16298 12724 16304 12736
rect 16356 12724 16362 12776
rect 16574 12773 16580 12776
rect 16568 12764 16580 12773
rect 16535 12736 16580 12764
rect 16568 12727 16580 12736
rect 16574 12724 16580 12727
rect 16632 12724 16638 12776
rect 16850 12724 16856 12776
rect 16908 12764 16914 12776
rect 17319 12764 17347 12804
rect 17494 12792 17500 12804
rect 17552 12792 17558 12844
rect 17862 12792 17868 12844
rect 17920 12832 17926 12844
rect 18601 12835 18659 12841
rect 18601 12832 18613 12835
rect 17920 12804 18613 12832
rect 17920 12792 17926 12804
rect 18601 12801 18613 12804
rect 18647 12801 18659 12835
rect 18601 12795 18659 12801
rect 18966 12792 18972 12844
rect 19024 12832 19030 12844
rect 19429 12835 19487 12841
rect 19024 12804 19380 12832
rect 19024 12792 19030 12804
rect 17773 12767 17831 12773
rect 17773 12764 17785 12767
rect 16908 12736 17347 12764
rect 17420 12736 17785 12764
rect 16908 12724 16914 12736
rect 12342 12696 12348 12708
rect 9876 12668 12348 12696
rect 9125 12659 9183 12665
rect 12342 12656 12348 12668
rect 12400 12656 12406 12708
rect 12618 12696 12624 12708
rect 12579 12668 12624 12696
rect 12618 12656 12624 12668
rect 12676 12656 12682 12708
rect 13256 12699 13314 12705
rect 13256 12665 13268 12699
rect 13302 12696 13314 12699
rect 15654 12696 15660 12708
rect 13302 12668 15660 12696
rect 13302 12665 13314 12668
rect 13256 12659 13314 12665
rect 15654 12656 15660 12668
rect 15712 12696 15718 12708
rect 17420 12696 17448 12736
rect 17773 12733 17785 12736
rect 17819 12733 17831 12767
rect 18417 12767 18475 12773
rect 18417 12764 18429 12767
rect 17773 12727 17831 12733
rect 17972 12736 18429 12764
rect 15712 12668 17448 12696
rect 15712 12656 15718 12668
rect 17494 12656 17500 12708
rect 17552 12696 17558 12708
rect 17972 12696 18000 12736
rect 18417 12733 18429 12736
rect 18463 12733 18475 12767
rect 18417 12727 18475 12733
rect 18874 12724 18880 12776
rect 18932 12764 18938 12776
rect 19245 12767 19303 12773
rect 19245 12764 19257 12767
rect 18932 12736 19257 12764
rect 18932 12724 18938 12736
rect 19245 12733 19257 12736
rect 19291 12733 19303 12767
rect 19352 12764 19380 12804
rect 19429 12801 19441 12835
rect 19475 12832 19487 12835
rect 19794 12832 19800 12844
rect 19475 12804 19800 12832
rect 19475 12801 19487 12804
rect 19429 12795 19487 12801
rect 19794 12792 19800 12804
rect 19852 12832 19858 12844
rect 20278 12841 20306 12940
rect 20990 12928 20996 12940
rect 21048 12968 21054 12980
rect 21358 12968 21364 12980
rect 21048 12940 21364 12968
rect 21048 12928 21054 12940
rect 21358 12928 21364 12940
rect 21416 12928 21422 12980
rect 21726 12968 21732 12980
rect 21687 12940 21732 12968
rect 21726 12928 21732 12940
rect 21784 12928 21790 12980
rect 20257 12835 20315 12841
rect 19852 12804 20208 12832
rect 19852 12792 19858 12804
rect 20180 12776 20208 12804
rect 20257 12801 20269 12835
rect 20303 12801 20315 12835
rect 22370 12832 22376 12844
rect 22331 12804 22376 12832
rect 20257 12795 20315 12801
rect 22370 12792 22376 12804
rect 22428 12792 22434 12844
rect 20073 12767 20131 12773
rect 20073 12764 20085 12767
rect 19352 12736 20085 12764
rect 19245 12727 19303 12733
rect 20073 12733 20085 12736
rect 20119 12733 20131 12767
rect 20073 12727 20131 12733
rect 20162 12724 20168 12776
rect 20220 12724 20226 12776
rect 20530 12773 20536 12776
rect 20513 12767 20536 12773
rect 20513 12733 20525 12767
rect 20513 12727 20536 12733
rect 20530 12724 20536 12727
rect 20588 12724 20594 12776
rect 18506 12696 18512 12708
rect 17552 12668 18000 12696
rect 18467 12668 18512 12696
rect 17552 12656 17558 12668
rect 18506 12656 18512 12668
rect 18564 12656 18570 12708
rect 19058 12656 19064 12708
rect 19116 12696 19122 12708
rect 19337 12699 19395 12705
rect 19337 12696 19349 12699
rect 19116 12668 19349 12696
rect 19116 12656 19122 12668
rect 19337 12665 19349 12668
rect 19383 12665 19395 12699
rect 22097 12699 22155 12705
rect 22097 12696 22109 12699
rect 19337 12659 19395 12665
rect 20364 12668 22109 12696
rect 8389 12631 8447 12637
rect 8389 12628 8401 12631
rect 8260 12600 8401 12628
rect 8260 12588 8266 12600
rect 8389 12597 8401 12600
rect 8435 12597 8447 12631
rect 9030 12628 9036 12640
rect 8991 12600 9036 12628
rect 8389 12591 8447 12597
rect 9030 12588 9036 12600
rect 9088 12588 9094 12640
rect 10137 12631 10195 12637
rect 10137 12597 10149 12631
rect 10183 12628 10195 12631
rect 10686 12628 10692 12640
rect 10183 12600 10692 12628
rect 10183 12597 10195 12600
rect 10137 12591 10195 12597
rect 10686 12588 10692 12600
rect 10744 12588 10750 12640
rect 12526 12588 12532 12640
rect 12584 12628 12590 12640
rect 12805 12631 12863 12637
rect 12805 12628 12817 12631
rect 12584 12600 12817 12628
rect 12584 12588 12590 12600
rect 12805 12597 12817 12600
rect 12851 12597 12863 12631
rect 12805 12591 12863 12597
rect 15378 12588 15384 12640
rect 15436 12628 15442 12640
rect 16025 12631 16083 12637
rect 16025 12628 16037 12631
rect 15436 12600 16037 12628
rect 15436 12588 15442 12600
rect 16025 12597 16037 12600
rect 16071 12628 16083 12631
rect 16850 12628 16856 12640
rect 16071 12600 16856 12628
rect 16071 12597 16083 12600
rect 16025 12591 16083 12597
rect 16850 12588 16856 12600
rect 16908 12588 16914 12640
rect 17678 12628 17684 12640
rect 17639 12600 17684 12628
rect 17678 12588 17684 12600
rect 17736 12588 17742 12640
rect 17773 12631 17831 12637
rect 17773 12597 17785 12631
rect 17819 12628 17831 12631
rect 20364 12628 20392 12668
rect 22097 12665 22109 12668
rect 22143 12665 22155 12699
rect 22097 12659 22155 12665
rect 17819 12600 20392 12628
rect 17819 12597 17831 12600
rect 17773 12591 17831 12597
rect 21266 12588 21272 12640
rect 21324 12628 21330 12640
rect 21637 12631 21695 12637
rect 21637 12628 21649 12631
rect 21324 12600 21649 12628
rect 21324 12588 21330 12600
rect 21637 12597 21649 12600
rect 21683 12597 21695 12631
rect 21637 12591 21695 12597
rect 22189 12631 22247 12637
rect 22189 12597 22201 12631
rect 22235 12628 22247 12631
rect 22278 12628 22284 12640
rect 22235 12600 22284 12628
rect 22235 12597 22247 12600
rect 22189 12591 22247 12597
rect 22278 12588 22284 12600
rect 22336 12588 22342 12640
rect 1104 12538 23276 12560
rect 1104 12486 8379 12538
rect 8431 12486 8443 12538
rect 8495 12486 8507 12538
rect 8559 12486 8571 12538
rect 8623 12486 15776 12538
rect 15828 12486 15840 12538
rect 15892 12486 15904 12538
rect 15956 12486 15968 12538
rect 16020 12486 23276 12538
rect 1104 12464 23276 12486
rect 2041 12427 2099 12433
rect 2041 12393 2053 12427
rect 2087 12424 2099 12427
rect 2130 12424 2136 12436
rect 2087 12396 2136 12424
rect 2087 12393 2099 12396
rect 2041 12387 2099 12393
rect 2130 12384 2136 12396
rect 2188 12384 2194 12436
rect 4249 12427 4307 12433
rect 4249 12393 4261 12427
rect 4295 12424 4307 12427
rect 4522 12424 4528 12436
rect 4295 12396 4528 12424
rect 4295 12393 4307 12396
rect 4249 12387 4307 12393
rect 4522 12384 4528 12396
rect 4580 12384 4586 12436
rect 5810 12384 5816 12436
rect 5868 12424 5874 12436
rect 5997 12427 6055 12433
rect 5997 12424 6009 12427
rect 5868 12396 6009 12424
rect 5868 12384 5874 12396
rect 5997 12393 6009 12396
rect 6043 12393 6055 12427
rect 8202 12424 8208 12436
rect 5997 12387 6055 12393
rect 7291 12396 8208 12424
rect 3142 12356 3148 12368
rect 3103 12328 3148 12356
rect 3142 12316 3148 12328
rect 3200 12316 3206 12368
rect 3234 12316 3240 12368
rect 3292 12356 3298 12368
rect 7291 12365 7319 12396
rect 8202 12384 8208 12396
rect 8260 12384 8266 12436
rect 8849 12427 8907 12433
rect 8849 12393 8861 12427
rect 8895 12393 8907 12427
rect 8849 12387 8907 12393
rect 9217 12427 9275 12433
rect 9217 12393 9229 12427
rect 9263 12424 9275 12427
rect 9674 12424 9680 12436
rect 9263 12396 9680 12424
rect 9263 12393 9275 12396
rect 9217 12387 9275 12393
rect 7276 12359 7334 12365
rect 3292 12328 4108 12356
rect 3292 12316 3298 12328
rect 2038 12248 2044 12300
rect 2096 12288 2102 12300
rect 2133 12291 2191 12297
rect 2133 12288 2145 12291
rect 2096 12260 2145 12288
rect 2096 12248 2102 12260
rect 2133 12257 2145 12260
rect 2179 12257 2191 12291
rect 2133 12251 2191 12257
rect 3053 12291 3111 12297
rect 3053 12257 3065 12291
rect 3099 12288 3111 12291
rect 3326 12288 3332 12300
rect 3099 12260 3332 12288
rect 3099 12257 3111 12260
rect 3053 12251 3111 12257
rect 3326 12248 3332 12260
rect 3384 12248 3390 12300
rect 4080 12297 4108 12328
rect 7276 12325 7288 12359
rect 7322 12325 7334 12359
rect 8864 12356 8892 12387
rect 9674 12384 9680 12396
rect 9732 12384 9738 12436
rect 9861 12427 9919 12433
rect 9861 12393 9873 12427
rect 9907 12424 9919 12427
rect 11514 12424 11520 12436
rect 9907 12396 11520 12424
rect 9907 12393 9919 12396
rect 9861 12387 9919 12393
rect 11514 12384 11520 12396
rect 11572 12384 11578 12436
rect 12342 12384 12348 12436
rect 12400 12424 12406 12436
rect 12713 12427 12771 12433
rect 12713 12424 12725 12427
rect 12400 12396 12725 12424
rect 12400 12384 12406 12396
rect 12713 12393 12725 12396
rect 12759 12393 12771 12427
rect 13446 12424 13452 12436
rect 12713 12387 12771 12393
rect 12912 12396 13452 12424
rect 12912 12356 12940 12396
rect 13446 12384 13452 12396
rect 13504 12384 13510 12436
rect 14921 12427 14979 12433
rect 14921 12393 14933 12427
rect 14967 12424 14979 12427
rect 15470 12424 15476 12436
rect 14967 12396 15476 12424
rect 14967 12393 14979 12396
rect 14921 12387 14979 12393
rect 15470 12384 15476 12396
rect 15528 12384 15534 12436
rect 15657 12427 15715 12433
rect 15657 12393 15669 12427
rect 15703 12424 15715 12427
rect 16206 12424 16212 12436
rect 15703 12396 16212 12424
rect 15703 12393 15715 12396
rect 15657 12387 15715 12393
rect 16206 12384 16212 12396
rect 16264 12384 16270 12436
rect 16298 12384 16304 12436
rect 16356 12424 16362 12436
rect 17126 12424 17132 12436
rect 16356 12396 17132 12424
rect 16356 12384 16362 12396
rect 17126 12384 17132 12396
rect 17184 12384 17190 12436
rect 17218 12384 17224 12436
rect 17276 12424 17282 12436
rect 17405 12427 17463 12433
rect 17405 12424 17417 12427
rect 17276 12396 17417 12424
rect 17276 12384 17282 12396
rect 17405 12393 17417 12396
rect 17451 12393 17463 12427
rect 17405 12387 17463 12393
rect 17492 12396 18175 12424
rect 13630 12356 13636 12368
rect 8864 12328 12940 12356
rect 12995 12328 13636 12356
rect 7276 12319 7334 12325
rect 4065 12291 4123 12297
rect 4065 12257 4077 12291
rect 4111 12257 4123 12291
rect 4065 12251 4123 12257
rect 4884 12291 4942 12297
rect 4884 12257 4896 12291
rect 4930 12288 4942 12291
rect 5810 12288 5816 12300
rect 4930 12260 5816 12288
rect 4930 12257 4942 12260
rect 4884 12251 4942 12257
rect 5810 12248 5816 12260
rect 5868 12248 5874 12300
rect 6457 12291 6515 12297
rect 6457 12257 6469 12291
rect 6503 12257 6515 12291
rect 7006 12288 7012 12300
rect 6967 12260 7012 12288
rect 6457 12251 6515 12257
rect 2317 12223 2375 12229
rect 2317 12189 2329 12223
rect 2363 12220 2375 12223
rect 3237 12223 3295 12229
rect 3237 12220 3249 12223
rect 2363 12192 3249 12220
rect 2363 12189 2375 12192
rect 2317 12183 2375 12189
rect 3237 12189 3249 12192
rect 3283 12220 3295 12223
rect 3878 12220 3884 12232
rect 3283 12192 3884 12220
rect 3283 12189 3295 12192
rect 3237 12183 3295 12189
rect 3878 12180 3884 12192
rect 3936 12180 3942 12232
rect 4154 12180 4160 12232
rect 4212 12220 4218 12232
rect 4617 12223 4675 12229
rect 4617 12220 4629 12223
rect 4212 12192 4629 12220
rect 4212 12180 4218 12192
rect 4617 12189 4629 12192
rect 4663 12189 4675 12223
rect 6472 12220 6500 12251
rect 7006 12248 7012 12260
rect 7064 12248 7070 12300
rect 8665 12291 8723 12297
rect 7116 12260 8616 12288
rect 7116 12220 7144 12260
rect 6472 12192 7144 12220
rect 8588 12220 8616 12260
rect 8665 12257 8677 12291
rect 8711 12288 8723 12291
rect 8846 12288 8852 12300
rect 8711 12260 8852 12288
rect 8711 12257 8723 12260
rect 8665 12251 8723 12257
rect 8846 12248 8852 12260
rect 8904 12248 8910 12300
rect 9122 12248 9128 12300
rect 9180 12288 9186 12300
rect 9401 12291 9459 12297
rect 9401 12288 9413 12291
rect 9180 12260 9413 12288
rect 9180 12248 9186 12260
rect 9401 12257 9413 12260
rect 9447 12257 9459 12291
rect 9401 12251 9459 12257
rect 9493 12291 9551 12297
rect 9493 12257 9505 12291
rect 9539 12288 9551 12291
rect 9677 12291 9735 12297
rect 9677 12288 9689 12291
rect 9539 12260 9689 12288
rect 9539 12257 9551 12260
rect 9493 12251 9551 12257
rect 9677 12257 9689 12260
rect 9723 12257 9735 12291
rect 9677 12251 9735 12257
rect 10413 12291 10471 12297
rect 10413 12257 10425 12291
rect 10459 12288 10471 12291
rect 10686 12288 10692 12300
rect 10459 12260 10692 12288
rect 10459 12257 10471 12260
rect 10413 12251 10471 12257
rect 10686 12248 10692 12260
rect 10744 12248 10750 12300
rect 11149 12291 11207 12297
rect 11149 12257 11161 12291
rect 11195 12288 11207 12291
rect 11333 12291 11391 12297
rect 11333 12288 11345 12291
rect 11195 12260 11345 12288
rect 11195 12257 11207 12260
rect 11149 12251 11207 12257
rect 11333 12257 11345 12260
rect 11379 12257 11391 12291
rect 11333 12251 11391 12257
rect 11425 12291 11483 12297
rect 11425 12257 11437 12291
rect 11471 12288 11483 12291
rect 11514 12288 11520 12300
rect 11471 12260 11520 12288
rect 11471 12257 11483 12260
rect 11425 12251 11483 12257
rect 11514 12248 11520 12260
rect 11572 12248 11578 12300
rect 12995 12220 13023 12328
rect 13630 12316 13636 12328
rect 13688 12316 13694 12368
rect 16316 12356 16344 12384
rect 16040 12328 16344 12356
rect 13532 12291 13590 12297
rect 13532 12257 13544 12291
rect 13578 12288 13590 12291
rect 13814 12288 13820 12300
rect 13578 12260 13820 12288
rect 13578 12257 13590 12260
rect 13532 12251 13590 12257
rect 13814 12248 13820 12260
rect 13872 12248 13878 12300
rect 14737 12291 14795 12297
rect 14737 12257 14749 12291
rect 14783 12257 14795 12291
rect 14737 12251 14795 12257
rect 15473 12291 15531 12297
rect 15473 12257 15485 12291
rect 15519 12288 15531 12291
rect 15562 12288 15568 12300
rect 15519 12260 15568 12288
rect 15519 12257 15531 12260
rect 15473 12251 15531 12257
rect 8588 12192 13023 12220
rect 13265 12223 13323 12229
rect 4617 12183 4675 12189
rect 13265 12189 13277 12223
rect 13311 12189 13323 12223
rect 13265 12183 13323 12189
rect 1673 12155 1731 12161
rect 1673 12121 1685 12155
rect 1719 12152 1731 12155
rect 6914 12152 6920 12164
rect 1719 12124 3004 12152
rect 1719 12121 1731 12124
rect 1673 12115 1731 12121
rect 1946 12044 1952 12096
rect 2004 12084 2010 12096
rect 2685 12087 2743 12093
rect 2685 12084 2697 12087
rect 2004 12056 2697 12084
rect 2004 12044 2010 12056
rect 2685 12053 2697 12056
rect 2731 12053 2743 12087
rect 2976 12084 3004 12124
rect 6564 12124 6920 12152
rect 3694 12084 3700 12096
rect 2976 12056 3700 12084
rect 2685 12047 2743 12053
rect 3694 12044 3700 12056
rect 3752 12044 3758 12096
rect 3878 12044 3884 12096
rect 3936 12084 3942 12096
rect 6564 12084 6592 12124
rect 6914 12112 6920 12124
rect 6972 12112 6978 12164
rect 8202 12112 8208 12164
rect 8260 12152 8266 12164
rect 9493 12155 9551 12161
rect 9493 12152 9505 12155
rect 8260 12124 9505 12152
rect 8260 12112 8266 12124
rect 9493 12121 9505 12124
rect 9539 12121 9551 12155
rect 9493 12115 9551 12121
rect 10965 12155 11023 12161
rect 10965 12121 10977 12155
rect 11011 12152 11023 12155
rect 12986 12152 12992 12164
rect 11011 12124 12992 12152
rect 11011 12121 11023 12124
rect 10965 12115 11023 12121
rect 12986 12112 12992 12124
rect 13044 12152 13050 12164
rect 13280 12152 13308 12183
rect 13044 12124 13308 12152
rect 13044 12112 13050 12124
rect 3936 12056 6592 12084
rect 6641 12087 6699 12093
rect 3936 12044 3942 12056
rect 6641 12053 6653 12087
rect 6687 12084 6699 12087
rect 8294 12084 8300 12096
rect 6687 12056 8300 12084
rect 6687 12053 6699 12056
rect 6641 12047 6699 12053
rect 8294 12044 8300 12056
rect 8352 12044 8358 12096
rect 8386 12044 8392 12096
rect 8444 12084 8450 12096
rect 9030 12084 9036 12096
rect 8444 12056 9036 12084
rect 8444 12044 8450 12056
rect 9030 12044 9036 12056
rect 9088 12044 9094 12096
rect 10042 12044 10048 12096
rect 10100 12084 10106 12096
rect 10229 12087 10287 12093
rect 10229 12084 10241 12087
rect 10100 12056 10241 12084
rect 10100 12044 10106 12056
rect 10229 12053 10241 12056
rect 10275 12053 10287 12087
rect 10229 12047 10287 12053
rect 11333 12087 11391 12093
rect 11333 12053 11345 12087
rect 11379 12084 11391 12087
rect 13262 12084 13268 12096
rect 11379 12056 13268 12084
rect 11379 12053 11391 12056
rect 11333 12047 11391 12053
rect 13262 12044 13268 12056
rect 13320 12044 13326 12096
rect 14642 12084 14648 12096
rect 14603 12056 14648 12084
rect 14642 12044 14648 12056
rect 14700 12044 14706 12096
rect 14752 12084 14780 12251
rect 15562 12248 15568 12260
rect 15620 12248 15626 12300
rect 16040 12297 16068 12328
rect 16758 12316 16764 12368
rect 16816 12356 16822 12368
rect 17492 12356 17520 12396
rect 18046 12365 18052 12368
rect 18040 12356 18052 12365
rect 16816 12328 17520 12356
rect 18007 12328 18052 12356
rect 16816 12316 16822 12328
rect 18040 12319 18052 12328
rect 18046 12316 18052 12319
rect 18104 12316 18110 12368
rect 18147 12356 18175 12396
rect 19058 12384 19064 12436
rect 19116 12424 19122 12436
rect 19153 12427 19211 12433
rect 19153 12424 19165 12427
rect 19116 12396 19165 12424
rect 19116 12384 19122 12396
rect 19153 12393 19165 12396
rect 19199 12424 19211 12427
rect 20806 12424 20812 12436
rect 19199 12396 20812 12424
rect 19199 12393 19211 12396
rect 19153 12387 19211 12393
rect 20806 12384 20812 12396
rect 20864 12384 20870 12436
rect 20898 12384 20904 12436
rect 20956 12424 20962 12436
rect 21174 12424 21180 12436
rect 20956 12396 21180 12424
rect 20956 12384 20962 12396
rect 21174 12384 21180 12396
rect 21232 12384 21238 12436
rect 21266 12365 21272 12368
rect 19889 12359 19947 12365
rect 19889 12356 19901 12359
rect 18147 12328 19901 12356
rect 19889 12325 19901 12328
rect 19935 12325 19947 12359
rect 21260 12356 21272 12365
rect 21227 12328 21272 12356
rect 19889 12319 19947 12325
rect 21260 12319 21272 12328
rect 21266 12316 21272 12319
rect 21324 12316 21330 12368
rect 16025 12291 16083 12297
rect 16025 12257 16037 12291
rect 16071 12257 16083 12291
rect 16025 12251 16083 12257
rect 16292 12291 16350 12297
rect 16292 12257 16304 12291
rect 16338 12288 16350 12291
rect 17586 12288 17592 12300
rect 16338 12260 17592 12288
rect 16338 12257 16350 12260
rect 16292 12251 16350 12257
rect 17586 12248 17592 12260
rect 17644 12248 17650 12300
rect 17773 12291 17831 12297
rect 17773 12288 17785 12291
rect 17696 12260 17785 12288
rect 17126 12180 17132 12232
rect 17184 12220 17190 12232
rect 17696 12220 17724 12260
rect 17773 12257 17785 12260
rect 17819 12257 17831 12291
rect 19610 12288 19616 12300
rect 17773 12251 17831 12257
rect 17880 12260 19616 12288
rect 17880 12220 17908 12260
rect 19610 12248 19616 12260
rect 19668 12248 19674 12300
rect 19794 12288 19800 12300
rect 19755 12260 19800 12288
rect 19794 12248 19800 12260
rect 19852 12248 19858 12300
rect 20162 12288 20168 12300
rect 19996 12260 20168 12288
rect 17184 12192 17724 12220
rect 17788 12192 17908 12220
rect 17184 12180 17190 12192
rect 17402 12152 17408 12164
rect 16960 12124 17408 12152
rect 16960 12084 16988 12124
rect 17402 12112 17408 12124
rect 17460 12112 17466 12164
rect 17678 12112 17684 12164
rect 17736 12152 17742 12164
rect 17788 12152 17816 12192
rect 18874 12180 18880 12232
rect 18932 12220 18938 12232
rect 19996 12229 20024 12260
rect 20162 12248 20168 12260
rect 20220 12248 20226 12300
rect 20990 12288 20996 12300
rect 20951 12260 20996 12288
rect 20990 12248 20996 12260
rect 21048 12248 21054 12300
rect 19981 12223 20039 12229
rect 19981 12220 19993 12223
rect 18932 12192 19993 12220
rect 18932 12180 18938 12192
rect 19981 12189 19993 12192
rect 20027 12189 20039 12223
rect 19981 12183 20039 12189
rect 17736 12124 17816 12152
rect 17736 12112 17742 12124
rect 14752 12056 16988 12084
rect 17954 12044 17960 12096
rect 18012 12084 18018 12096
rect 18138 12084 18144 12096
rect 18012 12056 18144 12084
rect 18012 12044 18018 12056
rect 18138 12044 18144 12056
rect 18196 12044 18202 12096
rect 19429 12087 19487 12093
rect 19429 12053 19441 12087
rect 19475 12084 19487 12087
rect 20254 12084 20260 12096
rect 19475 12056 20260 12084
rect 19475 12053 19487 12056
rect 19429 12047 19487 12053
rect 20254 12044 20260 12056
rect 20312 12044 20318 12096
rect 20990 12044 20996 12096
rect 21048 12084 21054 12096
rect 22373 12087 22431 12093
rect 22373 12084 22385 12087
rect 21048 12056 22385 12084
rect 21048 12044 21054 12056
rect 22373 12053 22385 12056
rect 22419 12053 22431 12087
rect 22373 12047 22431 12053
rect 1104 11994 23276 12016
rect 1104 11942 4680 11994
rect 4732 11942 4744 11994
rect 4796 11942 4808 11994
rect 4860 11942 4872 11994
rect 4924 11942 12078 11994
rect 12130 11942 12142 11994
rect 12194 11942 12206 11994
rect 12258 11942 12270 11994
rect 12322 11942 19475 11994
rect 19527 11942 19539 11994
rect 19591 11942 19603 11994
rect 19655 11942 19667 11994
rect 19719 11942 23276 11994
rect 1104 11920 23276 11942
rect 1489 11883 1547 11889
rect 1489 11849 1501 11883
rect 1535 11880 1547 11883
rect 3418 11880 3424 11892
rect 1535 11852 3424 11880
rect 1535 11849 1547 11852
rect 1489 11843 1547 11849
rect 3418 11840 3424 11852
rect 3476 11840 3482 11892
rect 3881 11883 3939 11889
rect 3881 11849 3893 11883
rect 3927 11880 3939 11883
rect 3973 11883 4031 11889
rect 3973 11880 3985 11883
rect 3927 11852 3985 11880
rect 3927 11849 3939 11852
rect 3881 11843 3939 11849
rect 3973 11849 3985 11852
rect 4019 11849 4031 11883
rect 5810 11880 5816 11892
rect 3973 11843 4031 11849
rect 4080 11852 5396 11880
rect 5771 11852 5816 11880
rect 3510 11772 3516 11824
rect 3568 11812 3574 11824
rect 4080 11812 4108 11852
rect 3568 11784 4108 11812
rect 4157 11815 4215 11821
rect 3568 11772 3574 11784
rect 4157 11781 4169 11815
rect 4203 11781 4215 11815
rect 5368 11812 5396 11852
rect 5810 11840 5816 11852
rect 5868 11840 5874 11892
rect 6365 11883 6423 11889
rect 6365 11849 6377 11883
rect 6411 11880 6423 11883
rect 7466 11880 7472 11892
rect 6411 11852 7472 11880
rect 6411 11849 6423 11852
rect 6365 11843 6423 11849
rect 7466 11840 7472 11852
rect 7524 11840 7530 11892
rect 7742 11840 7748 11892
rect 7800 11880 7806 11892
rect 8202 11880 8208 11892
rect 7800 11852 8208 11880
rect 7800 11840 7806 11852
rect 8202 11840 8208 11852
rect 8260 11840 8266 11892
rect 8294 11840 8300 11892
rect 8352 11880 8358 11892
rect 10962 11880 10968 11892
rect 8352 11852 10968 11880
rect 8352 11840 8358 11852
rect 10962 11840 10968 11852
rect 11020 11840 11026 11892
rect 11146 11840 11152 11892
rect 11204 11880 11210 11892
rect 11609 11883 11667 11889
rect 11609 11880 11621 11883
rect 11204 11852 11621 11880
rect 11204 11840 11210 11852
rect 11609 11849 11621 11852
rect 11655 11849 11667 11883
rect 11609 11843 11667 11849
rect 13814 11840 13820 11892
rect 13872 11880 13878 11892
rect 14185 11883 14243 11889
rect 14185 11880 14197 11883
rect 13872 11852 14197 11880
rect 13872 11840 13878 11852
rect 14185 11849 14197 11852
rect 14231 11880 14243 11883
rect 14231 11852 15608 11880
rect 14231 11849 14243 11852
rect 14185 11843 14243 11849
rect 5368 11784 6040 11812
rect 4157 11775 4215 11781
rect 1946 11744 1952 11756
rect 1907 11716 1952 11744
rect 1946 11704 1952 11716
rect 2004 11704 2010 11756
rect 2130 11744 2136 11756
rect 2091 11716 2136 11744
rect 2130 11704 2136 11716
rect 2188 11704 2194 11756
rect 3973 11747 4031 11753
rect 3973 11713 3985 11747
rect 4019 11744 4031 11747
rect 4062 11744 4068 11756
rect 4019 11716 4068 11744
rect 4019 11713 4031 11716
rect 3973 11707 4031 11713
rect 4062 11704 4068 11716
rect 4120 11704 4126 11756
rect 4172 11688 4200 11775
rect 4356 11716 4568 11744
rect 2501 11679 2559 11685
rect 2501 11645 2513 11679
rect 2547 11676 2559 11679
rect 4154 11676 4160 11688
rect 2547 11648 4160 11676
rect 2547 11645 2559 11648
rect 2501 11639 2559 11645
rect 1946 11568 1952 11620
rect 2004 11608 2010 11620
rect 2516 11608 2544 11639
rect 4154 11636 4160 11648
rect 4212 11676 4218 11688
rect 4356 11685 4384 11716
rect 4341 11679 4399 11685
rect 4212 11648 4292 11676
rect 4212 11636 4218 11648
rect 2004 11580 2544 11608
rect 2768 11611 2826 11617
rect 2004 11568 2010 11580
rect 2768 11577 2780 11611
rect 2814 11608 2826 11611
rect 3326 11608 3332 11620
rect 2814 11580 3332 11608
rect 2814 11577 2826 11580
rect 2768 11571 2826 11577
rect 3326 11568 3332 11580
rect 3384 11568 3390 11620
rect 4264 11608 4292 11648
rect 4341 11645 4353 11679
rect 4387 11645 4399 11679
rect 4341 11639 4399 11645
rect 4433 11679 4491 11685
rect 4433 11645 4445 11679
rect 4479 11645 4491 11679
rect 4540 11676 4568 11716
rect 5902 11676 5908 11688
rect 4540 11648 5908 11676
rect 4433 11639 4491 11645
rect 4448 11608 4476 11639
rect 5902 11636 5908 11648
rect 5960 11636 5966 11688
rect 4264 11580 4476 11608
rect 4700 11611 4758 11617
rect 4700 11577 4712 11611
rect 4746 11608 4758 11611
rect 5442 11608 5448 11620
rect 4746 11580 5448 11608
rect 4746 11577 4758 11580
rect 4700 11571 4758 11577
rect 5442 11568 5448 11580
rect 5500 11568 5506 11620
rect 6012 11608 6040 11784
rect 8110 11772 8116 11824
rect 8168 11812 8174 11824
rect 8481 11815 8539 11821
rect 8481 11812 8493 11815
rect 8168 11784 8493 11812
rect 8168 11772 8174 11784
rect 8481 11781 8493 11784
rect 8527 11781 8539 11815
rect 9950 11812 9956 11824
rect 8481 11775 8539 11781
rect 9054 11784 9956 11812
rect 9054 11744 9082 11784
rect 9950 11772 9956 11784
rect 10008 11772 10014 11824
rect 15580 11812 15608 11852
rect 15654 11840 15660 11892
rect 15712 11880 15718 11892
rect 15841 11883 15899 11889
rect 15841 11880 15853 11883
rect 15712 11852 15853 11880
rect 15712 11840 15718 11852
rect 15841 11849 15853 11852
rect 15887 11849 15899 11883
rect 19794 11880 19800 11892
rect 15841 11843 15899 11849
rect 15948 11852 19800 11880
rect 15948 11812 15976 11852
rect 19794 11840 19800 11852
rect 19852 11840 19858 11892
rect 20622 11840 20628 11892
rect 20680 11880 20686 11892
rect 22465 11883 22523 11889
rect 22465 11880 22477 11883
rect 20680 11852 22477 11880
rect 20680 11840 20686 11852
rect 22465 11849 22477 11852
rect 22511 11849 22523 11883
rect 22465 11843 22523 11849
rect 15580 11784 15976 11812
rect 16945 11815 17003 11821
rect 16945 11781 16957 11815
rect 16991 11812 17003 11815
rect 17678 11812 17684 11824
rect 16991 11784 17684 11812
rect 16991 11781 17003 11784
rect 16945 11775 17003 11781
rect 17678 11772 17684 11784
rect 17736 11772 17742 11824
rect 7852 11716 9082 11744
rect 9125 11747 9183 11753
rect 6181 11679 6239 11685
rect 6181 11645 6193 11679
rect 6227 11676 6239 11679
rect 6546 11676 6552 11688
rect 6227 11648 6552 11676
rect 6227 11645 6239 11648
rect 6181 11639 6239 11645
rect 6546 11636 6552 11648
rect 6604 11636 6610 11688
rect 6825 11679 6883 11685
rect 6825 11645 6837 11679
rect 6871 11676 6883 11679
rect 6914 11676 6920 11688
rect 6871 11648 6920 11676
rect 6871 11645 6883 11648
rect 6825 11639 6883 11645
rect 6914 11636 6920 11648
rect 6972 11636 6978 11688
rect 7852 11676 7880 11716
rect 9125 11713 9137 11747
rect 9171 11744 9183 11747
rect 9306 11744 9312 11756
rect 9171 11716 9312 11744
rect 9171 11713 9183 11716
rect 9125 11707 9183 11713
rect 9306 11704 9312 11716
rect 9364 11704 9370 11756
rect 10042 11704 10048 11756
rect 10100 11744 10106 11756
rect 10229 11747 10287 11753
rect 10229 11744 10241 11747
rect 10100 11716 10241 11744
rect 10100 11704 10106 11716
rect 10229 11713 10241 11716
rect 10275 11713 10287 11747
rect 10229 11707 10287 11713
rect 12618 11704 12624 11756
rect 12676 11744 12682 11756
rect 12805 11747 12863 11753
rect 12805 11744 12817 11747
rect 12676 11716 12817 11744
rect 12676 11704 12682 11716
rect 12805 11713 12817 11716
rect 12851 11713 12863 11747
rect 16758 11744 16764 11756
rect 12805 11707 12863 11713
rect 16132 11716 16764 11744
rect 7024 11648 7880 11676
rect 7024 11608 7052 11648
rect 8202 11636 8208 11688
rect 8260 11676 8266 11688
rect 8849 11679 8907 11685
rect 8849 11676 8861 11679
rect 8260 11648 8861 11676
rect 8260 11636 8266 11648
rect 8849 11645 8861 11648
rect 8895 11645 8907 11679
rect 8849 11639 8907 11645
rect 9674 11636 9680 11688
rect 9732 11676 9738 11688
rect 10502 11685 10508 11688
rect 10496 11676 10508 11685
rect 9732 11648 9777 11676
rect 10463 11648 10508 11676
rect 9732 11636 9738 11648
rect 10496 11639 10508 11648
rect 10502 11636 10508 11639
rect 10560 11636 10566 11688
rect 13998 11676 14004 11688
rect 13004 11648 14004 11676
rect 6012 11580 7052 11608
rect 7092 11611 7150 11617
rect 7092 11577 7104 11611
rect 7138 11608 7150 11611
rect 8386 11608 8392 11620
rect 7138 11580 8392 11608
rect 7138 11577 7150 11580
rect 7092 11571 7150 11577
rect 8386 11568 8392 11580
rect 8444 11568 8450 11620
rect 13004 11608 13032 11648
rect 13998 11636 14004 11648
rect 14056 11636 14062 11688
rect 14461 11679 14519 11685
rect 14461 11645 14473 11679
rect 14507 11676 14519 11679
rect 14550 11676 14556 11688
rect 14507 11648 14556 11676
rect 14507 11645 14519 11648
rect 14461 11639 14519 11645
rect 14550 11636 14556 11648
rect 14608 11636 14614 11688
rect 14734 11685 14740 11688
rect 14728 11676 14740 11685
rect 14695 11648 14740 11676
rect 14728 11639 14740 11648
rect 14734 11636 14740 11639
rect 14792 11636 14798 11688
rect 11164 11580 13032 11608
rect 13072 11611 13130 11617
rect 1857 11543 1915 11549
rect 1857 11509 1869 11543
rect 1903 11540 1915 11543
rect 3602 11540 3608 11552
rect 1903 11512 3608 11540
rect 1903 11509 1915 11512
rect 1857 11503 1915 11509
rect 3602 11500 3608 11512
rect 3660 11500 3666 11552
rect 3786 11500 3792 11552
rect 3844 11540 3850 11552
rect 4338 11540 4344 11552
rect 3844 11512 4344 11540
rect 3844 11500 3850 11512
rect 4338 11500 4344 11512
rect 4396 11540 4402 11552
rect 4522 11540 4528 11552
rect 4396 11512 4528 11540
rect 4396 11500 4402 11512
rect 4522 11500 4528 11512
rect 4580 11500 4586 11552
rect 7926 11500 7932 11552
rect 7984 11540 7990 11552
rect 8205 11543 8263 11549
rect 8205 11540 8217 11543
rect 7984 11512 8217 11540
rect 7984 11500 7990 11512
rect 8205 11509 8217 11512
rect 8251 11540 8263 11543
rect 8941 11543 8999 11549
rect 8941 11540 8953 11543
rect 8251 11512 8953 11540
rect 8251 11509 8263 11512
rect 8205 11503 8263 11509
rect 8941 11509 8953 11512
rect 8987 11509 8999 11543
rect 8941 11503 8999 11509
rect 9861 11543 9919 11549
rect 9861 11509 9873 11543
rect 9907 11540 9919 11543
rect 11164 11540 11192 11580
rect 13072 11577 13084 11611
rect 13118 11608 13130 11611
rect 16132 11608 16160 11716
rect 16758 11704 16764 11716
rect 16816 11704 16822 11756
rect 17402 11744 17408 11756
rect 17363 11716 17408 11744
rect 17402 11704 17408 11716
rect 17460 11704 17466 11756
rect 17589 11747 17647 11753
rect 17589 11713 17601 11747
rect 17635 11744 17647 11747
rect 17862 11744 17868 11756
rect 17635 11716 17868 11744
rect 17635 11713 17647 11716
rect 17589 11707 17647 11713
rect 17862 11704 17868 11716
rect 17920 11704 17926 11756
rect 19886 11704 19892 11756
rect 19944 11744 19950 11756
rect 20165 11747 20223 11753
rect 20165 11744 20177 11747
rect 19944 11716 20177 11744
rect 19944 11704 19950 11716
rect 20165 11713 20177 11716
rect 20211 11713 20223 11747
rect 20165 11707 20223 11713
rect 20346 11704 20352 11756
rect 20404 11744 20410 11756
rect 20628 11747 20686 11753
rect 20628 11744 20640 11747
rect 20404 11716 20640 11744
rect 20404 11704 20410 11716
rect 20628 11713 20640 11716
rect 20674 11713 20686 11747
rect 21910 11744 21916 11756
rect 20628 11707 20686 11713
rect 20824 11716 21916 11744
rect 16485 11679 16543 11685
rect 16485 11645 16497 11679
rect 16531 11676 16543 11679
rect 16853 11679 16911 11685
rect 16853 11676 16865 11679
rect 16531 11648 16865 11676
rect 16531 11645 16543 11648
rect 16485 11639 16543 11645
rect 16853 11645 16865 11648
rect 16899 11645 16911 11679
rect 16853 11639 16911 11645
rect 17310 11636 17316 11688
rect 17368 11676 17374 11688
rect 17368 11648 17413 11676
rect 17368 11636 17374 11648
rect 18138 11636 18144 11688
rect 18196 11676 18202 11688
rect 18233 11679 18291 11685
rect 18233 11676 18245 11679
rect 18196 11648 18245 11676
rect 18196 11636 18202 11648
rect 18233 11645 18245 11648
rect 18279 11645 18291 11679
rect 18233 11639 18291 11645
rect 18500 11679 18558 11685
rect 18500 11645 18512 11679
rect 18546 11676 18558 11679
rect 19058 11676 19064 11688
rect 18546 11648 19064 11676
rect 18546 11645 18558 11648
rect 18500 11639 18558 11645
rect 19058 11636 19064 11648
rect 19116 11636 19122 11688
rect 20824 11676 20852 11716
rect 21910 11704 21916 11716
rect 21968 11704 21974 11756
rect 20272 11648 20852 11676
rect 20901 11679 20959 11685
rect 13118 11580 16160 11608
rect 16301 11611 16359 11617
rect 13118 11577 13130 11580
rect 13072 11571 13130 11577
rect 14568 11552 14596 11580
rect 16301 11577 16313 11611
rect 16347 11608 16359 11611
rect 19334 11608 19340 11620
rect 16347 11580 19340 11608
rect 16347 11577 16359 11580
rect 16301 11571 16359 11577
rect 19334 11568 19340 11580
rect 19392 11568 19398 11620
rect 9907 11512 11192 11540
rect 11885 11543 11943 11549
rect 9907 11509 9919 11512
rect 9861 11503 9919 11509
rect 11885 11509 11897 11543
rect 11931 11540 11943 11543
rect 13814 11540 13820 11552
rect 11931 11512 13820 11540
rect 11931 11509 11943 11512
rect 11885 11503 11943 11509
rect 13814 11500 13820 11512
rect 13872 11500 13878 11552
rect 14550 11500 14556 11552
rect 14608 11500 14614 11552
rect 16206 11500 16212 11552
rect 16264 11540 16270 11552
rect 16669 11543 16727 11549
rect 16669 11540 16681 11543
rect 16264 11512 16681 11540
rect 16264 11500 16270 11512
rect 16669 11509 16681 11512
rect 16715 11509 16727 11543
rect 16669 11503 16727 11509
rect 16853 11543 16911 11549
rect 16853 11509 16865 11543
rect 16899 11540 16911 11543
rect 18046 11540 18052 11552
rect 16899 11512 18052 11540
rect 16899 11509 16911 11512
rect 16853 11503 16911 11509
rect 18046 11500 18052 11512
rect 18104 11500 18110 11552
rect 18322 11500 18328 11552
rect 18380 11540 18386 11552
rect 18966 11540 18972 11552
rect 18380 11512 18972 11540
rect 18380 11500 18386 11512
rect 18966 11500 18972 11512
rect 19024 11500 19030 11552
rect 19610 11540 19616 11552
rect 19523 11512 19616 11540
rect 19610 11500 19616 11512
rect 19668 11540 19674 11552
rect 20272 11540 20300 11648
rect 20901 11645 20913 11679
rect 20947 11676 20959 11679
rect 21266 11676 21272 11688
rect 20947 11648 21272 11676
rect 20947 11645 20959 11648
rect 20901 11639 20959 11645
rect 21266 11636 21272 11648
rect 21324 11636 21330 11688
rect 22278 11676 22284 11688
rect 22239 11648 22284 11676
rect 22278 11636 22284 11648
rect 22336 11636 22342 11688
rect 19668 11512 20300 11540
rect 19668 11500 19674 11512
rect 20530 11500 20536 11552
rect 20588 11540 20594 11552
rect 20631 11543 20689 11549
rect 20631 11540 20643 11543
rect 20588 11512 20643 11540
rect 20588 11500 20594 11512
rect 20631 11509 20643 11512
rect 20677 11509 20689 11543
rect 20631 11503 20689 11509
rect 20806 11500 20812 11552
rect 20864 11540 20870 11552
rect 22005 11543 22063 11549
rect 22005 11540 22017 11543
rect 20864 11512 22017 11540
rect 20864 11500 20870 11512
rect 22005 11509 22017 11512
rect 22051 11509 22063 11543
rect 22005 11503 22063 11509
rect 1104 11450 23276 11472
rect 1104 11398 8379 11450
rect 8431 11398 8443 11450
rect 8495 11398 8507 11450
rect 8559 11398 8571 11450
rect 8623 11398 15776 11450
rect 15828 11398 15840 11450
rect 15892 11398 15904 11450
rect 15956 11398 15968 11450
rect 16020 11398 23276 11450
rect 1104 11376 23276 11398
rect 1578 11336 1584 11348
rect 1539 11308 1584 11336
rect 1578 11296 1584 11308
rect 1636 11296 1642 11348
rect 2130 11296 2136 11348
rect 2188 11336 2194 11348
rect 3786 11336 3792 11348
rect 2188 11308 3792 11336
rect 2188 11296 2194 11308
rect 3786 11296 3792 11308
rect 3844 11296 3850 11348
rect 5442 11336 5448 11348
rect 3988 11308 4476 11336
rect 5403 11308 5448 11336
rect 2216 11271 2274 11277
rect 2216 11237 2228 11271
rect 2262 11268 2274 11271
rect 2774 11268 2780 11280
rect 2262 11240 2780 11268
rect 2262 11237 2274 11240
rect 2216 11231 2274 11237
rect 2774 11228 2780 11240
rect 2832 11268 2838 11280
rect 3142 11268 3148 11280
rect 2832 11240 3148 11268
rect 2832 11228 2838 11240
rect 3142 11228 3148 11240
rect 3200 11228 3206 11280
rect 1397 11203 1455 11209
rect 1397 11169 1409 11203
rect 1443 11200 1455 11203
rect 3988 11200 4016 11308
rect 4246 11228 4252 11280
rect 4304 11277 4310 11280
rect 4304 11271 4368 11277
rect 4304 11237 4322 11271
rect 4356 11237 4368 11271
rect 4304 11231 4368 11237
rect 4304 11228 4310 11231
rect 1443 11172 4016 11200
rect 4065 11203 4123 11209
rect 1443 11169 1455 11172
rect 1397 11163 1455 11169
rect 4065 11169 4077 11203
rect 4111 11200 4123 11203
rect 4154 11200 4160 11212
rect 4111 11172 4160 11200
rect 4111 11169 4123 11172
rect 4065 11163 4123 11169
rect 4154 11160 4160 11172
rect 4212 11160 4218 11212
rect 4448 11200 4476 11308
rect 5442 11296 5448 11308
rect 5500 11296 5506 11348
rect 5810 11296 5816 11348
rect 5868 11336 5874 11348
rect 6089 11339 6147 11345
rect 6089 11336 6101 11339
rect 5868 11308 6101 11336
rect 5868 11296 5874 11308
rect 6089 11305 6101 11308
rect 6135 11305 6147 11339
rect 9398 11336 9404 11348
rect 6089 11299 6147 11305
rect 6748 11308 9404 11336
rect 5460 11268 5488 11296
rect 6181 11271 6239 11277
rect 6181 11268 6193 11271
rect 5460 11240 6193 11268
rect 6181 11237 6193 11240
rect 6227 11237 6239 11271
rect 6181 11231 6239 11237
rect 6086 11200 6092 11212
rect 4448 11172 6092 11200
rect 6086 11160 6092 11172
rect 6144 11160 6150 11212
rect 6748 11200 6776 11308
rect 9398 11296 9404 11308
rect 9456 11296 9462 11348
rect 10502 11296 10508 11348
rect 10560 11336 10566 11348
rect 11333 11339 11391 11345
rect 11333 11336 11345 11339
rect 10560 11308 11345 11336
rect 10560 11296 10566 11308
rect 11333 11305 11345 11308
rect 11379 11305 11391 11339
rect 11333 11299 11391 11305
rect 11514 11296 11520 11348
rect 11572 11336 11578 11348
rect 19334 11336 19340 11348
rect 11572 11308 19340 11336
rect 11572 11296 11578 11308
rect 19334 11296 19340 11308
rect 19392 11296 19398 11348
rect 20162 11336 20168 11348
rect 19720 11308 20168 11336
rect 8941 11271 8999 11277
rect 8941 11237 8953 11271
rect 8987 11268 8999 11271
rect 9950 11268 9956 11280
rect 8987 11240 9956 11268
rect 8987 11237 8999 11240
rect 8941 11231 8999 11237
rect 9950 11228 9956 11240
rect 10008 11228 10014 11280
rect 14553 11271 14611 11277
rect 12176 11240 14504 11268
rect 6914 11200 6920 11212
rect 6196 11172 6776 11200
rect 6875 11172 6920 11200
rect 1946 11132 1952 11144
rect 1907 11104 1952 11132
rect 1946 11092 1952 11104
rect 2004 11092 2010 11144
rect 5534 11092 5540 11144
rect 5592 11132 5598 11144
rect 6196 11132 6224 11172
rect 6914 11160 6920 11172
rect 6972 11160 6978 11212
rect 7184 11203 7242 11209
rect 7184 11169 7196 11203
rect 7230 11200 7242 11203
rect 8202 11200 8208 11212
rect 7230 11172 8208 11200
rect 7230 11169 7242 11172
rect 7184 11163 7242 11169
rect 8202 11160 8208 11172
rect 8260 11160 8266 11212
rect 8754 11160 8760 11212
rect 8812 11200 8818 11212
rect 9582 11200 9588 11212
rect 8812 11172 9588 11200
rect 8812 11160 8818 11172
rect 9582 11160 9588 11172
rect 9640 11160 9646 11212
rect 10042 11200 10048 11212
rect 9968 11172 10048 11200
rect 6362 11132 6368 11144
rect 5592 11104 6224 11132
rect 6323 11104 6368 11132
rect 5592 11092 5598 11104
rect 6362 11092 6368 11104
rect 6420 11092 6426 11144
rect 9030 11132 9036 11144
rect 8991 11104 9036 11132
rect 9030 11092 9036 11104
rect 9088 11092 9094 11144
rect 9217 11135 9275 11141
rect 9217 11101 9229 11135
rect 9263 11132 9275 11135
rect 9306 11132 9312 11144
rect 9263 11104 9312 11132
rect 9263 11101 9275 11104
rect 9217 11095 9275 11101
rect 9306 11092 9312 11104
rect 9364 11092 9370 11144
rect 9968 11141 9996 11172
rect 10042 11160 10048 11172
rect 10100 11160 10106 11212
rect 10220 11203 10278 11209
rect 10220 11169 10232 11203
rect 10266 11200 10278 11203
rect 11146 11200 11152 11212
rect 10266 11172 11152 11200
rect 10266 11169 10278 11172
rect 10220 11163 10278 11169
rect 11146 11160 11152 11172
rect 11204 11160 11210 11212
rect 11606 11200 11612 11212
rect 11567 11172 11612 11200
rect 11606 11160 11612 11172
rect 11664 11160 11670 11212
rect 9953 11135 10011 11141
rect 9953 11101 9965 11135
rect 9999 11101 10011 11135
rect 9953 11095 10011 11101
rect 3326 11064 3332 11076
rect 3287 11036 3332 11064
rect 3326 11024 3332 11036
rect 3384 11024 3390 11076
rect 8573 11067 8631 11073
rect 5552 11036 5856 11064
rect 2590 10956 2596 11008
rect 2648 10996 2654 11008
rect 5552 10996 5580 11036
rect 5718 10996 5724 11008
rect 2648 10968 5580 10996
rect 5679 10968 5724 10996
rect 2648 10956 2654 10968
rect 5718 10956 5724 10968
rect 5776 10956 5782 11008
rect 5828 10996 5856 11036
rect 8128 11036 8432 11064
rect 8128 10996 8156 11036
rect 8294 10996 8300 11008
rect 5828 10968 8156 10996
rect 8255 10968 8300 10996
rect 8294 10956 8300 10968
rect 8352 10956 8358 11008
rect 8404 10996 8432 11036
rect 8573 11033 8585 11067
rect 8619 11064 8631 11067
rect 9858 11064 9864 11076
rect 8619 11036 9864 11064
rect 8619 11033 8631 11036
rect 8573 11027 8631 11033
rect 9858 11024 9864 11036
rect 9916 11024 9922 11076
rect 10962 11024 10968 11076
rect 11020 11064 11026 11076
rect 11793 11067 11851 11073
rect 11793 11064 11805 11067
rect 11020 11036 11805 11064
rect 11020 11024 11026 11036
rect 11793 11033 11805 11036
rect 11839 11033 11851 11067
rect 11793 11027 11851 11033
rect 12176 10996 12204 11240
rect 12434 11200 12440 11212
rect 12395 11172 12440 11200
rect 12434 11160 12440 11172
rect 12492 11160 12498 11212
rect 12529 11203 12587 11209
rect 12529 11169 12541 11203
rect 12575 11200 12587 11203
rect 12618 11200 12624 11212
rect 12575 11172 12624 11200
rect 12575 11169 12587 11172
rect 12529 11163 12587 11169
rect 12618 11160 12624 11172
rect 12676 11160 12682 11212
rect 12796 11203 12854 11209
rect 12796 11169 12808 11203
rect 12842 11200 12854 11203
rect 14274 11200 14280 11212
rect 12842 11172 14280 11200
rect 12842 11169 12854 11172
rect 12796 11163 12854 11169
rect 14274 11160 14280 11172
rect 14332 11160 14338 11212
rect 14476 11200 14504 11240
rect 14553 11237 14565 11271
rect 14599 11268 14611 11271
rect 15286 11268 15292 11280
rect 14599 11240 15292 11268
rect 14599 11237 14611 11240
rect 14553 11231 14611 11237
rect 15286 11228 15292 11240
rect 15344 11228 15350 11280
rect 15832 11271 15890 11277
rect 15488 11240 15792 11268
rect 15488 11200 15516 11240
rect 14476 11172 15516 11200
rect 15565 11203 15623 11209
rect 14642 11132 14648 11144
rect 14603 11104 14648 11132
rect 14642 11092 14648 11104
rect 14700 11092 14706 11144
rect 14752 11141 14780 11172
rect 15565 11169 15577 11203
rect 15611 11200 15623 11203
rect 15654 11200 15660 11212
rect 15611 11172 15660 11200
rect 15611 11169 15623 11172
rect 15565 11163 15623 11169
rect 15654 11160 15660 11172
rect 15712 11160 15718 11212
rect 15764 11200 15792 11240
rect 15832 11237 15844 11271
rect 15878 11268 15890 11271
rect 16482 11268 16488 11280
rect 15878 11240 16488 11268
rect 15878 11237 15890 11240
rect 15832 11231 15890 11237
rect 16482 11228 16488 11240
rect 16540 11228 16546 11280
rect 18138 11268 18144 11280
rect 17236 11240 18144 11268
rect 16666 11200 16672 11212
rect 15764 11172 16672 11200
rect 16666 11160 16672 11172
rect 16724 11160 16730 11212
rect 16758 11160 16764 11212
rect 16816 11200 16822 11212
rect 17236 11209 17264 11240
rect 18138 11228 18144 11240
rect 18196 11268 18202 11280
rect 19144 11271 19202 11277
rect 18196 11240 18920 11268
rect 18196 11228 18202 11240
rect 18892 11212 18920 11240
rect 19144 11237 19156 11271
rect 19190 11268 19202 11271
rect 19610 11268 19616 11280
rect 19190 11240 19616 11268
rect 19190 11237 19202 11240
rect 19144 11231 19202 11237
rect 19610 11228 19616 11240
rect 19668 11228 19674 11280
rect 17221 11203 17279 11209
rect 17221 11200 17233 11203
rect 16816 11172 17233 11200
rect 16816 11160 16822 11172
rect 17144 11144 17172 11172
rect 17221 11169 17233 11172
rect 17267 11169 17279 11203
rect 17221 11163 17279 11169
rect 17310 11160 17316 11212
rect 17368 11200 17374 11212
rect 17477 11203 17535 11209
rect 17477 11200 17489 11203
rect 17368 11172 17489 11200
rect 17368 11160 17374 11172
rect 17477 11169 17489 11172
rect 17523 11169 17535 11203
rect 18874 11200 18880 11212
rect 18787 11172 18880 11200
rect 17477 11163 17535 11169
rect 18874 11160 18880 11172
rect 18932 11160 18938 11212
rect 19720 11200 19748 11308
rect 20162 11296 20168 11308
rect 20220 11296 20226 11348
rect 20438 11296 20444 11348
rect 20496 11336 20502 11348
rect 20622 11336 20628 11348
rect 20496 11308 20628 11336
rect 20496 11296 20502 11308
rect 20622 11296 20628 11308
rect 20680 11296 20686 11348
rect 20901 11339 20959 11345
rect 20901 11305 20913 11339
rect 20947 11336 20959 11339
rect 22186 11336 22192 11348
rect 20947 11308 22192 11336
rect 20947 11305 20959 11308
rect 20901 11299 20959 11305
rect 22186 11296 22192 11308
rect 22244 11296 22250 11348
rect 18984 11172 19748 11200
rect 14737 11135 14795 11141
rect 14737 11101 14749 11135
rect 14783 11101 14795 11135
rect 14737 11095 14795 11101
rect 17126 11092 17132 11144
rect 17184 11092 17190 11144
rect 18322 11092 18328 11144
rect 18380 11132 18386 11144
rect 18984 11132 19012 11172
rect 20990 11160 20996 11212
rect 21048 11200 21054 11212
rect 21617 11203 21675 11209
rect 21617 11200 21629 11203
rect 21048 11172 21629 11200
rect 21048 11160 21054 11172
rect 21617 11169 21629 11172
rect 21663 11169 21675 11203
rect 21617 11163 21675 11169
rect 18380 11104 19012 11132
rect 18380 11092 18386 11104
rect 20254 11092 20260 11144
rect 20312 11132 20318 11144
rect 20622 11132 20628 11144
rect 20312 11104 20628 11132
rect 20312 11092 20318 11104
rect 20622 11092 20628 11104
rect 20680 11092 20686 11144
rect 20898 11092 20904 11144
rect 20956 11132 20962 11144
rect 21361 11135 21419 11141
rect 21361 11132 21373 11135
rect 20956 11104 21373 11132
rect 20956 11092 20962 11104
rect 21361 11101 21373 11104
rect 21407 11101 21419 11135
rect 21361 11095 21419 11101
rect 15010 11064 15016 11076
rect 13464 11036 15016 11064
rect 8404 10968 12204 10996
rect 12253 10999 12311 11005
rect 12253 10965 12265 10999
rect 12299 10996 12311 10999
rect 13464 10996 13492 11036
rect 15010 11024 15016 11036
rect 15068 11024 15074 11076
rect 18230 11024 18236 11076
rect 18288 11064 18294 11076
rect 18601 11067 18659 11073
rect 18601 11064 18613 11067
rect 18288 11036 18613 11064
rect 18288 11024 18294 11036
rect 18601 11033 18613 11036
rect 18647 11033 18659 11067
rect 18601 11027 18659 11033
rect 19978 11024 19984 11076
rect 20036 11064 20042 11076
rect 20438 11064 20444 11076
rect 20036 11036 20444 11064
rect 20036 11024 20042 11036
rect 20438 11024 20444 11036
rect 20496 11024 20502 11076
rect 22741 11067 22799 11073
rect 22741 11033 22753 11067
rect 22787 11064 22799 11067
rect 22830 11064 22836 11076
rect 22787 11036 22836 11064
rect 22787 11033 22799 11036
rect 22741 11027 22799 11033
rect 22830 11024 22836 11036
rect 22888 11024 22894 11076
rect 12299 10968 13492 10996
rect 12299 10965 12311 10968
rect 12253 10959 12311 10965
rect 13538 10956 13544 11008
rect 13596 10996 13602 11008
rect 13906 10996 13912 11008
rect 13596 10968 13912 10996
rect 13596 10956 13602 10968
rect 13906 10956 13912 10968
rect 13964 10956 13970 11008
rect 14182 10996 14188 11008
rect 14143 10968 14188 10996
rect 14182 10956 14188 10968
rect 14240 10956 14246 11008
rect 14366 10956 14372 11008
rect 14424 10996 14430 11008
rect 16945 10999 17003 11005
rect 16945 10996 16957 10999
rect 14424 10968 16957 10996
rect 14424 10956 14430 10968
rect 16945 10965 16957 10968
rect 16991 10996 17003 10999
rect 17494 10996 17500 11008
rect 16991 10968 17500 10996
rect 16991 10965 17003 10968
rect 16945 10959 17003 10965
rect 17494 10956 17500 10968
rect 17552 10956 17558 11008
rect 18782 10956 18788 11008
rect 18840 10996 18846 11008
rect 19058 10996 19064 11008
rect 18840 10968 19064 10996
rect 18840 10956 18846 10968
rect 19058 10956 19064 10968
rect 19116 10956 19122 11008
rect 20254 10996 20260 11008
rect 20215 10968 20260 10996
rect 20254 10956 20260 10968
rect 20312 10956 20318 11008
rect 1104 10906 23276 10928
rect 1104 10854 4680 10906
rect 4732 10854 4744 10906
rect 4796 10854 4808 10906
rect 4860 10854 4872 10906
rect 4924 10854 12078 10906
rect 12130 10854 12142 10906
rect 12194 10854 12206 10906
rect 12258 10854 12270 10906
rect 12322 10854 19475 10906
rect 19527 10854 19539 10906
rect 19591 10854 19603 10906
rect 19655 10854 19667 10906
rect 19719 10854 23276 10906
rect 1104 10832 23276 10854
rect 1486 10792 1492 10804
rect 1447 10764 1492 10792
rect 1486 10752 1492 10764
rect 1544 10752 1550 10804
rect 1762 10792 1768 10804
rect 1723 10764 1768 10792
rect 1762 10752 1768 10764
rect 1820 10752 1826 10804
rect 2133 10795 2191 10801
rect 2133 10761 2145 10795
rect 2179 10792 2191 10795
rect 2179 10764 4108 10792
rect 2179 10761 2191 10764
rect 2133 10755 2191 10761
rect 4080 10724 4108 10764
rect 4246 10752 4252 10804
rect 4304 10792 4310 10804
rect 4525 10795 4583 10801
rect 4525 10792 4537 10795
rect 4304 10764 4537 10792
rect 4304 10752 4310 10764
rect 4525 10761 4537 10764
rect 4571 10761 4583 10795
rect 4525 10755 4583 10761
rect 4801 10795 4859 10801
rect 4801 10761 4813 10795
rect 4847 10792 4859 10795
rect 5074 10792 5080 10804
rect 4847 10764 5080 10792
rect 4847 10761 4859 10764
rect 4801 10755 4859 10761
rect 5074 10752 5080 10764
rect 5132 10752 5138 10804
rect 5902 10792 5908 10804
rect 5863 10764 5908 10792
rect 5902 10752 5908 10764
rect 5960 10752 5966 10804
rect 7190 10792 7196 10804
rect 6012 10764 7196 10792
rect 4338 10724 4344 10736
rect 4080 10696 4344 10724
rect 4338 10684 4344 10696
rect 4396 10684 4402 10736
rect 4614 10684 4620 10736
rect 4672 10724 4678 10736
rect 6012 10724 6040 10764
rect 7190 10752 7196 10764
rect 7248 10752 7254 10804
rect 8202 10792 8208 10804
rect 8163 10764 8208 10792
rect 8202 10752 8208 10764
rect 8260 10752 8266 10804
rect 10870 10792 10876 10804
rect 8312 10764 10876 10792
rect 4672 10696 6040 10724
rect 4672 10684 4678 10696
rect 7834 10684 7840 10736
rect 7892 10724 7898 10736
rect 8312 10724 8340 10764
rect 10870 10752 10876 10764
rect 10928 10752 10934 10804
rect 11146 10792 11152 10804
rect 11107 10764 11152 10792
rect 11146 10752 11152 10764
rect 11204 10752 11210 10804
rect 11422 10752 11428 10804
rect 11480 10792 11486 10804
rect 11609 10795 11667 10801
rect 11609 10792 11621 10795
rect 11480 10764 11621 10792
rect 11480 10752 11486 10764
rect 11609 10761 11621 10764
rect 11655 10761 11667 10795
rect 17310 10792 17316 10804
rect 11609 10755 11667 10761
rect 12459 10764 17316 10792
rect 7892 10696 8340 10724
rect 8389 10727 8447 10733
rect 7892 10684 7898 10696
rect 8389 10693 8401 10727
rect 8435 10724 8447 10727
rect 9306 10724 9312 10736
rect 8435 10696 9312 10724
rect 8435 10693 8447 10696
rect 8389 10687 8447 10693
rect 9306 10684 9312 10696
rect 9364 10724 9370 10736
rect 9493 10727 9551 10733
rect 9493 10724 9505 10727
rect 9364 10696 9505 10724
rect 9364 10684 9370 10696
rect 9493 10693 9505 10696
rect 9539 10693 9551 10727
rect 9766 10724 9772 10736
rect 9493 10687 9551 10693
rect 9692 10696 9772 10724
rect 2777 10659 2835 10665
rect 2777 10625 2789 10659
rect 2823 10656 2835 10659
rect 2823 10628 3280 10656
rect 2823 10625 2835 10628
rect 2777 10619 2835 10625
rect 1486 10548 1492 10600
rect 1544 10588 1550 10600
rect 1581 10591 1639 10597
rect 1581 10588 1593 10591
rect 1544 10560 1593 10588
rect 1544 10548 1550 10560
rect 1581 10557 1593 10560
rect 1627 10557 1639 10591
rect 1581 10551 1639 10557
rect 1946 10548 1952 10600
rect 2004 10588 2010 10600
rect 3145 10591 3203 10597
rect 3145 10588 3157 10591
rect 2004 10560 3157 10588
rect 2004 10548 2010 10560
rect 3145 10557 3157 10560
rect 3191 10557 3203 10591
rect 3252 10588 3280 10628
rect 4522 10616 4528 10668
rect 4580 10656 4586 10668
rect 5353 10659 5411 10665
rect 5353 10656 5365 10659
rect 4580 10628 5365 10656
rect 4580 10616 4586 10628
rect 5353 10625 5365 10628
rect 5399 10625 5411 10659
rect 6641 10659 6699 10665
rect 6641 10656 6653 10659
rect 5353 10619 5411 10625
rect 6104 10628 6653 10656
rect 5166 10588 5172 10600
rect 3252 10560 4660 10588
rect 5127 10560 5172 10588
rect 3145 10551 3203 10557
rect 3412 10523 3470 10529
rect 3412 10489 3424 10523
rect 3458 10520 3470 10523
rect 4062 10520 4068 10532
rect 3458 10492 4068 10520
rect 3458 10489 3470 10492
rect 3412 10483 3470 10489
rect 4062 10480 4068 10492
rect 4120 10480 4126 10532
rect 2498 10452 2504 10464
rect 2459 10424 2504 10452
rect 2498 10412 2504 10424
rect 2556 10412 2562 10464
rect 2593 10455 2651 10461
rect 2593 10421 2605 10455
rect 2639 10452 2651 10455
rect 4522 10452 4528 10464
rect 2639 10424 4528 10452
rect 2639 10421 2651 10424
rect 2593 10415 2651 10421
rect 4522 10412 4528 10424
rect 4580 10412 4586 10464
rect 4632 10452 4660 10560
rect 5166 10548 5172 10560
rect 5224 10548 5230 10600
rect 5261 10591 5319 10597
rect 5261 10557 5273 10591
rect 5307 10588 5319 10591
rect 5718 10588 5724 10600
rect 5307 10560 5724 10588
rect 5307 10557 5319 10560
rect 5261 10551 5319 10557
rect 5718 10548 5724 10560
rect 5776 10548 5782 10600
rect 6104 10597 6132 10628
rect 6641 10625 6653 10628
rect 6687 10625 6699 10659
rect 6641 10619 6699 10625
rect 9125 10659 9183 10665
rect 9125 10625 9137 10659
rect 9171 10656 9183 10659
rect 9214 10656 9220 10668
rect 9171 10628 9220 10656
rect 9171 10625 9183 10628
rect 9125 10619 9183 10625
rect 9214 10616 9220 10628
rect 9272 10616 9278 10668
rect 6089 10591 6147 10597
rect 6089 10557 6101 10591
rect 6135 10557 6147 10591
rect 6089 10551 6147 10557
rect 6178 10548 6184 10600
rect 6236 10588 6242 10600
rect 6825 10591 6883 10597
rect 6236 10560 6281 10588
rect 6236 10548 6242 10560
rect 6825 10557 6837 10591
rect 6871 10588 6883 10591
rect 6914 10588 6920 10600
rect 6871 10560 6920 10588
rect 6871 10557 6883 10560
rect 6825 10551 6883 10557
rect 6914 10548 6920 10560
rect 6972 10548 6978 10600
rect 7092 10591 7150 10597
rect 7092 10557 7104 10591
rect 7138 10588 7150 10591
rect 7926 10588 7932 10600
rect 7138 10560 7932 10588
rect 7138 10557 7150 10560
rect 7092 10551 7150 10557
rect 7926 10548 7932 10560
rect 7984 10548 7990 10600
rect 9692 10597 9720 10696
rect 9766 10684 9772 10696
rect 9824 10684 9830 10736
rect 12459 10724 12487 10764
rect 17310 10752 17316 10764
rect 17368 10752 17374 10804
rect 17402 10752 17408 10804
rect 17460 10792 17466 10804
rect 18049 10795 18107 10801
rect 18049 10792 18061 10795
rect 17460 10764 18061 10792
rect 17460 10752 17466 10764
rect 18049 10761 18061 10764
rect 18095 10761 18107 10795
rect 18049 10755 18107 10761
rect 18874 10752 18880 10804
rect 18932 10792 18938 10804
rect 19061 10795 19119 10801
rect 19061 10792 19073 10795
rect 18932 10764 19073 10792
rect 18932 10752 18938 10764
rect 19061 10761 19073 10764
rect 19107 10761 19119 10795
rect 19061 10755 19119 10761
rect 19242 10752 19248 10804
rect 19300 10792 19306 10804
rect 21177 10795 21235 10801
rect 21177 10792 21189 10795
rect 19300 10764 21189 10792
rect 19300 10752 19306 10764
rect 21177 10761 21189 10764
rect 21223 10792 21235 10795
rect 21266 10792 21272 10804
rect 21223 10764 21272 10792
rect 21223 10761 21235 10764
rect 21177 10755 21235 10761
rect 21266 10752 21272 10764
rect 21324 10752 21330 10804
rect 23198 10792 23204 10804
rect 21376 10764 23204 10792
rect 11348 10696 12487 10724
rect 13817 10727 13875 10733
rect 9677 10591 9735 10597
rect 8036 10560 9628 10588
rect 5810 10480 5816 10532
rect 5868 10520 5874 10532
rect 8036 10520 8064 10560
rect 5868 10492 8064 10520
rect 5868 10480 5874 10492
rect 8294 10480 8300 10532
rect 8352 10520 8358 10532
rect 8941 10523 8999 10529
rect 8941 10520 8953 10523
rect 8352 10492 8953 10520
rect 8352 10480 8358 10492
rect 8941 10489 8953 10492
rect 8987 10489 8999 10523
rect 8941 10483 8999 10489
rect 6178 10452 6184 10464
rect 4632 10424 6184 10452
rect 6178 10412 6184 10424
rect 6236 10412 6242 10464
rect 6362 10452 6368 10464
rect 6323 10424 6368 10452
rect 6362 10412 6368 10424
rect 6420 10412 6426 10464
rect 6641 10455 6699 10461
rect 6641 10421 6653 10455
rect 6687 10452 6699 10455
rect 8389 10455 8447 10461
rect 8389 10452 8401 10455
rect 6687 10424 8401 10452
rect 6687 10421 6699 10424
rect 6641 10415 6699 10421
rect 8389 10421 8401 10424
rect 8435 10421 8447 10455
rect 8389 10415 8447 10421
rect 8481 10455 8539 10461
rect 8481 10421 8493 10455
rect 8527 10452 8539 10455
rect 8662 10452 8668 10464
rect 8527 10424 8668 10452
rect 8527 10421 8539 10424
rect 8481 10415 8539 10421
rect 8662 10412 8668 10424
rect 8720 10412 8726 10464
rect 8846 10452 8852 10464
rect 8807 10424 8852 10452
rect 8846 10412 8852 10424
rect 8904 10412 8910 10464
rect 9600 10452 9628 10560
rect 9677 10557 9689 10591
rect 9723 10557 9735 10591
rect 9677 10551 9735 10557
rect 9769 10591 9827 10597
rect 9769 10557 9781 10591
rect 9815 10588 9827 10591
rect 9858 10588 9864 10600
rect 9815 10560 9864 10588
rect 9815 10557 9827 10560
rect 9769 10551 9827 10557
rect 9858 10548 9864 10560
rect 9916 10548 9922 10600
rect 10502 10548 10508 10600
rect 10560 10588 10566 10600
rect 10962 10588 10968 10600
rect 10560 10560 10968 10588
rect 10560 10548 10566 10560
rect 10962 10548 10968 10560
rect 11020 10548 11026 10600
rect 10036 10523 10094 10529
rect 10036 10489 10048 10523
rect 10082 10520 10094 10523
rect 11054 10520 11060 10532
rect 10082 10492 11060 10520
rect 10082 10489 10094 10492
rect 10036 10483 10094 10489
rect 11054 10480 11060 10492
rect 11112 10480 11118 10532
rect 11348 10452 11376 10696
rect 13817 10693 13829 10727
rect 13863 10724 13875 10727
rect 14274 10724 14280 10736
rect 13863 10696 14280 10724
rect 13863 10693 13875 10696
rect 13817 10687 13875 10693
rect 14274 10684 14280 10696
rect 14332 10684 14338 10736
rect 16482 10684 16488 10736
rect 16540 10724 16546 10736
rect 16577 10727 16635 10733
rect 16577 10724 16589 10727
rect 16540 10696 16589 10724
rect 16540 10684 16546 10696
rect 16577 10693 16589 10696
rect 16623 10724 16635 10727
rect 18506 10724 18512 10736
rect 16623 10696 18512 10724
rect 16623 10693 16635 10696
rect 16577 10687 16635 10693
rect 18506 10684 18512 10696
rect 18564 10684 18570 10736
rect 14366 10656 14372 10668
rect 13832 10628 14372 10656
rect 11425 10591 11483 10597
rect 11425 10557 11437 10591
rect 11471 10557 11483 10591
rect 11425 10551 11483 10557
rect 11440 10520 11468 10551
rect 12434 10548 12440 10600
rect 12492 10588 12498 10600
rect 12704 10591 12762 10597
rect 12492 10560 12537 10588
rect 12492 10548 12498 10560
rect 12704 10557 12716 10591
rect 12750 10588 12762 10591
rect 13832 10588 13860 10628
rect 14366 10616 14372 10628
rect 14424 10616 14430 10668
rect 14734 10656 14740 10668
rect 14695 10628 14740 10656
rect 14734 10616 14740 10628
rect 14792 10616 14798 10668
rect 16206 10616 16212 10668
rect 16264 10656 16270 10668
rect 17494 10656 17500 10668
rect 16264 10628 17356 10656
rect 17455 10628 17500 10656
rect 16264 10616 16270 10628
rect 14553 10591 14611 10597
rect 14553 10588 14565 10591
rect 12750 10560 13860 10588
rect 13924 10560 14565 10588
rect 12750 10557 12762 10560
rect 12704 10551 12762 10557
rect 12526 10520 12532 10532
rect 11440 10492 12532 10520
rect 12526 10480 12532 10492
rect 12584 10480 12590 10532
rect 13814 10480 13820 10532
rect 13872 10520 13878 10532
rect 13924 10520 13952 10560
rect 14553 10557 14565 10560
rect 14599 10557 14611 10591
rect 14553 10551 14611 10557
rect 15197 10591 15255 10597
rect 15197 10557 15209 10591
rect 15243 10557 15255 10591
rect 15197 10551 15255 10557
rect 14645 10523 14703 10529
rect 14645 10520 14657 10523
rect 13872 10492 13952 10520
rect 14108 10492 14657 10520
rect 13872 10480 13878 10492
rect 14108 10464 14136 10492
rect 14645 10489 14657 10492
rect 14691 10489 14703 10523
rect 15212 10520 15240 10551
rect 15286 10548 15292 10600
rect 15344 10588 15350 10600
rect 15453 10591 15511 10597
rect 15453 10588 15465 10591
rect 15344 10560 15465 10588
rect 15344 10548 15350 10560
rect 15453 10557 15465 10560
rect 15499 10557 15511 10591
rect 16942 10588 16948 10600
rect 15453 10551 15511 10557
rect 16500 10560 16948 10588
rect 15654 10520 15660 10532
rect 15212 10492 15660 10520
rect 14645 10483 14703 10489
rect 15654 10480 15660 10492
rect 15712 10480 15718 10532
rect 9600 10424 11376 10452
rect 14090 10412 14096 10464
rect 14148 10412 14154 10464
rect 14185 10455 14243 10461
rect 14185 10421 14197 10455
rect 14231 10452 14243 10455
rect 14918 10452 14924 10464
rect 14231 10424 14924 10452
rect 14231 10421 14243 10424
rect 14185 10415 14243 10421
rect 14918 10412 14924 10424
rect 14976 10412 14982 10464
rect 15102 10412 15108 10464
rect 15160 10452 15166 10464
rect 16500 10452 16528 10560
rect 16942 10548 16948 10560
rect 17000 10548 17006 10600
rect 17328 10597 17356 10628
rect 17494 10616 17500 10628
rect 17552 10616 17558 10668
rect 17586 10616 17592 10668
rect 17644 10656 17650 10668
rect 18601 10659 18659 10665
rect 18601 10656 18613 10659
rect 17644 10628 18613 10656
rect 17644 10616 17650 10628
rect 18601 10625 18613 10628
rect 18647 10625 18659 10659
rect 18601 10619 18659 10625
rect 19610 10616 19616 10668
rect 19668 10656 19674 10668
rect 19800 10659 19858 10665
rect 19800 10656 19812 10659
rect 19668 10628 19812 10656
rect 19668 10616 19674 10628
rect 19800 10625 19812 10628
rect 19846 10656 19858 10659
rect 21376 10656 21404 10764
rect 23198 10752 23204 10764
rect 23256 10752 23262 10804
rect 19846 10628 21404 10656
rect 19846 10625 19858 10628
rect 19800 10619 19858 10625
rect 21542 10616 21548 10668
rect 21600 10656 21606 10668
rect 22189 10659 22247 10665
rect 22189 10656 22201 10659
rect 21600 10628 22201 10656
rect 21600 10616 21606 10628
rect 22189 10625 22201 10628
rect 22235 10625 22247 10659
rect 22189 10619 22247 10625
rect 17313 10591 17371 10597
rect 17313 10557 17325 10591
rect 17359 10557 17371 10591
rect 17313 10551 17371 10557
rect 18046 10548 18052 10600
rect 18104 10588 18110 10600
rect 19245 10591 19303 10597
rect 19245 10588 19257 10591
rect 18104 10560 19257 10588
rect 18104 10548 18110 10560
rect 19245 10557 19257 10560
rect 19291 10557 19303 10591
rect 19245 10551 19303 10557
rect 19337 10591 19395 10597
rect 19337 10557 19349 10591
rect 19383 10588 19395 10591
rect 19702 10588 19708 10600
rect 19383 10560 19708 10588
rect 19383 10557 19395 10560
rect 19337 10551 19395 10557
rect 19702 10548 19708 10560
rect 19760 10548 19766 10600
rect 19886 10548 19892 10600
rect 19944 10588 19950 10600
rect 20073 10591 20131 10597
rect 20073 10588 20085 10591
rect 19944 10560 20085 10588
rect 19944 10548 19950 10560
rect 20073 10557 20085 10560
rect 20119 10557 20131 10591
rect 20073 10551 20131 10557
rect 16666 10480 16672 10532
rect 16724 10520 16730 10532
rect 18138 10520 18144 10532
rect 16724 10492 18144 10520
rect 16724 10480 16730 10492
rect 18138 10480 18144 10492
rect 18196 10520 18202 10532
rect 18509 10523 18567 10529
rect 18509 10520 18521 10523
rect 18196 10492 18521 10520
rect 18196 10480 18202 10492
rect 18509 10489 18521 10492
rect 18555 10520 18567 10523
rect 18782 10520 18788 10532
rect 18555 10492 18788 10520
rect 18555 10489 18567 10492
rect 18509 10483 18567 10489
rect 18782 10480 18788 10492
rect 18840 10480 18846 10532
rect 21910 10480 21916 10532
rect 21968 10520 21974 10532
rect 22097 10523 22155 10529
rect 22097 10520 22109 10523
rect 21968 10492 22109 10520
rect 21968 10480 21974 10492
rect 22097 10489 22109 10492
rect 22143 10489 22155 10523
rect 22097 10483 22155 10489
rect 15160 10424 16528 10452
rect 15160 10412 15166 10424
rect 16574 10412 16580 10464
rect 16632 10452 16638 10464
rect 16850 10452 16856 10464
rect 16632 10424 16856 10452
rect 16632 10412 16638 10424
rect 16850 10412 16856 10424
rect 16908 10452 16914 10464
rect 16945 10455 17003 10461
rect 16945 10452 16957 10455
rect 16908 10424 16957 10452
rect 16908 10412 16914 10424
rect 16945 10421 16957 10424
rect 16991 10421 17003 10455
rect 16945 10415 17003 10421
rect 17402 10412 17408 10464
rect 17460 10452 17466 10464
rect 17460 10424 17505 10452
rect 17460 10412 17466 10424
rect 17954 10412 17960 10464
rect 18012 10452 18018 10464
rect 18417 10455 18475 10461
rect 18417 10452 18429 10455
rect 18012 10424 18429 10452
rect 18012 10412 18018 10424
rect 18417 10421 18429 10424
rect 18463 10421 18475 10455
rect 18417 10415 18475 10421
rect 19242 10412 19248 10464
rect 19300 10452 19306 10464
rect 19803 10455 19861 10461
rect 19803 10452 19815 10455
rect 19300 10424 19815 10452
rect 19300 10412 19306 10424
rect 19803 10421 19815 10424
rect 19849 10452 19861 10455
rect 20438 10452 20444 10464
rect 19849 10424 20444 10452
rect 19849 10421 19861 10424
rect 19803 10415 19861 10421
rect 20438 10412 20444 10424
rect 20496 10412 20502 10464
rect 21266 10412 21272 10464
rect 21324 10452 21330 10464
rect 21637 10455 21695 10461
rect 21637 10452 21649 10455
rect 21324 10424 21649 10452
rect 21324 10412 21330 10424
rect 21637 10421 21649 10424
rect 21683 10452 21695 10455
rect 21818 10452 21824 10464
rect 21683 10424 21824 10452
rect 21683 10421 21695 10424
rect 21637 10415 21695 10421
rect 21818 10412 21824 10424
rect 21876 10412 21882 10464
rect 22002 10452 22008 10464
rect 21963 10424 22008 10452
rect 22002 10412 22008 10424
rect 22060 10412 22066 10464
rect 1104 10362 23276 10384
rect 1104 10310 8379 10362
rect 8431 10310 8443 10362
rect 8495 10310 8507 10362
rect 8559 10310 8571 10362
rect 8623 10310 15776 10362
rect 15828 10310 15840 10362
rect 15892 10310 15904 10362
rect 15956 10310 15968 10362
rect 16020 10310 23276 10362
rect 1104 10288 23276 10310
rect 2590 10248 2596 10260
rect 2551 10220 2596 10248
rect 2590 10208 2596 10220
rect 2648 10208 2654 10260
rect 4065 10251 4123 10257
rect 4065 10217 4077 10251
rect 4111 10217 4123 10251
rect 4065 10211 4123 10217
rect 3329 10183 3387 10189
rect 3329 10149 3341 10183
rect 3375 10180 3387 10183
rect 3694 10180 3700 10192
rect 3375 10152 3700 10180
rect 3375 10149 3387 10152
rect 3329 10143 3387 10149
rect 3694 10140 3700 10152
rect 3752 10140 3758 10192
rect 4080 10180 4108 10211
rect 4246 10208 4252 10260
rect 4304 10248 4310 10260
rect 4433 10251 4491 10257
rect 4433 10248 4445 10251
rect 4304 10220 4445 10248
rect 4304 10208 4310 10220
rect 4433 10217 4445 10220
rect 4479 10217 4491 10251
rect 4433 10211 4491 10217
rect 4525 10251 4583 10257
rect 4525 10217 4537 10251
rect 4571 10248 4583 10251
rect 4614 10248 4620 10260
rect 4571 10220 4620 10248
rect 4571 10217 4583 10220
rect 4525 10211 4583 10217
rect 4614 10208 4620 10220
rect 4672 10208 4678 10260
rect 5445 10251 5503 10257
rect 5445 10217 5457 10251
rect 5491 10248 5503 10251
rect 7834 10248 7840 10260
rect 5491 10220 7840 10248
rect 5491 10217 5503 10220
rect 5445 10211 5503 10217
rect 7834 10208 7840 10220
rect 7892 10208 7898 10260
rect 8481 10251 8539 10257
rect 8481 10217 8493 10251
rect 8527 10248 8539 10251
rect 8846 10248 8852 10260
rect 8527 10220 8852 10248
rect 8527 10217 8539 10220
rect 8481 10211 8539 10217
rect 8846 10208 8852 10220
rect 8904 10208 8910 10260
rect 9217 10251 9275 10257
rect 9217 10217 9229 10251
rect 9263 10248 9275 10251
rect 9401 10251 9459 10257
rect 9401 10248 9413 10251
rect 9263 10220 9413 10248
rect 9263 10217 9275 10220
rect 9217 10211 9275 10217
rect 9401 10217 9413 10220
rect 9447 10217 9459 10251
rect 9401 10211 9459 10217
rect 9493 10251 9551 10257
rect 9493 10217 9505 10251
rect 9539 10248 9551 10251
rect 9674 10248 9680 10260
rect 9539 10220 9680 10248
rect 9539 10217 9551 10220
rect 9493 10211 9551 10217
rect 9674 10208 9680 10220
rect 9732 10208 9738 10260
rect 11054 10248 11060 10260
rect 9784 10220 10079 10248
rect 11015 10220 11060 10248
rect 5537 10183 5595 10189
rect 4080 10152 5488 10180
rect 1857 10115 1915 10121
rect 1857 10081 1869 10115
rect 1903 10081 1915 10115
rect 1857 10075 1915 10081
rect 2409 10115 2467 10121
rect 2409 10081 2421 10115
rect 2455 10112 2467 10115
rect 2682 10112 2688 10124
rect 2455 10084 2688 10112
rect 2455 10081 2467 10084
rect 2409 10075 2467 10081
rect 1872 10044 1900 10075
rect 2682 10072 2688 10084
rect 2740 10072 2746 10124
rect 3421 10115 3479 10121
rect 3421 10081 3433 10115
rect 3467 10112 3479 10115
rect 4154 10112 4160 10124
rect 3467 10084 4160 10112
rect 3467 10081 3479 10084
rect 3421 10075 3479 10081
rect 3436 10044 3464 10075
rect 4154 10072 4160 10084
rect 4212 10072 4218 10124
rect 5460 10112 5488 10152
rect 5537 10149 5549 10183
rect 5583 10180 5595 10183
rect 7190 10180 7196 10192
rect 5583 10152 7196 10180
rect 5583 10149 5595 10152
rect 5537 10143 5595 10149
rect 7190 10140 7196 10152
rect 7248 10140 7254 10192
rect 7368 10183 7426 10189
rect 7368 10149 7380 10183
rect 7414 10180 7426 10183
rect 8202 10180 8208 10192
rect 7414 10152 8208 10180
rect 7414 10149 7426 10152
rect 7368 10143 7426 10149
rect 8202 10140 8208 10152
rect 8260 10140 8266 10192
rect 9784 10180 9812 10220
rect 10051 10192 10079 10220
rect 11054 10208 11060 10220
rect 11112 10248 11118 10260
rect 11793 10251 11851 10257
rect 11793 10248 11805 10251
rect 11112 10220 11805 10248
rect 11112 10208 11118 10220
rect 11793 10217 11805 10220
rect 11839 10217 11851 10251
rect 11793 10211 11851 10217
rect 11974 10208 11980 10260
rect 12032 10248 12038 10260
rect 15102 10248 15108 10260
rect 12032 10220 15108 10248
rect 12032 10208 12038 10220
rect 15102 10208 15108 10220
rect 15160 10208 15166 10260
rect 15286 10208 15292 10260
rect 15344 10248 15350 10260
rect 16669 10251 16727 10257
rect 16669 10248 16681 10251
rect 15344 10220 16681 10248
rect 15344 10208 15350 10220
rect 16669 10217 16681 10220
rect 16715 10217 16727 10251
rect 16669 10211 16727 10217
rect 17310 10208 17316 10260
rect 17368 10248 17374 10260
rect 18417 10251 18475 10257
rect 18417 10248 18429 10251
rect 17368 10220 18429 10248
rect 17368 10208 17374 10220
rect 18417 10217 18429 10220
rect 18463 10217 18475 10251
rect 19334 10248 19340 10260
rect 18417 10211 18475 10217
rect 18616 10220 19340 10248
rect 8956 10152 9812 10180
rect 6362 10112 6368 10124
rect 5460 10084 6368 10112
rect 6362 10072 6368 10084
rect 6420 10072 6426 10124
rect 6457 10115 6515 10121
rect 6457 10081 6469 10115
rect 6503 10081 6515 10115
rect 6457 10075 6515 10081
rect 6549 10115 6607 10121
rect 6549 10081 6561 10115
rect 6595 10112 6607 10115
rect 8956 10112 8984 10152
rect 9858 10140 9864 10192
rect 9916 10189 9922 10192
rect 9916 10183 9980 10189
rect 9916 10149 9934 10183
rect 9968 10149 9980 10183
rect 9916 10143 9980 10149
rect 9916 10140 9922 10143
rect 10033 10140 10039 10192
rect 10091 10140 10097 10192
rect 11146 10140 11152 10192
rect 11204 10180 11210 10192
rect 11701 10183 11759 10189
rect 11701 10180 11713 10183
rect 11204 10152 11713 10180
rect 11204 10140 11210 10152
rect 11701 10149 11713 10152
rect 11747 10149 11759 10183
rect 15194 10180 15200 10192
rect 11701 10143 11759 10149
rect 12636 10152 14320 10180
rect 6595 10084 8984 10112
rect 9033 10115 9091 10121
rect 6595 10081 6607 10084
rect 6549 10075 6607 10081
rect 9033 10081 9045 10115
rect 9079 10112 9091 10115
rect 9493 10115 9551 10121
rect 9493 10112 9505 10115
rect 9079 10084 9505 10112
rect 9079 10081 9091 10084
rect 9033 10075 9091 10081
rect 9493 10081 9505 10084
rect 9539 10081 9551 10115
rect 9493 10075 9551 10081
rect 3602 10044 3608 10056
rect 1872 10016 3464 10044
rect 3563 10016 3608 10044
rect 3602 10004 3608 10016
rect 3660 10004 3666 10056
rect 4709 10047 4767 10053
rect 4709 10013 4721 10047
rect 4755 10044 4767 10047
rect 5258 10044 5264 10056
rect 4755 10016 5264 10044
rect 4755 10013 4767 10016
rect 4709 10007 4767 10013
rect 5258 10004 5264 10016
rect 5316 10004 5322 10056
rect 5721 10047 5779 10053
rect 5721 10013 5733 10047
rect 5767 10044 5779 10047
rect 5810 10044 5816 10056
rect 5767 10016 5816 10044
rect 5767 10013 5779 10016
rect 5721 10007 5779 10013
rect 5810 10004 5816 10016
rect 5868 10004 5874 10056
rect 6472 10044 6500 10075
rect 9582 10072 9588 10124
rect 9640 10112 9646 10124
rect 12636 10121 12664 10152
rect 9677 10115 9735 10121
rect 9677 10112 9689 10115
rect 9640 10084 9689 10112
rect 9640 10072 9646 10084
rect 9677 10081 9689 10084
rect 9723 10081 9735 10115
rect 12621 10115 12679 10121
rect 9677 10075 9735 10081
rect 9784 10084 11928 10112
rect 6733 10047 6791 10053
rect 6472 10016 6592 10044
rect 6564 9988 6592 10016
rect 6733 10013 6745 10047
rect 6779 10013 6791 10047
rect 6733 10007 6791 10013
rect 4246 9936 4252 9988
rect 4304 9976 4310 9988
rect 4304 9948 6500 9976
rect 4304 9936 4310 9948
rect 2041 9911 2099 9917
rect 2041 9877 2053 9911
rect 2087 9908 2099 9911
rect 2130 9908 2136 9920
rect 2087 9880 2136 9908
rect 2087 9877 2099 9880
rect 2041 9871 2099 9877
rect 2130 9868 2136 9880
rect 2188 9868 2194 9920
rect 2961 9911 3019 9917
rect 2961 9877 2973 9911
rect 3007 9908 3019 9911
rect 3050 9908 3056 9920
rect 3007 9880 3056 9908
rect 3007 9877 3019 9880
rect 2961 9871 3019 9877
rect 3050 9868 3056 9880
rect 3108 9868 3114 9920
rect 5077 9911 5135 9917
rect 5077 9877 5089 9911
rect 5123 9908 5135 9911
rect 5626 9908 5632 9920
rect 5123 9880 5632 9908
rect 5123 9877 5135 9880
rect 5077 9871 5135 9877
rect 5626 9868 5632 9880
rect 5684 9868 5690 9920
rect 6086 9908 6092 9920
rect 6047 9880 6092 9908
rect 6086 9868 6092 9880
rect 6144 9868 6150 9920
rect 6472 9908 6500 9948
rect 6546 9936 6552 9988
rect 6604 9936 6610 9988
rect 6748 9976 6776 10007
rect 6914 10004 6920 10056
rect 6972 10044 6978 10056
rect 7101 10047 7159 10053
rect 7101 10044 7113 10047
rect 6972 10016 7113 10044
rect 6972 10004 6978 10016
rect 7101 10013 7113 10016
rect 7147 10013 7159 10047
rect 7101 10007 7159 10013
rect 9214 10004 9220 10056
rect 9272 10044 9278 10056
rect 9784 10044 9812 10084
rect 11900 10053 11928 10084
rect 12621 10081 12633 10115
rect 12667 10081 12679 10115
rect 12621 10075 12679 10081
rect 12980 10115 13038 10121
rect 12980 10081 12992 10115
rect 13026 10112 13038 10115
rect 13538 10112 13544 10124
rect 13026 10084 13544 10112
rect 13026 10081 13038 10084
rect 12980 10075 13038 10081
rect 13538 10072 13544 10084
rect 13596 10072 13602 10124
rect 14292 10056 14320 10152
rect 14384 10152 15200 10180
rect 14384 10121 14412 10152
rect 15194 10140 15200 10152
rect 15252 10140 15258 10192
rect 15654 10180 15660 10192
rect 15304 10152 15660 10180
rect 14369 10115 14427 10121
rect 14369 10081 14381 10115
rect 14415 10081 14427 10115
rect 14369 10075 14427 10081
rect 14550 10072 14556 10124
rect 14608 10072 14614 10124
rect 15010 10072 15016 10124
rect 15068 10112 15074 10124
rect 15304 10121 15332 10152
rect 15654 10140 15660 10152
rect 15712 10180 15718 10192
rect 16482 10180 16488 10192
rect 15712 10152 16488 10180
rect 15712 10140 15718 10152
rect 16482 10140 16488 10152
rect 16540 10140 16546 10192
rect 16942 10140 16948 10192
rect 17000 10180 17006 10192
rect 18616 10180 18644 10220
rect 19334 10208 19340 10220
rect 19392 10208 19398 10260
rect 20533 10251 20591 10257
rect 20533 10217 20545 10251
rect 20579 10217 20591 10251
rect 20533 10211 20591 10217
rect 17000 10152 18644 10180
rect 18693 10183 18751 10189
rect 17000 10140 17006 10152
rect 18693 10149 18705 10183
rect 18739 10180 18751 10183
rect 20438 10180 20444 10192
rect 18739 10152 20444 10180
rect 18739 10149 18751 10152
rect 18693 10143 18751 10149
rect 20438 10140 20444 10152
rect 20496 10140 20502 10192
rect 20548 10180 20576 10211
rect 21450 10208 21456 10260
rect 21508 10248 21514 10260
rect 21818 10248 21824 10260
rect 21508 10220 21824 10248
rect 21508 10208 21514 10220
rect 21818 10208 21824 10220
rect 21876 10208 21882 10260
rect 22462 10208 22468 10260
rect 22520 10248 22526 10260
rect 22557 10251 22615 10257
rect 22557 10248 22569 10251
rect 22520 10220 22569 10248
rect 22520 10208 22526 10220
rect 22557 10217 22569 10220
rect 22603 10217 22615 10251
rect 22557 10211 22615 10217
rect 21168 10183 21226 10189
rect 21168 10180 21180 10183
rect 20548 10152 21180 10180
rect 21168 10149 21180 10152
rect 21214 10180 21226 10183
rect 23014 10180 23020 10192
rect 21214 10152 23020 10180
rect 21214 10149 21226 10152
rect 21168 10143 21226 10149
rect 23014 10140 23020 10152
rect 23072 10140 23078 10192
rect 15105 10115 15163 10121
rect 15105 10112 15117 10115
rect 15068 10084 15117 10112
rect 15068 10072 15074 10084
rect 15105 10081 15117 10084
rect 15151 10081 15163 10115
rect 15289 10115 15347 10121
rect 15289 10112 15301 10115
rect 15105 10075 15163 10081
rect 15212 10084 15301 10112
rect 9272 10016 9812 10044
rect 11885 10047 11943 10053
rect 9272 10004 9278 10016
rect 11885 10013 11897 10047
rect 11931 10013 11943 10047
rect 12710 10044 12716 10056
rect 12671 10016 12716 10044
rect 11885 10007 11943 10013
rect 12710 10004 12716 10016
rect 12768 10004 12774 10056
rect 14274 10004 14280 10056
rect 14332 10004 14338 10056
rect 14568 10044 14596 10072
rect 14476 10016 14596 10044
rect 7006 9976 7012 9988
rect 6748 9948 7012 9976
rect 7006 9936 7012 9948
rect 7064 9936 7070 9988
rect 9401 9979 9459 9985
rect 9401 9945 9413 9979
rect 9447 9976 9459 9979
rect 9582 9976 9588 9988
rect 9447 9948 9588 9976
rect 9447 9945 9459 9948
rect 9401 9939 9459 9945
rect 9582 9936 9588 9948
rect 9640 9936 9646 9988
rect 10686 9936 10692 9988
rect 10744 9976 10750 9988
rect 11333 9979 11391 9985
rect 11333 9976 11345 9979
rect 10744 9948 11345 9976
rect 10744 9936 10750 9948
rect 11333 9945 11345 9948
rect 11379 9945 11391 9979
rect 11333 9939 11391 9945
rect 14093 9979 14151 9985
rect 14093 9945 14105 9979
rect 14139 9976 14151 9979
rect 14476 9976 14504 10016
rect 14642 10004 14648 10056
rect 14700 10044 14706 10056
rect 15212 10044 15240 10084
rect 15289 10081 15301 10084
rect 15335 10081 15347 10115
rect 15289 10075 15347 10081
rect 15378 10072 15384 10124
rect 15436 10112 15442 10124
rect 15545 10115 15603 10121
rect 15545 10112 15557 10115
rect 15436 10084 15557 10112
rect 15436 10072 15442 10084
rect 15545 10081 15557 10084
rect 15591 10081 15603 10115
rect 15545 10075 15603 10081
rect 17037 10115 17095 10121
rect 17037 10081 17049 10115
rect 17083 10112 17095 10115
rect 17126 10112 17132 10124
rect 17083 10084 17132 10112
rect 17083 10081 17095 10084
rect 17037 10075 17095 10081
rect 17126 10072 17132 10084
rect 17184 10072 17190 10124
rect 17310 10121 17316 10124
rect 17304 10075 17316 10121
rect 17368 10112 17374 10124
rect 18230 10112 18236 10124
rect 17368 10084 18236 10112
rect 17310 10072 17316 10075
rect 17368 10072 17374 10084
rect 18230 10072 18236 10084
rect 18288 10072 18294 10124
rect 18598 10072 18604 10124
rect 18656 10112 18662 10124
rect 18874 10112 18880 10124
rect 18656 10084 18880 10112
rect 18656 10072 18662 10084
rect 18874 10072 18880 10084
rect 18932 10112 18938 10124
rect 19426 10121 19432 10124
rect 19153 10115 19211 10121
rect 19153 10112 19165 10115
rect 18932 10084 19165 10112
rect 18932 10072 18938 10084
rect 19153 10081 19165 10084
rect 19199 10081 19211 10115
rect 19420 10112 19432 10121
rect 19339 10084 19432 10112
rect 19153 10075 19211 10081
rect 19420 10075 19432 10084
rect 19484 10112 19490 10124
rect 20254 10112 20260 10124
rect 19484 10084 20260 10112
rect 14700 10016 15240 10044
rect 14700 10004 14706 10016
rect 14139 9948 14504 9976
rect 14553 9979 14611 9985
rect 14139 9945 14151 9948
rect 14093 9939 14151 9945
rect 14553 9945 14565 9979
rect 14599 9976 14611 9979
rect 14599 9948 15332 9976
rect 14599 9945 14611 9948
rect 14553 9939 14611 9945
rect 11974 9908 11980 9920
rect 6472 9880 11980 9908
rect 11974 9868 11980 9880
rect 12032 9868 12038 9920
rect 12434 9868 12440 9920
rect 12492 9908 12498 9920
rect 12618 9908 12624 9920
rect 12492 9880 12624 9908
rect 12492 9868 12498 9880
rect 12618 9868 12624 9880
rect 12676 9868 12682 9920
rect 14921 9911 14979 9917
rect 14921 9877 14933 9911
rect 14967 9908 14979 9911
rect 15010 9908 15016 9920
rect 14967 9880 15016 9908
rect 14967 9877 14979 9880
rect 14921 9871 14979 9877
rect 15010 9868 15016 9880
rect 15068 9868 15074 9920
rect 15304 9908 15332 9948
rect 18874 9936 18880 9988
rect 18932 9976 18938 9988
rect 19058 9976 19064 9988
rect 18932 9948 19064 9976
rect 18932 9936 18938 9948
rect 19058 9936 19064 9948
rect 19116 9936 19122 9988
rect 16022 9908 16028 9920
rect 15304 9880 16028 9908
rect 16022 9868 16028 9880
rect 16080 9868 16086 9920
rect 18322 9868 18328 9920
rect 18380 9908 18386 9920
rect 18690 9908 18696 9920
rect 18380 9880 18696 9908
rect 18380 9868 18386 9880
rect 18690 9868 18696 9880
rect 18748 9868 18754 9920
rect 19168 9908 19196 10075
rect 19426 10072 19432 10075
rect 19484 10072 19490 10084
rect 20254 10072 20260 10084
rect 20312 10072 20318 10124
rect 20898 10044 20904 10056
rect 20732 10016 20904 10044
rect 20732 9908 20760 10016
rect 20898 10004 20904 10016
rect 20956 10004 20962 10056
rect 22186 9936 22192 9988
rect 22244 9976 22250 9988
rect 22281 9979 22339 9985
rect 22281 9976 22293 9979
rect 22244 9948 22293 9976
rect 22244 9936 22250 9948
rect 22281 9945 22293 9948
rect 22327 9976 22339 9979
rect 22922 9976 22928 9988
rect 22327 9948 22928 9976
rect 22327 9945 22339 9948
rect 22281 9939 22339 9945
rect 22922 9936 22928 9948
rect 22980 9936 22986 9988
rect 19168 9880 20760 9908
rect 1104 9818 23276 9840
rect 1104 9766 4680 9818
rect 4732 9766 4744 9818
rect 4796 9766 4808 9818
rect 4860 9766 4872 9818
rect 4924 9766 12078 9818
rect 12130 9766 12142 9818
rect 12194 9766 12206 9818
rect 12258 9766 12270 9818
rect 12322 9766 19475 9818
rect 19527 9766 19539 9818
rect 19591 9766 19603 9818
rect 19655 9766 19667 9818
rect 19719 9766 23276 9818
rect 1104 9744 23276 9766
rect 4522 9704 4528 9716
rect 4483 9676 4528 9704
rect 4522 9664 4528 9676
rect 4580 9664 4586 9716
rect 7006 9704 7012 9716
rect 5460 9676 7012 9704
rect 2774 9596 2780 9648
rect 2832 9636 2838 9648
rect 3329 9639 3387 9645
rect 2832 9608 2877 9636
rect 2832 9596 2838 9608
rect 3329 9605 3341 9639
rect 3375 9636 3387 9639
rect 5460 9636 5488 9676
rect 7006 9664 7012 9676
rect 7064 9664 7070 9716
rect 9766 9704 9772 9716
rect 7760 9676 9260 9704
rect 6270 9636 6276 9648
rect 3375 9608 5488 9636
rect 6196 9608 6276 9636
rect 3375 9605 3387 9608
rect 3329 9599 3387 9605
rect 4246 9568 4252 9580
rect 4207 9540 4252 9568
rect 4246 9528 4252 9540
rect 4304 9528 4310 9580
rect 5169 9571 5227 9577
rect 5169 9537 5181 9571
rect 5215 9568 5227 9571
rect 5258 9568 5264 9580
rect 5215 9540 5264 9568
rect 5215 9537 5227 9540
rect 5169 9531 5227 9537
rect 5258 9528 5264 9540
rect 5316 9528 5322 9580
rect 6196 9577 6224 9608
rect 6270 9596 6276 9608
rect 6328 9596 6334 9648
rect 7760 9577 7788 9676
rect 9030 9596 9036 9648
rect 9088 9636 9094 9648
rect 9125 9639 9183 9645
rect 9125 9636 9137 9639
rect 9088 9608 9137 9636
rect 9088 9596 9094 9608
rect 9125 9605 9137 9608
rect 9171 9605 9183 9639
rect 9232 9636 9260 9676
rect 9416 9676 9772 9704
rect 9416 9636 9444 9676
rect 9766 9664 9772 9676
rect 9824 9664 9830 9716
rect 10042 9664 10048 9716
rect 10100 9704 10106 9716
rect 10781 9707 10839 9713
rect 10781 9704 10793 9707
rect 10100 9676 10793 9704
rect 10100 9664 10106 9676
rect 10781 9673 10793 9676
rect 10827 9673 10839 9707
rect 10781 9667 10839 9673
rect 11808 9676 15424 9704
rect 9232 9608 9444 9636
rect 9125 9599 9183 9605
rect 6181 9571 6239 9577
rect 6181 9537 6193 9571
rect 6227 9537 6239 9571
rect 6181 9531 6239 9537
rect 6365 9571 6423 9577
rect 6365 9537 6377 9571
rect 6411 9568 6423 9571
rect 7745 9571 7803 9577
rect 6411 9540 7696 9568
rect 6411 9537 6423 9540
rect 6365 9531 6423 9537
rect 1397 9503 1455 9509
rect 1397 9469 1409 9503
rect 1443 9500 1455 9503
rect 1946 9500 1952 9512
rect 1443 9472 1952 9500
rect 1443 9469 1455 9472
rect 1397 9463 1455 9469
rect 1946 9460 1952 9472
rect 2004 9460 2010 9512
rect 2866 9460 2872 9512
rect 2924 9500 2930 9512
rect 3145 9503 3203 9509
rect 3145 9500 3157 9503
rect 2924 9472 3157 9500
rect 2924 9460 2930 9472
rect 3145 9469 3157 9472
rect 3191 9469 3203 9503
rect 4890 9500 4896 9512
rect 4851 9472 4896 9500
rect 3145 9463 3203 9469
rect 4890 9460 4896 9472
rect 4948 9460 4954 9512
rect 4985 9503 5043 9509
rect 4985 9469 4997 9503
rect 5031 9500 5043 9503
rect 5350 9500 5356 9512
rect 5031 9472 5356 9500
rect 5031 9469 5043 9472
rect 4985 9463 5043 9469
rect 5350 9460 5356 9472
rect 5408 9460 5414 9512
rect 5629 9503 5687 9509
rect 5629 9469 5641 9503
rect 5675 9500 5687 9503
rect 5994 9500 6000 9512
rect 5675 9472 6000 9500
rect 5675 9469 5687 9472
rect 5629 9463 5687 9469
rect 5994 9460 6000 9472
rect 6052 9500 6058 9512
rect 6089 9503 6147 9509
rect 6089 9500 6101 9503
rect 6052 9472 6101 9500
rect 6052 9460 6058 9472
rect 6089 9469 6101 9472
rect 6135 9469 6147 9503
rect 7190 9500 7196 9512
rect 7151 9472 7196 9500
rect 6089 9463 6147 9469
rect 7190 9460 7196 9472
rect 7248 9460 7254 9512
rect 1486 9392 1492 9444
rect 1544 9432 1550 9444
rect 1642 9435 1700 9441
rect 1642 9432 1654 9435
rect 1544 9404 1654 9432
rect 1544 9392 1550 9404
rect 1642 9401 1654 9404
rect 1688 9401 1700 9435
rect 1642 9395 1700 9401
rect 4157 9435 4215 9441
rect 4157 9401 4169 9435
rect 4203 9432 4215 9435
rect 5074 9432 5080 9444
rect 4203 9404 5080 9432
rect 4203 9401 4215 9404
rect 4157 9395 4215 9401
rect 5074 9392 5080 9404
rect 5132 9392 5138 9444
rect 7668 9432 7696 9540
rect 7745 9537 7757 9571
rect 7791 9537 7803 9571
rect 9140 9568 9168 9599
rect 9416 9577 9444 9608
rect 10410 9596 10416 9648
rect 10468 9636 10474 9648
rect 11333 9639 11391 9645
rect 11333 9636 11345 9639
rect 10468 9608 11345 9636
rect 10468 9596 10474 9608
rect 11333 9605 11345 9608
rect 11379 9605 11391 9639
rect 11333 9599 11391 9605
rect 9401 9571 9459 9577
rect 9140 9540 9352 9568
rect 7745 9531 7803 9537
rect 8012 9503 8070 9509
rect 8012 9469 8024 9503
rect 8058 9500 8070 9503
rect 8846 9500 8852 9512
rect 8058 9472 8852 9500
rect 8058 9469 8070 9472
rect 8012 9463 8070 9469
rect 8846 9460 8852 9472
rect 8904 9460 8910 9512
rect 8938 9460 8944 9512
rect 8996 9500 9002 9512
rect 9324 9500 9352 9540
rect 9401 9537 9413 9571
rect 9447 9537 9459 9571
rect 11808 9568 11836 9676
rect 13449 9639 13507 9645
rect 13449 9605 13461 9639
rect 13495 9636 13507 9639
rect 14090 9636 14096 9648
rect 13495 9608 14096 9636
rect 13495 9605 13507 9608
rect 13449 9599 13507 9605
rect 14090 9596 14096 9608
rect 14148 9596 14154 9648
rect 15396 9636 15424 9676
rect 15470 9664 15476 9716
rect 15528 9704 15534 9716
rect 15841 9707 15899 9713
rect 15841 9704 15853 9707
rect 15528 9676 15853 9704
rect 15528 9664 15534 9676
rect 15841 9673 15853 9676
rect 15887 9673 15899 9707
rect 15841 9667 15899 9673
rect 16025 9707 16083 9713
rect 16025 9673 16037 9707
rect 16071 9704 16083 9707
rect 17310 9704 17316 9716
rect 16071 9676 17316 9704
rect 16071 9673 16083 9676
rect 16025 9667 16083 9673
rect 17310 9664 17316 9676
rect 17368 9664 17374 9716
rect 18230 9664 18236 9716
rect 18288 9704 18294 9716
rect 18288 9676 19472 9704
rect 18288 9664 18294 9676
rect 16117 9639 16175 9645
rect 15396 9608 15516 9636
rect 9401 9531 9459 9537
rect 10704 9540 11836 9568
rect 9657 9503 9715 9509
rect 9657 9500 9669 9503
rect 8996 9472 9168 9500
rect 9324 9472 9669 9500
rect 8996 9460 9002 9472
rect 9140 9432 9168 9472
rect 9657 9469 9669 9472
rect 9703 9469 9715 9503
rect 9657 9463 9715 9469
rect 10704 9432 10732 9540
rect 11882 9528 11888 9580
rect 11940 9568 11946 9580
rect 12618 9568 12624 9580
rect 11940 9540 11985 9568
rect 12084 9540 12624 9568
rect 11940 9528 11946 9540
rect 11701 9503 11759 9509
rect 11701 9469 11713 9503
rect 11747 9500 11759 9503
rect 12084 9500 12112 9540
rect 12618 9528 12624 9540
rect 12676 9528 12682 9580
rect 13081 9571 13139 9577
rect 13081 9537 13093 9571
rect 13127 9537 13139 9571
rect 13998 9568 14004 9580
rect 13959 9540 14004 9568
rect 13081 9531 13139 9537
rect 13096 9500 13124 9531
rect 13998 9528 14004 9540
rect 14056 9528 14062 9580
rect 15488 9568 15516 9608
rect 16117 9605 16129 9639
rect 16163 9636 16175 9639
rect 17402 9636 17408 9648
rect 16163 9608 17408 9636
rect 16163 9605 16175 9608
rect 16117 9599 16175 9605
rect 17402 9596 17408 9608
rect 17460 9596 17466 9648
rect 19444 9636 19472 9676
rect 19981 9639 20039 9645
rect 19981 9636 19993 9639
rect 19444 9608 19993 9636
rect 19981 9605 19993 9608
rect 20027 9605 20039 9639
rect 19981 9599 20039 9605
rect 20165 9639 20223 9645
rect 20165 9605 20177 9639
rect 20211 9605 20223 9639
rect 20165 9599 20223 9605
rect 16574 9568 16580 9580
rect 15488 9540 16580 9568
rect 16574 9528 16580 9540
rect 16632 9528 16638 9580
rect 16758 9568 16764 9580
rect 16719 9540 16764 9568
rect 16758 9528 16764 9540
rect 16816 9528 16822 9580
rect 18230 9528 18236 9580
rect 18288 9568 18294 9580
rect 18512 9571 18570 9577
rect 18512 9568 18524 9571
rect 18288 9540 18524 9568
rect 18288 9528 18294 9540
rect 18512 9537 18524 9540
rect 18558 9537 18570 9571
rect 18782 9568 18788 9580
rect 18743 9540 18788 9568
rect 18512 9531 18570 9537
rect 18782 9528 18788 9540
rect 18840 9528 18846 9580
rect 19426 9528 19432 9580
rect 19484 9568 19490 9580
rect 20180 9568 20208 9599
rect 19484 9540 20208 9568
rect 19484 9528 19490 9540
rect 20254 9528 20260 9580
rect 20312 9568 20318 9580
rect 20717 9571 20775 9577
rect 20717 9568 20729 9571
rect 20312 9540 20729 9568
rect 20312 9528 20318 9540
rect 20717 9537 20729 9540
rect 20763 9537 20775 9571
rect 20717 9531 20775 9537
rect 20898 9528 20904 9580
rect 20956 9568 20962 9580
rect 21361 9571 21419 9577
rect 21361 9568 21373 9571
rect 20956 9540 21373 9568
rect 20956 9528 20962 9540
rect 21361 9537 21373 9540
rect 21407 9537 21419 9571
rect 21361 9531 21419 9537
rect 13538 9500 13544 9512
rect 11747 9472 12112 9500
rect 12176 9472 12940 9500
rect 13096 9472 13544 9500
rect 11747 9469 11759 9472
rect 11701 9463 11759 9469
rect 12176 9432 12204 9472
rect 12802 9432 12808 9444
rect 7668 9404 9076 9432
rect 9140 9404 10732 9432
rect 11716 9404 12204 9432
rect 12763 9404 12808 9432
rect 3694 9364 3700 9376
rect 3655 9336 3700 9364
rect 3694 9324 3700 9336
rect 3752 9324 3758 9376
rect 4062 9364 4068 9376
rect 4023 9336 4068 9364
rect 4062 9324 4068 9336
rect 4120 9324 4126 9376
rect 5718 9364 5724 9376
rect 5679 9336 5724 9364
rect 5718 9324 5724 9336
rect 5776 9324 5782 9376
rect 7377 9367 7435 9373
rect 7377 9333 7389 9367
rect 7423 9364 7435 9367
rect 7466 9364 7472 9376
rect 7423 9336 7472 9364
rect 7423 9333 7435 9336
rect 7377 9327 7435 9333
rect 7466 9324 7472 9336
rect 7524 9324 7530 9376
rect 7834 9324 7840 9376
rect 7892 9364 7898 9376
rect 8938 9364 8944 9376
rect 7892 9336 8944 9364
rect 7892 9324 7898 9336
rect 8938 9324 8944 9336
rect 8996 9324 9002 9376
rect 9048 9364 9076 9404
rect 11716 9364 11744 9404
rect 12802 9392 12808 9404
rect 12860 9392 12866 9444
rect 12912 9432 12940 9472
rect 13538 9460 13544 9472
rect 13596 9460 13602 9512
rect 13630 9460 13636 9512
rect 13688 9500 13694 9512
rect 14461 9503 14519 9509
rect 14461 9500 14473 9503
rect 13688 9472 14473 9500
rect 13688 9460 13694 9472
rect 14461 9469 14473 9472
rect 14507 9500 14519 9503
rect 14550 9500 14556 9512
rect 14507 9472 14556 9500
rect 14507 9469 14519 9472
rect 14461 9463 14519 9469
rect 14550 9460 14556 9472
rect 14608 9460 14614 9512
rect 14734 9509 14740 9512
rect 14728 9500 14740 9509
rect 14695 9472 14740 9500
rect 14728 9463 14740 9472
rect 14734 9460 14740 9463
rect 14792 9460 14798 9512
rect 15010 9460 15016 9512
rect 15068 9500 15074 9512
rect 15068 9472 16611 9500
rect 15068 9460 15074 9472
rect 12912 9404 15240 9432
rect 9048 9336 11744 9364
rect 11793 9367 11851 9373
rect 11793 9333 11805 9367
rect 11839 9364 11851 9367
rect 12437 9367 12495 9373
rect 12437 9364 12449 9367
rect 11839 9336 12449 9364
rect 11839 9333 11851 9336
rect 11793 9327 11851 9333
rect 12437 9333 12449 9336
rect 12483 9333 12495 9367
rect 12894 9364 12900 9376
rect 12855 9336 12900 9364
rect 12437 9327 12495 9333
rect 12894 9324 12900 9336
rect 12952 9324 12958 9376
rect 13814 9364 13820 9376
rect 13775 9336 13820 9364
rect 13814 9324 13820 9336
rect 13872 9324 13878 9376
rect 13909 9367 13967 9373
rect 13909 9333 13921 9367
rect 13955 9364 13967 9367
rect 15102 9364 15108 9376
rect 13955 9336 15108 9364
rect 13955 9333 13967 9336
rect 13909 9327 13967 9333
rect 15102 9324 15108 9336
rect 15160 9324 15166 9376
rect 15212 9364 15240 9404
rect 15378 9392 15384 9444
rect 15436 9432 15442 9444
rect 16485 9435 16543 9441
rect 16485 9432 16497 9435
rect 15436 9404 16497 9432
rect 15436 9392 15442 9404
rect 16485 9401 16497 9404
rect 16531 9401 16543 9435
rect 16583 9432 16611 9472
rect 17034 9460 17040 9512
rect 17092 9500 17098 9512
rect 17129 9503 17187 9509
rect 17129 9500 17141 9503
rect 17092 9472 17141 9500
rect 17092 9460 17098 9472
rect 17129 9469 17141 9472
rect 17175 9469 17187 9503
rect 17129 9463 17187 9469
rect 17865 9503 17923 9509
rect 17865 9469 17877 9503
rect 17911 9469 17923 9503
rect 17865 9463 17923 9469
rect 18049 9503 18107 9509
rect 18049 9469 18061 9503
rect 18095 9500 18107 9503
rect 18372 9503 18430 9509
rect 18095 9472 18184 9500
rect 18095 9469 18107 9472
rect 18049 9463 18107 9469
rect 17880 9432 17908 9463
rect 16583 9404 17908 9432
rect 16485 9395 16543 9401
rect 16025 9367 16083 9373
rect 16025 9364 16037 9367
rect 15212 9336 16037 9364
rect 16025 9333 16037 9336
rect 16071 9333 16083 9367
rect 16574 9364 16580 9376
rect 16535 9336 16580 9364
rect 16025 9327 16083 9333
rect 16574 9324 16580 9336
rect 16632 9324 16638 9376
rect 17310 9364 17316 9376
rect 17271 9336 17316 9364
rect 17310 9324 17316 9336
rect 17368 9324 17374 9376
rect 17681 9367 17739 9373
rect 17681 9333 17693 9367
rect 17727 9364 17739 9367
rect 18046 9364 18052 9376
rect 17727 9336 18052 9364
rect 17727 9333 17739 9336
rect 17681 9327 17739 9333
rect 18046 9324 18052 9336
rect 18104 9324 18110 9376
rect 18156 9364 18184 9472
rect 18372 9469 18384 9503
rect 18418 9500 18430 9503
rect 19242 9500 19248 9512
rect 18418 9472 19248 9500
rect 18418 9469 18430 9472
rect 18372 9463 18430 9469
rect 19242 9460 19248 9472
rect 19300 9460 19306 9512
rect 20438 9460 20444 9512
rect 20496 9500 20502 9512
rect 20533 9503 20591 9509
rect 20533 9500 20545 9503
rect 20496 9472 20545 9500
rect 20496 9460 20502 9472
rect 20533 9469 20545 9472
rect 20579 9469 20591 9503
rect 20533 9463 20591 9469
rect 21628 9503 21686 9509
rect 21628 9469 21640 9503
rect 21674 9500 21686 9503
rect 22186 9500 22192 9512
rect 21674 9472 22192 9500
rect 21674 9469 21686 9472
rect 21628 9463 21686 9469
rect 22186 9460 22192 9472
rect 22244 9460 22250 9512
rect 20625 9435 20683 9441
rect 20625 9432 20637 9435
rect 19444 9404 20637 9432
rect 18506 9364 18512 9376
rect 18156 9336 18512 9364
rect 18506 9324 18512 9336
rect 18564 9324 18570 9376
rect 18782 9324 18788 9376
rect 18840 9364 18846 9376
rect 19444 9364 19472 9404
rect 20625 9401 20637 9404
rect 20671 9401 20683 9435
rect 20625 9395 20683 9401
rect 19886 9364 19892 9376
rect 18840 9336 19472 9364
rect 19847 9336 19892 9364
rect 18840 9324 18846 9336
rect 19886 9324 19892 9336
rect 19944 9324 19950 9376
rect 19981 9367 20039 9373
rect 19981 9333 19993 9367
rect 20027 9364 20039 9367
rect 22741 9367 22799 9373
rect 22741 9364 22753 9367
rect 20027 9336 22753 9364
rect 20027 9333 20039 9336
rect 19981 9327 20039 9333
rect 22741 9333 22753 9336
rect 22787 9333 22799 9367
rect 22741 9327 22799 9333
rect 1104 9274 23276 9296
rect 1104 9222 8379 9274
rect 8431 9222 8443 9274
rect 8495 9222 8507 9274
rect 8559 9222 8571 9274
rect 8623 9222 15776 9274
rect 15828 9222 15840 9274
rect 15892 9222 15904 9274
rect 15956 9222 15968 9274
rect 16020 9222 23276 9274
rect 1104 9200 23276 9222
rect 2961 9163 3019 9169
rect 2961 9129 2973 9163
rect 3007 9160 3019 9163
rect 3510 9160 3516 9172
rect 3007 9132 3516 9160
rect 3007 9129 3019 9132
rect 2961 9123 3019 9129
rect 3510 9120 3516 9132
rect 3568 9120 3574 9172
rect 4154 9120 4160 9172
rect 4212 9160 4218 9172
rect 4709 9163 4767 9169
rect 4709 9160 4721 9163
rect 4212 9132 4721 9160
rect 4212 9120 4218 9132
rect 4709 9129 4721 9132
rect 4755 9129 4767 9163
rect 4709 9123 4767 9129
rect 5626 9120 5632 9172
rect 5684 9160 5690 9172
rect 6181 9163 6239 9169
rect 6181 9160 6193 9163
rect 5684 9132 6193 9160
rect 5684 9120 5690 9132
rect 6181 9129 6193 9132
rect 6227 9129 6239 9163
rect 6181 9123 6239 9129
rect 6546 9120 6552 9172
rect 6604 9160 6610 9172
rect 6733 9163 6791 9169
rect 6733 9160 6745 9163
rect 6604 9132 6745 9160
rect 6604 9120 6610 9132
rect 6733 9129 6745 9132
rect 6779 9129 6791 9163
rect 6733 9123 6791 9129
rect 7101 9163 7159 9169
rect 7101 9129 7113 9163
rect 7147 9160 7159 9163
rect 7282 9160 7288 9172
rect 7147 9132 7288 9160
rect 7147 9129 7159 9132
rect 7101 9123 7159 9129
rect 7282 9120 7288 9132
rect 7340 9120 7346 9172
rect 7742 9160 7748 9172
rect 7703 9132 7748 9160
rect 7742 9120 7748 9132
rect 7800 9120 7806 9172
rect 8113 9163 8171 9169
rect 8113 9129 8125 9163
rect 8159 9160 8171 9163
rect 8662 9160 8668 9172
rect 8159 9132 8668 9160
rect 8159 9129 8171 9132
rect 8113 9123 8171 9129
rect 8662 9120 8668 9132
rect 8720 9120 8726 9172
rect 8757 9163 8815 9169
rect 8757 9129 8769 9163
rect 8803 9160 8815 9163
rect 9674 9160 9680 9172
rect 8803 9132 9536 9160
rect 9635 9132 9680 9160
rect 8803 9129 8815 9132
rect 8757 9123 8815 9129
rect 5077 9095 5135 9101
rect 5077 9061 5089 9095
rect 5123 9092 5135 9095
rect 6914 9092 6920 9104
rect 5123 9064 6920 9092
rect 5123 9061 5135 9064
rect 5077 9055 5135 9061
rect 6914 9052 6920 9064
rect 6972 9052 6978 9104
rect 7193 9095 7251 9101
rect 7193 9061 7205 9095
rect 7239 9092 7251 9095
rect 7466 9092 7472 9104
rect 7239 9064 7472 9092
rect 7239 9061 7251 9064
rect 7193 9055 7251 9061
rect 7466 9052 7472 9064
rect 7524 9052 7530 9104
rect 9306 9092 9312 9104
rect 8964 9064 9312 9092
rect 3421 9027 3479 9033
rect 3421 8993 3433 9027
rect 3467 9024 3479 9027
rect 3970 9024 3976 9036
rect 3467 8996 3976 9024
rect 3467 8993 3479 8996
rect 3421 8987 3479 8993
rect 3970 8984 3976 8996
rect 4028 8984 4034 9036
rect 4157 9027 4215 9033
rect 4157 8993 4169 9027
rect 4203 9024 4215 9027
rect 4430 9024 4436 9036
rect 4203 8996 4436 9024
rect 4203 8993 4215 8996
rect 4157 8987 4215 8993
rect 4430 8984 4436 8996
rect 4488 8984 4494 9036
rect 5169 9027 5227 9033
rect 5169 8993 5181 9027
rect 5215 9024 5227 9027
rect 5350 9024 5356 9036
rect 5215 8996 5356 9024
rect 5215 8993 5227 8996
rect 5169 8987 5227 8993
rect 5350 8984 5356 8996
rect 5408 8984 5414 9036
rect 6089 9027 6147 9033
rect 6089 8993 6101 9027
rect 6135 9024 6147 9027
rect 7650 9024 7656 9036
rect 6135 8996 6868 9024
rect 6135 8993 6147 8996
rect 6089 8987 6147 8993
rect 5261 8959 5319 8965
rect 5261 8925 5273 8959
rect 5307 8925 5319 8959
rect 5261 8919 5319 8925
rect 6365 8959 6423 8965
rect 6365 8925 6377 8959
rect 6411 8925 6423 8959
rect 6840 8956 6868 8996
rect 7208 8996 7656 9024
rect 7208 8956 7236 8996
rect 7650 8984 7656 8996
rect 7708 8984 7714 9036
rect 8110 8984 8116 9036
rect 8168 9024 8174 9036
rect 8964 9033 8992 9064
rect 9306 9052 9312 9064
rect 9364 9052 9370 9104
rect 9508 9092 9536 9132
rect 9674 9120 9680 9132
rect 9732 9120 9738 9172
rect 10045 9163 10103 9169
rect 10045 9129 10057 9163
rect 10091 9160 10103 9163
rect 10686 9160 10692 9172
rect 10091 9132 10692 9160
rect 10091 9129 10103 9132
rect 10045 9123 10103 9129
rect 10686 9120 10692 9132
rect 10744 9120 10750 9172
rect 10962 9120 10968 9172
rect 11020 9160 11026 9172
rect 12621 9163 12679 9169
rect 12621 9160 12633 9163
rect 11020 9132 12633 9160
rect 11020 9120 11026 9132
rect 12621 9129 12633 9132
rect 12667 9160 12679 9163
rect 12894 9160 12900 9172
rect 12667 9132 12900 9160
rect 12667 9129 12679 9132
rect 12621 9123 12679 9129
rect 12894 9120 12900 9132
rect 12952 9120 12958 9172
rect 13173 9163 13231 9169
rect 13173 9129 13185 9163
rect 13219 9160 13231 9163
rect 13722 9160 13728 9172
rect 13219 9132 13728 9160
rect 13219 9129 13231 9132
rect 13173 9123 13231 9129
rect 13722 9120 13728 9132
rect 13780 9120 13786 9172
rect 14734 9120 14740 9172
rect 14792 9160 14798 9172
rect 14921 9163 14979 9169
rect 14921 9160 14933 9163
rect 14792 9132 14933 9160
rect 14792 9120 14798 9132
rect 14921 9129 14933 9132
rect 14967 9129 14979 9163
rect 14921 9123 14979 9129
rect 15102 9120 15108 9172
rect 15160 9160 15166 9172
rect 15286 9160 15292 9172
rect 15160 9132 15292 9160
rect 15160 9120 15166 9132
rect 15286 9120 15292 9132
rect 15344 9120 15350 9172
rect 15378 9120 15384 9172
rect 15436 9160 15442 9172
rect 15657 9163 15715 9169
rect 15657 9160 15669 9163
rect 15436 9132 15669 9160
rect 15436 9120 15442 9132
rect 15657 9129 15669 9132
rect 15703 9129 15715 9163
rect 15657 9123 15715 9129
rect 16390 9120 16396 9172
rect 16448 9160 16454 9172
rect 16485 9163 16543 9169
rect 16485 9160 16497 9163
rect 16448 9132 16497 9160
rect 16448 9120 16454 9132
rect 16485 9129 16497 9132
rect 16531 9129 16543 9163
rect 16485 9123 16543 9129
rect 16666 9120 16672 9172
rect 16724 9160 16730 9172
rect 19334 9160 19340 9172
rect 16724 9132 19340 9160
rect 16724 9120 16730 9132
rect 19334 9120 19340 9132
rect 19392 9120 19398 9172
rect 21910 9160 21916 9172
rect 21871 9132 21916 9160
rect 21910 9120 21916 9132
rect 21968 9120 21974 9172
rect 10594 9092 10600 9104
rect 9508 9064 10600 9092
rect 10594 9052 10600 9064
rect 10652 9092 10658 9104
rect 11422 9092 11428 9104
rect 10652 9064 11428 9092
rect 10652 9052 10658 9064
rect 11422 9052 11428 9064
rect 11480 9052 11486 9104
rect 11606 9052 11612 9104
rect 11664 9092 11670 9104
rect 11664 9064 12655 9092
rect 11664 9052 11670 9064
rect 8205 9027 8263 9033
rect 8205 9024 8217 9027
rect 8168 8996 8217 9024
rect 8168 8984 8174 8996
rect 8205 8993 8217 8996
rect 8251 8993 8263 9027
rect 8205 8987 8263 8993
rect 8949 9027 9007 9033
rect 8949 8993 8961 9027
rect 8995 8993 9007 9027
rect 8949 8987 9007 8993
rect 9036 8984 9042 9036
rect 9094 9033 9100 9036
rect 9094 9027 9116 9033
rect 9104 8993 9116 9027
rect 9094 8987 9116 8993
rect 9094 8984 9100 8987
rect 9858 8984 9864 9036
rect 9916 9024 9922 9036
rect 10137 9027 10195 9033
rect 10137 9024 10149 9027
rect 9916 8996 10149 9024
rect 9916 8984 9922 8996
rect 10137 8993 10149 8996
rect 10183 8993 10195 9027
rect 10137 8987 10195 8993
rect 10689 9027 10747 9033
rect 10689 8993 10701 9027
rect 10735 9024 10747 9027
rect 10870 9024 10876 9036
rect 10735 8996 10876 9024
rect 10735 8993 10747 8996
rect 10689 8987 10747 8993
rect 10870 8984 10876 8996
rect 10928 8984 10934 9036
rect 11508 9027 11566 9033
rect 11508 8993 11520 9027
rect 11554 9024 11566 9027
rect 11554 8996 12572 9024
rect 11554 8993 11566 8996
rect 11508 8987 11566 8993
rect 6840 8928 7236 8956
rect 7377 8959 7435 8965
rect 6365 8919 6423 8925
rect 7377 8925 7389 8959
rect 7423 8956 7435 8959
rect 7834 8956 7840 8968
rect 7423 8928 7840 8956
rect 7423 8925 7435 8928
rect 7377 8919 7435 8925
rect 3605 8891 3663 8897
rect 3605 8857 3617 8891
rect 3651 8888 3663 8891
rect 4246 8888 4252 8900
rect 3651 8860 4252 8888
rect 3651 8857 3663 8860
rect 3605 8851 3663 8857
rect 4246 8848 4252 8860
rect 4304 8888 4310 8900
rect 5276 8888 5304 8919
rect 4304 8860 5304 8888
rect 6380 8888 6408 8919
rect 7834 8916 7840 8928
rect 7892 8916 7898 8968
rect 8389 8959 8447 8965
rect 8389 8925 8401 8959
rect 8435 8956 8447 8959
rect 10229 8959 10287 8965
rect 10229 8956 10241 8959
rect 8435 8928 10241 8956
rect 8435 8925 8447 8928
rect 8389 8919 8447 8925
rect 10229 8925 10241 8928
rect 10275 8956 10287 8959
rect 10502 8956 10508 8968
rect 10275 8928 10508 8956
rect 10275 8925 10287 8928
rect 10229 8919 10287 8925
rect 10502 8916 10508 8928
rect 10560 8916 10566 8968
rect 10594 8916 10600 8968
rect 10652 8956 10658 8968
rect 11241 8959 11299 8965
rect 11241 8956 11253 8959
rect 10652 8928 11253 8956
rect 10652 8916 10658 8928
rect 11241 8925 11253 8928
rect 11287 8925 11299 8959
rect 11241 8919 11299 8925
rect 8202 8888 8208 8900
rect 6380 8860 8208 8888
rect 4304 8848 4310 8860
rect 8202 8848 8208 8860
rect 8260 8848 8266 8900
rect 9490 8848 9496 8900
rect 9548 8888 9554 8900
rect 11146 8888 11152 8900
rect 9548 8860 11152 8888
rect 9548 8848 9554 8860
rect 11146 8848 11152 8860
rect 11204 8848 11210 8900
rect 12544 8888 12572 8996
rect 12627 8956 12655 9064
rect 12710 9052 12716 9104
rect 12768 9092 12774 9104
rect 12768 9064 13584 9092
rect 12768 9052 12774 9064
rect 12989 9027 13047 9033
rect 12989 8993 13001 9027
rect 13035 9024 13047 9027
rect 13078 9024 13084 9036
rect 13035 8996 13084 9024
rect 13035 8993 13047 8996
rect 12989 8987 13047 8993
rect 13078 8984 13084 8996
rect 13136 8984 13142 9036
rect 13556 9033 13584 9064
rect 13998 9052 14004 9104
rect 14056 9052 14062 9104
rect 14458 9052 14464 9104
rect 14516 9092 14522 9104
rect 17212 9095 17270 9101
rect 14516 9064 16344 9092
rect 14516 9052 14522 9064
rect 13541 9027 13599 9033
rect 13541 8993 13553 9027
rect 13587 9024 13599 9027
rect 13630 9024 13636 9036
rect 13587 8996 13636 9024
rect 13587 8993 13599 8996
rect 13541 8987 13599 8993
rect 13630 8984 13636 8996
rect 13688 8984 13694 9036
rect 13808 9027 13866 9033
rect 13808 8993 13820 9027
rect 13854 9024 13866 9027
rect 14016 9024 14044 9052
rect 13854 8996 14587 9024
rect 13854 8993 13866 8996
rect 13808 8987 13866 8993
rect 13170 8956 13176 8968
rect 12627 8928 13176 8956
rect 13170 8916 13176 8928
rect 13228 8916 13234 8968
rect 14559 8888 14587 8996
rect 14642 8984 14648 9036
rect 14700 9024 14706 9036
rect 16316 9033 16344 9064
rect 17212 9061 17224 9095
rect 17258 9092 17270 9095
rect 17586 9092 17592 9104
rect 17258 9064 17592 9092
rect 17258 9061 17270 9064
rect 17212 9055 17270 9061
rect 17586 9052 17592 9064
rect 17644 9052 17650 9104
rect 18874 9052 18880 9104
rect 18932 9092 18938 9104
rect 21269 9095 21327 9101
rect 21269 9092 21281 9095
rect 18932 9064 21281 9092
rect 18932 9052 18938 9064
rect 21269 9061 21281 9064
rect 21315 9061 21327 9095
rect 21269 9055 21327 9061
rect 21726 9052 21732 9104
rect 21784 9092 21790 9104
rect 22373 9095 22431 9101
rect 22373 9092 22385 9095
rect 21784 9064 22385 9092
rect 21784 9052 21790 9064
rect 22373 9061 22385 9064
rect 22419 9061 22431 9095
rect 22373 9055 22431 9061
rect 16301 9027 16359 9033
rect 14700 8996 15976 9024
rect 14700 8984 14706 8996
rect 15746 8956 15752 8968
rect 15707 8928 15752 8956
rect 15746 8916 15752 8928
rect 15804 8916 15810 8968
rect 15841 8959 15899 8965
rect 15841 8925 15853 8959
rect 15887 8925 15899 8959
rect 15948 8956 15976 8996
rect 16301 8993 16313 9027
rect 16347 8993 16359 9027
rect 16301 8987 16359 8993
rect 16482 8984 16488 9036
rect 16540 9024 16546 9036
rect 16945 9027 17003 9033
rect 16945 9024 16957 9027
rect 16540 8996 16957 9024
rect 16540 8984 16546 8996
rect 16945 8993 16957 8996
rect 16991 8993 17003 9027
rect 17954 9024 17960 9036
rect 16945 8987 17003 8993
rect 17052 8996 17960 9024
rect 16390 8956 16396 8968
rect 15948 8928 16396 8956
rect 15841 8919 15899 8925
rect 15470 8888 15476 8900
rect 12544 8860 13584 8888
rect 14559 8860 15476 8888
rect 4341 8823 4399 8829
rect 4341 8789 4353 8823
rect 4387 8820 4399 8823
rect 5442 8820 5448 8832
rect 4387 8792 5448 8820
rect 4387 8789 4399 8792
rect 4341 8783 4399 8789
rect 5442 8780 5448 8792
rect 5500 8780 5506 8832
rect 5721 8823 5779 8829
rect 5721 8789 5733 8823
rect 5767 8820 5779 8823
rect 8570 8820 8576 8832
rect 5767 8792 8576 8820
rect 5767 8789 5779 8792
rect 5721 8783 5779 8789
rect 8570 8780 8576 8792
rect 8628 8780 8634 8832
rect 9217 8823 9275 8829
rect 9217 8789 9229 8823
rect 9263 8820 9275 8823
rect 10686 8820 10692 8832
rect 9263 8792 10692 8820
rect 9263 8789 9275 8792
rect 9217 8783 9275 8789
rect 10686 8780 10692 8792
rect 10744 8780 10750 8832
rect 10873 8823 10931 8829
rect 10873 8789 10885 8823
rect 10919 8820 10931 8823
rect 13446 8820 13452 8832
rect 10919 8792 13452 8820
rect 10919 8789 10931 8792
rect 10873 8783 10931 8789
rect 13446 8780 13452 8792
rect 13504 8780 13510 8832
rect 13556 8820 13584 8860
rect 15470 8848 15476 8860
rect 15528 8848 15534 8900
rect 15654 8848 15660 8900
rect 15712 8888 15718 8900
rect 15856 8888 15884 8919
rect 16390 8916 16396 8928
rect 16448 8916 16454 8968
rect 17052 8956 17080 8996
rect 17954 8984 17960 8996
rect 18012 8984 18018 9036
rect 18322 8984 18328 9036
rect 18380 9024 18386 9036
rect 19041 9027 19099 9033
rect 19041 9024 19053 9027
rect 18380 8996 19053 9024
rect 18380 8984 18386 8996
rect 19041 8993 19053 8996
rect 19087 8993 19099 9027
rect 19041 8987 19099 8993
rect 20346 8984 20352 9036
rect 20404 9024 20410 9036
rect 22281 9027 22339 9033
rect 22281 9024 22293 9027
rect 20404 8996 22293 9024
rect 20404 8984 20410 8996
rect 22281 8993 22293 8996
rect 22327 8993 22339 9027
rect 22281 8987 22339 8993
rect 16500 8928 17080 8956
rect 16500 8900 16528 8928
rect 18598 8916 18604 8968
rect 18656 8956 18662 8968
rect 18785 8959 18843 8965
rect 18785 8956 18797 8959
rect 18656 8928 18797 8956
rect 18656 8916 18662 8928
rect 18785 8925 18797 8928
rect 18831 8925 18843 8959
rect 18785 8919 18843 8925
rect 20622 8916 20628 8968
rect 20680 8956 20686 8968
rect 21361 8959 21419 8965
rect 21361 8956 21373 8959
rect 20680 8928 21373 8956
rect 20680 8916 20686 8928
rect 21361 8925 21373 8928
rect 21407 8925 21419 8959
rect 21361 8919 21419 8925
rect 21450 8916 21456 8968
rect 21508 8956 21514 8968
rect 22462 8956 22468 8968
rect 21508 8928 21553 8956
rect 22423 8928 22468 8956
rect 21508 8916 21514 8928
rect 22462 8916 22468 8928
rect 22520 8916 22526 8968
rect 15712 8860 15884 8888
rect 15712 8848 15718 8860
rect 16482 8848 16488 8900
rect 16540 8848 16546 8900
rect 17880 8860 18460 8888
rect 17880 8820 17908 8860
rect 13556 8792 17908 8820
rect 17954 8780 17960 8832
rect 18012 8820 18018 8832
rect 18325 8823 18383 8829
rect 18325 8820 18337 8823
rect 18012 8792 18337 8820
rect 18012 8780 18018 8792
rect 18325 8789 18337 8792
rect 18371 8789 18383 8823
rect 18432 8820 18460 8860
rect 20165 8823 20223 8829
rect 20165 8820 20177 8823
rect 18432 8792 20177 8820
rect 18325 8783 18383 8789
rect 20165 8789 20177 8792
rect 20211 8820 20223 8823
rect 20254 8820 20260 8832
rect 20211 8792 20260 8820
rect 20211 8789 20223 8792
rect 20165 8783 20223 8789
rect 20254 8780 20260 8792
rect 20312 8780 20318 8832
rect 20901 8823 20959 8829
rect 20901 8789 20913 8823
rect 20947 8820 20959 8823
rect 22278 8820 22284 8832
rect 20947 8792 22284 8820
rect 20947 8789 20959 8792
rect 20901 8783 20959 8789
rect 22278 8780 22284 8792
rect 22336 8780 22342 8832
rect 1104 8730 23276 8752
rect 1104 8678 4680 8730
rect 4732 8678 4744 8730
rect 4796 8678 4808 8730
rect 4860 8678 4872 8730
rect 4924 8678 12078 8730
rect 12130 8678 12142 8730
rect 12194 8678 12206 8730
rect 12258 8678 12270 8730
rect 12322 8678 19475 8730
rect 19527 8678 19539 8730
rect 19591 8678 19603 8730
rect 19655 8678 19667 8730
rect 19719 8678 23276 8730
rect 1104 8656 23276 8678
rect 4062 8576 4068 8628
rect 4120 8616 4126 8628
rect 4341 8619 4399 8625
rect 4341 8616 4353 8619
rect 4120 8588 4353 8616
rect 4120 8576 4126 8588
rect 4341 8585 4353 8588
rect 4387 8585 4399 8619
rect 4341 8579 4399 8585
rect 7009 8619 7067 8625
rect 7009 8585 7021 8619
rect 7055 8616 7067 8619
rect 10321 8619 10379 8625
rect 7055 8588 9444 8616
rect 7055 8585 7067 8588
rect 7009 8579 7067 8585
rect 4706 8548 4712 8560
rect 4667 8520 4712 8548
rect 4706 8508 4712 8520
rect 4764 8508 4770 8560
rect 5721 8551 5779 8557
rect 5721 8517 5733 8551
rect 5767 8517 5779 8551
rect 5721 8511 5779 8517
rect 7377 8551 7435 8557
rect 7377 8517 7389 8551
rect 7423 8548 7435 8551
rect 8386 8548 8392 8560
rect 7423 8520 8392 8548
rect 7423 8517 7435 8520
rect 7377 8511 7435 8517
rect 1854 8440 1860 8492
rect 1912 8480 1918 8492
rect 1949 8483 2007 8489
rect 1949 8480 1961 8483
rect 1912 8452 1961 8480
rect 1912 8440 1918 8452
rect 1949 8449 1961 8452
rect 1995 8449 2007 8483
rect 5350 8480 5356 8492
rect 5311 8452 5356 8480
rect 1949 8443 2007 8449
rect 5350 8440 5356 8452
rect 5408 8440 5414 8492
rect 1762 8412 1768 8424
rect 1723 8384 1768 8412
rect 1762 8372 1768 8384
rect 1820 8372 1826 8424
rect 4157 8415 4215 8421
rect 4157 8381 4169 8415
rect 4203 8412 4215 8415
rect 5736 8412 5764 8511
rect 8386 8508 8392 8520
rect 8444 8508 8450 8560
rect 6270 8480 6276 8492
rect 6231 8452 6276 8480
rect 6270 8440 6276 8452
rect 6328 8440 6334 8492
rect 7926 8480 7932 8492
rect 7887 8452 7932 8480
rect 7926 8440 7932 8452
rect 7984 8440 7990 8492
rect 9416 8480 9444 8588
rect 10321 8585 10333 8619
rect 10367 8616 10379 8619
rect 11698 8616 11704 8628
rect 10367 8588 11704 8616
rect 10367 8585 10379 8588
rect 10321 8579 10379 8585
rect 11698 8576 11704 8588
rect 11756 8576 11762 8628
rect 11790 8576 11796 8628
rect 11848 8616 11854 8628
rect 12069 8619 12127 8625
rect 12069 8616 12081 8619
rect 11848 8588 12081 8616
rect 11848 8576 11854 8588
rect 12069 8585 12081 8588
rect 12115 8616 12127 8619
rect 12802 8616 12808 8628
rect 12115 8588 12808 8616
rect 12115 8585 12127 8588
rect 12069 8579 12127 8585
rect 12802 8576 12808 8588
rect 12860 8576 12866 8628
rect 13170 8576 13176 8628
rect 13228 8616 13234 8628
rect 15470 8616 15476 8628
rect 13228 8588 15148 8616
rect 15431 8588 15476 8616
rect 13228 8576 13234 8588
rect 10597 8551 10655 8557
rect 10597 8548 10609 8551
rect 9692 8520 10609 8548
rect 9692 8480 9720 8520
rect 10597 8517 10609 8520
rect 10643 8517 10655 8551
rect 10597 8511 10655 8517
rect 13446 8508 13452 8560
rect 13504 8548 13510 8560
rect 13817 8551 13875 8557
rect 13817 8548 13829 8551
rect 13504 8520 13829 8548
rect 13504 8508 13510 8520
rect 13817 8517 13829 8520
rect 13863 8517 13875 8551
rect 13817 8511 13875 8517
rect 9416 8452 9720 8480
rect 10060 8452 10640 8480
rect 6822 8412 6828 8424
rect 4203 8384 5764 8412
rect 6012 8384 6684 8412
rect 6783 8384 6828 8412
rect 4203 8381 4215 8384
rect 4157 8375 4215 8381
rect 5169 8347 5227 8353
rect 5169 8313 5181 8347
rect 5215 8344 5227 8347
rect 6012 8344 6040 8384
rect 6178 8344 6184 8356
rect 5215 8316 6040 8344
rect 6139 8316 6184 8344
rect 5215 8313 5227 8316
rect 5169 8307 5227 8313
rect 6178 8304 6184 8316
rect 6236 8304 6242 8356
rect 6656 8344 6684 8384
rect 6822 8372 6828 8384
rect 6880 8372 6886 8424
rect 8389 8415 8447 8421
rect 8389 8381 8401 8415
rect 8435 8412 8447 8415
rect 10060 8412 10088 8452
rect 10612 8424 10640 8452
rect 12434 8440 12440 8492
rect 12492 8480 12498 8492
rect 12492 8452 12537 8480
rect 12492 8440 12498 8452
rect 13630 8440 13636 8492
rect 13688 8480 13694 8492
rect 14093 8483 14151 8489
rect 14093 8480 14105 8483
rect 13688 8452 14105 8480
rect 13688 8440 13694 8452
rect 14093 8449 14105 8452
rect 14139 8449 14151 8483
rect 15120 8480 15148 8588
rect 15470 8576 15476 8588
rect 15528 8576 15534 8628
rect 18230 8616 18236 8628
rect 15571 8588 18236 8616
rect 15286 8508 15292 8560
rect 15344 8548 15350 8560
rect 15571 8548 15599 8588
rect 18230 8576 18236 8588
rect 18288 8576 18294 8628
rect 18874 8616 18880 8628
rect 18835 8588 18880 8616
rect 18874 8576 18880 8588
rect 18932 8576 18938 8628
rect 19150 8616 19156 8628
rect 18984 8588 19156 8616
rect 15344 8520 15599 8548
rect 17681 8551 17739 8557
rect 15344 8508 15350 8520
rect 17681 8517 17693 8551
rect 17727 8548 17739 8551
rect 18138 8548 18144 8560
rect 17727 8520 18144 8548
rect 17727 8517 17739 8520
rect 17681 8511 17739 8517
rect 18138 8508 18144 8520
rect 18196 8508 18202 8560
rect 18785 8551 18843 8557
rect 18340 8520 18736 8548
rect 15120 8452 15424 8480
rect 14093 8443 14151 8449
rect 8435 8384 10088 8412
rect 10137 8415 10195 8421
rect 8435 8381 8447 8384
rect 8389 8375 8447 8381
rect 10137 8381 10149 8415
rect 10183 8412 10195 8415
rect 10410 8412 10416 8424
rect 10183 8384 10416 8412
rect 10183 8381 10195 8384
rect 10137 8375 10195 8381
rect 10410 8372 10416 8384
rect 10468 8372 10474 8424
rect 10594 8372 10600 8424
rect 10652 8412 10658 8424
rect 10689 8415 10747 8421
rect 10689 8412 10701 8415
rect 10652 8384 10701 8412
rect 10652 8372 10658 8384
rect 10689 8381 10701 8384
rect 10735 8381 10747 8415
rect 10689 8375 10747 8381
rect 10888 8384 11192 8412
rect 7650 8344 7656 8356
rect 6656 8316 7656 8344
rect 7650 8304 7656 8316
rect 7708 8304 7714 8356
rect 7837 8347 7895 8353
rect 7837 8313 7849 8347
rect 7883 8344 7895 8347
rect 8656 8347 8714 8353
rect 7883 8316 8616 8344
rect 7883 8313 7895 8316
rect 7837 8307 7895 8313
rect 5077 8279 5135 8285
rect 5077 8245 5089 8279
rect 5123 8276 5135 8279
rect 5258 8276 5264 8288
rect 5123 8248 5264 8276
rect 5123 8245 5135 8248
rect 5077 8239 5135 8245
rect 5258 8236 5264 8248
rect 5316 8236 5322 8288
rect 6089 8279 6147 8285
rect 6089 8245 6101 8279
rect 6135 8276 6147 8279
rect 7006 8276 7012 8288
rect 6135 8248 7012 8276
rect 6135 8245 6147 8248
rect 6089 8239 6147 8245
rect 7006 8236 7012 8248
rect 7064 8236 7070 8288
rect 7745 8279 7803 8285
rect 7745 8245 7757 8279
rect 7791 8276 7803 8279
rect 8202 8276 8208 8288
rect 7791 8248 8208 8276
rect 7791 8245 7803 8248
rect 7745 8239 7803 8245
rect 8202 8236 8208 8248
rect 8260 8236 8266 8288
rect 8588 8276 8616 8316
rect 8656 8313 8668 8347
rect 8702 8344 8714 8347
rect 10888 8344 10916 8384
rect 10962 8353 10968 8356
rect 8702 8316 10916 8344
rect 8702 8313 8714 8316
rect 8656 8307 8714 8313
rect 10956 8307 10968 8353
rect 11020 8344 11026 8356
rect 11164 8344 11192 8384
rect 11238 8372 11244 8424
rect 11296 8412 11302 8424
rect 15286 8412 15292 8424
rect 11296 8384 15292 8412
rect 11296 8372 11302 8384
rect 15286 8372 15292 8384
rect 15344 8372 15350 8424
rect 15396 8412 15424 8452
rect 15470 8440 15476 8492
rect 15528 8480 15534 8492
rect 15841 8483 15899 8489
rect 15841 8480 15853 8483
rect 15528 8452 15853 8480
rect 15528 8440 15534 8452
rect 15841 8449 15853 8452
rect 15887 8480 15899 8483
rect 16114 8480 16120 8492
rect 15887 8452 16120 8480
rect 15887 8449 15899 8452
rect 15841 8443 15899 8449
rect 16114 8440 16120 8452
rect 16172 8440 16178 8492
rect 16304 8483 16362 8489
rect 16304 8449 16316 8483
rect 16350 8480 16362 8483
rect 16482 8480 16488 8492
rect 16350 8452 16488 8480
rect 16350 8449 16362 8452
rect 16304 8443 16362 8449
rect 16482 8440 16488 8452
rect 16540 8440 16546 8492
rect 16574 8440 16580 8492
rect 16632 8480 16638 8492
rect 18340 8480 18368 8520
rect 16632 8452 16677 8480
rect 16767 8452 18368 8480
rect 16632 8440 16638 8452
rect 16767 8412 16795 8452
rect 18414 8440 18420 8492
rect 18472 8480 18478 8492
rect 18708 8480 18736 8520
rect 18785 8517 18797 8551
rect 18831 8548 18843 8551
rect 18984 8548 19012 8588
rect 19150 8576 19156 8588
rect 19208 8576 19214 8628
rect 19242 8576 19248 8628
rect 19300 8616 19306 8628
rect 19705 8619 19763 8625
rect 19705 8616 19717 8619
rect 19300 8588 19717 8616
rect 19300 8576 19306 8588
rect 19705 8585 19717 8588
rect 19751 8585 19763 8619
rect 19705 8579 19763 8585
rect 22646 8576 22652 8628
rect 22704 8616 22710 8628
rect 22922 8616 22928 8628
rect 22704 8588 22928 8616
rect 22704 8576 22710 8588
rect 22922 8576 22928 8588
rect 22980 8576 22986 8628
rect 19886 8548 19892 8560
rect 18831 8520 19012 8548
rect 19056 8520 19892 8548
rect 18831 8517 18843 8520
rect 18785 8511 18843 8517
rect 19056 8480 19084 8520
rect 19886 8508 19892 8520
rect 19944 8508 19950 8560
rect 18472 8452 18517 8480
rect 18708 8452 19084 8480
rect 18472 8440 18478 8452
rect 19150 8440 19156 8492
rect 19208 8480 19214 8492
rect 19337 8483 19395 8489
rect 19337 8480 19349 8483
rect 19208 8452 19349 8480
rect 19208 8440 19214 8452
rect 19337 8449 19349 8452
rect 19383 8449 19395 8483
rect 19337 8443 19395 8449
rect 19426 8440 19432 8492
rect 19484 8480 19490 8492
rect 19702 8480 19708 8492
rect 19484 8452 19529 8480
rect 19615 8452 19708 8480
rect 19484 8440 19490 8452
rect 19702 8440 19708 8452
rect 19760 8480 19766 8492
rect 20212 8483 20270 8489
rect 20212 8480 20224 8483
rect 19760 8452 20224 8480
rect 19760 8440 19766 8452
rect 20212 8449 20224 8452
rect 20258 8449 20270 8483
rect 20212 8443 20270 8449
rect 20346 8440 20352 8492
rect 20404 8480 20410 8492
rect 20622 8480 20628 8492
rect 20404 8452 20449 8480
rect 20583 8452 20628 8480
rect 20404 8440 20410 8452
rect 20622 8440 20628 8452
rect 20680 8440 20686 8492
rect 22278 8440 22284 8492
rect 22336 8480 22342 8492
rect 22465 8483 22523 8489
rect 22465 8480 22477 8483
rect 22336 8452 22477 8480
rect 22336 8440 22342 8452
rect 22465 8449 22477 8452
rect 22511 8449 22523 8483
rect 22646 8480 22652 8492
rect 22607 8452 22652 8480
rect 22465 8443 22523 8449
rect 22646 8440 22652 8452
rect 22704 8440 22710 8492
rect 15396 8384 16795 8412
rect 17218 8372 17224 8424
rect 17276 8412 17282 8424
rect 17862 8412 17868 8424
rect 17276 8384 17868 8412
rect 17276 8372 17282 8384
rect 17862 8372 17868 8384
rect 17920 8372 17926 8424
rect 18141 8415 18199 8421
rect 18141 8412 18153 8415
rect 17972 8384 18153 8412
rect 11020 8316 11056 8344
rect 11164 8316 12480 8344
rect 10962 8304 10968 8307
rect 11020 8304 11026 8316
rect 9582 8276 9588 8288
rect 8588 8248 9588 8276
rect 9582 8236 9588 8248
rect 9640 8236 9646 8288
rect 9769 8279 9827 8285
rect 9769 8245 9781 8279
rect 9815 8276 9827 8279
rect 10134 8276 10140 8288
rect 9815 8248 10140 8276
rect 9815 8245 9827 8248
rect 9769 8239 9827 8245
rect 10134 8236 10140 8248
rect 10192 8236 10198 8288
rect 10597 8279 10655 8285
rect 10597 8245 10609 8279
rect 10643 8276 10655 8279
rect 12342 8276 12348 8288
rect 10643 8248 12348 8276
rect 10643 8245 10655 8248
rect 10597 8239 10655 8245
rect 12342 8236 12348 8248
rect 12400 8236 12406 8288
rect 12452 8276 12480 8316
rect 12526 8304 12532 8356
rect 12584 8344 12590 8356
rect 12682 8347 12740 8353
rect 12682 8344 12694 8347
rect 12584 8316 12694 8344
rect 12584 8304 12590 8316
rect 12682 8313 12694 8316
rect 12728 8313 12740 8347
rect 12682 8307 12740 8313
rect 14360 8347 14418 8353
rect 14360 8313 14372 8347
rect 14406 8344 14418 8347
rect 15746 8344 15752 8356
rect 14406 8316 15752 8344
rect 14406 8313 14418 8316
rect 14360 8307 14418 8313
rect 15746 8304 15752 8316
rect 15804 8304 15810 8356
rect 15838 8304 15844 8356
rect 15896 8304 15902 8356
rect 13446 8276 13452 8288
rect 12452 8248 13452 8276
rect 13446 8236 13452 8248
rect 13504 8236 13510 8288
rect 15102 8236 15108 8288
rect 15160 8276 15166 8288
rect 15856 8276 15884 8304
rect 15160 8248 15884 8276
rect 15160 8236 15166 8248
rect 16298 8236 16304 8288
rect 16356 8285 16362 8288
rect 16356 8276 16365 8285
rect 17310 8276 17316 8288
rect 16356 8248 17316 8276
rect 16356 8239 16365 8248
rect 16356 8236 16362 8239
rect 17310 8236 17316 8248
rect 17368 8236 17374 8288
rect 17862 8236 17868 8288
rect 17920 8276 17926 8288
rect 17972 8276 18000 8384
rect 18141 8381 18153 8384
rect 18187 8381 18199 8415
rect 18141 8375 18199 8381
rect 18230 8372 18236 8424
rect 18288 8412 18294 8424
rect 18785 8415 18843 8421
rect 18785 8412 18797 8415
rect 18288 8384 18797 8412
rect 18288 8372 18294 8384
rect 18785 8381 18797 8384
rect 18831 8381 18843 8415
rect 18785 8375 18843 8381
rect 19794 8372 19800 8424
rect 19852 8412 19858 8424
rect 19889 8415 19947 8421
rect 19889 8412 19901 8415
rect 19852 8384 19901 8412
rect 19852 8372 19858 8384
rect 19889 8381 19901 8384
rect 19935 8381 19947 8415
rect 19889 8375 19947 8381
rect 18874 8344 18880 8356
rect 18156 8316 18880 8344
rect 18156 8288 18184 8316
rect 18874 8304 18880 8316
rect 18932 8304 18938 8356
rect 22373 8347 22431 8353
rect 22373 8313 22385 8347
rect 22419 8344 22431 8347
rect 22554 8344 22560 8356
rect 22419 8316 22560 8344
rect 22419 8313 22431 8316
rect 22373 8307 22431 8313
rect 22554 8304 22560 8316
rect 22612 8304 22618 8356
rect 17920 8248 18000 8276
rect 17920 8236 17926 8248
rect 18138 8236 18144 8288
rect 18196 8236 18202 8288
rect 18414 8236 18420 8288
rect 18472 8276 18478 8288
rect 19245 8279 19303 8285
rect 19245 8276 19257 8279
rect 18472 8248 19257 8276
rect 18472 8236 18478 8248
rect 19245 8245 19257 8248
rect 19291 8245 19303 8279
rect 21726 8276 21732 8288
rect 21687 8248 21732 8276
rect 19245 8239 19303 8245
rect 21726 8236 21732 8248
rect 21784 8236 21790 8288
rect 22005 8279 22063 8285
rect 22005 8245 22017 8279
rect 22051 8276 22063 8279
rect 22922 8276 22928 8288
rect 22051 8248 22928 8276
rect 22051 8245 22063 8248
rect 22005 8239 22063 8245
rect 22922 8236 22928 8248
rect 22980 8236 22986 8288
rect 1104 8186 23276 8208
rect 1104 8134 8379 8186
rect 8431 8134 8443 8186
rect 8495 8134 8507 8186
rect 8559 8134 8571 8186
rect 8623 8134 15776 8186
rect 15828 8134 15840 8186
rect 15892 8134 15904 8186
rect 15956 8134 15968 8186
rect 16020 8134 23276 8186
rect 1104 8112 23276 8134
rect 4617 8075 4675 8081
rect 4617 8041 4629 8075
rect 4663 8072 4675 8075
rect 4982 8072 4988 8084
rect 4663 8044 4988 8072
rect 4663 8041 4675 8044
rect 4617 8035 4675 8041
rect 4982 8032 4988 8044
rect 5040 8032 5046 8084
rect 5074 8032 5080 8084
rect 5132 8072 5138 8084
rect 5537 8075 5595 8081
rect 5132 8044 5177 8072
rect 5132 8032 5138 8044
rect 5537 8041 5549 8075
rect 5583 8072 5595 8075
rect 5997 8075 6055 8081
rect 5997 8072 6009 8075
rect 5583 8044 6009 8072
rect 5583 8041 5595 8044
rect 5537 8035 5595 8041
rect 5997 8041 6009 8044
rect 6043 8072 6055 8075
rect 6730 8072 6736 8084
rect 6043 8044 6736 8072
rect 6043 8041 6055 8044
rect 5997 8035 6055 8041
rect 6730 8032 6736 8044
rect 6788 8032 6794 8084
rect 7837 8075 7895 8081
rect 7837 8041 7849 8075
rect 7883 8072 7895 8075
rect 9493 8075 9551 8081
rect 9493 8072 9505 8075
rect 7883 8044 9505 8072
rect 7883 8041 7895 8044
rect 7837 8035 7895 8041
rect 9493 8041 9505 8044
rect 9539 8041 9551 8075
rect 9493 8035 9551 8041
rect 9582 8032 9588 8084
rect 9640 8072 9646 8084
rect 9677 8075 9735 8081
rect 9677 8072 9689 8075
rect 9640 8044 9689 8072
rect 9640 8032 9646 8044
rect 9677 8041 9689 8044
rect 9723 8041 9735 8075
rect 12526 8072 12532 8084
rect 9677 8035 9735 8041
rect 10152 8044 12204 8072
rect 12487 8044 12532 8072
rect 1762 7964 1768 8016
rect 1820 8004 1826 8016
rect 6089 8007 6147 8013
rect 1820 7976 5028 8004
rect 1820 7964 1826 7976
rect 4338 7896 4344 7948
rect 4396 7936 4402 7948
rect 4893 7939 4951 7945
rect 4893 7936 4905 7939
rect 4396 7908 4905 7936
rect 4396 7896 4402 7908
rect 4893 7905 4905 7908
rect 4939 7905 4951 7939
rect 5000 7936 5028 7976
rect 6089 7973 6101 8007
rect 6135 8004 6147 8007
rect 7282 8004 7288 8016
rect 6135 7976 7288 8004
rect 6135 7973 6147 7976
rect 6089 7967 6147 7973
rect 7282 7964 7288 7976
rect 7340 7964 7346 8016
rect 10152 8004 10180 8044
rect 10962 8004 10968 8016
rect 7392 7976 10180 8004
rect 10244 7976 10968 8004
rect 6822 7936 6828 7948
rect 5000 7908 6828 7936
rect 4893 7899 4951 7905
rect 6822 7896 6828 7908
rect 6880 7896 6886 7948
rect 6273 7871 6331 7877
rect 6273 7837 6285 7871
rect 6319 7868 6331 7871
rect 7392 7868 7420 7976
rect 7469 7939 7527 7945
rect 7469 7905 7481 7939
rect 7515 7936 7527 7939
rect 7837 7939 7895 7945
rect 7837 7936 7849 7939
rect 7515 7908 7849 7936
rect 7515 7905 7527 7908
rect 7469 7899 7527 7905
rect 7837 7905 7849 7908
rect 7883 7905 7895 7939
rect 7837 7899 7895 7905
rect 8196 7939 8254 7945
rect 8196 7905 8208 7939
rect 8242 7936 8254 7939
rect 9950 7936 9956 7948
rect 8242 7908 9956 7936
rect 8242 7905 8254 7908
rect 8196 7899 8254 7905
rect 9950 7896 9956 7908
rect 10008 7936 10014 7948
rect 10045 7939 10103 7945
rect 10045 7936 10057 7939
rect 10008 7908 10057 7936
rect 10008 7896 10014 7908
rect 10045 7905 10057 7908
rect 10091 7905 10103 7939
rect 10045 7899 10103 7905
rect 7926 7868 7932 7880
rect 6319 7840 7420 7868
rect 7887 7840 7932 7868
rect 6319 7837 6331 7840
rect 6273 7831 6331 7837
rect 7926 7828 7932 7840
rect 7984 7828 7990 7880
rect 9493 7871 9551 7877
rect 9493 7837 9505 7871
rect 9539 7868 9551 7871
rect 9858 7868 9864 7880
rect 9539 7840 9864 7868
rect 9539 7837 9551 7840
rect 9493 7831 9551 7837
rect 9858 7828 9864 7840
rect 9916 7828 9922 7880
rect 10134 7868 10140 7880
rect 10095 7840 10140 7868
rect 10134 7828 10140 7840
rect 10192 7828 10198 7880
rect 10244 7877 10272 7976
rect 10962 7964 10968 7976
rect 11020 7964 11026 8016
rect 11416 8007 11474 8013
rect 11416 7973 11428 8007
rect 11462 8004 11474 8007
rect 11790 8004 11796 8016
rect 11462 7976 11796 8004
rect 11462 7973 11474 7976
rect 11416 7967 11474 7973
rect 11790 7964 11796 7976
rect 11848 7964 11854 8016
rect 12176 8004 12204 8044
rect 12526 8032 12532 8044
rect 12584 8072 12590 8084
rect 13265 8075 13323 8081
rect 13265 8072 13277 8075
rect 12584 8044 13277 8072
rect 12584 8032 12590 8044
rect 13265 8041 13277 8044
rect 13311 8041 13323 8075
rect 13265 8035 13323 8041
rect 13354 8032 13360 8084
rect 13412 8072 13418 8084
rect 14185 8075 14243 8081
rect 14185 8072 14197 8075
rect 13412 8044 14197 8072
rect 13412 8032 13418 8044
rect 14185 8041 14197 8044
rect 14231 8041 14243 8075
rect 14185 8035 14243 8041
rect 14366 8032 14372 8084
rect 14424 8072 14430 8084
rect 14826 8072 14832 8084
rect 14424 8044 14832 8072
rect 14424 8032 14430 8044
rect 14826 8032 14832 8044
rect 14884 8032 14890 8084
rect 15378 8032 15384 8084
rect 15436 8072 15442 8084
rect 15755 8075 15813 8081
rect 15755 8072 15767 8075
rect 15436 8044 15767 8072
rect 15436 8032 15442 8044
rect 15755 8041 15767 8044
rect 15801 8072 15813 8075
rect 16298 8072 16304 8084
rect 15801 8044 16304 8072
rect 15801 8041 15813 8044
rect 15755 8035 15813 8041
rect 16298 8032 16304 8044
rect 16356 8032 16362 8084
rect 16482 8032 16488 8084
rect 16540 8072 16546 8084
rect 17129 8075 17187 8081
rect 17129 8072 17141 8075
rect 16540 8044 17141 8072
rect 16540 8032 16546 8044
rect 17129 8041 17141 8044
rect 17175 8041 17187 8075
rect 17129 8035 17187 8041
rect 17957 8075 18015 8081
rect 17957 8041 17969 8075
rect 18003 8072 18015 8075
rect 20441 8075 20499 8081
rect 18003 8044 20024 8072
rect 18003 8041 18015 8044
rect 17957 8035 18015 8041
rect 12986 8004 12992 8016
rect 12176 7976 12992 8004
rect 12986 7964 12992 7976
rect 13044 7964 13050 8016
rect 14277 8007 14335 8013
rect 14277 8004 14289 8007
rect 13096 7976 14289 8004
rect 10318 7896 10324 7948
rect 10376 7936 10382 7948
rect 10594 7936 10600 7948
rect 10376 7908 10600 7936
rect 10376 7896 10382 7908
rect 10594 7896 10600 7908
rect 10652 7936 10658 7948
rect 11149 7939 11207 7945
rect 11149 7936 11161 7939
rect 10652 7908 11161 7936
rect 10652 7896 10658 7908
rect 11149 7905 11161 7908
rect 11195 7905 11207 7939
rect 11149 7899 11207 7905
rect 11698 7896 11704 7948
rect 11756 7936 11762 7948
rect 13096 7936 13124 7976
rect 14277 7973 14289 7976
rect 14323 7973 14335 8007
rect 14277 7967 14335 7973
rect 17310 7964 17316 8016
rect 17368 8004 17374 8016
rect 17368 7976 18716 8004
rect 17368 7964 17374 7976
rect 11756 7908 13124 7936
rect 13173 7939 13231 7945
rect 11756 7896 11762 7908
rect 13173 7905 13185 7939
rect 13219 7936 13231 7939
rect 13446 7936 13452 7948
rect 13219 7908 13452 7936
rect 13219 7905 13231 7908
rect 13173 7899 13231 7905
rect 13446 7896 13452 7908
rect 13504 7896 13510 7948
rect 13814 7896 13820 7948
rect 13872 7936 13878 7948
rect 15010 7936 15016 7948
rect 13872 7908 14872 7936
rect 14971 7908 15016 7936
rect 13872 7896 13878 7908
rect 10229 7871 10287 7877
rect 10229 7837 10241 7871
rect 10275 7837 10287 7871
rect 10229 7831 10287 7837
rect 10689 7871 10747 7877
rect 10689 7837 10701 7871
rect 10735 7837 10747 7871
rect 10689 7831 10747 7837
rect 5626 7800 5632 7812
rect 5587 7772 5632 7800
rect 5626 7760 5632 7772
rect 5684 7760 5690 7812
rect 8956 7772 9628 7800
rect 8294 7692 8300 7744
rect 8352 7732 8358 7744
rect 8956 7732 8984 7772
rect 8352 7704 8984 7732
rect 8352 7692 8358 7704
rect 9030 7692 9036 7744
rect 9088 7732 9094 7744
rect 9309 7735 9367 7741
rect 9309 7732 9321 7735
rect 9088 7704 9321 7732
rect 9088 7692 9094 7704
rect 9309 7701 9321 7704
rect 9355 7701 9367 7735
rect 9600 7732 9628 7772
rect 9674 7760 9680 7812
rect 9732 7800 9738 7812
rect 10244 7800 10272 7831
rect 9732 7772 10272 7800
rect 9732 7760 9738 7772
rect 10318 7732 10324 7744
rect 9600 7704 10324 7732
rect 9309 7695 9367 7701
rect 10318 7692 10324 7704
rect 10376 7692 10382 7744
rect 10704 7732 10732 7831
rect 12342 7828 12348 7880
rect 12400 7868 12406 7880
rect 13357 7871 13415 7877
rect 12400 7840 13308 7868
rect 12400 7828 12406 7840
rect 12158 7760 12164 7812
rect 12216 7800 12222 7812
rect 12216 7772 12572 7800
rect 12216 7760 12222 7772
rect 12434 7732 12440 7744
rect 10704 7704 12440 7732
rect 12434 7692 12440 7704
rect 12492 7692 12498 7744
rect 12544 7732 12572 7772
rect 12618 7760 12624 7812
rect 12676 7800 12682 7812
rect 12805 7803 12863 7809
rect 12805 7800 12817 7803
rect 12676 7772 12817 7800
rect 12676 7760 12682 7772
rect 12805 7769 12817 7772
rect 12851 7769 12863 7803
rect 13280 7800 13308 7840
rect 13357 7837 13369 7871
rect 13403 7868 13415 7871
rect 13538 7868 13544 7880
rect 13403 7840 13544 7868
rect 13403 7837 13415 7840
rect 13357 7831 13415 7837
rect 13538 7828 13544 7840
rect 13596 7828 13602 7880
rect 14369 7871 14427 7877
rect 14369 7837 14381 7871
rect 14415 7837 14427 7871
rect 14844 7868 14872 7908
rect 15010 7896 15016 7908
rect 15068 7896 15074 7948
rect 15286 7936 15292 7948
rect 15247 7908 15292 7936
rect 15286 7896 15292 7908
rect 15344 7896 15350 7948
rect 16025 7939 16083 7945
rect 16025 7936 16037 7939
rect 15396 7908 16037 7936
rect 15396 7868 15424 7908
rect 16025 7905 16037 7908
rect 16071 7936 16083 7939
rect 17954 7936 17960 7948
rect 16071 7908 17960 7936
rect 16071 7905 16083 7908
rect 16025 7899 16083 7905
rect 17954 7896 17960 7908
rect 18012 7896 18018 7948
rect 18049 7939 18107 7945
rect 18049 7905 18061 7939
rect 18095 7936 18107 7939
rect 18138 7936 18144 7948
rect 18095 7908 18144 7936
rect 18095 7905 18107 7908
rect 18049 7899 18107 7905
rect 18138 7896 18144 7908
rect 18196 7896 18202 7948
rect 18506 7896 18512 7948
rect 18564 7936 18570 7948
rect 18601 7939 18659 7945
rect 18601 7936 18613 7939
rect 18564 7908 18613 7936
rect 18564 7896 18570 7908
rect 18601 7905 18613 7908
rect 18647 7905 18659 7939
rect 18688 7936 18716 7976
rect 18874 7936 18880 7948
rect 18688 7908 18880 7936
rect 18601 7899 18659 7905
rect 18874 7896 18880 7908
rect 18932 7945 18938 7948
rect 18932 7939 18982 7945
rect 18932 7905 18936 7939
rect 18970 7905 18982 7939
rect 18932 7899 18982 7905
rect 19337 7939 19395 7945
rect 19337 7905 19349 7939
rect 19383 7936 19395 7939
rect 19996 7936 20024 8044
rect 20441 8041 20453 8075
rect 20487 8072 20499 8075
rect 20622 8072 20628 8084
rect 20487 8044 20628 8072
rect 20487 8041 20499 8044
rect 20441 8035 20499 8041
rect 20622 8032 20628 8044
rect 20680 8032 20686 8084
rect 21536 8007 21594 8013
rect 21536 7973 21548 8007
rect 21582 8004 21594 8007
rect 22462 8004 22468 8016
rect 21582 7976 22468 8004
rect 21582 7973 21594 7976
rect 21536 7967 21594 7973
rect 22462 7964 22468 7976
rect 22520 7964 22526 8016
rect 20070 7936 20076 7948
rect 19383 7908 20076 7936
rect 19383 7905 19395 7908
rect 19337 7899 19395 7905
rect 18932 7896 18938 7899
rect 20070 7896 20076 7908
rect 20128 7896 20134 7948
rect 20898 7896 20904 7948
rect 20956 7936 20962 7948
rect 21269 7939 21327 7945
rect 21269 7936 21281 7939
rect 20956 7908 21281 7936
rect 20956 7896 20962 7908
rect 21269 7905 21281 7908
rect 21315 7905 21327 7939
rect 21269 7899 21327 7905
rect 14844 7840 15424 7868
rect 14369 7831 14427 7837
rect 13998 7800 14004 7812
rect 13280 7772 14004 7800
rect 12805 7763 12863 7769
rect 13998 7760 14004 7772
rect 14056 7800 14062 7812
rect 14384 7800 14412 7831
rect 15746 7828 15752 7880
rect 15804 7868 15810 7880
rect 15804 7840 15849 7868
rect 15804 7828 15810 7840
rect 16114 7828 16120 7880
rect 16172 7868 16178 7880
rect 18233 7871 18291 7877
rect 16172 7840 18184 7868
rect 16172 7828 16178 7840
rect 14056 7772 14412 7800
rect 14056 7760 14062 7772
rect 16666 7760 16672 7812
rect 16724 7800 16730 7812
rect 17678 7800 17684 7812
rect 16724 7772 17684 7800
rect 16724 7760 16730 7772
rect 17678 7760 17684 7772
rect 17736 7760 17742 7812
rect 18156 7800 18184 7840
rect 18233 7837 18245 7871
rect 18279 7868 18291 7871
rect 18322 7868 18328 7880
rect 18279 7840 18328 7868
rect 18279 7837 18291 7840
rect 18233 7831 18291 7837
rect 18322 7828 18328 7840
rect 18380 7828 18386 7880
rect 19107 7871 19165 7877
rect 19107 7837 19119 7871
rect 19153 7868 19165 7871
rect 19518 7868 19524 7880
rect 19153 7840 19524 7868
rect 19153 7837 19165 7840
rect 19107 7831 19165 7837
rect 19518 7828 19524 7840
rect 19576 7828 19582 7880
rect 20714 7828 20720 7880
rect 20772 7868 20778 7880
rect 20990 7868 20996 7880
rect 20772 7840 20996 7868
rect 20772 7828 20778 7840
rect 20990 7828 20996 7840
rect 21048 7828 21054 7880
rect 18506 7800 18512 7812
rect 18156 7772 18512 7800
rect 18506 7760 18512 7772
rect 18564 7760 18570 7812
rect 21174 7800 21180 7812
rect 20916 7772 21180 7800
rect 13170 7732 13176 7744
rect 12544 7704 13176 7732
rect 13170 7692 13176 7704
rect 13228 7692 13234 7744
rect 13817 7735 13875 7741
rect 13817 7701 13829 7735
rect 13863 7732 13875 7735
rect 14458 7732 14464 7744
rect 13863 7704 14464 7732
rect 13863 7701 13875 7704
rect 13817 7695 13875 7701
rect 14458 7692 14464 7704
rect 14516 7692 14522 7744
rect 14550 7692 14556 7744
rect 14608 7732 14614 7744
rect 16942 7732 16948 7744
rect 14608 7704 16948 7732
rect 14608 7692 14614 7704
rect 16942 7692 16948 7704
rect 17000 7692 17006 7744
rect 17589 7735 17647 7741
rect 17589 7701 17601 7735
rect 17635 7732 17647 7735
rect 18782 7732 18788 7744
rect 17635 7704 18788 7732
rect 17635 7701 17647 7704
rect 17589 7695 17647 7701
rect 18782 7692 18788 7704
rect 18840 7692 18846 7744
rect 18874 7692 18880 7744
rect 18932 7732 18938 7744
rect 20916 7732 20944 7772
rect 21174 7760 21180 7772
rect 21232 7760 21238 7812
rect 18932 7704 20944 7732
rect 18932 7692 18938 7704
rect 22370 7692 22376 7744
rect 22428 7732 22434 7744
rect 22649 7735 22707 7741
rect 22649 7732 22661 7735
rect 22428 7704 22661 7732
rect 22428 7692 22434 7704
rect 22649 7701 22661 7704
rect 22695 7701 22707 7735
rect 22649 7695 22707 7701
rect 1104 7642 23276 7664
rect 1104 7590 4680 7642
rect 4732 7590 4744 7642
rect 4796 7590 4808 7642
rect 4860 7590 4872 7642
rect 4924 7590 12078 7642
rect 12130 7590 12142 7642
rect 12194 7590 12206 7642
rect 12258 7590 12270 7642
rect 12322 7590 19475 7642
rect 19527 7590 19539 7642
rect 19591 7590 19603 7642
rect 19655 7590 19667 7642
rect 19719 7590 23276 7642
rect 1104 7568 23276 7590
rect 5442 7488 5448 7540
rect 5500 7528 5506 7540
rect 6365 7531 6423 7537
rect 6365 7528 6377 7531
rect 5500 7500 6377 7528
rect 5500 7488 5506 7500
rect 6365 7497 6377 7500
rect 6411 7497 6423 7531
rect 6365 7491 6423 7497
rect 7193 7531 7251 7537
rect 7193 7497 7205 7531
rect 7239 7528 7251 7531
rect 7374 7528 7380 7540
rect 7239 7500 7380 7528
rect 7239 7497 7251 7500
rect 7193 7491 7251 7497
rect 7374 7488 7380 7500
rect 7432 7488 7438 7540
rect 7561 7531 7619 7537
rect 7561 7497 7573 7531
rect 7607 7528 7619 7531
rect 8294 7528 8300 7540
rect 7607 7500 8300 7528
rect 7607 7497 7619 7500
rect 7561 7491 7619 7497
rect 8294 7488 8300 7500
rect 8352 7488 8358 7540
rect 9950 7528 9956 7540
rect 8588 7500 9812 7528
rect 9911 7500 9956 7528
rect 8588 7460 8616 7500
rect 7024 7432 8616 7460
rect 9784 7460 9812 7500
rect 9950 7488 9956 7500
rect 10008 7488 10014 7540
rect 11974 7528 11980 7540
rect 10244 7500 11980 7528
rect 10244 7460 10272 7500
rect 11974 7488 11980 7500
rect 12032 7488 12038 7540
rect 15654 7528 15660 7540
rect 13648 7500 15516 7528
rect 15615 7500 15660 7528
rect 9784 7432 10272 7460
rect 5534 7284 5540 7336
rect 5592 7324 5598 7336
rect 5629 7327 5687 7333
rect 5629 7324 5641 7327
rect 5592 7296 5641 7324
rect 5592 7284 5598 7296
rect 5629 7293 5641 7296
rect 5675 7293 5687 7327
rect 5629 7287 5687 7293
rect 6181 7327 6239 7333
rect 6181 7293 6193 7327
rect 6227 7324 6239 7327
rect 6914 7324 6920 7336
rect 6227 7296 6920 7324
rect 6227 7293 6239 7296
rect 6181 7287 6239 7293
rect 6914 7284 6920 7296
rect 6972 7284 6978 7336
rect 7024 7333 7052 7432
rect 11882 7420 11888 7472
rect 11940 7420 11946 7472
rect 7377 7395 7435 7401
rect 7377 7361 7389 7395
rect 7423 7392 7435 7395
rect 8110 7392 8116 7404
rect 7423 7364 8116 7392
rect 7423 7361 7435 7364
rect 7377 7355 7435 7361
rect 8110 7352 8116 7364
rect 8168 7352 8174 7404
rect 9674 7352 9680 7404
rect 9732 7392 9738 7404
rect 10226 7392 10232 7404
rect 9732 7364 10232 7392
rect 9732 7352 9738 7364
rect 10226 7352 10232 7364
rect 10284 7352 10290 7404
rect 11238 7352 11244 7404
rect 11296 7392 11302 7404
rect 11900 7392 11928 7420
rect 12989 7395 13047 7401
rect 12989 7392 13001 7395
rect 11296 7364 13001 7392
rect 11296 7352 11302 7364
rect 12989 7361 13001 7364
rect 13035 7361 13047 7395
rect 12989 7355 13047 7361
rect 7009 7327 7067 7333
rect 7009 7293 7021 7327
rect 7055 7293 7067 7327
rect 7009 7287 7067 7293
rect 7926 7284 7932 7336
rect 7984 7324 7990 7336
rect 8573 7327 8631 7333
rect 8573 7324 8585 7327
rect 7984 7296 8585 7324
rect 7984 7284 7990 7296
rect 8573 7293 8585 7296
rect 8619 7293 8631 7327
rect 8573 7287 8631 7293
rect 8840 7327 8898 7333
rect 8840 7293 8852 7327
rect 8886 7324 8898 7327
rect 10134 7324 10140 7336
rect 8886 7296 10140 7324
rect 8886 7293 8898 7296
rect 8840 7287 8898 7293
rect 6362 7216 6368 7268
rect 6420 7256 6426 7268
rect 8021 7259 8079 7265
rect 8021 7256 8033 7259
rect 6420 7228 8033 7256
rect 6420 7216 6426 7228
rect 8021 7225 8033 7228
rect 8067 7225 8079 7259
rect 8588 7256 8616 7287
rect 10134 7284 10140 7296
rect 10192 7284 10198 7336
rect 10318 7284 10324 7336
rect 10376 7324 10382 7336
rect 11790 7324 11796 7336
rect 10376 7296 11796 7324
rect 10376 7284 10382 7296
rect 11790 7284 11796 7296
rect 11848 7284 11854 7336
rect 11885 7327 11943 7333
rect 11885 7293 11897 7327
rect 11931 7324 11943 7327
rect 13354 7324 13360 7336
rect 11931 7296 13360 7324
rect 11931 7293 11943 7296
rect 11885 7287 11943 7293
rect 13354 7284 13360 7296
rect 13412 7284 13418 7336
rect 13648 7333 13676 7500
rect 14274 7460 14280 7472
rect 13740 7432 14280 7460
rect 13740 7333 13768 7432
rect 14274 7420 14280 7432
rect 14332 7420 14338 7472
rect 15488 7460 15516 7500
rect 15654 7488 15660 7500
rect 15712 7488 15718 7540
rect 16316 7500 17540 7528
rect 16316 7460 16344 7500
rect 15488 7432 16344 7460
rect 17512 7460 17540 7500
rect 17586 7488 17592 7540
rect 17644 7528 17650 7540
rect 17681 7531 17739 7537
rect 17681 7528 17693 7531
rect 17644 7500 17693 7528
rect 17644 7488 17650 7500
rect 17681 7497 17693 7500
rect 17727 7497 17739 7531
rect 17681 7491 17739 7497
rect 18322 7488 18328 7540
rect 18380 7528 18386 7540
rect 20165 7531 20223 7537
rect 20165 7528 20177 7531
rect 18380 7500 20177 7528
rect 18380 7488 18386 7500
rect 20165 7497 20177 7500
rect 20211 7497 20223 7531
rect 20165 7491 20223 7497
rect 22462 7488 22468 7540
rect 22520 7528 22526 7540
rect 22557 7531 22615 7537
rect 22557 7528 22569 7531
rect 22520 7500 22569 7528
rect 22520 7488 22526 7500
rect 22557 7497 22569 7500
rect 22603 7497 22615 7531
rect 22557 7491 22615 7497
rect 18046 7460 18052 7472
rect 17512 7432 18052 7460
rect 18046 7420 18052 7432
rect 18104 7420 18110 7472
rect 18417 7463 18475 7469
rect 18417 7429 18429 7463
rect 18463 7429 18475 7463
rect 18417 7423 18475 7429
rect 18432 7392 18460 7423
rect 19886 7420 19892 7472
rect 19944 7460 19950 7472
rect 20898 7460 20904 7472
rect 19944 7432 20904 7460
rect 19944 7420 19950 7432
rect 18432 7364 18920 7392
rect 13633 7327 13691 7333
rect 13633 7293 13645 7327
rect 13679 7293 13691 7327
rect 13633 7287 13691 7293
rect 13725 7327 13783 7333
rect 13725 7293 13737 7327
rect 13771 7293 13783 7327
rect 14274 7324 14280 7336
rect 14235 7296 14280 7324
rect 13725 7287 13783 7293
rect 14274 7284 14280 7296
rect 14332 7284 14338 7336
rect 14826 7284 14832 7336
rect 14884 7324 14890 7336
rect 16117 7327 16175 7333
rect 16117 7324 16129 7327
rect 14884 7296 16129 7324
rect 14884 7284 14890 7296
rect 16117 7293 16129 7296
rect 16163 7293 16175 7327
rect 16117 7287 16175 7293
rect 16209 7327 16267 7333
rect 16209 7293 16221 7327
rect 16255 7324 16267 7327
rect 16301 7327 16359 7333
rect 16301 7324 16313 7327
rect 16255 7296 16313 7324
rect 16255 7293 16267 7296
rect 16209 7287 16267 7293
rect 16301 7293 16313 7296
rect 16347 7293 16359 7327
rect 18138 7324 18144 7336
rect 16301 7287 16359 7293
rect 16500 7296 18144 7324
rect 8754 7256 8760 7268
rect 8588 7228 8760 7256
rect 8021 7219 8079 7225
rect 8754 7216 8760 7228
rect 8812 7216 8818 7268
rect 9030 7216 9036 7268
rect 9088 7256 9094 7268
rect 10474 7259 10532 7265
rect 10474 7256 10486 7259
rect 9088 7228 10486 7256
rect 9088 7216 9094 7228
rect 10474 7225 10486 7228
rect 10520 7225 10532 7259
rect 10474 7219 10532 7225
rect 12250 7216 12256 7268
rect 12308 7256 12314 7268
rect 12897 7259 12955 7265
rect 12897 7256 12909 7259
rect 12308 7228 12909 7256
rect 12308 7216 12314 7228
rect 12897 7225 12909 7228
rect 12943 7225 12955 7259
rect 12897 7219 12955 7225
rect 14544 7259 14602 7265
rect 14544 7225 14556 7259
rect 14590 7256 14602 7259
rect 15286 7256 15292 7268
rect 14590 7228 15292 7256
rect 14590 7225 14602 7228
rect 14544 7219 14602 7225
rect 15286 7216 15292 7228
rect 15344 7216 15350 7268
rect 16500 7256 16528 7296
rect 18138 7284 18144 7296
rect 18196 7284 18202 7336
rect 18233 7327 18291 7333
rect 18233 7293 18245 7327
rect 18279 7293 18291 7327
rect 18233 7287 18291 7293
rect 15856 7228 16528 7256
rect 16568 7259 16626 7265
rect 5813 7191 5871 7197
rect 5813 7157 5825 7191
rect 5859 7188 5871 7191
rect 6270 7188 6276 7200
rect 5859 7160 6276 7188
rect 5859 7157 5871 7160
rect 5813 7151 5871 7157
rect 6270 7148 6276 7160
rect 6328 7188 6334 7200
rect 7377 7191 7435 7197
rect 7377 7188 7389 7191
rect 6328 7160 7389 7188
rect 6328 7148 6334 7160
rect 7377 7157 7389 7160
rect 7423 7157 7435 7191
rect 7377 7151 7435 7157
rect 7929 7191 7987 7197
rect 7929 7157 7941 7191
rect 7975 7188 7987 7191
rect 8846 7188 8852 7200
rect 7975 7160 8852 7188
rect 7975 7157 7987 7160
rect 7929 7151 7987 7157
rect 8846 7148 8852 7160
rect 8904 7148 8910 7200
rect 8938 7148 8944 7200
rect 8996 7188 9002 7200
rect 11609 7191 11667 7197
rect 11609 7188 11621 7191
rect 8996 7160 11621 7188
rect 8996 7148 9002 7160
rect 11609 7157 11621 7160
rect 11655 7157 11667 7191
rect 11609 7151 11667 7157
rect 12434 7148 12440 7200
rect 12492 7188 12498 7200
rect 12802 7188 12808 7200
rect 12492 7160 12537 7188
rect 12763 7160 12808 7188
rect 12492 7148 12498 7160
rect 12802 7148 12808 7160
rect 12860 7148 12866 7200
rect 13449 7191 13507 7197
rect 13449 7157 13461 7191
rect 13495 7188 13507 7191
rect 13814 7188 13820 7200
rect 13495 7160 13820 7188
rect 13495 7157 13507 7160
rect 13449 7151 13507 7157
rect 13814 7148 13820 7160
rect 13872 7148 13878 7200
rect 13909 7191 13967 7197
rect 13909 7157 13921 7191
rect 13955 7188 13967 7191
rect 15856 7188 15884 7228
rect 16568 7225 16580 7259
rect 16614 7256 16626 7259
rect 17494 7256 17500 7268
rect 16614 7228 17500 7256
rect 16614 7225 16626 7228
rect 16568 7219 16626 7225
rect 17494 7216 17500 7228
rect 17552 7216 17558 7268
rect 18248 7256 18276 7287
rect 18598 7284 18604 7336
rect 18656 7324 18662 7336
rect 18785 7327 18843 7333
rect 18785 7324 18797 7327
rect 18656 7296 18797 7324
rect 18656 7284 18662 7296
rect 18785 7293 18797 7296
rect 18831 7293 18843 7327
rect 18892 7324 18920 7364
rect 20346 7324 20352 7336
rect 18892 7296 20352 7324
rect 18785 7287 18843 7293
rect 20346 7284 20352 7296
rect 20404 7284 20410 7336
rect 20456 7333 20484 7432
rect 20898 7420 20904 7432
rect 20956 7420 20962 7472
rect 20530 7352 20536 7404
rect 20588 7392 20594 7404
rect 20717 7395 20775 7401
rect 20717 7392 20729 7395
rect 20588 7364 20729 7392
rect 20588 7352 20594 7364
rect 20717 7361 20729 7364
rect 20763 7361 20775 7395
rect 20717 7355 20775 7361
rect 20441 7327 20499 7333
rect 20441 7293 20453 7327
rect 20487 7293 20499 7327
rect 20441 7287 20499 7293
rect 20898 7284 20904 7336
rect 20956 7324 20962 7336
rect 21177 7327 21235 7333
rect 21177 7324 21189 7327
rect 20956 7296 21189 7324
rect 20956 7284 20962 7296
rect 21177 7293 21189 7296
rect 21223 7293 21235 7327
rect 21177 7287 21235 7293
rect 21444 7327 21502 7333
rect 21444 7293 21456 7327
rect 21490 7324 21502 7327
rect 22646 7324 22652 7336
rect 21490 7296 22652 7324
rect 21490 7293 21502 7296
rect 21444 7287 21502 7293
rect 22646 7284 22652 7296
rect 22704 7284 22710 7336
rect 19052 7259 19110 7265
rect 18248 7228 19012 7256
rect 13955 7160 15884 7188
rect 15933 7191 15991 7197
rect 13955 7157 13967 7160
rect 13909 7151 13967 7157
rect 15933 7157 15945 7191
rect 15979 7188 15991 7191
rect 16114 7188 16120 7200
rect 15979 7160 16120 7188
rect 15979 7157 15991 7160
rect 15933 7151 15991 7157
rect 16114 7148 16120 7160
rect 16172 7188 16178 7200
rect 16209 7191 16267 7197
rect 16209 7188 16221 7191
rect 16172 7160 16221 7188
rect 16172 7148 16178 7160
rect 16209 7157 16221 7160
rect 16255 7157 16267 7191
rect 18984 7188 19012 7228
rect 19052 7225 19064 7259
rect 19098 7256 19110 7259
rect 21542 7256 21548 7268
rect 19098 7228 21548 7256
rect 19098 7225 19110 7228
rect 19052 7219 19110 7225
rect 21542 7216 21548 7228
rect 21600 7256 21606 7268
rect 22370 7256 22376 7268
rect 21600 7228 22376 7256
rect 21600 7216 21606 7228
rect 22370 7216 22376 7228
rect 22428 7216 22434 7268
rect 19334 7188 19340 7200
rect 18984 7160 19340 7188
rect 16209 7151 16267 7157
rect 19334 7148 19340 7160
rect 19392 7148 19398 7200
rect 19794 7148 19800 7200
rect 19852 7188 19858 7200
rect 21818 7188 21824 7200
rect 19852 7160 21824 7188
rect 19852 7148 19858 7160
rect 21818 7148 21824 7160
rect 21876 7148 21882 7200
rect 1104 7098 23276 7120
rect 1104 7046 8379 7098
rect 8431 7046 8443 7098
rect 8495 7046 8507 7098
rect 8559 7046 8571 7098
rect 8623 7046 15776 7098
rect 15828 7046 15840 7098
rect 15892 7046 15904 7098
rect 15956 7046 15968 7098
rect 16020 7046 23276 7098
rect 1104 7024 23276 7046
rect 7469 6987 7527 6993
rect 7469 6953 7481 6987
rect 7515 6984 7527 6987
rect 7558 6984 7564 6996
rect 7515 6956 7564 6984
rect 7515 6953 7527 6956
rect 7469 6947 7527 6953
rect 7558 6944 7564 6956
rect 7616 6944 7622 6996
rect 9582 6944 9588 6996
rect 9640 6984 9646 6996
rect 13262 6984 13268 6996
rect 9640 6956 13268 6984
rect 9640 6944 9646 6956
rect 13262 6944 13268 6956
rect 13320 6944 13326 6996
rect 13725 6987 13783 6993
rect 13725 6984 13737 6987
rect 13372 6956 13737 6984
rect 6454 6848 6460 6860
rect 6415 6820 6460 6848
rect 6454 6808 6460 6820
rect 6512 6808 6518 6860
rect 6825 6851 6883 6857
rect 6825 6817 6837 6851
rect 6871 6817 6883 6851
rect 7576 6848 7604 6944
rect 9030 6916 9036 6928
rect 8991 6888 9036 6916
rect 9030 6876 9036 6888
rect 9088 6876 9094 6928
rect 10962 6876 10968 6928
rect 11020 6916 11026 6928
rect 12710 6916 12716 6928
rect 11020 6888 11836 6916
rect 12671 6888 12716 6916
rect 11020 6876 11026 6888
rect 7929 6851 7987 6857
rect 7929 6848 7941 6851
rect 7576 6820 7941 6848
rect 6825 6811 6883 6817
rect 7929 6817 7941 6820
rect 7975 6817 7987 6851
rect 7929 6811 7987 6817
rect 8021 6851 8079 6857
rect 8021 6817 8033 6851
rect 8067 6848 8079 6851
rect 8938 6848 8944 6860
rect 8067 6820 8800 6848
rect 8899 6820 8944 6848
rect 8067 6817 8079 6820
rect 8021 6811 8079 6817
rect 3694 6740 3700 6792
rect 3752 6780 3758 6792
rect 6840 6780 6868 6811
rect 3752 6752 6868 6780
rect 8205 6783 8263 6789
rect 3752 6740 3758 6752
rect 8205 6749 8217 6783
rect 8251 6780 8263 6783
rect 8294 6780 8300 6792
rect 8251 6752 8300 6780
rect 8251 6749 8263 6752
rect 8205 6743 8263 6749
rect 8294 6740 8300 6752
rect 8352 6740 8358 6792
rect 8772 6780 8800 6820
rect 8938 6808 8944 6820
rect 8996 6808 9002 6860
rect 9766 6848 9772 6860
rect 9048 6820 9772 6848
rect 9048 6780 9076 6820
rect 9766 6808 9772 6820
rect 9824 6808 9830 6860
rect 9950 6857 9956 6860
rect 9944 6811 9956 6857
rect 10008 6848 10014 6860
rect 10008 6820 10044 6848
rect 9950 6808 9956 6811
rect 10008 6808 10014 6820
rect 11606 6808 11612 6860
rect 11664 6848 11670 6860
rect 11701 6851 11759 6857
rect 11701 6848 11713 6851
rect 11664 6820 11713 6848
rect 11664 6808 11670 6820
rect 11701 6817 11713 6820
rect 11747 6817 11759 6851
rect 11808 6848 11836 6888
rect 12710 6876 12716 6888
rect 12768 6876 12774 6928
rect 12894 6876 12900 6928
rect 12952 6916 12958 6928
rect 13372 6916 13400 6956
rect 13725 6953 13737 6956
rect 13771 6953 13783 6987
rect 13725 6947 13783 6953
rect 16942 6944 16948 6996
rect 17000 6984 17006 6996
rect 19153 6987 19211 6993
rect 17000 6956 17540 6984
rect 17000 6944 17006 6956
rect 12952 6888 13400 6916
rect 12952 6876 12958 6888
rect 13814 6876 13820 6928
rect 13872 6916 13878 6928
rect 16298 6916 16304 6928
rect 13872 6888 16304 6916
rect 13872 6876 13878 6888
rect 16298 6876 16304 6888
rect 16356 6916 16362 6928
rect 16356 6888 16620 6916
rect 16356 6876 16362 6888
rect 13538 6848 13544 6860
rect 11808 6820 13544 6848
rect 11701 6811 11759 6817
rect 8772 6752 9076 6780
rect 9217 6783 9275 6789
rect 9217 6749 9229 6783
rect 9263 6780 9275 6783
rect 9490 6780 9496 6792
rect 9263 6752 9496 6780
rect 9263 6749 9275 6752
rect 9217 6743 9275 6749
rect 9490 6740 9496 6752
rect 9548 6740 9554 6792
rect 9674 6780 9680 6792
rect 9635 6752 9680 6780
rect 9674 6740 9680 6752
rect 9732 6740 9738 6792
rect 10686 6740 10692 6792
rect 10744 6780 10750 6792
rect 11054 6780 11060 6792
rect 10744 6752 11060 6780
rect 10744 6740 10750 6752
rect 11054 6740 11060 6752
rect 11112 6740 11118 6792
rect 11146 6740 11152 6792
rect 11204 6780 11210 6792
rect 11900 6789 11928 6820
rect 11793 6783 11851 6789
rect 11793 6780 11805 6783
rect 11204 6752 11805 6780
rect 11204 6740 11210 6752
rect 11793 6749 11805 6752
rect 11839 6749 11851 6783
rect 11793 6743 11851 6749
rect 11885 6783 11943 6789
rect 11885 6749 11897 6783
rect 11931 6749 11943 6783
rect 11885 6743 11943 6749
rect 11992 6752 12388 6780
rect 7558 6712 7564 6724
rect 7519 6684 7564 6712
rect 7558 6672 7564 6684
rect 7616 6672 7622 6724
rect 8478 6712 8484 6724
rect 8128 6684 8484 6712
rect 5350 6604 5356 6656
rect 5408 6644 5414 6656
rect 6638 6644 6644 6656
rect 5408 6616 6644 6644
rect 5408 6604 5414 6616
rect 6638 6604 6644 6616
rect 6696 6604 6702 6656
rect 7009 6647 7067 6653
rect 7009 6613 7021 6647
rect 7055 6644 7067 6647
rect 8128 6644 8156 6684
rect 8478 6672 8484 6684
rect 8536 6672 8542 6724
rect 8573 6715 8631 6721
rect 8573 6681 8585 6715
rect 8619 6712 8631 6715
rect 8662 6712 8668 6724
rect 8619 6684 8668 6712
rect 8619 6681 8631 6684
rect 8573 6675 8631 6681
rect 8662 6672 8668 6684
rect 8720 6672 8726 6724
rect 8754 6672 8760 6724
rect 8812 6712 8818 6724
rect 9692 6712 9720 6740
rect 11992 6712 12020 6752
rect 8812 6684 9720 6712
rect 10888 6684 12020 6712
rect 8812 6672 8818 6684
rect 7055 6616 8156 6644
rect 7055 6613 7067 6616
rect 7009 6607 7067 6613
rect 8202 6604 8208 6656
rect 8260 6644 8266 6656
rect 10888 6644 10916 6684
rect 12250 6672 12256 6724
rect 12308 6672 12314 6724
rect 12360 6712 12388 6752
rect 12618 6740 12624 6792
rect 12676 6780 12682 6792
rect 13004 6789 13032 6820
rect 13538 6808 13544 6820
rect 13596 6808 13602 6860
rect 14185 6851 14243 6857
rect 14185 6817 14197 6851
rect 14231 6848 14243 6851
rect 14369 6851 14427 6857
rect 14369 6848 14381 6851
rect 14231 6820 14381 6848
rect 14231 6817 14243 6820
rect 14185 6811 14243 6817
rect 14369 6817 14381 6820
rect 14415 6817 14427 6851
rect 14550 6848 14556 6860
rect 14511 6820 14556 6848
rect 14369 6811 14427 6817
rect 14550 6808 14556 6820
rect 14608 6808 14614 6860
rect 15562 6857 15568 6860
rect 15556 6848 15568 6857
rect 15523 6820 15568 6848
rect 15556 6811 15568 6820
rect 15562 6808 15568 6811
rect 15620 6808 15626 6860
rect 12805 6783 12863 6789
rect 12805 6780 12817 6783
rect 12676 6752 12817 6780
rect 12676 6740 12682 6752
rect 12805 6749 12817 6752
rect 12851 6749 12863 6783
rect 12805 6743 12863 6749
rect 12989 6783 13047 6789
rect 12989 6749 13001 6783
rect 13035 6749 13047 6783
rect 12989 6743 13047 6749
rect 13078 6740 13084 6792
rect 13136 6780 13142 6792
rect 13817 6783 13875 6789
rect 13817 6780 13829 6783
rect 13136 6752 13829 6780
rect 13136 6740 13142 6752
rect 13817 6749 13829 6752
rect 13863 6749 13875 6783
rect 13998 6780 14004 6792
rect 13959 6752 14004 6780
rect 13817 6743 13875 6749
rect 13998 6740 14004 6752
rect 14056 6740 14062 6792
rect 15010 6740 15016 6792
rect 15068 6780 15074 6792
rect 15289 6783 15347 6789
rect 15289 6780 15301 6783
rect 15068 6752 15301 6780
rect 15068 6740 15074 6752
rect 15289 6749 15301 6752
rect 15335 6749 15347 6783
rect 16592 6780 16620 6888
rect 16666 6876 16672 6928
rect 16724 6916 16730 6928
rect 17402 6916 17408 6928
rect 16724 6888 17408 6916
rect 16724 6876 16730 6888
rect 17402 6876 17408 6888
rect 17460 6876 17466 6928
rect 17512 6916 17540 6956
rect 19153 6953 19165 6987
rect 19199 6984 19211 6987
rect 19334 6984 19340 6996
rect 19199 6956 19340 6984
rect 19199 6953 19211 6956
rect 19153 6947 19211 6953
rect 19334 6944 19340 6956
rect 19392 6984 19398 6996
rect 19797 6987 19855 6993
rect 19797 6984 19809 6987
rect 19392 6956 19809 6984
rect 19392 6944 19398 6956
rect 19797 6953 19809 6956
rect 19843 6953 19855 6987
rect 19797 6947 19855 6953
rect 22281 6987 22339 6993
rect 22281 6953 22293 6987
rect 22327 6984 22339 6987
rect 22646 6984 22652 6996
rect 22327 6956 22652 6984
rect 22327 6953 22339 6956
rect 22281 6947 22339 6953
rect 22646 6944 22652 6956
rect 22704 6944 22710 6996
rect 20254 6916 20260 6928
rect 17512 6888 20260 6916
rect 20254 6876 20260 6888
rect 20312 6876 20318 6928
rect 16758 6808 16764 6860
rect 16816 6848 16822 6860
rect 17201 6851 17259 6857
rect 17201 6848 17213 6851
rect 16816 6820 17213 6848
rect 16816 6808 16822 6820
rect 17201 6817 17213 6820
rect 17247 6817 17259 6851
rect 17201 6811 17259 6817
rect 17494 6808 17500 6860
rect 17552 6848 17558 6860
rect 20162 6848 20168 6860
rect 17552 6820 19380 6848
rect 20123 6820 20168 6848
rect 17552 6808 17558 6820
rect 16945 6783 17003 6789
rect 16945 6780 16957 6783
rect 16592 6752 16957 6780
rect 15289 6743 15347 6749
rect 16945 6749 16957 6752
rect 16991 6749 17003 6783
rect 16945 6743 17003 6749
rect 18598 6740 18604 6792
rect 18656 6780 18662 6792
rect 19352 6789 19380 6820
rect 20162 6808 20168 6820
rect 20220 6808 20226 6860
rect 21168 6851 21226 6857
rect 21168 6817 21180 6851
rect 21214 6848 21226 6851
rect 21450 6848 21456 6860
rect 21214 6820 21456 6848
rect 21214 6817 21226 6820
rect 21168 6811 21226 6817
rect 21450 6808 21456 6820
rect 21508 6808 21514 6860
rect 22554 6848 22560 6860
rect 22515 6820 22560 6848
rect 22554 6808 22560 6820
rect 22612 6808 22618 6860
rect 23382 6848 23388 6860
rect 23343 6820 23388 6848
rect 23382 6808 23388 6820
rect 23440 6808 23446 6860
rect 19245 6783 19303 6789
rect 19245 6780 19257 6783
rect 18656 6752 19257 6780
rect 18656 6740 18662 6752
rect 19245 6749 19257 6752
rect 19291 6749 19303 6783
rect 19245 6743 19303 6749
rect 19337 6783 19395 6789
rect 19337 6749 19349 6783
rect 19383 6749 19395 6783
rect 20254 6780 20260 6792
rect 20215 6752 20260 6780
rect 19337 6743 19395 6749
rect 20254 6740 20260 6752
rect 20312 6740 20318 6792
rect 20349 6783 20407 6789
rect 20349 6749 20361 6783
rect 20395 6749 20407 6783
rect 20898 6780 20904 6792
rect 20859 6752 20904 6780
rect 20349 6743 20407 6749
rect 14737 6715 14795 6721
rect 14737 6712 14749 6715
rect 12360 6684 14749 6712
rect 14737 6681 14749 6684
rect 14783 6681 14795 6715
rect 14737 6675 14795 6681
rect 16669 6715 16727 6721
rect 16669 6681 16681 6715
rect 16715 6712 16727 6715
rect 16758 6712 16764 6724
rect 16715 6684 16764 6712
rect 16715 6681 16727 6684
rect 16669 6675 16727 6681
rect 16758 6672 16764 6684
rect 16816 6672 16822 6724
rect 17954 6672 17960 6724
rect 18012 6712 18018 6724
rect 18012 6684 19012 6712
rect 18012 6672 18018 6684
rect 11054 6644 11060 6656
rect 8260 6616 10916 6644
rect 11015 6616 11060 6644
rect 8260 6604 8266 6616
rect 11054 6604 11060 6616
rect 11112 6604 11118 6656
rect 11330 6644 11336 6656
rect 11291 6616 11336 6644
rect 11330 6604 11336 6616
rect 11388 6604 11394 6656
rect 12268 6644 12296 6672
rect 12345 6647 12403 6653
rect 12345 6644 12357 6647
rect 12268 6616 12357 6644
rect 12345 6613 12357 6616
rect 12391 6613 12403 6647
rect 13354 6644 13360 6656
rect 13315 6616 13360 6644
rect 12345 6607 12403 6613
rect 13354 6604 13360 6616
rect 13412 6644 13418 6656
rect 14090 6644 14096 6656
rect 13412 6616 14096 6644
rect 13412 6604 13418 6616
rect 14090 6604 14096 6616
rect 14148 6604 14154 6656
rect 14185 6647 14243 6653
rect 14185 6613 14197 6647
rect 14231 6644 14243 6647
rect 17126 6644 17132 6656
rect 14231 6616 17132 6644
rect 14231 6613 14243 6616
rect 14185 6607 14243 6613
rect 17126 6604 17132 6616
rect 17184 6604 17190 6656
rect 17586 6604 17592 6656
rect 17644 6644 17650 6656
rect 18325 6647 18383 6653
rect 18325 6644 18337 6647
rect 17644 6616 18337 6644
rect 17644 6604 17650 6616
rect 18325 6613 18337 6616
rect 18371 6613 18383 6647
rect 18782 6644 18788 6656
rect 18743 6616 18788 6644
rect 18325 6607 18383 6613
rect 18782 6604 18788 6616
rect 18840 6604 18846 6656
rect 18984 6644 19012 6684
rect 19058 6672 19064 6724
rect 19116 6712 19122 6724
rect 20364 6712 20392 6743
rect 20898 6740 20904 6752
rect 20956 6740 20962 6792
rect 19116 6684 20392 6712
rect 19116 6672 19122 6684
rect 20714 6644 20720 6656
rect 18984 6616 20720 6644
rect 20714 6604 20720 6616
rect 20772 6604 20778 6656
rect 1104 6554 23276 6576
rect 1104 6502 4680 6554
rect 4732 6502 4744 6554
rect 4796 6502 4808 6554
rect 4860 6502 4872 6554
rect 4924 6502 12078 6554
rect 12130 6502 12142 6554
rect 12194 6502 12206 6554
rect 12258 6502 12270 6554
rect 12322 6502 19475 6554
rect 19527 6502 19539 6554
rect 19591 6502 19603 6554
rect 19655 6502 19667 6554
rect 19719 6502 23276 6554
rect 1104 6480 23276 6502
rect 7098 6400 7104 6452
rect 7156 6440 7162 6452
rect 7837 6443 7895 6449
rect 7837 6440 7849 6443
rect 7156 6412 7849 6440
rect 7156 6400 7162 6412
rect 7837 6409 7849 6412
rect 7883 6409 7895 6443
rect 7837 6403 7895 6409
rect 8294 6400 8300 6452
rect 8352 6440 8358 6452
rect 8352 6412 9720 6440
rect 8352 6400 8358 6412
rect 8389 6375 8447 6381
rect 8389 6341 8401 6375
rect 8435 6372 8447 6375
rect 8662 6372 8668 6384
rect 8435 6344 8668 6372
rect 8435 6341 8447 6344
rect 8389 6335 8447 6341
rect 8662 6332 8668 6344
rect 8720 6332 8726 6384
rect 9692 6372 9720 6412
rect 9950 6400 9956 6452
rect 10008 6440 10014 6452
rect 10137 6443 10195 6449
rect 10137 6440 10149 6443
rect 10008 6412 10149 6440
rect 10008 6400 10014 6412
rect 10137 6409 10149 6412
rect 10183 6440 10195 6443
rect 10183 6412 10824 6440
rect 10183 6409 10195 6412
rect 10137 6403 10195 6409
rect 10594 6372 10600 6384
rect 9692 6344 10600 6372
rect 10594 6332 10600 6344
rect 10652 6332 10658 6384
rect 8754 6304 8760 6316
rect 8715 6276 8760 6304
rect 8754 6264 8760 6276
rect 8812 6264 8818 6316
rect 10796 6304 10824 6412
rect 10870 6400 10876 6452
rect 10928 6440 10934 6452
rect 14277 6443 14335 6449
rect 10928 6412 14228 6440
rect 10928 6400 10934 6412
rect 10873 6307 10931 6313
rect 10873 6304 10885 6307
rect 10796 6276 10885 6304
rect 10873 6273 10885 6276
rect 10919 6273 10931 6307
rect 10873 6267 10931 6273
rect 10962 6264 10968 6316
rect 11020 6304 11026 6316
rect 11020 6276 11065 6304
rect 11020 6264 11026 6276
rect 12342 6264 12348 6316
rect 12400 6304 12406 6316
rect 12897 6307 12955 6313
rect 12897 6304 12909 6307
rect 12400 6276 12909 6304
rect 12400 6264 12406 6276
rect 12897 6273 12909 6276
rect 12943 6273 12955 6307
rect 12897 6267 12955 6273
rect 7653 6239 7711 6245
rect 7653 6205 7665 6239
rect 7699 6205 7711 6239
rect 8202 6236 8208 6248
rect 8163 6208 8208 6236
rect 7653 6199 7711 6205
rect 7668 6168 7696 6199
rect 8202 6196 8208 6208
rect 8260 6196 8266 6248
rect 10410 6236 10416 6248
rect 8864 6208 10416 6236
rect 8864 6168 8892 6208
rect 10410 6196 10416 6208
rect 10468 6196 10474 6248
rect 10781 6239 10839 6245
rect 10781 6205 10793 6239
rect 10827 6236 10839 6239
rect 11054 6236 11060 6248
rect 10827 6208 11060 6236
rect 10827 6205 10839 6208
rect 10781 6199 10839 6205
rect 11054 6196 11060 6208
rect 11112 6196 11118 6248
rect 11514 6196 11520 6248
rect 11572 6236 11578 6248
rect 11609 6239 11667 6245
rect 11609 6236 11621 6239
rect 11572 6208 11621 6236
rect 11572 6196 11578 6208
rect 11609 6205 11621 6208
rect 11655 6205 11667 6239
rect 11609 6199 11667 6205
rect 11793 6239 11851 6245
rect 11793 6205 11805 6239
rect 11839 6236 11851 6239
rect 12250 6236 12256 6248
rect 11839 6208 12256 6236
rect 11839 6205 11851 6208
rect 11793 6199 11851 6205
rect 12250 6196 12256 6208
rect 12308 6196 12314 6248
rect 12437 6239 12495 6245
rect 12437 6205 12449 6239
rect 12483 6236 12495 6239
rect 12483 6208 13860 6236
rect 12483 6205 12495 6208
rect 12437 6199 12495 6205
rect 13832 6180 13860 6208
rect 7668 6140 8892 6168
rect 8938 6128 8944 6180
rect 8996 6177 9002 6180
rect 8996 6171 9060 6177
rect 8996 6137 9014 6171
rect 9048 6137 9060 6171
rect 8996 6131 9060 6137
rect 13164 6171 13222 6177
rect 13164 6137 13176 6171
rect 13210 6168 13222 6171
rect 13354 6168 13360 6180
rect 13210 6140 13360 6168
rect 13210 6137 13222 6140
rect 13164 6131 13222 6137
rect 8996 6128 9002 6131
rect 13354 6128 13360 6140
rect 13412 6168 13418 6180
rect 13722 6168 13728 6180
rect 13412 6140 13728 6168
rect 13412 6128 13418 6140
rect 13722 6128 13728 6140
rect 13780 6128 13786 6180
rect 13814 6128 13820 6180
rect 13872 6128 13878 6180
rect 14200 6168 14228 6412
rect 14277 6409 14289 6443
rect 14323 6440 14335 6443
rect 14550 6440 14556 6452
rect 14323 6412 14556 6440
rect 14323 6409 14335 6412
rect 14277 6403 14335 6409
rect 14550 6400 14556 6412
rect 14608 6400 14614 6452
rect 15286 6400 15292 6452
rect 15344 6440 15350 6452
rect 15654 6440 15660 6452
rect 15344 6412 15660 6440
rect 15344 6400 15350 6412
rect 15654 6400 15660 6412
rect 15712 6440 15718 6452
rect 15933 6443 15991 6449
rect 15933 6440 15945 6443
rect 15712 6412 15945 6440
rect 15712 6400 15718 6412
rect 15933 6409 15945 6412
rect 15979 6409 15991 6443
rect 15933 6403 15991 6409
rect 16945 6443 17003 6449
rect 16945 6409 16957 6443
rect 16991 6440 17003 6443
rect 18230 6440 18236 6452
rect 16991 6412 18236 6440
rect 16991 6409 17003 6412
rect 16945 6403 17003 6409
rect 18230 6400 18236 6412
rect 18288 6400 18294 6452
rect 20438 6440 20444 6452
rect 18616 6412 20444 6440
rect 14568 6304 14596 6400
rect 18616 6372 18644 6412
rect 20438 6400 20444 6412
rect 20496 6400 20502 6452
rect 20901 6443 20959 6449
rect 20901 6409 20913 6443
rect 20947 6440 20959 6443
rect 21450 6440 21456 6452
rect 20947 6412 21456 6440
rect 20947 6409 20959 6412
rect 20901 6403 20959 6409
rect 21450 6400 21456 6412
rect 21508 6400 21514 6452
rect 15580 6344 18644 6372
rect 14568 6276 14688 6304
rect 14366 6196 14372 6248
rect 14424 6236 14430 6248
rect 14553 6239 14611 6245
rect 14553 6236 14565 6239
rect 14424 6208 14565 6236
rect 14424 6196 14430 6208
rect 14553 6205 14565 6208
rect 14599 6205 14611 6239
rect 14660 6236 14688 6276
rect 14809 6239 14867 6245
rect 14809 6236 14821 6239
rect 14660 6208 14821 6236
rect 14553 6199 14611 6205
rect 14809 6205 14821 6208
rect 14855 6205 14867 6239
rect 14809 6199 14867 6205
rect 15580 6168 15608 6344
rect 18690 6332 18696 6384
rect 18748 6372 18754 6384
rect 18748 6344 19564 6372
rect 18748 6332 18754 6344
rect 17402 6304 17408 6316
rect 14200 6140 15608 6168
rect 15856 6276 17408 6304
rect 10410 6100 10416 6112
rect 10371 6072 10416 6100
rect 10410 6060 10416 6072
rect 10468 6060 10474 6112
rect 11238 6060 11244 6112
rect 11296 6100 11302 6112
rect 11425 6103 11483 6109
rect 11425 6100 11437 6103
rect 11296 6072 11437 6100
rect 11296 6060 11302 6072
rect 11425 6069 11437 6072
rect 11471 6069 11483 6103
rect 11425 6063 11483 6069
rect 11977 6103 12035 6109
rect 11977 6069 11989 6103
rect 12023 6100 12035 6103
rect 15856 6100 15884 6276
rect 17402 6264 17408 6276
rect 17460 6264 17466 6316
rect 17589 6307 17647 6313
rect 17589 6273 17601 6307
rect 17635 6304 17647 6307
rect 17635 6276 18092 6304
rect 17635 6273 17647 6276
rect 17589 6267 17647 6273
rect 16393 6239 16451 6245
rect 16393 6205 16405 6239
rect 16439 6236 16451 6239
rect 17678 6236 17684 6248
rect 16439 6208 17684 6236
rect 16439 6205 16451 6208
rect 16393 6199 16451 6205
rect 17678 6196 17684 6208
rect 17736 6196 17742 6248
rect 18064 6236 18092 6276
rect 18138 6264 18144 6316
rect 18196 6304 18202 6316
rect 19058 6304 19064 6316
rect 18196 6276 19064 6304
rect 18196 6264 18202 6276
rect 19058 6264 19064 6276
rect 19116 6264 19122 6316
rect 19536 6313 19564 6344
rect 19521 6307 19579 6313
rect 19521 6273 19533 6307
rect 19567 6273 19579 6307
rect 19521 6267 19579 6273
rect 19536 6236 19564 6267
rect 21818 6264 21824 6316
rect 21876 6304 21882 6316
rect 22097 6307 22155 6313
rect 22097 6304 22109 6307
rect 21876 6276 22109 6304
rect 21876 6264 21882 6276
rect 22097 6273 22109 6276
rect 22143 6273 22155 6307
rect 22097 6267 22155 6273
rect 20898 6236 20904 6248
rect 18064 6208 19104 6236
rect 19536 6208 20904 6236
rect 19076 6180 19104 6208
rect 20898 6196 20904 6208
rect 20956 6196 20962 6248
rect 22002 6196 22008 6248
rect 22060 6236 22066 6248
rect 22557 6239 22615 6245
rect 22557 6236 22569 6239
rect 22060 6208 22569 6236
rect 22060 6196 22066 6208
rect 22557 6205 22569 6208
rect 22603 6205 22615 6239
rect 22557 6199 22615 6205
rect 18969 6171 19027 6177
rect 18969 6168 18981 6171
rect 16592 6140 18981 6168
rect 16592 6109 16620 6140
rect 18969 6137 18981 6140
rect 19015 6137 19027 6171
rect 18969 6131 19027 6137
rect 19058 6128 19064 6180
rect 19116 6128 19122 6180
rect 19242 6128 19248 6180
rect 19300 6168 19306 6180
rect 19766 6171 19824 6177
rect 19766 6168 19778 6171
rect 19300 6140 19778 6168
rect 19300 6128 19306 6140
rect 19766 6137 19778 6140
rect 19812 6137 19824 6171
rect 21910 6168 21916 6180
rect 21871 6140 21916 6168
rect 19766 6131 19824 6137
rect 21910 6128 21916 6140
rect 21968 6128 21974 6180
rect 12023 6072 15884 6100
rect 16577 6103 16635 6109
rect 12023 6069 12035 6072
rect 11977 6063 12035 6069
rect 16577 6069 16589 6103
rect 16623 6069 16635 6103
rect 17310 6100 17316 6112
rect 17271 6072 17316 6100
rect 16577 6063 16635 6069
rect 17310 6060 17316 6072
rect 17368 6060 17374 6112
rect 17405 6103 17463 6109
rect 17405 6069 17417 6103
rect 17451 6100 17463 6103
rect 17954 6100 17960 6112
rect 17451 6072 17960 6100
rect 17451 6069 17463 6072
rect 17405 6063 17463 6069
rect 17954 6060 17960 6072
rect 18012 6060 18018 6112
rect 18049 6103 18107 6109
rect 18049 6069 18061 6103
rect 18095 6100 18107 6103
rect 18414 6100 18420 6112
rect 18095 6072 18420 6100
rect 18095 6069 18107 6072
rect 18049 6063 18107 6069
rect 18414 6060 18420 6072
rect 18472 6060 18478 6112
rect 18509 6103 18567 6109
rect 18509 6069 18521 6103
rect 18555 6100 18567 6103
rect 18598 6100 18604 6112
rect 18555 6072 18604 6100
rect 18555 6069 18567 6072
rect 18509 6063 18567 6069
rect 18598 6060 18604 6072
rect 18656 6060 18662 6112
rect 18874 6100 18880 6112
rect 18835 6072 18880 6100
rect 18874 6060 18880 6072
rect 18932 6060 18938 6112
rect 20990 6060 20996 6112
rect 21048 6100 21054 6112
rect 21545 6103 21603 6109
rect 21545 6100 21557 6103
rect 21048 6072 21557 6100
rect 21048 6060 21054 6072
rect 21545 6069 21557 6072
rect 21591 6069 21603 6103
rect 22002 6100 22008 6112
rect 21963 6072 22008 6100
rect 21545 6063 21603 6069
rect 22002 6060 22008 6072
rect 22060 6060 22066 6112
rect 1104 6010 23276 6032
rect 1104 5958 8379 6010
rect 8431 5958 8443 6010
rect 8495 5958 8507 6010
rect 8559 5958 8571 6010
rect 8623 5958 15776 6010
rect 15828 5958 15840 6010
rect 15892 5958 15904 6010
rect 15956 5958 15968 6010
rect 16020 5958 23276 6010
rect 1104 5936 23276 5958
rect 8018 5856 8024 5908
rect 8076 5896 8082 5908
rect 8113 5899 8171 5905
rect 8113 5896 8125 5899
rect 8076 5868 8125 5896
rect 8076 5856 8082 5868
rect 8113 5865 8125 5868
rect 8159 5865 8171 5899
rect 8113 5859 8171 5865
rect 9401 5899 9459 5905
rect 9401 5865 9413 5899
rect 9447 5896 9459 5899
rect 9447 5868 11836 5896
rect 9447 5865 9459 5868
rect 9401 5859 9459 5865
rect 8941 5831 8999 5837
rect 8941 5797 8953 5831
rect 8987 5828 8999 5831
rect 11808 5828 11836 5868
rect 12342 5856 12348 5908
rect 12400 5896 12406 5908
rect 12897 5899 12955 5905
rect 12897 5896 12909 5899
rect 12400 5868 12909 5896
rect 12400 5856 12406 5868
rect 12897 5865 12909 5868
rect 12943 5865 12955 5899
rect 13630 5896 13636 5908
rect 12897 5859 12955 5865
rect 13096 5868 13636 5896
rect 13096 5828 13124 5868
rect 13630 5856 13636 5868
rect 13688 5856 13694 5908
rect 13722 5856 13728 5908
rect 13780 5896 13786 5908
rect 14369 5899 14427 5905
rect 14369 5896 14381 5899
rect 13780 5868 14381 5896
rect 13780 5856 13786 5868
rect 14369 5865 14381 5868
rect 14415 5865 14427 5899
rect 17218 5896 17224 5908
rect 14369 5859 14427 5865
rect 15488 5868 17224 5896
rect 8987 5800 11744 5828
rect 11808 5800 13124 5828
rect 8987 5797 8999 5800
rect 8941 5791 8999 5797
rect 6638 5720 6644 5772
rect 6696 5760 6702 5772
rect 9766 5760 9772 5772
rect 6696 5732 9772 5760
rect 6696 5720 6702 5732
rect 9766 5720 9772 5732
rect 9824 5720 9830 5772
rect 9944 5763 10002 5769
rect 9944 5729 9956 5763
rect 9990 5760 10002 5763
rect 11054 5760 11060 5772
rect 9990 5732 11060 5760
rect 9990 5729 10002 5732
rect 9944 5723 10002 5729
rect 11054 5720 11060 5732
rect 11112 5720 11118 5772
rect 11606 5769 11612 5772
rect 11600 5760 11612 5769
rect 11567 5732 11612 5760
rect 11600 5723 11612 5732
rect 11606 5720 11612 5723
rect 11664 5720 11670 5772
rect 11716 5760 11744 5800
rect 12526 5760 12532 5772
rect 11716 5732 12532 5760
rect 12526 5720 12532 5732
rect 12584 5720 12590 5772
rect 12897 5763 12955 5769
rect 12897 5729 12909 5763
rect 12943 5760 12955 5763
rect 12989 5763 13047 5769
rect 12989 5760 13001 5763
rect 12943 5732 13001 5760
rect 12943 5729 12955 5732
rect 12897 5723 12955 5729
rect 12989 5729 13001 5732
rect 13035 5729 13047 5763
rect 12989 5723 13047 5729
rect 13256 5763 13314 5769
rect 13256 5729 13268 5763
rect 13302 5760 13314 5763
rect 13722 5760 13728 5772
rect 13302 5732 13728 5760
rect 13302 5729 13314 5732
rect 13256 5723 13314 5729
rect 13722 5720 13728 5732
rect 13780 5720 13786 5772
rect 14645 5763 14703 5769
rect 14645 5729 14657 5763
rect 14691 5760 14703 5763
rect 15488 5760 15516 5868
rect 17218 5856 17224 5868
rect 17276 5856 17282 5908
rect 17494 5896 17500 5908
rect 17407 5868 17500 5896
rect 17494 5856 17500 5868
rect 17552 5896 17558 5908
rect 18233 5899 18291 5905
rect 18233 5896 18245 5899
rect 17552 5868 18245 5896
rect 17552 5856 17558 5868
rect 18233 5865 18245 5868
rect 18279 5865 18291 5899
rect 18233 5859 18291 5865
rect 19242 5856 19248 5908
rect 19300 5896 19306 5908
rect 20165 5899 20223 5905
rect 20165 5896 20177 5899
rect 19300 5868 20177 5896
rect 19300 5856 19306 5868
rect 20165 5865 20177 5868
rect 20211 5865 20223 5899
rect 23385 5899 23443 5905
rect 23385 5896 23397 5899
rect 20165 5859 20223 5865
rect 22112 5868 23397 5896
rect 15580 5800 19840 5828
rect 15580 5769 15608 5800
rect 14691 5732 15516 5760
rect 15565 5763 15623 5769
rect 14691 5729 14703 5732
rect 14645 5723 14703 5729
rect 15565 5729 15577 5763
rect 15611 5729 15623 5763
rect 15565 5723 15623 5729
rect 16384 5763 16442 5769
rect 16384 5729 16396 5763
rect 16430 5760 16442 5763
rect 16430 5732 17172 5760
rect 16430 5729 16442 5732
rect 16384 5723 16442 5729
rect 9033 5695 9091 5701
rect 9033 5661 9045 5695
rect 9079 5661 9091 5695
rect 9033 5655 9091 5661
rect 9217 5695 9275 5701
rect 9217 5661 9229 5695
rect 9263 5692 9275 5695
rect 9401 5695 9459 5701
rect 9401 5692 9413 5695
rect 9263 5664 9413 5692
rect 9263 5661 9275 5664
rect 9217 5655 9275 5661
rect 9401 5661 9413 5664
rect 9447 5661 9459 5695
rect 9674 5692 9680 5704
rect 9635 5664 9680 5692
rect 9401 5655 9459 5661
rect 7650 5584 7656 5636
rect 7708 5624 7714 5636
rect 8573 5627 8631 5633
rect 8573 5624 8585 5627
rect 7708 5596 8585 5624
rect 7708 5584 7714 5596
rect 8573 5593 8585 5596
rect 8619 5593 8631 5627
rect 8573 5587 8631 5593
rect 9048 5556 9076 5655
rect 9674 5652 9680 5664
rect 9732 5652 9738 5704
rect 11238 5652 11244 5704
rect 11296 5692 11302 5704
rect 11333 5695 11391 5701
rect 11333 5692 11345 5695
rect 11296 5664 11345 5692
rect 11296 5652 11302 5664
rect 11333 5661 11345 5664
rect 11379 5661 11391 5695
rect 16114 5692 16120 5704
rect 16075 5664 16120 5692
rect 11333 5655 11391 5661
rect 16114 5652 16120 5664
rect 16172 5652 16178 5704
rect 17144 5692 17172 5732
rect 17678 5720 17684 5772
rect 17736 5760 17742 5772
rect 18141 5763 18199 5769
rect 18141 5760 18153 5763
rect 17736 5732 18153 5760
rect 17736 5720 17742 5732
rect 18141 5729 18153 5732
rect 18187 5729 18199 5763
rect 18141 5723 18199 5729
rect 18690 5720 18696 5772
rect 18748 5760 18754 5772
rect 19058 5769 19064 5772
rect 18785 5763 18843 5769
rect 18785 5760 18797 5763
rect 18748 5732 18797 5760
rect 18748 5720 18754 5732
rect 18785 5729 18797 5732
rect 18831 5729 18843 5763
rect 19052 5760 19064 5769
rect 19019 5732 19064 5760
rect 18785 5723 18843 5729
rect 19052 5723 19064 5732
rect 19058 5720 19064 5723
rect 19116 5720 19122 5772
rect 19812 5760 19840 5800
rect 20438 5788 20444 5840
rect 20496 5828 20502 5840
rect 22112 5828 22140 5868
rect 23385 5865 23397 5868
rect 23431 5865 23443 5899
rect 23385 5859 23443 5865
rect 22554 5828 22560 5840
rect 20496 5800 22324 5828
rect 22515 5800 22560 5828
rect 20496 5788 20502 5800
rect 20898 5760 20904 5772
rect 19812 5732 20904 5760
rect 20898 5720 20904 5732
rect 20956 5720 20962 5772
rect 21542 5720 21548 5772
rect 21600 5760 21606 5772
rect 22296 5769 22324 5800
rect 22554 5788 22560 5800
rect 22612 5788 22618 5840
rect 21637 5763 21695 5769
rect 21637 5760 21649 5763
rect 21600 5732 21649 5760
rect 21600 5720 21606 5732
rect 21637 5729 21649 5732
rect 21683 5729 21695 5763
rect 21637 5723 21695 5729
rect 22281 5763 22339 5769
rect 22281 5729 22293 5763
rect 22327 5729 22339 5763
rect 22281 5723 22339 5729
rect 17770 5692 17776 5704
rect 17144 5664 17776 5692
rect 17770 5652 17776 5664
rect 17828 5652 17834 5704
rect 18322 5692 18328 5704
rect 18283 5664 18328 5692
rect 18322 5652 18328 5664
rect 18380 5652 18386 5704
rect 21726 5692 21732 5704
rect 21687 5664 21732 5692
rect 21726 5652 21732 5664
rect 21784 5652 21790 5704
rect 21818 5652 21824 5704
rect 21876 5692 21882 5704
rect 21876 5664 21969 5692
rect 21876 5652 21882 5664
rect 11057 5627 11115 5633
rect 11057 5593 11069 5627
rect 11103 5624 11115 5627
rect 11146 5624 11152 5636
rect 11103 5596 11152 5624
rect 11103 5593 11115 5596
rect 11057 5587 11115 5593
rect 11146 5584 11152 5596
rect 11204 5584 11210 5636
rect 12618 5584 12624 5636
rect 12676 5624 12682 5636
rect 12713 5627 12771 5633
rect 12713 5624 12725 5627
rect 12676 5596 12725 5624
rect 12676 5584 12682 5596
rect 12713 5593 12725 5596
rect 12759 5593 12771 5627
rect 12713 5587 12771 5593
rect 14090 5584 14096 5636
rect 14148 5624 14154 5636
rect 14550 5624 14556 5636
rect 14148 5596 14556 5624
rect 14148 5584 14154 5596
rect 14550 5584 14556 5596
rect 14608 5584 14614 5636
rect 14829 5627 14887 5633
rect 14829 5593 14841 5627
rect 14875 5624 14887 5627
rect 16022 5624 16028 5636
rect 14875 5596 16028 5624
rect 14875 5593 14887 5596
rect 14829 5587 14887 5593
rect 16022 5584 16028 5596
rect 16080 5584 16086 5636
rect 17696 5596 18644 5624
rect 11974 5556 11980 5568
rect 9048 5528 11980 5556
rect 11974 5516 11980 5528
rect 12032 5516 12038 5568
rect 12526 5516 12532 5568
rect 12584 5556 12590 5568
rect 12897 5559 12955 5565
rect 12897 5556 12909 5559
rect 12584 5528 12909 5556
rect 12584 5516 12590 5528
rect 12897 5525 12909 5528
rect 12943 5556 12955 5559
rect 14366 5556 14372 5568
rect 12943 5528 14372 5556
rect 12943 5525 12955 5528
rect 12897 5519 12955 5525
rect 14366 5516 14372 5528
rect 14424 5516 14430 5568
rect 15749 5559 15807 5565
rect 15749 5525 15761 5559
rect 15795 5556 15807 5559
rect 17696 5556 17724 5596
rect 15795 5528 17724 5556
rect 17773 5559 17831 5565
rect 15795 5525 15807 5528
rect 15749 5519 15807 5525
rect 17773 5525 17785 5559
rect 17819 5556 17831 5559
rect 18506 5556 18512 5568
rect 17819 5528 18512 5556
rect 17819 5525 17831 5528
rect 17773 5519 17831 5525
rect 18506 5516 18512 5528
rect 18564 5516 18570 5568
rect 18616 5556 18644 5596
rect 20438 5584 20444 5636
rect 20496 5624 20502 5636
rect 21836 5624 21864 5652
rect 20496 5596 21864 5624
rect 20496 5584 20502 5596
rect 20162 5556 20168 5568
rect 18616 5528 20168 5556
rect 20162 5516 20168 5528
rect 20220 5516 20226 5568
rect 20806 5516 20812 5568
rect 20864 5556 20870 5568
rect 21269 5559 21327 5565
rect 21269 5556 21281 5559
rect 20864 5528 21281 5556
rect 20864 5516 20870 5528
rect 21269 5525 21281 5528
rect 21315 5525 21327 5559
rect 21269 5519 21327 5525
rect 1104 5466 23276 5488
rect 1104 5414 4680 5466
rect 4732 5414 4744 5466
rect 4796 5414 4808 5466
rect 4860 5414 4872 5466
rect 4924 5414 12078 5466
rect 12130 5414 12142 5466
rect 12194 5414 12206 5466
rect 12258 5414 12270 5466
rect 12322 5414 19475 5466
rect 19527 5414 19539 5466
rect 19591 5414 19603 5466
rect 19655 5414 19667 5466
rect 19719 5414 23276 5466
rect 1104 5392 23276 5414
rect 9585 5355 9643 5361
rect 9585 5321 9597 5355
rect 9631 5352 9643 5355
rect 11333 5355 11391 5361
rect 9631 5324 11008 5352
rect 9631 5321 9643 5324
rect 9585 5315 9643 5321
rect 10980 5216 11008 5324
rect 11333 5321 11345 5355
rect 11379 5352 11391 5355
rect 11606 5352 11612 5364
rect 11379 5324 11612 5352
rect 11379 5321 11391 5324
rect 11333 5315 11391 5321
rect 11606 5312 11612 5324
rect 11664 5312 11670 5364
rect 15102 5352 15108 5364
rect 15063 5324 15108 5352
rect 15102 5312 15108 5324
rect 15160 5312 15166 5364
rect 16022 5312 16028 5364
rect 16080 5352 16086 5364
rect 17678 5352 17684 5364
rect 16080 5324 17540 5352
rect 17639 5324 17684 5352
rect 16080 5312 16086 5324
rect 13722 5244 13728 5296
rect 13780 5284 13786 5296
rect 13817 5287 13875 5293
rect 13817 5284 13829 5287
rect 13780 5256 13829 5284
rect 13780 5244 13786 5256
rect 13817 5253 13829 5256
rect 13863 5253 13875 5287
rect 13817 5247 13875 5253
rect 14366 5244 14372 5296
rect 14424 5284 14430 5296
rect 14424 5256 14688 5284
rect 14424 5244 14430 5256
rect 10980 5188 12572 5216
rect 9398 5148 9404 5160
rect 9359 5120 9404 5148
rect 9398 5108 9404 5120
rect 9456 5108 9462 5160
rect 9674 5108 9680 5160
rect 9732 5148 9738 5160
rect 9953 5151 10011 5157
rect 9953 5148 9965 5151
rect 9732 5120 9965 5148
rect 9732 5108 9738 5120
rect 9953 5117 9965 5120
rect 9999 5117 10011 5151
rect 9953 5111 10011 5117
rect 10220 5151 10278 5157
rect 10220 5117 10232 5151
rect 10266 5148 10278 5151
rect 11146 5148 11152 5160
rect 10266 5120 11152 5148
rect 10266 5117 10278 5120
rect 10220 5111 10278 5117
rect 9968 5080 9996 5111
rect 11146 5108 11152 5120
rect 11204 5108 11210 5160
rect 11793 5151 11851 5157
rect 11793 5117 11805 5151
rect 11839 5148 11851 5151
rect 12250 5148 12256 5160
rect 11839 5120 12256 5148
rect 11839 5117 11851 5120
rect 11793 5111 11851 5117
rect 12250 5108 12256 5120
rect 12308 5108 12314 5160
rect 12437 5151 12495 5157
rect 12437 5117 12449 5151
rect 12483 5117 12495 5151
rect 12437 5111 12495 5117
rect 11238 5080 11244 5092
rect 9968 5052 11244 5080
rect 11238 5040 11244 5052
rect 11296 5040 11302 5092
rect 8938 5012 8944 5024
rect 8899 4984 8944 5012
rect 8938 4972 8944 4984
rect 8996 4972 9002 5024
rect 11977 5015 12035 5021
rect 11977 4981 11989 5015
rect 12023 5012 12035 5015
rect 12342 5012 12348 5024
rect 12023 4984 12348 5012
rect 12023 4981 12035 4984
rect 11977 4975 12035 4981
rect 12342 4972 12348 4984
rect 12400 4972 12406 5024
rect 12452 5012 12480 5111
rect 12544 5080 12572 5188
rect 13906 5176 13912 5228
rect 13964 5216 13970 5228
rect 14458 5216 14464 5228
rect 13964 5188 14464 5216
rect 13964 5176 13970 5188
rect 14458 5176 14464 5188
rect 14516 5216 14522 5228
rect 14660 5225 14688 5256
rect 14553 5219 14611 5225
rect 14553 5216 14565 5219
rect 14516 5188 14565 5216
rect 14516 5176 14522 5188
rect 14553 5185 14565 5188
rect 14599 5185 14611 5219
rect 14553 5179 14611 5185
rect 14645 5219 14703 5225
rect 14645 5185 14657 5219
rect 14691 5185 14703 5219
rect 15654 5216 15660 5228
rect 15615 5188 15660 5216
rect 14645 5179 14703 5185
rect 15654 5176 15660 5188
rect 15712 5176 15718 5228
rect 16298 5216 16304 5228
rect 16259 5188 16304 5216
rect 16298 5176 16304 5188
rect 16356 5176 16362 5228
rect 17512 5216 17540 5324
rect 17678 5312 17684 5324
rect 17736 5312 17742 5364
rect 18046 5352 18052 5364
rect 18007 5324 18052 5352
rect 18046 5312 18052 5324
rect 18104 5312 18110 5364
rect 18138 5312 18144 5364
rect 18196 5352 18202 5364
rect 19794 5352 19800 5364
rect 18196 5324 19800 5352
rect 18196 5312 18202 5324
rect 19794 5312 19800 5324
rect 19852 5312 19858 5364
rect 20349 5355 20407 5361
rect 20349 5321 20361 5355
rect 20395 5352 20407 5355
rect 20898 5352 20904 5364
rect 20395 5324 20904 5352
rect 20395 5321 20407 5324
rect 20349 5315 20407 5321
rect 20898 5312 20904 5324
rect 20956 5312 20962 5364
rect 17586 5244 17592 5296
rect 17644 5284 17650 5296
rect 19245 5287 19303 5293
rect 19245 5284 19257 5287
rect 17644 5256 19257 5284
rect 17644 5244 17650 5256
rect 19245 5253 19257 5256
rect 19291 5253 19303 5287
rect 19245 5247 19303 5253
rect 18322 5216 18328 5228
rect 17512 5188 18328 5216
rect 18322 5176 18328 5188
rect 18380 5176 18386 5228
rect 18506 5216 18512 5228
rect 18467 5188 18512 5216
rect 18506 5176 18512 5188
rect 18564 5176 18570 5228
rect 18601 5219 18659 5225
rect 18601 5185 18613 5219
rect 18647 5216 18659 5219
rect 19610 5216 19616 5228
rect 18647 5188 19616 5216
rect 18647 5185 18659 5188
rect 18601 5179 18659 5185
rect 12710 5157 12716 5160
rect 12704 5148 12716 5157
rect 12671 5120 12716 5148
rect 12704 5111 12716 5120
rect 12710 5108 12716 5111
rect 12768 5108 12774 5160
rect 13814 5108 13820 5160
rect 13872 5148 13878 5160
rect 16390 5148 16396 5160
rect 13872 5120 16396 5148
rect 13872 5108 13878 5120
rect 16390 5108 16396 5120
rect 16448 5108 16454 5160
rect 16568 5151 16626 5157
rect 16568 5117 16580 5151
rect 16614 5148 16626 5151
rect 17494 5148 17500 5160
rect 16614 5120 17500 5148
rect 16614 5117 16626 5120
rect 16568 5111 16626 5117
rect 17494 5108 17500 5120
rect 17552 5108 17558 5160
rect 17862 5108 17868 5160
rect 17920 5148 17926 5160
rect 18616 5148 18644 5179
rect 19610 5176 19616 5188
rect 19668 5216 19674 5228
rect 19797 5219 19855 5225
rect 19797 5216 19809 5219
rect 19668 5188 19809 5216
rect 19668 5176 19674 5188
rect 19797 5185 19809 5188
rect 19843 5185 19855 5219
rect 20806 5216 20812 5228
rect 20767 5188 20812 5216
rect 19797 5179 19855 5185
rect 20806 5176 20812 5188
rect 20864 5176 20870 5228
rect 20898 5176 20904 5228
rect 20956 5216 20962 5228
rect 20956 5188 21001 5216
rect 20956 5176 20962 5188
rect 17920 5120 18644 5148
rect 17920 5108 17926 5120
rect 18690 5108 18696 5160
rect 18748 5148 18754 5160
rect 20622 5148 20628 5160
rect 18748 5120 20628 5148
rect 18748 5108 18754 5120
rect 20622 5108 20628 5120
rect 20680 5108 20686 5160
rect 20717 5151 20775 5157
rect 20717 5117 20729 5151
rect 20763 5148 20775 5151
rect 20990 5148 20996 5160
rect 20763 5120 20996 5148
rect 20763 5117 20775 5120
rect 20717 5111 20775 5117
rect 20990 5108 20996 5120
rect 21048 5108 21054 5160
rect 21174 5108 21180 5160
rect 21232 5148 21238 5160
rect 21361 5151 21419 5157
rect 21361 5148 21373 5151
rect 21232 5120 21373 5148
rect 21232 5108 21238 5120
rect 21361 5117 21373 5120
rect 21407 5117 21419 5151
rect 21361 5111 21419 5117
rect 13078 5080 13084 5092
rect 12544 5052 13084 5080
rect 13078 5040 13084 5052
rect 13136 5040 13142 5092
rect 14182 5040 14188 5092
rect 14240 5080 14246 5092
rect 15473 5083 15531 5089
rect 15473 5080 15485 5083
rect 14240 5052 15485 5080
rect 14240 5040 14246 5052
rect 15473 5049 15485 5052
rect 15519 5049 15531 5083
rect 15473 5043 15531 5049
rect 15654 5040 15660 5092
rect 15712 5080 15718 5092
rect 18874 5080 18880 5092
rect 15712 5052 18880 5080
rect 15712 5040 15718 5052
rect 18874 5040 18880 5052
rect 18932 5040 18938 5092
rect 19058 5040 19064 5092
rect 19116 5080 19122 5092
rect 19116 5052 19932 5080
rect 19116 5040 19122 5052
rect 12526 5012 12532 5024
rect 12452 4984 12532 5012
rect 12526 4972 12532 4984
rect 12584 4972 12590 5024
rect 13814 4972 13820 5024
rect 13872 5012 13878 5024
rect 14093 5015 14151 5021
rect 14093 5012 14105 5015
rect 13872 4984 14105 5012
rect 13872 4972 13878 4984
rect 14093 4981 14105 4984
rect 14139 4981 14151 5015
rect 14458 5012 14464 5024
rect 14419 4984 14464 5012
rect 14093 4975 14151 4981
rect 14458 4972 14464 4984
rect 14516 4972 14522 5024
rect 14550 4972 14556 5024
rect 14608 5012 14614 5024
rect 15565 5015 15623 5021
rect 15565 5012 15577 5015
rect 14608 4984 15577 5012
rect 14608 4972 14614 4984
rect 15565 4981 15577 4984
rect 15611 4981 15623 5015
rect 18414 5012 18420 5024
rect 18375 4984 18420 5012
rect 15565 4975 15623 4981
rect 18414 4972 18420 4984
rect 18472 4972 18478 5024
rect 19610 5012 19616 5024
rect 19571 4984 19616 5012
rect 19610 4972 19616 4984
rect 19668 4972 19674 5024
rect 19705 5015 19763 5021
rect 19705 4981 19717 5015
rect 19751 5012 19763 5015
rect 19794 5012 19800 5024
rect 19751 4984 19800 5012
rect 19751 4981 19763 4984
rect 19705 4975 19763 4981
rect 19794 4972 19800 4984
rect 19852 4972 19858 5024
rect 19904 5012 19932 5052
rect 20898 5040 20904 5092
rect 20956 5080 20962 5092
rect 21634 5089 21640 5092
rect 21606 5083 21640 5089
rect 21606 5080 21618 5083
rect 20956 5052 21618 5080
rect 20956 5040 20962 5052
rect 21606 5049 21618 5052
rect 21692 5080 21698 5092
rect 21692 5052 21754 5080
rect 21606 5043 21640 5049
rect 21634 5040 21640 5043
rect 21692 5040 21698 5052
rect 22741 5015 22799 5021
rect 22741 5012 22753 5015
rect 19904 4984 22753 5012
rect 22741 4981 22753 4984
rect 22787 4981 22799 5015
rect 22741 4975 22799 4981
rect 1104 4922 23276 4944
rect 1104 4870 8379 4922
rect 8431 4870 8443 4922
rect 8495 4870 8507 4922
rect 8559 4870 8571 4922
rect 8623 4870 15776 4922
rect 15828 4870 15840 4922
rect 15892 4870 15904 4922
rect 15956 4870 15968 4922
rect 16020 4870 23276 4922
rect 1104 4848 23276 4870
rect 9398 4768 9404 4820
rect 9456 4808 9462 4820
rect 10137 4811 10195 4817
rect 10137 4808 10149 4811
rect 9456 4780 10149 4808
rect 9456 4768 9462 4780
rect 10137 4777 10149 4780
rect 10183 4777 10195 4811
rect 10137 4771 10195 4777
rect 10410 4768 10416 4820
rect 10468 4808 10474 4820
rect 10597 4811 10655 4817
rect 10597 4808 10609 4811
rect 10468 4780 10609 4808
rect 10468 4768 10474 4780
rect 10597 4777 10609 4780
rect 10643 4777 10655 4811
rect 10597 4771 10655 4777
rect 11514 4768 11520 4820
rect 11572 4768 11578 4820
rect 12710 4808 12716 4820
rect 12671 4780 12716 4808
rect 12710 4768 12716 4780
rect 12768 4768 12774 4820
rect 12802 4768 12808 4820
rect 12860 4808 12866 4820
rect 12989 4811 13047 4817
rect 12989 4808 13001 4811
rect 12860 4780 13001 4808
rect 12860 4768 12866 4780
rect 12989 4777 13001 4780
rect 13035 4777 13047 4811
rect 13354 4808 13360 4820
rect 13315 4780 13360 4808
rect 12989 4771 13047 4777
rect 13354 4768 13360 4780
rect 13412 4768 13418 4820
rect 13449 4811 13507 4817
rect 13449 4777 13461 4811
rect 13495 4808 13507 4811
rect 13722 4808 13728 4820
rect 13495 4780 13728 4808
rect 13495 4777 13507 4780
rect 13449 4771 13507 4777
rect 13722 4768 13728 4780
rect 13780 4768 13786 4820
rect 14366 4808 14372 4820
rect 14327 4780 14372 4808
rect 14366 4768 14372 4780
rect 14424 4768 14430 4820
rect 15473 4811 15531 4817
rect 15473 4777 15485 4811
rect 15519 4808 15531 4811
rect 15654 4808 15660 4820
rect 15519 4780 15660 4808
rect 15519 4777 15531 4780
rect 15473 4771 15531 4777
rect 15654 4768 15660 4780
rect 15712 4768 15718 4820
rect 17218 4808 17224 4820
rect 16040 4780 17224 4808
rect 10505 4743 10563 4749
rect 10505 4709 10517 4743
rect 10551 4740 10563 4743
rect 11330 4740 11336 4752
rect 10551 4712 11336 4740
rect 10551 4709 10563 4712
rect 10505 4703 10563 4709
rect 11330 4700 11336 4712
rect 11388 4700 11394 4752
rect 11532 4672 11560 4768
rect 11600 4743 11658 4749
rect 11600 4709 11612 4743
rect 11646 4740 11658 4743
rect 12618 4740 12624 4752
rect 11646 4712 12624 4740
rect 11646 4709 11658 4712
rect 11600 4703 11658 4709
rect 12618 4700 12624 4712
rect 12676 4700 12682 4752
rect 16040 4740 16068 4780
rect 17218 4768 17224 4780
rect 17276 4768 17282 4820
rect 17497 4811 17555 4817
rect 17497 4777 17509 4811
rect 17543 4808 17555 4811
rect 18414 4808 18420 4820
rect 17543 4780 18420 4808
rect 17543 4777 17555 4780
rect 17497 4771 17555 4777
rect 18414 4768 18420 4780
rect 18472 4768 18478 4820
rect 19610 4768 19616 4820
rect 19668 4808 19674 4820
rect 19705 4811 19763 4817
rect 19705 4808 19717 4811
rect 19668 4780 19717 4808
rect 19668 4768 19674 4780
rect 19705 4777 19717 4780
rect 19751 4777 19763 4811
rect 19705 4771 19763 4777
rect 21634 4768 21640 4820
rect 21692 4808 21698 4820
rect 22741 4811 22799 4817
rect 22741 4808 22753 4811
rect 21692 4780 22753 4808
rect 21692 4768 21698 4780
rect 22741 4777 22753 4780
rect 22787 4777 22799 4811
rect 22741 4771 22799 4777
rect 15120 4712 16068 4740
rect 16108 4743 16166 4749
rect 15120 4672 15148 4712
rect 16108 4709 16120 4743
rect 16154 4740 16166 4743
rect 17678 4740 17684 4752
rect 16154 4712 17684 4740
rect 16154 4709 16166 4712
rect 16108 4703 16166 4709
rect 17678 4700 17684 4712
rect 17736 4700 17742 4752
rect 18322 4700 18328 4752
rect 18380 4740 18386 4752
rect 18966 4740 18972 4752
rect 18380 4712 18972 4740
rect 18380 4700 18386 4712
rect 18966 4700 18972 4712
rect 19024 4740 19030 4752
rect 19024 4712 19104 4740
rect 19024 4700 19030 4712
rect 15286 4672 15292 4684
rect 10796 4644 11560 4672
rect 14476 4644 15148 4672
rect 15247 4644 15292 4672
rect 10796 4613 10824 4644
rect 10781 4607 10839 4613
rect 10781 4573 10793 4607
rect 10827 4573 10839 4607
rect 10781 4567 10839 4573
rect 11238 4564 11244 4616
rect 11296 4604 11302 4616
rect 11333 4607 11391 4613
rect 11333 4604 11345 4607
rect 11296 4576 11345 4604
rect 11296 4564 11302 4576
rect 11333 4573 11345 4576
rect 11379 4573 11391 4607
rect 11333 4567 11391 4573
rect 12342 4564 12348 4616
rect 12400 4604 12406 4616
rect 13446 4604 13452 4616
rect 12400 4576 13452 4604
rect 12400 4564 12406 4576
rect 13446 4564 13452 4576
rect 13504 4564 13510 4616
rect 13538 4564 13544 4616
rect 13596 4604 13602 4616
rect 14476 4613 14504 4644
rect 15286 4632 15292 4644
rect 15344 4632 15350 4684
rect 15930 4672 15936 4684
rect 15856 4644 15936 4672
rect 14461 4607 14519 4613
rect 13596 4576 13641 4604
rect 13596 4564 13602 4576
rect 14461 4573 14473 4607
rect 14507 4573 14519 4607
rect 14642 4604 14648 4616
rect 14603 4576 14648 4604
rect 14461 4567 14519 4573
rect 14642 4564 14648 4576
rect 14700 4564 14706 4616
rect 15654 4564 15660 4616
rect 15712 4604 15718 4616
rect 15856 4613 15884 4644
rect 15930 4632 15936 4644
rect 15988 4632 15994 4684
rect 17126 4632 17132 4684
rect 17184 4672 17190 4684
rect 17865 4675 17923 4681
rect 17865 4672 17877 4675
rect 17184 4644 17877 4672
rect 17184 4632 17190 4644
rect 17865 4641 17877 4644
rect 17911 4641 17923 4675
rect 17865 4635 17923 4641
rect 18138 4632 18144 4684
rect 18196 4672 18202 4684
rect 18877 4675 18935 4681
rect 18877 4672 18889 4675
rect 18196 4644 18889 4672
rect 18196 4632 18202 4644
rect 18877 4641 18889 4644
rect 18923 4641 18935 4675
rect 18877 4635 18935 4641
rect 15841 4607 15899 4613
rect 15841 4604 15853 4607
rect 15712 4576 15853 4604
rect 15712 4564 15718 4576
rect 15841 4573 15853 4576
rect 15887 4573 15899 4607
rect 17957 4607 18015 4613
rect 17957 4604 17969 4607
rect 15841 4567 15899 4573
rect 17236 4576 17969 4604
rect 13170 4496 13176 4548
rect 13228 4536 13234 4548
rect 14001 4539 14059 4545
rect 14001 4536 14013 4539
rect 13228 4508 14013 4536
rect 13228 4496 13234 4508
rect 14001 4505 14013 4508
rect 14047 4505 14059 4539
rect 14001 4499 14059 4505
rect 8938 4428 8944 4480
rect 8996 4468 9002 4480
rect 13354 4468 13360 4480
rect 8996 4440 13360 4468
rect 8996 4428 9002 4440
rect 13354 4428 13360 4440
rect 13412 4428 13418 4480
rect 16574 4428 16580 4480
rect 16632 4468 16638 4480
rect 17236 4477 17264 4576
rect 17957 4573 17969 4576
rect 18003 4573 18015 4607
rect 17957 4567 18015 4573
rect 18049 4607 18107 4613
rect 18049 4573 18061 4607
rect 18095 4604 18107 4607
rect 18322 4604 18328 4616
rect 18095 4576 18328 4604
rect 18095 4573 18107 4576
rect 18049 4567 18107 4573
rect 18322 4564 18328 4576
rect 18380 4564 18386 4616
rect 19076 4613 19104 4712
rect 20714 4700 20720 4752
rect 20772 4740 20778 4752
rect 20901 4743 20959 4749
rect 20901 4740 20913 4743
rect 20772 4712 20913 4740
rect 20772 4700 20778 4712
rect 20901 4709 20913 4712
rect 20947 4709 20959 4743
rect 20901 4703 20959 4709
rect 20073 4675 20131 4681
rect 20073 4641 20085 4675
rect 20119 4672 20131 4675
rect 20806 4672 20812 4684
rect 20119 4644 20812 4672
rect 20119 4641 20131 4644
rect 20073 4635 20131 4641
rect 20806 4632 20812 4644
rect 20864 4632 20870 4684
rect 21628 4675 21686 4681
rect 21628 4641 21640 4675
rect 21674 4672 21686 4675
rect 21910 4672 21916 4684
rect 21674 4644 21916 4672
rect 21674 4641 21686 4644
rect 21628 4635 21686 4641
rect 21910 4632 21916 4644
rect 21968 4632 21974 4684
rect 18969 4607 19027 4613
rect 18969 4573 18981 4607
rect 19015 4573 19027 4607
rect 18969 4567 19027 4573
rect 19061 4607 19119 4613
rect 19061 4573 19073 4607
rect 19107 4573 19119 4607
rect 20162 4604 20168 4616
rect 20123 4576 20168 4604
rect 19061 4567 19119 4573
rect 17402 4496 17408 4548
rect 17460 4536 17466 4548
rect 18984 4536 19012 4567
rect 17460 4508 19012 4536
rect 19076 4536 19104 4567
rect 20162 4564 20168 4576
rect 20220 4564 20226 4616
rect 20257 4607 20315 4613
rect 20257 4573 20269 4607
rect 20303 4573 20315 4607
rect 20257 4567 20315 4573
rect 20272 4536 20300 4567
rect 20990 4564 20996 4616
rect 21048 4604 21054 4616
rect 21174 4604 21180 4616
rect 21048 4576 21180 4604
rect 21048 4564 21054 4576
rect 21174 4564 21180 4576
rect 21232 4604 21238 4616
rect 21361 4607 21419 4613
rect 21361 4604 21373 4607
rect 21232 4576 21373 4604
rect 21232 4564 21238 4576
rect 21361 4573 21373 4576
rect 21407 4573 21419 4607
rect 21361 4567 21419 4573
rect 20346 4536 20352 4548
rect 19076 4508 20352 4536
rect 17460 4496 17466 4508
rect 20346 4496 20352 4508
rect 20404 4496 20410 4548
rect 17221 4471 17279 4477
rect 17221 4468 17233 4471
rect 16632 4440 17233 4468
rect 16632 4428 16638 4440
rect 17221 4437 17233 4440
rect 17267 4437 17279 4471
rect 17221 4431 17279 4437
rect 17954 4428 17960 4480
rect 18012 4468 18018 4480
rect 18509 4471 18567 4477
rect 18509 4468 18521 4471
rect 18012 4440 18521 4468
rect 18012 4428 18018 4440
rect 18509 4437 18521 4440
rect 18555 4437 18567 4471
rect 18509 4431 18567 4437
rect 18690 4428 18696 4480
rect 18748 4468 18754 4480
rect 20622 4468 20628 4480
rect 18748 4440 20628 4468
rect 18748 4428 18754 4440
rect 20622 4428 20628 4440
rect 20680 4428 20686 4480
rect 1104 4378 23276 4400
rect 1104 4326 4680 4378
rect 4732 4326 4744 4378
rect 4796 4326 4808 4378
rect 4860 4326 4872 4378
rect 4924 4326 12078 4378
rect 12130 4326 12142 4378
rect 12194 4326 12206 4378
rect 12258 4326 12270 4378
rect 12322 4326 19475 4378
rect 19527 4326 19539 4378
rect 19591 4326 19603 4378
rect 19655 4326 19667 4378
rect 19719 4326 23276 4378
rect 1104 4304 23276 4326
rect 8110 4224 8116 4276
rect 8168 4264 8174 4276
rect 8168 4236 13308 4264
rect 8168 4224 8174 4236
rect 11422 4156 11428 4208
rect 11480 4196 11486 4208
rect 11480 4168 11928 4196
rect 11480 4156 11486 4168
rect 6914 4088 6920 4140
rect 6972 4128 6978 4140
rect 11900 4137 11928 4168
rect 13280 4137 13308 4236
rect 13354 4224 13360 4276
rect 13412 4264 13418 4276
rect 13725 4267 13783 4273
rect 13725 4264 13737 4267
rect 13412 4236 13737 4264
rect 13412 4224 13418 4236
rect 13725 4233 13737 4236
rect 13771 4233 13783 4267
rect 17126 4264 17132 4276
rect 13725 4227 13783 4233
rect 15304 4236 16988 4264
rect 17087 4236 17132 4264
rect 13446 4156 13452 4208
rect 13504 4196 13510 4208
rect 15304 4196 15332 4236
rect 13504 4168 15332 4196
rect 16960 4196 16988 4236
rect 17126 4224 17132 4236
rect 17184 4224 17190 4276
rect 17218 4224 17224 4276
rect 17276 4264 17282 4276
rect 19058 4264 19064 4276
rect 17276 4236 19064 4264
rect 17276 4224 17282 4236
rect 19058 4224 19064 4236
rect 19116 4224 19122 4276
rect 19705 4267 19763 4273
rect 19705 4233 19717 4267
rect 19751 4264 19763 4267
rect 19794 4264 19800 4276
rect 19751 4236 19800 4264
rect 19751 4233 19763 4236
rect 19705 4227 19763 4233
rect 19794 4224 19800 4236
rect 19852 4224 19858 4276
rect 17862 4196 17868 4208
rect 16960 4168 17868 4196
rect 13504 4156 13510 4168
rect 11885 4131 11943 4137
rect 6972 4100 11836 4128
rect 6972 4088 6978 4100
rect 10778 4060 10784 4072
rect 10739 4032 10784 4060
rect 10778 4020 10784 4032
rect 10836 4020 10842 4072
rect 11698 4060 11704 4072
rect 11659 4032 11704 4060
rect 11698 4020 11704 4032
rect 11756 4020 11762 4072
rect 11808 4060 11836 4100
rect 11885 4097 11897 4131
rect 11931 4097 11943 4131
rect 11885 4091 11943 4097
rect 13265 4131 13323 4137
rect 13265 4097 13277 4131
rect 13311 4097 13323 4131
rect 14274 4128 14280 4140
rect 14235 4100 14280 4128
rect 13265 4091 13323 4097
rect 14274 4088 14280 4100
rect 14332 4088 14338 4140
rect 14645 4131 14703 4137
rect 14645 4097 14657 4131
rect 14691 4128 14703 4131
rect 15010 4128 15016 4140
rect 14691 4100 15016 4128
rect 14691 4097 14703 4100
rect 14645 4091 14703 4097
rect 15010 4088 15016 4100
rect 15068 4088 15074 4140
rect 15304 4137 15332 4168
rect 17862 4156 17868 4168
rect 17920 4156 17926 4208
rect 20346 4196 20352 4208
rect 20272 4168 20352 4196
rect 20272 4137 20300 4168
rect 20346 4156 20352 4168
rect 20404 4156 20410 4208
rect 15289 4131 15347 4137
rect 15289 4097 15301 4131
rect 15335 4097 15347 4131
rect 20257 4131 20315 4137
rect 15289 4091 15347 4097
rect 17420 4100 18184 4128
rect 13170 4060 13176 4072
rect 11808 4032 11928 4060
rect 13131 4032 13176 4060
rect 7282 3952 7288 4004
rect 7340 3992 7346 4004
rect 7340 3964 11376 3992
rect 7340 3952 7346 3964
rect 5166 3884 5172 3936
rect 5224 3924 5230 3936
rect 11348 3933 11376 3964
rect 11606 3952 11612 4004
rect 11664 3992 11670 4004
rect 11793 3995 11851 4001
rect 11793 3992 11805 3995
rect 11664 3964 11805 3992
rect 11664 3952 11670 3964
rect 11793 3961 11805 3964
rect 11839 3961 11851 3995
rect 11793 3955 11851 3961
rect 10965 3927 11023 3933
rect 10965 3924 10977 3927
rect 5224 3896 10977 3924
rect 5224 3884 5230 3896
rect 10965 3893 10977 3896
rect 11011 3893 11023 3927
rect 10965 3887 11023 3893
rect 11333 3927 11391 3933
rect 11333 3893 11345 3927
rect 11379 3893 11391 3927
rect 11900 3924 11928 4032
rect 13170 4020 13176 4032
rect 13228 4020 13234 4072
rect 14185 4063 14243 4069
rect 14185 4029 14197 4063
rect 14231 4060 14243 4063
rect 14734 4060 14740 4072
rect 14231 4032 14740 4060
rect 14231 4029 14243 4032
rect 14185 4023 14243 4029
rect 14734 4020 14740 4032
rect 14792 4020 14798 4072
rect 15105 4063 15163 4069
rect 15105 4029 15117 4063
rect 15151 4060 15163 4063
rect 15194 4060 15200 4072
rect 15151 4032 15200 4060
rect 15151 4029 15163 4032
rect 15105 4023 15163 4029
rect 15194 4020 15200 4032
rect 15252 4020 15258 4072
rect 15654 4020 15660 4072
rect 15712 4060 15718 4072
rect 15749 4063 15807 4069
rect 15749 4060 15761 4063
rect 15712 4032 15761 4060
rect 15712 4020 15718 4032
rect 15749 4029 15761 4032
rect 15795 4029 15807 4063
rect 15749 4023 15807 4029
rect 16016 4063 16074 4069
rect 16016 4029 16028 4063
rect 16062 4060 16074 4063
rect 16574 4060 16580 4072
rect 16062 4032 16580 4060
rect 16062 4029 16074 4032
rect 16016 4023 16074 4029
rect 16574 4020 16580 4032
rect 16632 4020 16638 4072
rect 17420 4069 17448 4100
rect 17405 4063 17463 4069
rect 17405 4029 17417 4063
rect 17451 4029 17463 4063
rect 17405 4023 17463 4029
rect 17494 4020 17500 4072
rect 17552 4060 17558 4072
rect 17770 4060 17776 4072
rect 17552 4032 17776 4060
rect 17552 4020 17558 4032
rect 17770 4020 17776 4032
rect 17828 4060 17834 4072
rect 18049 4063 18107 4069
rect 18049 4060 18061 4063
rect 17828 4032 18061 4060
rect 17828 4020 17834 4032
rect 18049 4029 18061 4032
rect 18095 4029 18107 4063
rect 18156 4060 18184 4100
rect 20257 4097 20269 4131
rect 20303 4097 20315 4131
rect 20257 4091 20315 4097
rect 18598 4060 18604 4072
rect 18156 4032 18604 4060
rect 18049 4023 18107 4029
rect 12802 3952 12808 4004
rect 12860 3992 12866 4004
rect 14550 3992 14556 4004
rect 12860 3964 14556 3992
rect 12860 3952 12866 3964
rect 14550 3952 14556 3964
rect 14608 3952 14614 4004
rect 15286 3992 15292 4004
rect 14752 3964 15292 3992
rect 12713 3927 12771 3933
rect 12713 3924 12725 3927
rect 11900 3896 12725 3924
rect 11333 3887 11391 3893
rect 12713 3893 12725 3896
rect 12759 3893 12771 3927
rect 12713 3887 12771 3893
rect 13081 3927 13139 3933
rect 13081 3893 13093 3927
rect 13127 3924 13139 3927
rect 13170 3924 13176 3936
rect 13127 3896 13176 3924
rect 13127 3893 13139 3896
rect 13081 3887 13139 3893
rect 13170 3884 13176 3896
rect 13228 3884 13234 3936
rect 14752 3933 14780 3964
rect 15286 3952 15292 3964
rect 15344 3952 15350 4004
rect 17954 3992 17960 4004
rect 16868 3964 17960 3992
rect 14093 3927 14151 3933
rect 14093 3893 14105 3927
rect 14139 3924 14151 3927
rect 14645 3927 14703 3933
rect 14645 3924 14657 3927
rect 14139 3896 14657 3924
rect 14139 3893 14151 3896
rect 14093 3887 14151 3893
rect 14645 3893 14657 3896
rect 14691 3893 14703 3927
rect 14645 3887 14703 3893
rect 14737 3927 14795 3933
rect 14737 3893 14749 3927
rect 14783 3893 14795 3927
rect 14737 3887 14795 3893
rect 15197 3927 15255 3933
rect 15197 3893 15209 3927
rect 15243 3924 15255 3927
rect 16868 3924 16896 3964
rect 17954 3952 17960 3964
rect 18012 3952 18018 4004
rect 15243 3896 16896 3924
rect 15243 3893 15255 3896
rect 15197 3887 15255 3893
rect 17310 3884 17316 3936
rect 17368 3924 17374 3936
rect 17589 3927 17647 3933
rect 17589 3924 17601 3927
rect 17368 3896 17601 3924
rect 17368 3884 17374 3896
rect 17589 3893 17601 3896
rect 17635 3893 17647 3927
rect 18064 3924 18092 4023
rect 18598 4020 18604 4032
rect 18656 4020 18662 4072
rect 19242 4020 19248 4072
rect 19300 4060 19306 4072
rect 19300 4032 20300 4060
rect 19300 4020 19306 4032
rect 18316 3995 18374 4001
rect 18316 3961 18328 3995
rect 18362 3992 18374 3995
rect 18874 3992 18880 4004
rect 18362 3964 18880 3992
rect 18362 3961 18374 3964
rect 18316 3955 18374 3961
rect 18874 3952 18880 3964
rect 18932 3952 18938 4004
rect 20165 3995 20223 4001
rect 20165 3992 20177 3995
rect 19444 3964 20177 3992
rect 19444 3936 19472 3964
rect 20165 3961 20177 3964
rect 20211 3961 20223 3995
rect 20272 3992 20300 4032
rect 20530 4020 20536 4072
rect 20588 4060 20594 4072
rect 20717 4063 20775 4069
rect 20717 4060 20729 4063
rect 20588 4032 20729 4060
rect 20588 4020 20594 4032
rect 20717 4029 20729 4032
rect 20763 4029 20775 4063
rect 20898 4060 20904 4072
rect 20859 4032 20904 4060
rect 20717 4023 20775 4029
rect 20898 4020 20904 4032
rect 20956 4020 20962 4072
rect 20990 4020 20996 4072
rect 21048 4060 21054 4072
rect 21361 4063 21419 4069
rect 21361 4060 21373 4063
rect 21048 4032 21373 4060
rect 21048 4020 21054 4032
rect 21361 4029 21373 4032
rect 21407 4029 21419 4063
rect 21361 4023 21419 4029
rect 21628 4063 21686 4069
rect 21628 4029 21640 4063
rect 21674 4060 21686 4063
rect 22002 4060 22008 4072
rect 21674 4032 22008 4060
rect 21674 4029 21686 4032
rect 21628 4023 21686 4029
rect 21836 4004 21864 4032
rect 22002 4020 22008 4032
rect 22060 4020 22066 4072
rect 21085 3995 21143 4001
rect 21085 3992 21097 3995
rect 20272 3964 21097 3992
rect 20165 3955 20223 3961
rect 21085 3961 21097 3964
rect 21131 3961 21143 3995
rect 21085 3955 21143 3961
rect 21818 3952 21824 4004
rect 21876 3952 21882 4004
rect 19058 3924 19064 3936
rect 18064 3896 19064 3924
rect 17589 3887 17647 3893
rect 19058 3884 19064 3896
rect 19116 3884 19122 3936
rect 19426 3924 19432 3936
rect 19339 3896 19432 3924
rect 19426 3884 19432 3896
rect 19484 3884 19490 3936
rect 20073 3927 20131 3933
rect 20073 3893 20085 3927
rect 20119 3924 20131 3927
rect 20438 3924 20444 3936
rect 20119 3896 20444 3924
rect 20119 3893 20131 3896
rect 20073 3887 20131 3893
rect 20438 3884 20444 3896
rect 20496 3884 20502 3936
rect 21910 3884 21916 3936
rect 21968 3924 21974 3936
rect 22741 3927 22799 3933
rect 22741 3924 22753 3927
rect 21968 3896 22753 3924
rect 21968 3884 21974 3896
rect 22741 3893 22753 3896
rect 22787 3893 22799 3927
rect 22741 3887 22799 3893
rect 1104 3834 23276 3856
rect 1104 3782 8379 3834
rect 8431 3782 8443 3834
rect 8495 3782 8507 3834
rect 8559 3782 8571 3834
rect 8623 3782 15776 3834
rect 15828 3782 15840 3834
rect 15892 3782 15904 3834
rect 15956 3782 15968 3834
rect 16020 3782 23276 3834
rect 1104 3760 23276 3782
rect 10318 3720 10324 3732
rect 2516 3692 10324 3720
rect 2516 3593 2544 3692
rect 10318 3680 10324 3692
rect 10376 3680 10382 3732
rect 12802 3720 12808 3732
rect 12763 3692 12808 3720
rect 12802 3680 12808 3692
rect 12860 3680 12866 3732
rect 16942 3720 16948 3732
rect 14200 3692 16948 3720
rect 3237 3655 3295 3661
rect 3237 3621 3249 3655
rect 3283 3652 3295 3655
rect 3878 3652 3884 3664
rect 3283 3624 3884 3652
rect 3283 3621 3295 3624
rect 3237 3615 3295 3621
rect 3878 3612 3884 3624
rect 3936 3612 3942 3664
rect 13630 3652 13636 3664
rect 12636 3624 13636 3652
rect 2501 3587 2559 3593
rect 2501 3553 2513 3587
rect 2547 3553 2559 3587
rect 2501 3547 2559 3553
rect 11977 3587 12035 3593
rect 11977 3553 11989 3587
rect 12023 3584 12035 3587
rect 12434 3584 12440 3596
rect 12023 3556 12440 3584
rect 12023 3553 12035 3556
rect 11977 3547 12035 3553
rect 1762 3476 1768 3528
rect 1820 3516 1826 3528
rect 2516 3516 2544 3547
rect 12434 3544 12440 3556
rect 12492 3544 12498 3596
rect 12636 3593 12664 3624
rect 13630 3612 13636 3624
rect 13688 3612 13694 3664
rect 12621 3587 12679 3593
rect 12621 3553 12633 3587
rect 12667 3553 12679 3587
rect 13538 3584 13544 3596
rect 13499 3556 13544 3584
rect 12621 3547 12679 3553
rect 13538 3544 13544 3556
rect 13596 3544 13602 3596
rect 1820 3488 2544 3516
rect 1820 3476 1826 3488
rect 12066 3476 12072 3528
rect 12124 3516 12130 3528
rect 13630 3516 13636 3528
rect 12124 3488 12940 3516
rect 13591 3488 13636 3516
rect 12124 3476 12130 3488
rect 12161 3451 12219 3457
rect 12161 3417 12173 3451
rect 12207 3448 12219 3451
rect 12802 3448 12808 3460
rect 12207 3420 12808 3448
rect 12207 3417 12219 3420
rect 12161 3411 12219 3417
rect 12802 3408 12808 3420
rect 12860 3408 12866 3460
rect 2498 3340 2504 3392
rect 2556 3380 2562 3392
rect 11606 3380 11612 3392
rect 2556 3352 11612 3380
rect 2556 3340 2562 3352
rect 11606 3340 11612 3352
rect 11664 3380 11670 3392
rect 11974 3380 11980 3392
rect 11664 3352 11980 3380
rect 11664 3340 11670 3352
rect 11974 3340 11980 3352
rect 12032 3340 12038 3392
rect 12912 3380 12940 3488
rect 13630 3476 13636 3488
rect 13688 3476 13694 3528
rect 13817 3519 13875 3525
rect 13817 3485 13829 3519
rect 13863 3516 13875 3519
rect 14200 3516 14228 3692
rect 16942 3680 16948 3692
rect 17000 3680 17006 3732
rect 18874 3720 18880 3732
rect 18835 3692 18880 3720
rect 18874 3680 18880 3692
rect 18932 3680 18938 3732
rect 21542 3680 21548 3732
rect 21600 3720 21606 3732
rect 22281 3723 22339 3729
rect 22281 3720 22293 3723
rect 21600 3692 22293 3720
rect 21600 3680 21606 3692
rect 22281 3689 22293 3692
rect 22327 3689 22339 3723
rect 22281 3683 22339 3689
rect 14645 3655 14703 3661
rect 14645 3621 14657 3655
rect 14691 3652 14703 3655
rect 14918 3652 14924 3664
rect 14691 3624 14924 3652
rect 14691 3621 14703 3624
rect 14645 3615 14703 3621
rect 14918 3612 14924 3624
rect 14976 3612 14982 3664
rect 16108 3655 16166 3661
rect 16108 3621 16120 3655
rect 16154 3652 16166 3655
rect 17126 3652 17132 3664
rect 16154 3624 17132 3652
rect 16154 3621 16166 3624
rect 16108 3615 16166 3621
rect 17126 3612 17132 3624
rect 17184 3612 17190 3664
rect 19426 3661 19432 3664
rect 19420 3652 19432 3661
rect 19387 3624 19432 3652
rect 19420 3615 19432 3624
rect 19426 3612 19432 3615
rect 19484 3612 19490 3664
rect 21168 3655 21226 3661
rect 21168 3621 21180 3655
rect 21214 3652 21226 3655
rect 21726 3652 21732 3664
rect 21214 3624 21732 3652
rect 21214 3621 21226 3624
rect 21168 3615 21226 3621
rect 21726 3612 21732 3624
rect 21784 3612 21790 3664
rect 14553 3587 14611 3593
rect 14553 3553 14565 3587
rect 14599 3584 14611 3587
rect 14826 3584 14832 3596
rect 14599 3556 14832 3584
rect 14599 3553 14611 3556
rect 14553 3547 14611 3553
rect 14826 3544 14832 3556
rect 14884 3544 14890 3596
rect 15289 3587 15347 3593
rect 15289 3553 15301 3587
rect 15335 3584 15347 3587
rect 17586 3584 17592 3596
rect 15335 3556 17592 3584
rect 15335 3553 15347 3556
rect 15289 3547 15347 3553
rect 17586 3544 17592 3556
rect 17644 3544 17650 3596
rect 17770 3593 17776 3596
rect 17764 3547 17776 3593
rect 17828 3584 17834 3596
rect 17828 3556 17864 3584
rect 17770 3544 17776 3547
rect 17828 3544 17834 3556
rect 19058 3544 19064 3596
rect 19116 3584 19122 3596
rect 19153 3587 19211 3593
rect 19153 3584 19165 3587
rect 19116 3556 19165 3584
rect 19116 3544 19122 3556
rect 19153 3553 19165 3556
rect 19199 3553 19211 3587
rect 19153 3547 19211 3553
rect 13863 3488 14228 3516
rect 13863 3485 13875 3488
rect 13817 3479 13875 3485
rect 14274 3476 14280 3528
rect 14332 3516 14338 3528
rect 14737 3519 14795 3525
rect 14737 3516 14749 3519
rect 14332 3488 14749 3516
rect 14332 3476 14338 3488
rect 14737 3485 14749 3488
rect 14783 3516 14795 3519
rect 15562 3516 15568 3528
rect 14783 3488 15568 3516
rect 14783 3485 14795 3488
rect 14737 3479 14795 3485
rect 15562 3476 15568 3488
rect 15620 3476 15626 3528
rect 15654 3476 15660 3528
rect 15712 3516 15718 3528
rect 15841 3519 15899 3525
rect 15841 3516 15853 3519
rect 15712 3488 15853 3516
rect 15712 3476 15718 3488
rect 15841 3485 15853 3488
rect 15887 3485 15899 3519
rect 17494 3516 17500 3528
rect 17455 3488 17500 3516
rect 15841 3479 15899 3485
rect 17494 3476 17500 3488
rect 17552 3476 17558 3528
rect 20898 3516 20904 3528
rect 20859 3488 20904 3516
rect 20898 3476 20904 3488
rect 20956 3476 20962 3528
rect 12986 3408 12992 3460
rect 13044 3448 13050 3460
rect 14185 3451 14243 3457
rect 14185 3448 14197 3451
rect 13044 3420 14197 3448
rect 13044 3408 13050 3420
rect 14185 3417 14197 3420
rect 14231 3417 14243 3451
rect 14185 3411 14243 3417
rect 17221 3451 17279 3457
rect 17221 3417 17233 3451
rect 17267 3448 17279 3451
rect 17402 3448 17408 3460
rect 17267 3420 17408 3448
rect 17267 3417 17279 3420
rect 17221 3411 17279 3417
rect 17402 3408 17408 3420
rect 17460 3408 17466 3460
rect 13173 3383 13231 3389
rect 13173 3380 13185 3383
rect 12912 3352 13185 3380
rect 13173 3349 13185 3352
rect 13219 3380 13231 3383
rect 14366 3380 14372 3392
rect 13219 3352 14372 3380
rect 13219 3349 13231 3352
rect 13173 3343 13231 3349
rect 14366 3340 14372 3352
rect 14424 3340 14430 3392
rect 15473 3383 15531 3389
rect 15473 3349 15485 3383
rect 15519 3380 15531 3383
rect 20254 3380 20260 3392
rect 15519 3352 20260 3380
rect 15519 3349 15531 3352
rect 15473 3343 15531 3349
rect 20254 3340 20260 3352
rect 20312 3340 20318 3392
rect 20438 3340 20444 3392
rect 20496 3380 20502 3392
rect 20533 3383 20591 3389
rect 20533 3380 20545 3383
rect 20496 3352 20545 3380
rect 20496 3340 20502 3352
rect 20533 3349 20545 3352
rect 20579 3349 20591 3383
rect 20533 3343 20591 3349
rect 1104 3290 23276 3312
rect 1104 3238 4680 3290
rect 4732 3238 4744 3290
rect 4796 3238 4808 3290
rect 4860 3238 4872 3290
rect 4924 3238 12078 3290
rect 12130 3238 12142 3290
rect 12194 3238 12206 3290
rect 12258 3238 12270 3290
rect 12322 3238 19475 3290
rect 19527 3238 19539 3290
rect 19591 3238 19603 3290
rect 19655 3238 19667 3290
rect 19719 3238 23276 3290
rect 1104 3216 23276 3238
rect 13078 3176 13084 3188
rect 13039 3148 13084 3176
rect 13078 3136 13084 3148
rect 13136 3136 13142 3188
rect 13630 3136 13636 3188
rect 13688 3176 13694 3188
rect 14001 3179 14059 3185
rect 14001 3176 14013 3179
rect 13688 3148 14013 3176
rect 13688 3136 13694 3148
rect 14001 3145 14013 3148
rect 14047 3145 14059 3179
rect 16390 3176 16396 3188
rect 14001 3139 14059 3145
rect 16040 3148 16396 3176
rect 2590 3068 2596 3120
rect 2648 3108 2654 3120
rect 15013 3111 15071 3117
rect 15013 3108 15025 3111
rect 2648 3080 15025 3108
rect 2648 3068 2654 3080
rect 15013 3077 15025 3080
rect 15059 3077 15071 3111
rect 15013 3071 15071 3077
rect 1946 3040 1952 3052
rect 1907 3012 1952 3040
rect 1946 3000 1952 3012
rect 2004 3000 2010 3052
rect 14645 3043 14703 3049
rect 14645 3009 14657 3043
rect 14691 3040 14703 3043
rect 15470 3040 15476 3052
rect 14691 3012 15476 3040
rect 14691 3009 14703 3012
rect 14645 3003 14703 3009
rect 15470 3000 15476 3012
rect 15528 3000 15534 3052
rect 15562 3000 15568 3052
rect 15620 3040 15626 3052
rect 16040 3049 16068 3148
rect 16390 3136 16396 3148
rect 16448 3176 16454 3188
rect 17405 3179 17463 3185
rect 16448 3148 16988 3176
rect 16448 3136 16454 3148
rect 16960 3108 16988 3148
rect 17405 3145 17417 3179
rect 17451 3176 17463 3179
rect 18138 3176 18144 3188
rect 17451 3148 18144 3176
rect 17451 3145 17463 3148
rect 17405 3139 17463 3145
rect 18138 3136 18144 3148
rect 18196 3136 18202 3188
rect 20162 3136 20168 3188
rect 20220 3176 20226 3188
rect 20257 3179 20315 3185
rect 20257 3176 20269 3179
rect 20220 3148 20269 3176
rect 20220 3136 20226 3148
rect 20257 3145 20269 3148
rect 20303 3145 20315 3179
rect 20257 3139 20315 3145
rect 21726 3136 21732 3188
rect 21784 3176 21790 3188
rect 21913 3179 21971 3185
rect 21913 3176 21925 3179
rect 21784 3148 21925 3176
rect 21784 3136 21790 3148
rect 21913 3145 21925 3148
rect 21959 3145 21971 3179
rect 21913 3139 21971 3145
rect 17494 3108 17500 3120
rect 16960 3080 17500 3108
rect 17494 3068 17500 3080
rect 17552 3068 17558 3120
rect 18046 3068 18052 3120
rect 18104 3108 18110 3120
rect 18509 3111 18567 3117
rect 18509 3108 18521 3111
rect 18104 3080 18521 3108
rect 18104 3068 18110 3080
rect 18509 3077 18521 3080
rect 18555 3077 18567 3111
rect 18509 3071 18567 3077
rect 16025 3043 16083 3049
rect 15620 3012 15665 3040
rect 15620 3000 15626 3012
rect 16025 3009 16037 3043
rect 16071 3009 16083 3043
rect 16025 3003 16083 3009
rect 1762 2972 1768 2984
rect 1723 2944 1768 2972
rect 1762 2932 1768 2944
rect 1820 2932 1826 2984
rect 2498 2972 2504 2984
rect 2459 2944 2504 2972
rect 2498 2932 2504 2944
rect 2556 2932 2562 2984
rect 5074 2972 5080 2984
rect 5035 2944 5080 2972
rect 5074 2932 5080 2944
rect 5132 2932 5138 2984
rect 11882 2932 11888 2984
rect 11940 2972 11946 2984
rect 12897 2975 12955 2981
rect 12897 2972 12909 2975
rect 11940 2944 12909 2972
rect 11940 2932 11946 2944
rect 12897 2941 12909 2944
rect 12943 2941 12955 2975
rect 12897 2935 12955 2941
rect 13449 2975 13507 2981
rect 13449 2941 13461 2975
rect 13495 2972 13507 2975
rect 13906 2972 13912 2984
rect 13495 2944 13912 2972
rect 13495 2941 13507 2944
rect 13449 2935 13507 2941
rect 13906 2932 13912 2944
rect 13964 2932 13970 2984
rect 15381 2975 15439 2981
rect 15381 2941 15393 2975
rect 15427 2972 15439 2975
rect 16114 2972 16120 2984
rect 15427 2944 16120 2972
rect 15427 2941 15439 2944
rect 15381 2935 15439 2941
rect 16114 2932 16120 2944
rect 16172 2932 16178 2984
rect 16292 2975 16350 2981
rect 16292 2941 16304 2975
rect 16338 2972 16350 2975
rect 17402 2972 17408 2984
rect 16338 2944 17408 2972
rect 16338 2941 16350 2944
rect 16292 2935 16350 2941
rect 17402 2932 17408 2944
rect 17460 2932 17466 2984
rect 18325 2975 18383 2981
rect 18325 2941 18337 2975
rect 18371 2972 18383 2975
rect 18782 2972 18788 2984
rect 18371 2944 18788 2972
rect 18371 2941 18383 2944
rect 18325 2935 18383 2941
rect 18782 2932 18788 2944
rect 18840 2932 18846 2984
rect 18877 2975 18935 2981
rect 18877 2941 18889 2975
rect 18923 2941 18935 2975
rect 18877 2935 18935 2941
rect 19144 2975 19202 2981
rect 19144 2941 19156 2975
rect 19190 2972 19202 2975
rect 20438 2972 20444 2984
rect 19190 2944 20444 2972
rect 19190 2941 19202 2944
rect 19144 2935 19202 2941
rect 2130 2864 2136 2916
rect 2188 2904 2194 2916
rect 14369 2907 14427 2913
rect 14369 2904 14381 2907
rect 2188 2876 14381 2904
rect 2188 2864 2194 2876
rect 14369 2873 14381 2876
rect 14415 2873 14427 2907
rect 14369 2867 14427 2873
rect 15473 2907 15531 2913
rect 15473 2873 15485 2907
rect 15519 2904 15531 2907
rect 17034 2904 17040 2916
rect 15519 2876 17040 2904
rect 15519 2873 15531 2876
rect 15473 2867 15531 2873
rect 17034 2864 17040 2876
rect 17092 2864 17098 2916
rect 18892 2904 18920 2935
rect 20438 2932 20444 2944
rect 20496 2932 20502 2984
rect 20806 2981 20812 2984
rect 20533 2975 20591 2981
rect 20533 2941 20545 2975
rect 20579 2941 20591 2975
rect 20800 2972 20812 2981
rect 20767 2944 20812 2972
rect 20533 2935 20591 2941
rect 20800 2935 20812 2944
rect 19058 2904 19064 2916
rect 18892 2876 19064 2904
rect 19058 2864 19064 2876
rect 19116 2904 19122 2916
rect 20548 2904 20576 2935
rect 20806 2932 20812 2935
rect 20864 2932 20870 2984
rect 22094 2932 22100 2984
rect 22152 2972 22158 2984
rect 22189 2975 22247 2981
rect 22189 2972 22201 2975
rect 22152 2944 22201 2972
rect 22152 2932 22158 2944
rect 22189 2941 22201 2944
rect 22235 2941 22247 2975
rect 22189 2935 22247 2941
rect 20898 2904 20904 2916
rect 19116 2876 20904 2904
rect 19116 2864 19122 2876
rect 20898 2864 20904 2876
rect 20956 2864 20962 2916
rect 22465 2907 22523 2913
rect 22465 2873 22477 2907
rect 22511 2904 22523 2907
rect 22554 2904 22560 2916
rect 22511 2876 22560 2904
rect 22511 2873 22523 2876
rect 22465 2867 22523 2873
rect 22554 2864 22560 2876
rect 22612 2864 22618 2916
rect 1670 2796 1676 2848
rect 1728 2836 1734 2848
rect 2685 2839 2743 2845
rect 2685 2836 2697 2839
rect 1728 2808 2697 2836
rect 1728 2796 1734 2808
rect 2685 2805 2697 2808
rect 2731 2805 2743 2839
rect 2685 2799 2743 2805
rect 7006 2796 7012 2848
rect 7064 2836 7070 2848
rect 12986 2836 12992 2848
rect 7064 2808 12992 2836
rect 7064 2796 7070 2808
rect 12986 2796 12992 2808
rect 13044 2796 13050 2848
rect 13633 2839 13691 2845
rect 13633 2805 13645 2839
rect 13679 2836 13691 2839
rect 14182 2836 14188 2848
rect 13679 2808 14188 2836
rect 13679 2805 13691 2808
rect 13633 2799 13691 2805
rect 14182 2796 14188 2808
rect 14240 2796 14246 2848
rect 14458 2796 14464 2848
rect 14516 2836 14522 2848
rect 14516 2808 14561 2836
rect 14516 2796 14522 2808
rect 17678 2796 17684 2848
rect 17736 2836 17742 2848
rect 22738 2836 22744 2848
rect 17736 2808 22744 2836
rect 17736 2796 17742 2808
rect 22738 2796 22744 2808
rect 22796 2796 22802 2848
rect 1104 2746 23276 2768
rect 1104 2694 8379 2746
rect 8431 2694 8443 2746
rect 8495 2694 8507 2746
rect 8559 2694 8571 2746
rect 8623 2694 15776 2746
rect 15828 2694 15840 2746
rect 15892 2694 15904 2746
rect 15956 2694 15968 2746
rect 16020 2694 23276 2746
rect 1104 2672 23276 2694
rect 14001 2635 14059 2641
rect 14001 2601 14013 2635
rect 14047 2601 14059 2635
rect 14001 2595 14059 2601
rect 14016 2564 14044 2595
rect 14366 2592 14372 2644
rect 14424 2632 14430 2644
rect 14737 2635 14795 2641
rect 14737 2632 14749 2635
rect 14424 2604 14749 2632
rect 14424 2592 14430 2604
rect 14737 2601 14749 2604
rect 14783 2601 14795 2635
rect 14737 2595 14795 2601
rect 15841 2635 15899 2641
rect 15841 2601 15853 2635
rect 15887 2632 15899 2635
rect 15887 2604 16712 2632
rect 15887 2601 15899 2604
rect 15841 2595 15899 2601
rect 14458 2564 14464 2576
rect 14016 2536 14464 2564
rect 14458 2524 14464 2536
rect 14516 2524 14522 2576
rect 15562 2524 15568 2576
rect 15620 2564 15626 2576
rect 15620 2536 16068 2564
rect 15620 2524 15626 2536
rect 3050 2456 3056 2508
rect 3108 2496 3114 2508
rect 13817 2499 13875 2505
rect 13817 2496 13829 2499
rect 3108 2468 13829 2496
rect 3108 2456 3114 2468
rect 13817 2465 13829 2468
rect 13863 2465 13875 2499
rect 15930 2496 15936 2508
rect 15891 2468 15936 2496
rect 13817 2459 13875 2465
rect 15930 2456 15936 2468
rect 15988 2456 15994 2508
rect 14826 2428 14832 2440
rect 14787 2400 14832 2428
rect 14826 2388 14832 2400
rect 14884 2388 14890 2440
rect 15010 2428 15016 2440
rect 14971 2400 15016 2428
rect 15010 2388 15016 2400
rect 15068 2388 15074 2440
rect 16040 2437 16068 2536
rect 16390 2456 16396 2508
rect 16448 2496 16454 2508
rect 16485 2499 16543 2505
rect 16485 2496 16497 2499
rect 16448 2468 16497 2496
rect 16448 2456 16454 2468
rect 16485 2465 16497 2468
rect 16531 2465 16543 2499
rect 16684 2496 16712 2604
rect 17770 2592 17776 2644
rect 17828 2632 17834 2644
rect 17865 2635 17923 2641
rect 17865 2632 17877 2635
rect 17828 2604 17877 2632
rect 17828 2592 17834 2604
rect 17865 2601 17877 2604
rect 17911 2632 17923 2635
rect 18693 2635 18751 2641
rect 17911 2604 18276 2632
rect 17911 2601 17923 2604
rect 17865 2595 17923 2601
rect 16752 2567 16810 2573
rect 16752 2533 16764 2567
rect 16798 2564 16810 2567
rect 18138 2564 18144 2576
rect 16798 2536 18144 2564
rect 16798 2533 16810 2536
rect 16752 2527 16810 2533
rect 18138 2524 18144 2536
rect 18196 2524 18202 2576
rect 18248 2564 18276 2604
rect 18693 2601 18705 2635
rect 18739 2632 18751 2635
rect 18874 2632 18880 2644
rect 18739 2604 18880 2632
rect 18739 2601 18751 2604
rect 18693 2595 18751 2601
rect 18874 2592 18880 2604
rect 18932 2592 18938 2644
rect 20717 2635 20775 2641
rect 18984 2604 20300 2632
rect 18785 2567 18843 2573
rect 18785 2564 18797 2567
rect 18248 2536 18797 2564
rect 18785 2533 18797 2536
rect 18831 2533 18843 2567
rect 18785 2527 18843 2533
rect 18984 2496 19012 2604
rect 19604 2567 19662 2573
rect 19604 2533 19616 2567
rect 19650 2564 19662 2567
rect 20162 2564 20168 2576
rect 19650 2536 20168 2564
rect 19650 2533 19662 2536
rect 19604 2527 19662 2533
rect 20162 2524 20168 2536
rect 20220 2524 20226 2576
rect 20272 2564 20300 2604
rect 20717 2601 20729 2635
rect 20763 2632 20775 2635
rect 20806 2632 20812 2644
rect 20763 2604 20812 2632
rect 20763 2601 20775 2604
rect 20717 2595 20775 2601
rect 20806 2592 20812 2604
rect 20864 2592 20870 2644
rect 21818 2592 21824 2644
rect 21876 2632 21882 2644
rect 22557 2635 22615 2641
rect 22557 2632 22569 2635
rect 21876 2604 22569 2632
rect 21876 2592 21882 2604
rect 22557 2601 22569 2604
rect 22603 2601 22615 2635
rect 22557 2595 22615 2601
rect 21082 2564 21088 2576
rect 20272 2536 21088 2564
rect 21082 2524 21088 2536
rect 21140 2524 21146 2576
rect 21444 2567 21502 2573
rect 21444 2533 21456 2567
rect 21490 2564 21502 2567
rect 21634 2564 21640 2576
rect 21490 2536 21640 2564
rect 21490 2533 21502 2536
rect 21444 2527 21502 2533
rect 21634 2524 21640 2536
rect 21692 2524 21698 2576
rect 16684 2468 19012 2496
rect 16485 2459 16543 2465
rect 19058 2456 19064 2508
rect 19116 2496 19122 2508
rect 19337 2499 19395 2505
rect 19337 2496 19349 2499
rect 19116 2468 19349 2496
rect 19116 2456 19122 2468
rect 19337 2465 19349 2468
rect 19383 2465 19395 2499
rect 19337 2459 19395 2465
rect 20898 2456 20904 2508
rect 20956 2496 20962 2508
rect 21177 2499 21235 2505
rect 21177 2496 21189 2499
rect 20956 2468 21189 2496
rect 20956 2456 20962 2468
rect 21177 2465 21189 2468
rect 21223 2465 21235 2499
rect 21177 2459 21235 2465
rect 16025 2431 16083 2437
rect 16025 2397 16037 2431
rect 16071 2397 16083 2431
rect 18966 2428 18972 2440
rect 18927 2400 18972 2428
rect 16025 2391 16083 2397
rect 18966 2388 18972 2400
rect 19024 2388 19030 2440
rect 6178 2320 6184 2372
rect 6236 2360 6242 2372
rect 15473 2363 15531 2369
rect 15473 2360 15485 2363
rect 6236 2332 15485 2360
rect 6236 2320 6242 2332
rect 15473 2329 15485 2332
rect 15519 2329 15531 2363
rect 15473 2323 15531 2329
rect 9858 2252 9864 2304
rect 9916 2292 9922 2304
rect 14369 2295 14427 2301
rect 14369 2292 14381 2295
rect 9916 2264 14381 2292
rect 9916 2252 9922 2264
rect 14369 2261 14381 2264
rect 14415 2261 14427 2295
rect 14369 2255 14427 2261
rect 15194 2252 15200 2304
rect 15252 2292 15258 2304
rect 18325 2295 18383 2301
rect 18325 2292 18337 2295
rect 15252 2264 18337 2292
rect 15252 2252 15258 2264
rect 18325 2261 18337 2264
rect 18371 2261 18383 2295
rect 18325 2255 18383 2261
rect 1104 2202 23276 2224
rect 1104 2150 4680 2202
rect 4732 2150 4744 2202
rect 4796 2150 4808 2202
rect 4860 2150 4872 2202
rect 4924 2150 12078 2202
rect 12130 2150 12142 2202
rect 12194 2150 12206 2202
rect 12258 2150 12270 2202
rect 12322 2150 19475 2202
rect 19527 2150 19539 2202
rect 19591 2150 19603 2202
rect 19655 2150 19667 2202
rect 19719 2150 23276 2202
rect 1104 2128 23276 2150
rect 14826 2048 14832 2100
rect 14884 2088 14890 2100
rect 19978 2088 19984 2100
rect 14884 2060 19984 2088
rect 14884 2048 14890 2060
rect 19978 2048 19984 2060
rect 20036 2048 20042 2100
rect 15010 1980 15016 2032
rect 15068 2020 15074 2032
rect 21450 2020 21456 2032
rect 15068 1992 21456 2020
rect 15068 1980 15074 1992
rect 21450 1980 21456 1992
rect 21508 1980 21514 2032
rect 16850 1912 16856 1964
rect 16908 1952 16914 1964
rect 19886 1952 19892 1964
rect 16908 1924 19892 1952
rect 16908 1912 16914 1924
rect 19886 1912 19892 1924
rect 19944 1912 19950 1964
<< via1 >>
rect 8576 22856 8628 22908
rect 9496 22856 9548 22908
rect 15384 22856 15436 22908
rect 19432 22856 19484 22908
rect 17684 22584 17736 22636
rect 19340 22584 19392 22636
rect 18328 22312 18380 22364
rect 19800 22312 19852 22364
rect 9220 22108 9272 22160
rect 10968 22108 11020 22160
rect 7932 22040 7984 22092
rect 9404 22040 9456 22092
rect 9680 22040 9732 22092
rect 21640 22040 21692 22092
rect 8760 21972 8812 22024
rect 12716 21972 12768 22024
rect 16948 21972 17000 22024
rect 2044 21904 2096 21956
rect 10048 21904 10100 21956
rect 13452 21904 13504 21956
rect 19156 21904 19208 21956
rect 19616 21904 19668 21956
rect 6644 21836 6696 21888
rect 7748 21836 7800 21888
rect 8208 21836 8260 21888
rect 11612 21836 11664 21888
rect 14188 21836 14240 21888
rect 19800 21836 19852 21888
rect 20628 21836 20680 21888
rect 4680 21734 4732 21786
rect 4744 21734 4796 21786
rect 4808 21734 4860 21786
rect 4872 21734 4924 21786
rect 12078 21734 12130 21786
rect 12142 21734 12194 21786
rect 12206 21734 12258 21786
rect 12270 21734 12322 21786
rect 19475 21734 19527 21786
rect 19539 21734 19591 21786
rect 19603 21734 19655 21786
rect 19667 21734 19719 21786
rect 10048 21675 10100 21684
rect 10048 21641 10057 21675
rect 10057 21641 10091 21675
rect 10091 21641 10100 21675
rect 10048 21632 10100 21641
rect 3056 21496 3108 21548
rect 5632 21564 5684 21616
rect 8392 21564 8444 21616
rect 17592 21632 17644 21684
rect 18972 21632 19024 21684
rect 5264 21496 5316 21548
rect 6644 21496 6696 21548
rect 6736 21496 6788 21548
rect 7656 21496 7708 21548
rect 8668 21496 8720 21548
rect 11336 21564 11388 21616
rect 11428 21564 11480 21616
rect 11888 21564 11940 21616
rect 11520 21496 11572 21548
rect 11612 21539 11664 21548
rect 11612 21505 11621 21539
rect 11621 21505 11655 21539
rect 11655 21505 11664 21539
rect 11612 21496 11664 21505
rect 11980 21496 12032 21548
rect 14188 21539 14240 21548
rect 14188 21505 14197 21539
rect 14197 21505 14231 21539
rect 14231 21505 14240 21539
rect 14188 21496 14240 21505
rect 2872 21428 2924 21480
rect 1584 21360 1636 21412
rect 1400 21292 1452 21344
rect 2228 21335 2280 21344
rect 2228 21301 2237 21335
rect 2237 21301 2271 21335
rect 2271 21301 2280 21335
rect 2228 21292 2280 21301
rect 6092 21471 6144 21480
rect 6092 21437 6101 21471
rect 6101 21437 6135 21471
rect 6135 21437 6144 21471
rect 6092 21428 6144 21437
rect 6276 21428 6328 21480
rect 8392 21471 8444 21480
rect 8392 21437 8401 21471
rect 8401 21437 8435 21471
rect 8435 21437 8444 21471
rect 8392 21428 8444 21437
rect 8944 21471 8996 21480
rect 8944 21437 8953 21471
rect 8953 21437 8987 21471
rect 8987 21437 8996 21471
rect 8944 21428 8996 21437
rect 9036 21428 9088 21480
rect 14648 21428 14700 21480
rect 15108 21428 15160 21480
rect 16212 21496 16264 21548
rect 16764 21428 16816 21480
rect 16856 21428 16908 21480
rect 3148 21335 3200 21344
rect 3148 21301 3157 21335
rect 3157 21301 3191 21335
rect 3191 21301 3200 21335
rect 3148 21292 3200 21301
rect 3240 21335 3292 21344
rect 3240 21301 3249 21335
rect 3249 21301 3283 21335
rect 3283 21301 3292 21335
rect 3240 21292 3292 21301
rect 4344 21292 4396 21344
rect 4528 21335 4580 21344
rect 4528 21301 4537 21335
rect 4537 21301 4571 21335
rect 4571 21301 4580 21335
rect 4528 21292 4580 21301
rect 5540 21292 5592 21344
rect 12532 21360 12584 21412
rect 6920 21292 6972 21344
rect 7380 21335 7432 21344
rect 7380 21301 7389 21335
rect 7389 21301 7423 21335
rect 7423 21301 7432 21335
rect 7380 21292 7432 21301
rect 9772 21292 9824 21344
rect 11244 21292 11296 21344
rect 11428 21335 11480 21344
rect 11428 21301 11437 21335
rect 11437 21301 11471 21335
rect 11471 21301 11480 21335
rect 11428 21292 11480 21301
rect 11612 21292 11664 21344
rect 12072 21335 12124 21344
rect 12072 21301 12081 21335
rect 12081 21301 12115 21335
rect 12115 21301 12124 21335
rect 12072 21292 12124 21301
rect 14464 21360 14516 21412
rect 20536 21564 20588 21616
rect 20628 21564 20680 21616
rect 24032 21632 24084 21684
rect 21640 21564 21692 21616
rect 19340 21496 19392 21548
rect 19892 21496 19944 21548
rect 22008 21496 22060 21548
rect 22928 21496 22980 21548
rect 17408 21428 17460 21480
rect 18236 21428 18288 21480
rect 20352 21428 20404 21480
rect 21272 21428 21324 21480
rect 19156 21403 19208 21412
rect 19156 21369 19165 21403
rect 19165 21369 19199 21403
rect 19199 21369 19208 21403
rect 19156 21360 19208 21369
rect 12992 21335 13044 21344
rect 12992 21301 13001 21335
rect 13001 21301 13035 21335
rect 13035 21301 13044 21335
rect 12992 21292 13044 21301
rect 13084 21335 13136 21344
rect 13084 21301 13093 21335
rect 13093 21301 13127 21335
rect 13127 21301 13136 21335
rect 13084 21292 13136 21301
rect 13820 21292 13872 21344
rect 14004 21335 14056 21344
rect 14004 21301 14013 21335
rect 14013 21301 14047 21335
rect 14047 21301 14056 21335
rect 14004 21292 14056 21301
rect 15476 21335 15528 21344
rect 15476 21301 15485 21335
rect 15485 21301 15519 21335
rect 15519 21301 15528 21335
rect 15476 21292 15528 21301
rect 16488 21335 16540 21344
rect 16488 21301 16497 21335
rect 16497 21301 16531 21335
rect 16531 21301 16540 21335
rect 16488 21292 16540 21301
rect 17776 21292 17828 21344
rect 18052 21292 18104 21344
rect 19432 21292 19484 21344
rect 19800 21292 19852 21344
rect 20076 21335 20128 21344
rect 20076 21301 20085 21335
rect 20085 21301 20119 21335
rect 20119 21301 20128 21335
rect 20076 21292 20128 21301
rect 20628 21335 20680 21344
rect 20628 21301 20637 21335
rect 20637 21301 20671 21335
rect 20671 21301 20680 21335
rect 20628 21292 20680 21301
rect 21180 21335 21232 21344
rect 21180 21301 21189 21335
rect 21189 21301 21223 21335
rect 21223 21301 21232 21335
rect 21180 21292 21232 21301
rect 21732 21292 21784 21344
rect 23204 21292 23256 21344
rect 8379 21190 8431 21242
rect 8443 21190 8495 21242
rect 8507 21190 8559 21242
rect 8571 21190 8623 21242
rect 15776 21190 15828 21242
rect 15840 21190 15892 21242
rect 15904 21190 15956 21242
rect 15968 21190 16020 21242
rect 296 21088 348 21140
rect 3148 21088 3200 21140
rect 3516 21131 3568 21140
rect 3516 21097 3525 21131
rect 3525 21097 3559 21131
rect 3559 21097 3568 21131
rect 3516 21088 3568 21097
rect 5172 21020 5224 21072
rect 5540 21088 5592 21140
rect 7840 21088 7892 21140
rect 6736 21020 6788 21072
rect 7196 21020 7248 21072
rect 7380 21020 7432 21072
rect 7472 21020 7524 21072
rect 12072 21088 12124 21140
rect 13360 21088 13412 21140
rect 14464 21131 14516 21140
rect 2044 20952 2096 21004
rect 3240 20952 3292 21004
rect 4344 20995 4396 21004
rect 4344 20961 4378 20995
rect 4378 20961 4396 20995
rect 4344 20952 4396 20961
rect 6552 20952 6604 21004
rect 8024 20952 8076 21004
rect 3332 20884 3384 20936
rect 5080 20884 5132 20936
rect 6460 20884 6512 20936
rect 7840 20884 7892 20936
rect 9036 20927 9088 20936
rect 5264 20816 5316 20868
rect 5448 20816 5500 20868
rect 2780 20748 2832 20800
rect 4436 20748 4488 20800
rect 5816 20748 5868 20800
rect 8668 20816 8720 20868
rect 9036 20893 9045 20927
rect 9045 20893 9079 20927
rect 9079 20893 9088 20927
rect 9036 20884 9088 20893
rect 10232 20952 10284 21004
rect 11520 21020 11572 21072
rect 12532 21020 12584 21072
rect 11980 20952 12032 21004
rect 14096 20952 14148 21004
rect 9588 20816 9640 20868
rect 8576 20791 8628 20800
rect 8576 20757 8585 20791
rect 8585 20757 8619 20791
rect 8619 20757 8628 20791
rect 8576 20748 8628 20757
rect 8852 20748 8904 20800
rect 9956 20748 10008 20800
rect 12440 20816 12492 20868
rect 12900 20816 12952 20868
rect 14464 21097 14473 21131
rect 14473 21097 14507 21131
rect 14507 21097 14516 21131
rect 14464 21088 14516 21097
rect 14648 21088 14700 21140
rect 15200 21088 15252 21140
rect 15476 21088 15528 21140
rect 20076 21088 20128 21140
rect 20628 21088 20680 21140
rect 15568 21063 15620 21072
rect 15568 21029 15602 21063
rect 15602 21029 15620 21063
rect 15568 21020 15620 21029
rect 18788 21020 18840 21072
rect 14372 20884 14424 20936
rect 19892 20952 19944 21004
rect 20260 21020 20312 21072
rect 20352 21020 20404 21072
rect 17408 20927 17460 20936
rect 17408 20893 17417 20927
rect 17417 20893 17451 20927
rect 17451 20893 17460 20927
rect 17408 20884 17460 20893
rect 17592 20927 17644 20936
rect 17592 20893 17601 20927
rect 17601 20893 17635 20927
rect 17635 20893 17644 20927
rect 17592 20884 17644 20893
rect 17960 20884 18012 20936
rect 22468 20952 22520 21004
rect 22652 20995 22704 21004
rect 22652 20961 22661 20995
rect 22661 20961 22695 20995
rect 22695 20961 22704 20995
rect 22652 20952 22704 20961
rect 21364 20927 21416 20936
rect 11060 20791 11112 20800
rect 11060 20757 11069 20791
rect 11069 20757 11103 20791
rect 11103 20757 11112 20791
rect 11060 20748 11112 20757
rect 11244 20748 11296 20800
rect 11980 20748 12032 20800
rect 12532 20748 12584 20800
rect 19156 20816 19208 20868
rect 21364 20893 21373 20927
rect 21373 20893 21407 20927
rect 21407 20893 21416 20927
rect 21364 20884 21416 20893
rect 21088 20816 21140 20868
rect 23020 20884 23072 20936
rect 14372 20748 14424 20800
rect 15476 20748 15528 20800
rect 16488 20748 16540 20800
rect 16580 20748 16632 20800
rect 19800 20748 19852 20800
rect 20904 20791 20956 20800
rect 20904 20757 20913 20791
rect 20913 20757 20947 20791
rect 20947 20757 20956 20791
rect 20904 20748 20956 20757
rect 21180 20748 21232 20800
rect 22836 20791 22888 20800
rect 22836 20757 22845 20791
rect 22845 20757 22879 20791
rect 22879 20757 22888 20791
rect 22836 20748 22888 20757
rect 4680 20646 4732 20698
rect 4744 20646 4796 20698
rect 4808 20646 4860 20698
rect 4872 20646 4924 20698
rect 12078 20646 12130 20698
rect 12142 20646 12194 20698
rect 12206 20646 12258 20698
rect 12270 20646 12322 20698
rect 19475 20646 19527 20698
rect 19539 20646 19591 20698
rect 19603 20646 19655 20698
rect 19667 20646 19719 20698
rect 848 20544 900 20596
rect 3056 20544 3108 20596
rect 3240 20544 3292 20596
rect 4344 20544 4396 20596
rect 5264 20544 5316 20596
rect 2780 20340 2832 20392
rect 3332 20340 3384 20392
rect 3516 20340 3568 20392
rect 3976 20340 4028 20392
rect 6000 20476 6052 20528
rect 5724 20451 5776 20460
rect 5724 20417 5733 20451
rect 5733 20417 5767 20451
rect 5767 20417 5776 20451
rect 5724 20408 5776 20417
rect 8116 20544 8168 20596
rect 8576 20544 8628 20596
rect 10232 20587 10284 20596
rect 10232 20553 10241 20587
rect 10241 20553 10275 20587
rect 10275 20553 10284 20587
rect 10232 20544 10284 20553
rect 11520 20544 11572 20596
rect 14096 20587 14148 20596
rect 12440 20476 12492 20528
rect 14096 20553 14105 20587
rect 14105 20553 14139 20587
rect 14139 20553 14148 20587
rect 14096 20544 14148 20553
rect 15108 20544 15160 20596
rect 6460 20340 6512 20392
rect 8852 20383 8904 20392
rect 8852 20349 8861 20383
rect 8861 20349 8895 20383
rect 8895 20349 8904 20383
rect 8852 20340 8904 20349
rect 9956 20408 10008 20460
rect 10232 20408 10284 20460
rect 10416 20340 10468 20392
rect 2964 20272 3016 20324
rect 4160 20272 4212 20324
rect 7104 20315 7156 20324
rect 2136 20204 2188 20256
rect 3608 20204 3660 20256
rect 4344 20204 4396 20256
rect 5448 20247 5500 20256
rect 5448 20213 5457 20247
rect 5457 20213 5491 20247
rect 5491 20213 5500 20247
rect 5448 20204 5500 20213
rect 5632 20204 5684 20256
rect 7104 20281 7138 20315
rect 7138 20281 7156 20315
rect 7104 20272 7156 20281
rect 9312 20272 9364 20324
rect 9496 20272 9548 20324
rect 12440 20340 12492 20392
rect 11060 20272 11112 20324
rect 11704 20272 11756 20324
rect 11980 20272 12032 20324
rect 13912 20340 13964 20392
rect 14004 20272 14056 20324
rect 14372 20451 14424 20460
rect 14372 20417 14381 20451
rect 14381 20417 14415 20451
rect 14415 20417 14424 20451
rect 14372 20408 14424 20417
rect 14464 20340 14516 20392
rect 14924 20340 14976 20392
rect 19340 20544 19392 20596
rect 19892 20544 19944 20596
rect 20352 20544 20404 20596
rect 21364 20544 21416 20596
rect 20904 20476 20956 20528
rect 23388 20476 23440 20528
rect 20720 20408 20772 20460
rect 16120 20340 16172 20392
rect 17960 20340 18012 20392
rect 18144 20340 18196 20392
rect 19156 20340 19208 20392
rect 19708 20383 19760 20392
rect 19708 20349 19717 20383
rect 19717 20349 19751 20383
rect 19751 20349 19760 20383
rect 19708 20340 19760 20349
rect 19800 20340 19852 20392
rect 9864 20204 9916 20256
rect 11152 20204 11204 20256
rect 11612 20204 11664 20256
rect 15568 20204 15620 20256
rect 16580 20272 16632 20324
rect 19892 20272 19944 20324
rect 20076 20272 20128 20324
rect 21916 20272 21968 20324
rect 16764 20204 16816 20256
rect 20720 20204 20772 20256
rect 21088 20247 21140 20256
rect 21088 20213 21097 20247
rect 21097 20213 21131 20247
rect 21131 20213 21140 20247
rect 21088 20204 21140 20213
rect 21548 20247 21600 20256
rect 21548 20213 21557 20247
rect 21557 20213 21591 20247
rect 21591 20213 21600 20247
rect 21548 20204 21600 20213
rect 22376 20247 22428 20256
rect 22376 20213 22385 20247
rect 22385 20213 22419 20247
rect 22419 20213 22428 20247
rect 22376 20204 22428 20213
rect 8379 20102 8431 20154
rect 8443 20102 8495 20154
rect 8507 20102 8559 20154
rect 8571 20102 8623 20154
rect 15776 20102 15828 20154
rect 15840 20102 15892 20154
rect 15904 20102 15956 20154
rect 15968 20102 16020 20154
rect 2964 20043 3016 20052
rect 2964 20009 2973 20043
rect 2973 20009 3007 20043
rect 3007 20009 3016 20043
rect 2964 20000 3016 20009
rect 3056 20000 3108 20052
rect 4528 20000 4580 20052
rect 1860 19975 1912 19984
rect 1860 19941 1894 19975
rect 1894 19941 1912 19975
rect 1860 19932 1912 19941
rect 4620 19932 4672 19984
rect 6460 20000 6512 20052
rect 5816 19932 5868 19984
rect 1676 19864 1728 19916
rect 3424 19864 3476 19916
rect 4252 19864 4304 19916
rect 4804 19864 4856 19916
rect 3884 19796 3936 19848
rect 4068 19728 4120 19780
rect 6368 19864 6420 19916
rect 8668 20000 8720 20052
rect 9680 20000 9732 20052
rect 9864 20043 9916 20052
rect 9864 20009 9873 20043
rect 9873 20009 9907 20043
rect 9907 20009 9916 20043
rect 9864 20000 9916 20009
rect 10600 20000 10652 20052
rect 14004 20000 14056 20052
rect 18144 20000 18196 20052
rect 18236 20000 18288 20052
rect 20812 20000 20864 20052
rect 21456 20000 21508 20052
rect 7472 19975 7524 19984
rect 7472 19941 7506 19975
rect 7506 19941 7524 19975
rect 7472 19932 7524 19941
rect 7748 19932 7800 19984
rect 7012 19864 7064 19916
rect 7840 19864 7892 19916
rect 9220 19864 9272 19916
rect 9680 19907 9732 19916
rect 9680 19873 9689 19907
rect 9689 19873 9723 19907
rect 9723 19873 9732 19907
rect 9680 19864 9732 19873
rect 12716 19932 12768 19984
rect 12900 19932 12952 19984
rect 13176 19932 13228 19984
rect 14648 19932 14700 19984
rect 15568 19932 15620 19984
rect 16764 19975 16816 19984
rect 16764 19941 16798 19975
rect 16798 19941 16816 19975
rect 10416 19728 10468 19780
rect 11428 19796 11480 19848
rect 14004 19796 14056 19848
rect 15016 19864 15068 19916
rect 16764 19932 16816 19941
rect 17960 19932 18012 19984
rect 18604 19932 18656 19984
rect 21088 19932 21140 19984
rect 16028 19864 16080 19916
rect 21456 19907 21508 19916
rect 16120 19796 16172 19848
rect 18236 19796 18288 19848
rect 18696 19839 18748 19848
rect 18696 19805 18705 19839
rect 18705 19805 18739 19839
rect 18739 19805 18748 19839
rect 18696 19796 18748 19805
rect 16212 19728 16264 19780
rect 17500 19728 17552 19780
rect 21456 19873 21490 19907
rect 21490 19873 21508 19907
rect 21456 19864 21508 19873
rect 21824 19864 21876 19916
rect 7104 19660 7156 19712
rect 8116 19660 8168 19712
rect 8300 19660 8352 19712
rect 8760 19660 8812 19712
rect 10232 19703 10284 19712
rect 10232 19669 10241 19703
rect 10241 19669 10275 19703
rect 10275 19669 10284 19703
rect 10232 19660 10284 19669
rect 11060 19660 11112 19712
rect 14464 19660 14516 19712
rect 17408 19660 17460 19712
rect 17776 19660 17828 19712
rect 18420 19660 18472 19712
rect 18880 19660 18932 19712
rect 20536 19796 20588 19848
rect 20996 19796 21048 19848
rect 19800 19660 19852 19712
rect 22560 19703 22612 19712
rect 22560 19669 22569 19703
rect 22569 19669 22603 19703
rect 22603 19669 22612 19703
rect 22560 19660 22612 19669
rect 22836 19703 22888 19712
rect 22836 19669 22845 19703
rect 22845 19669 22879 19703
rect 22879 19669 22888 19703
rect 22836 19660 22888 19669
rect 4680 19558 4732 19610
rect 4744 19558 4796 19610
rect 4808 19558 4860 19610
rect 4872 19558 4924 19610
rect 12078 19558 12130 19610
rect 12142 19558 12194 19610
rect 12206 19558 12258 19610
rect 12270 19558 12322 19610
rect 19475 19558 19527 19610
rect 19539 19558 19591 19610
rect 19603 19558 19655 19610
rect 19667 19558 19719 19610
rect 4160 19456 4212 19508
rect 4988 19456 5040 19508
rect 1492 19388 1544 19440
rect 3056 19388 3108 19440
rect 3884 19388 3936 19440
rect 3148 19363 3200 19372
rect 3148 19329 3157 19363
rect 3157 19329 3191 19363
rect 3191 19329 3200 19363
rect 3148 19320 3200 19329
rect 3332 19320 3384 19372
rect 4620 19388 4672 19440
rect 2228 19252 2280 19304
rect 4528 19320 4580 19372
rect 3148 19184 3200 19236
rect 1584 19159 1636 19168
rect 1584 19125 1593 19159
rect 1593 19125 1627 19159
rect 1627 19125 1636 19159
rect 1584 19116 1636 19125
rect 1952 19159 2004 19168
rect 1952 19125 1961 19159
rect 1961 19125 1995 19159
rect 1995 19125 2004 19159
rect 1952 19116 2004 19125
rect 2872 19116 2924 19168
rect 3516 19116 3568 19168
rect 5172 19252 5224 19304
rect 3884 19184 3936 19236
rect 6276 19295 6328 19304
rect 6276 19261 6285 19295
rect 6285 19261 6319 19295
rect 6319 19261 6328 19295
rect 6276 19252 6328 19261
rect 13176 19456 13228 19508
rect 9128 19388 9180 19440
rect 9404 19388 9456 19440
rect 7748 19320 7800 19372
rect 7932 19320 7984 19372
rect 11796 19388 11848 19440
rect 14096 19456 14148 19508
rect 14188 19456 14240 19508
rect 13728 19388 13780 19440
rect 14556 19388 14608 19440
rect 4068 19159 4120 19168
rect 4068 19125 4077 19159
rect 4077 19125 4111 19159
rect 4111 19125 4120 19159
rect 4068 19116 4120 19125
rect 5816 19116 5868 19168
rect 7104 19116 7156 19168
rect 7656 19252 7708 19304
rect 8208 19252 8260 19304
rect 9128 19252 9180 19304
rect 9036 19184 9088 19236
rect 9680 19252 9732 19304
rect 9588 19116 9640 19168
rect 11704 19320 11756 19372
rect 10324 19252 10376 19304
rect 10508 19252 10560 19304
rect 12532 19252 12584 19304
rect 15660 19388 15712 19440
rect 16580 19456 16632 19508
rect 20076 19499 20128 19508
rect 17500 19388 17552 19440
rect 20076 19465 20085 19499
rect 20085 19465 20119 19499
rect 20119 19465 20128 19499
rect 20076 19456 20128 19465
rect 21640 19456 21692 19508
rect 22100 19456 22152 19508
rect 15200 19320 15252 19372
rect 16212 19320 16264 19372
rect 17592 19320 17644 19372
rect 18512 19363 18564 19372
rect 18512 19329 18524 19363
rect 18524 19329 18558 19363
rect 18558 19329 18564 19363
rect 18512 19320 18564 19329
rect 18788 19320 18840 19372
rect 19800 19320 19852 19372
rect 11060 19184 11112 19236
rect 11336 19184 11388 19236
rect 9864 19116 9916 19168
rect 11704 19116 11756 19168
rect 11980 19116 12032 19168
rect 12716 19116 12768 19168
rect 12992 19116 13044 19168
rect 13084 19116 13136 19168
rect 13544 19116 13596 19168
rect 17960 19252 18012 19304
rect 14832 19159 14884 19168
rect 14832 19125 14841 19159
rect 14841 19125 14875 19159
rect 14875 19125 14884 19159
rect 14832 19116 14884 19125
rect 15292 19116 15344 19168
rect 15568 19116 15620 19168
rect 16120 19116 16172 19168
rect 16212 19116 16264 19168
rect 18144 19116 18196 19168
rect 18788 19116 18840 19168
rect 19064 19116 19116 19168
rect 21640 19184 21692 19236
rect 20076 19116 20128 19168
rect 20352 19116 20404 19168
rect 20904 19116 20956 19168
rect 22192 19116 22244 19168
rect 8379 19014 8431 19066
rect 8443 19014 8495 19066
rect 8507 19014 8559 19066
rect 8571 19014 8623 19066
rect 15776 19014 15828 19066
rect 15840 19014 15892 19066
rect 15904 19014 15956 19066
rect 15968 19014 16020 19066
rect 2780 18912 2832 18964
rect 3056 18912 3108 18964
rect 3516 18912 3568 18964
rect 3700 18912 3752 18964
rect 5448 18912 5500 18964
rect 5632 18912 5684 18964
rect 14004 18955 14056 18964
rect 1952 18844 2004 18896
rect 1676 18776 1728 18828
rect 3056 18776 3108 18828
rect 5264 18844 5316 18896
rect 3516 18776 3568 18828
rect 6092 18776 6144 18828
rect 7656 18844 7708 18896
rect 8024 18844 8076 18896
rect 6460 18776 6512 18828
rect 3424 18708 3476 18760
rect 4620 18708 4672 18760
rect 5816 18751 5868 18760
rect 5816 18717 5825 18751
rect 5825 18717 5859 18751
rect 5859 18717 5868 18751
rect 7380 18776 7432 18828
rect 7472 18776 7524 18828
rect 5816 18708 5868 18717
rect 7932 18708 7984 18760
rect 9496 18708 9548 18760
rect 6368 18615 6420 18624
rect 6368 18581 6377 18615
rect 6377 18581 6411 18615
rect 6411 18581 6420 18615
rect 6368 18572 6420 18581
rect 8760 18640 8812 18692
rect 8208 18615 8260 18624
rect 8208 18581 8217 18615
rect 8217 18581 8251 18615
rect 8251 18581 8260 18615
rect 8484 18615 8536 18624
rect 8208 18572 8260 18581
rect 8484 18581 8493 18615
rect 8493 18581 8527 18615
rect 8527 18581 8536 18615
rect 8484 18572 8536 18581
rect 11704 18844 11756 18896
rect 13544 18844 13596 18896
rect 14004 18921 14013 18955
rect 14013 18921 14047 18955
rect 14047 18921 14056 18955
rect 14004 18912 14056 18921
rect 14372 18912 14424 18964
rect 16120 18912 16172 18964
rect 18144 18912 18196 18964
rect 19984 18912 20036 18964
rect 20168 18912 20220 18964
rect 21180 18912 21232 18964
rect 21732 18912 21784 18964
rect 14280 18844 14332 18896
rect 9680 18819 9732 18828
rect 9680 18785 9689 18819
rect 9689 18785 9723 18819
rect 9723 18785 9732 18819
rect 9680 18776 9732 18785
rect 10324 18776 10376 18828
rect 11060 18776 11112 18828
rect 11152 18776 11204 18828
rect 10048 18708 10100 18760
rect 10140 18751 10192 18760
rect 10140 18717 10152 18751
rect 10152 18717 10186 18751
rect 10186 18717 10192 18751
rect 12716 18776 12768 18828
rect 15568 18844 15620 18896
rect 20536 18844 20588 18896
rect 15108 18776 15160 18828
rect 10140 18708 10192 18717
rect 11704 18640 11756 18692
rect 12072 18640 12124 18692
rect 11796 18572 11848 18624
rect 16488 18776 16540 18828
rect 16580 18776 16632 18828
rect 16856 18776 16908 18828
rect 17500 18776 17552 18828
rect 17960 18819 18012 18828
rect 17960 18785 17994 18819
rect 17994 18785 18012 18819
rect 17960 18776 18012 18785
rect 18328 18776 18380 18828
rect 18512 18776 18564 18828
rect 19800 18776 19852 18828
rect 19892 18776 19944 18828
rect 21180 18776 21232 18828
rect 15752 18751 15804 18760
rect 12900 18572 12952 18624
rect 15752 18717 15761 18751
rect 15761 18717 15795 18751
rect 15795 18717 15804 18751
rect 15752 18708 15804 18717
rect 19248 18708 19300 18760
rect 18696 18640 18748 18692
rect 17040 18572 17092 18624
rect 17132 18615 17184 18624
rect 17132 18581 17141 18615
rect 17141 18581 17175 18615
rect 17175 18581 17184 18615
rect 17408 18615 17460 18624
rect 17132 18572 17184 18581
rect 17408 18581 17417 18615
rect 17417 18581 17451 18615
rect 17451 18581 17460 18615
rect 17408 18572 17460 18581
rect 18604 18572 18656 18624
rect 19156 18615 19208 18624
rect 19156 18581 19165 18615
rect 19165 18581 19199 18615
rect 19199 18581 19208 18615
rect 20168 18615 20220 18624
rect 19156 18572 19208 18581
rect 20168 18581 20177 18615
rect 20177 18581 20211 18615
rect 20211 18581 20220 18615
rect 20812 18708 20864 18760
rect 20996 18640 21048 18692
rect 22008 18708 22060 18760
rect 21364 18615 21416 18624
rect 20168 18572 20220 18581
rect 21364 18581 21373 18615
rect 21373 18581 21407 18615
rect 21407 18581 21416 18615
rect 21364 18572 21416 18581
rect 22100 18572 22152 18624
rect 4680 18470 4732 18522
rect 4744 18470 4796 18522
rect 4808 18470 4860 18522
rect 4872 18470 4924 18522
rect 12078 18470 12130 18522
rect 12142 18470 12194 18522
rect 12206 18470 12258 18522
rect 12270 18470 12322 18522
rect 19475 18470 19527 18522
rect 19539 18470 19591 18522
rect 19603 18470 19655 18522
rect 19667 18470 19719 18522
rect 3056 18411 3108 18420
rect 3056 18377 3065 18411
rect 3065 18377 3099 18411
rect 3099 18377 3108 18411
rect 3056 18368 3108 18377
rect 8852 18368 8904 18420
rect 9128 18411 9180 18420
rect 9128 18377 9137 18411
rect 9137 18377 9171 18411
rect 9171 18377 9180 18411
rect 9128 18368 9180 18377
rect 11520 18368 11572 18420
rect 15568 18368 15620 18420
rect 4988 18300 5040 18352
rect 6552 18300 6604 18352
rect 5816 18275 5868 18284
rect 5816 18241 5825 18275
rect 5825 18241 5859 18275
rect 5859 18241 5868 18275
rect 5816 18232 5868 18241
rect 7104 18232 7156 18284
rect 7656 18232 7708 18284
rect 12900 18300 12952 18352
rect 18788 18368 18840 18420
rect 18880 18368 18932 18420
rect 19248 18368 19300 18420
rect 20352 18368 20404 18420
rect 1768 18164 1820 18216
rect 3332 18207 3384 18216
rect 3332 18173 3341 18207
rect 3341 18173 3375 18207
rect 3375 18173 3384 18207
rect 3332 18164 3384 18173
rect 4068 18164 4120 18216
rect 4528 18164 4580 18216
rect 6920 18164 6972 18216
rect 8024 18207 8076 18216
rect 8024 18173 8033 18207
rect 8033 18173 8067 18207
rect 8067 18173 8076 18207
rect 8024 18164 8076 18173
rect 8116 18164 8168 18216
rect 3148 18096 3200 18148
rect 5172 18096 5224 18148
rect 5724 18139 5776 18148
rect 5724 18105 5733 18139
rect 5733 18105 5767 18139
rect 5767 18105 5776 18139
rect 5724 18096 5776 18105
rect 9680 18164 9732 18216
rect 9772 18207 9824 18216
rect 9772 18173 9781 18207
rect 9781 18173 9815 18207
rect 9815 18173 9824 18207
rect 9772 18164 9824 18173
rect 14924 18232 14976 18284
rect 15200 18275 15252 18284
rect 15200 18241 15209 18275
rect 15209 18241 15243 18275
rect 15243 18241 15252 18275
rect 15200 18232 15252 18241
rect 10508 18207 10560 18216
rect 10508 18173 10517 18207
rect 10517 18173 10551 18207
rect 10551 18173 10560 18207
rect 10508 18164 10560 18173
rect 3884 18028 3936 18080
rect 5632 18071 5684 18080
rect 5632 18037 5641 18071
rect 5641 18037 5675 18071
rect 5675 18037 5684 18071
rect 5632 18028 5684 18037
rect 7104 18028 7156 18080
rect 10048 18096 10100 18148
rect 11244 18096 11296 18148
rect 12808 18164 12860 18216
rect 14372 18164 14424 18216
rect 16028 18232 16080 18284
rect 17868 18232 17920 18284
rect 18052 18275 18104 18284
rect 18052 18241 18061 18275
rect 18061 18241 18095 18275
rect 18095 18241 18104 18275
rect 18052 18232 18104 18241
rect 19524 18300 19576 18352
rect 15568 18096 15620 18148
rect 11888 18028 11940 18080
rect 12440 18071 12492 18080
rect 12440 18037 12449 18071
rect 12449 18037 12483 18071
rect 12483 18037 12492 18071
rect 12440 18028 12492 18037
rect 12808 18028 12860 18080
rect 16488 18164 16540 18216
rect 18512 18207 18564 18216
rect 18512 18173 18521 18207
rect 18521 18173 18555 18207
rect 18555 18173 18564 18207
rect 18512 18164 18564 18173
rect 21916 18232 21968 18284
rect 20076 18164 20128 18216
rect 20904 18164 20956 18216
rect 17408 18096 17460 18148
rect 18052 18096 18104 18148
rect 19156 18096 19208 18148
rect 19248 18028 19300 18080
rect 20352 18096 20404 18148
rect 21640 18028 21692 18080
rect 22008 18028 22060 18080
rect 22284 18071 22336 18080
rect 22284 18037 22293 18071
rect 22293 18037 22327 18071
rect 22327 18037 22336 18071
rect 22284 18028 22336 18037
rect 22376 18071 22428 18080
rect 22376 18037 22385 18071
rect 22385 18037 22419 18071
rect 22419 18037 22428 18071
rect 22376 18028 22428 18037
rect 8379 17926 8431 17978
rect 8443 17926 8495 17978
rect 8507 17926 8559 17978
rect 8571 17926 8623 17978
rect 15776 17926 15828 17978
rect 15840 17926 15892 17978
rect 15904 17926 15956 17978
rect 15968 17926 16020 17978
rect 3148 17867 3200 17876
rect 3148 17833 3157 17867
rect 3157 17833 3191 17867
rect 3191 17833 3200 17867
rect 3148 17824 3200 17833
rect 3608 17867 3660 17876
rect 3608 17833 3617 17867
rect 3617 17833 3651 17867
rect 3651 17833 3660 17867
rect 3608 17824 3660 17833
rect 4252 17867 4304 17876
rect 4252 17833 4261 17867
rect 4261 17833 4295 17867
rect 4295 17833 4304 17867
rect 4252 17824 4304 17833
rect 5264 17824 5316 17876
rect 7472 17824 7524 17876
rect 7564 17824 7616 17876
rect 8852 17867 8904 17876
rect 8852 17833 8861 17867
rect 8861 17833 8895 17867
rect 8895 17833 8904 17867
rect 8852 17824 8904 17833
rect 10508 17824 10560 17876
rect 10600 17824 10652 17876
rect 11428 17867 11480 17876
rect 3884 17756 3936 17808
rect 8760 17799 8812 17808
rect 8760 17765 8769 17799
rect 8769 17765 8803 17799
rect 8803 17765 8812 17799
rect 8760 17756 8812 17765
rect 1860 17688 1912 17740
rect 3792 17688 3844 17740
rect 4896 17688 4948 17740
rect 3332 17620 3384 17672
rect 1768 17484 1820 17536
rect 5264 17484 5316 17536
rect 5724 17484 5776 17536
rect 8116 17688 8168 17740
rect 6644 17620 6696 17672
rect 7748 17620 7800 17672
rect 9864 17756 9916 17808
rect 9128 17688 9180 17740
rect 11152 17756 11204 17808
rect 11428 17833 11437 17867
rect 11437 17833 11471 17867
rect 11471 17833 11480 17867
rect 11428 17824 11480 17833
rect 12440 17824 12492 17876
rect 14188 17824 14240 17876
rect 14372 17867 14424 17876
rect 14372 17833 14381 17867
rect 14381 17833 14415 17867
rect 14415 17833 14424 17867
rect 14372 17824 14424 17833
rect 15384 17824 15436 17876
rect 14924 17756 14976 17808
rect 15200 17756 15252 17808
rect 15292 17756 15344 17808
rect 11060 17688 11112 17740
rect 8944 17620 8996 17672
rect 9312 17620 9364 17672
rect 9496 17620 9548 17672
rect 11980 17663 12032 17672
rect 8392 17527 8444 17536
rect 8392 17493 8401 17527
rect 8401 17493 8435 17527
rect 8435 17493 8444 17527
rect 8392 17484 8444 17493
rect 11980 17629 11989 17663
rect 11989 17629 12023 17663
rect 12023 17629 12032 17663
rect 11980 17620 12032 17629
rect 12532 17688 12584 17740
rect 13084 17688 13136 17740
rect 13820 17688 13872 17740
rect 14648 17731 14700 17740
rect 14648 17697 14657 17731
rect 14657 17697 14691 17731
rect 14691 17697 14700 17731
rect 14648 17688 14700 17697
rect 14832 17688 14884 17740
rect 17040 17824 17092 17876
rect 19340 17824 19392 17876
rect 20260 17867 20312 17876
rect 20260 17833 20269 17867
rect 20269 17833 20303 17867
rect 20303 17833 20312 17867
rect 20260 17824 20312 17833
rect 21456 17824 21508 17876
rect 16764 17756 16816 17808
rect 16856 17688 16908 17740
rect 17040 17688 17092 17740
rect 17316 17731 17368 17740
rect 17316 17697 17325 17731
rect 17325 17697 17359 17731
rect 17359 17697 17368 17731
rect 17316 17688 17368 17697
rect 18604 17756 18656 17808
rect 18788 17756 18840 17808
rect 19064 17756 19116 17808
rect 20996 17756 21048 17808
rect 21088 17756 21140 17808
rect 22192 17756 22244 17808
rect 12532 17552 12584 17604
rect 12716 17552 12768 17604
rect 12900 17552 12952 17604
rect 15108 17620 15160 17672
rect 16396 17620 16448 17672
rect 17592 17663 17644 17672
rect 17592 17629 17601 17663
rect 17601 17629 17635 17663
rect 17635 17629 17644 17663
rect 17592 17620 17644 17629
rect 18052 17620 18104 17672
rect 19248 17620 19300 17672
rect 20536 17620 20588 17672
rect 20904 17663 20956 17672
rect 20904 17629 20913 17663
rect 20913 17629 20947 17663
rect 20947 17629 20956 17663
rect 20904 17620 20956 17629
rect 22836 17620 22888 17672
rect 11244 17484 11296 17536
rect 13728 17484 13780 17536
rect 17408 17484 17460 17536
rect 19156 17484 19208 17536
rect 20168 17484 20220 17536
rect 22744 17484 22796 17536
rect 4680 17382 4732 17434
rect 4744 17382 4796 17434
rect 4808 17382 4860 17434
rect 4872 17382 4924 17434
rect 12078 17382 12130 17434
rect 12142 17382 12194 17434
rect 12206 17382 12258 17434
rect 12270 17382 12322 17434
rect 19475 17382 19527 17434
rect 19539 17382 19591 17434
rect 19603 17382 19655 17434
rect 19667 17382 19719 17434
rect 8392 17280 8444 17332
rect 9404 17323 9456 17332
rect 9404 17289 9413 17323
rect 9413 17289 9447 17323
rect 9447 17289 9456 17323
rect 9404 17280 9456 17289
rect 9864 17280 9916 17332
rect 11060 17323 11112 17332
rect 4068 17212 4120 17264
rect 4252 17212 4304 17264
rect 7748 17212 7800 17264
rect 5908 17144 5960 17196
rect 7196 17144 7248 17196
rect 1860 17076 1912 17128
rect 3516 17076 3568 17128
rect 4160 17076 4212 17128
rect 4988 17076 5040 17128
rect 5172 17119 5224 17128
rect 5172 17085 5206 17119
rect 5206 17085 5224 17119
rect 5172 17076 5224 17085
rect 7012 17076 7064 17128
rect 11060 17289 11069 17323
rect 11069 17289 11103 17323
rect 11103 17289 11112 17323
rect 11060 17280 11112 17289
rect 11152 17280 11204 17332
rect 12900 17280 12952 17332
rect 22100 17280 22152 17332
rect 8300 17119 8352 17128
rect 8300 17085 8323 17119
rect 8323 17085 8352 17119
rect 2136 16940 2188 16992
rect 3332 16940 3384 16992
rect 4528 16983 4580 16992
rect 4528 16949 4537 16983
rect 4537 16949 4571 16983
rect 4571 16949 4580 16983
rect 4528 16940 4580 16949
rect 7932 17008 7984 17060
rect 8300 17076 8352 17085
rect 9496 17076 9548 17128
rect 13820 17212 13872 17264
rect 15016 17212 15068 17264
rect 19064 17212 19116 17264
rect 14832 17144 14884 17196
rect 16304 17144 16356 17196
rect 16764 17144 16816 17196
rect 11980 17076 12032 17128
rect 12440 17076 12492 17128
rect 13268 17076 13320 17128
rect 9956 17051 10008 17060
rect 9956 17017 9990 17051
rect 9990 17017 10008 17051
rect 11704 17051 11756 17060
rect 9956 17008 10008 17017
rect 11704 17017 11713 17051
rect 11713 17017 11747 17051
rect 11747 17017 11756 17051
rect 11704 17008 11756 17017
rect 13360 17008 13412 17060
rect 16672 17076 16724 17128
rect 17224 17076 17276 17128
rect 18052 17119 18104 17128
rect 18052 17085 18061 17119
rect 18061 17085 18095 17119
rect 18095 17085 18104 17119
rect 18052 17076 18104 17085
rect 19340 17144 19392 17196
rect 20168 17187 20220 17196
rect 19892 17076 19944 17128
rect 20168 17153 20177 17187
rect 20177 17153 20211 17187
rect 20211 17153 20220 17187
rect 20168 17144 20220 17153
rect 20260 17187 20312 17196
rect 20260 17153 20269 17187
rect 20269 17153 20303 17187
rect 20303 17153 20312 17187
rect 20260 17144 20312 17153
rect 20904 17144 20956 17196
rect 20720 17119 20772 17128
rect 20720 17085 20729 17119
rect 20729 17085 20763 17119
rect 20763 17085 20772 17119
rect 20720 17076 20772 17085
rect 14004 17008 14056 17060
rect 18144 17008 18196 17060
rect 6276 16983 6328 16992
rect 6276 16949 6285 16983
rect 6285 16949 6319 16983
rect 6319 16949 6328 16983
rect 6276 16940 6328 16949
rect 7104 16940 7156 16992
rect 7472 16983 7524 16992
rect 7472 16949 7481 16983
rect 7481 16949 7515 16983
rect 7515 16949 7524 16983
rect 7472 16940 7524 16949
rect 8116 16940 8168 16992
rect 11336 16983 11388 16992
rect 11336 16949 11345 16983
rect 11345 16949 11379 16983
rect 11379 16949 11388 16983
rect 11336 16940 11388 16949
rect 12348 16940 12400 16992
rect 12716 16940 12768 16992
rect 12900 16983 12952 16992
rect 12900 16949 12909 16983
rect 12909 16949 12943 16983
rect 12943 16949 12952 16983
rect 12900 16940 12952 16949
rect 13728 16940 13780 16992
rect 15108 16940 15160 16992
rect 15292 16940 15344 16992
rect 16304 16940 16356 16992
rect 16488 16983 16540 16992
rect 16488 16949 16497 16983
rect 16497 16949 16531 16983
rect 16531 16949 16540 16983
rect 16488 16940 16540 16949
rect 16948 16983 17000 16992
rect 16948 16949 16957 16983
rect 16957 16949 16991 16983
rect 16991 16949 17000 16983
rect 16948 16940 17000 16949
rect 17040 16940 17092 16992
rect 17868 16940 17920 16992
rect 18512 16940 18564 16992
rect 19064 16940 19116 16992
rect 19248 16940 19300 16992
rect 19892 16940 19944 16992
rect 21180 17076 21232 17128
rect 22192 17076 22244 17128
rect 21180 16940 21232 16992
rect 21456 16940 21508 16992
rect 21640 17051 21692 17060
rect 21640 17017 21674 17051
rect 21674 17017 21692 17051
rect 21640 17008 21692 17017
rect 22560 17008 22612 17060
rect 21732 16940 21784 16992
rect 8379 16838 8431 16890
rect 8443 16838 8495 16890
rect 8507 16838 8559 16890
rect 8571 16838 8623 16890
rect 15776 16838 15828 16890
rect 15840 16838 15892 16890
rect 15904 16838 15956 16890
rect 15968 16838 16020 16890
rect 1768 16779 1820 16788
rect 1768 16745 1777 16779
rect 1777 16745 1811 16779
rect 1811 16745 1820 16779
rect 1768 16736 1820 16745
rect 3516 16779 3568 16788
rect 3516 16745 3525 16779
rect 3525 16745 3559 16779
rect 3559 16745 3568 16779
rect 3516 16736 3568 16745
rect 5908 16736 5960 16788
rect 6092 16736 6144 16788
rect 3424 16668 3476 16720
rect 4344 16668 4396 16720
rect 5632 16668 5684 16720
rect 6276 16668 6328 16720
rect 7288 16736 7340 16788
rect 8208 16736 8260 16788
rect 14924 16736 14976 16788
rect 16488 16736 16540 16788
rect 20904 16779 20956 16788
rect 20904 16745 20913 16779
rect 20913 16745 20947 16779
rect 20947 16745 20956 16779
rect 20904 16736 20956 16745
rect 20996 16736 21048 16788
rect 4436 16600 4488 16652
rect 7012 16600 7064 16652
rect 7932 16600 7984 16652
rect 8208 16600 8260 16652
rect 8760 16643 8812 16652
rect 8760 16609 8769 16643
rect 8769 16609 8803 16643
rect 8803 16609 8812 16643
rect 8760 16600 8812 16609
rect 9496 16643 9548 16652
rect 1492 16532 1544 16584
rect 2136 16575 2188 16584
rect 2136 16541 2145 16575
rect 2145 16541 2179 16575
rect 2179 16541 2188 16575
rect 2136 16532 2188 16541
rect 4804 16575 4856 16584
rect 4804 16541 4813 16575
rect 4813 16541 4847 16575
rect 4847 16541 4856 16575
rect 4804 16532 4856 16541
rect 6920 16532 6972 16584
rect 9496 16609 9505 16643
rect 9505 16609 9539 16643
rect 9539 16609 9548 16643
rect 9496 16600 9548 16609
rect 10048 16668 10100 16720
rect 10140 16600 10192 16652
rect 10324 16600 10376 16652
rect 10416 16532 10468 16584
rect 10692 16575 10744 16584
rect 10692 16541 10704 16575
rect 10704 16541 10738 16575
rect 10738 16541 10744 16575
rect 10968 16575 11020 16584
rect 10692 16532 10744 16541
rect 10968 16541 10977 16575
rect 10977 16541 11011 16575
rect 11011 16541 11020 16575
rect 10968 16532 11020 16541
rect 11244 16600 11296 16652
rect 14188 16668 14240 16720
rect 16028 16668 16080 16720
rect 16948 16668 17000 16720
rect 12992 16600 13044 16652
rect 14832 16600 14884 16652
rect 15108 16600 15160 16652
rect 12348 16575 12400 16584
rect 12348 16541 12357 16575
rect 12357 16541 12391 16575
rect 12391 16541 12400 16575
rect 12348 16532 12400 16541
rect 4528 16396 4580 16448
rect 9220 16396 9272 16448
rect 12256 16464 12308 16516
rect 14004 16507 14056 16516
rect 11888 16396 11940 16448
rect 12716 16396 12768 16448
rect 13728 16439 13780 16448
rect 13728 16405 13737 16439
rect 13737 16405 13771 16439
rect 13771 16405 13780 16439
rect 13728 16396 13780 16405
rect 14004 16473 14013 16507
rect 14013 16473 14047 16507
rect 14047 16473 14056 16507
rect 14004 16464 14056 16473
rect 14188 16464 14240 16516
rect 14740 16532 14792 16584
rect 16488 16600 16540 16652
rect 16764 16600 16816 16652
rect 17224 16643 17276 16652
rect 17224 16609 17258 16643
rect 17258 16609 17276 16643
rect 17224 16600 17276 16609
rect 18144 16668 18196 16720
rect 18052 16600 18104 16652
rect 16948 16575 17000 16584
rect 16948 16541 16957 16575
rect 16957 16541 16991 16575
rect 16991 16541 17000 16575
rect 16948 16532 17000 16541
rect 18972 16600 19024 16652
rect 16672 16507 16724 16516
rect 16672 16473 16681 16507
rect 16681 16473 16715 16507
rect 16715 16473 16724 16507
rect 16672 16464 16724 16473
rect 16764 16464 16816 16516
rect 17868 16396 17920 16448
rect 18144 16396 18196 16448
rect 20076 16668 20128 16720
rect 22100 16668 22152 16720
rect 21364 16643 21416 16652
rect 21364 16609 21373 16643
rect 21373 16609 21407 16643
rect 21407 16609 21416 16643
rect 21364 16600 21416 16609
rect 23112 16600 23164 16652
rect 20168 16532 20220 16584
rect 21456 16575 21508 16584
rect 21456 16541 21465 16575
rect 21465 16541 21499 16575
rect 21499 16541 21508 16575
rect 21456 16532 21508 16541
rect 20260 16464 20312 16516
rect 4680 16294 4732 16346
rect 4744 16294 4796 16346
rect 4808 16294 4860 16346
rect 4872 16294 4924 16346
rect 12078 16294 12130 16346
rect 12142 16294 12194 16346
rect 12206 16294 12258 16346
rect 12270 16294 12322 16346
rect 19475 16294 19527 16346
rect 19539 16294 19591 16346
rect 19603 16294 19655 16346
rect 19667 16294 19719 16346
rect 2780 16192 2832 16244
rect 3700 16192 3752 16244
rect 4160 16192 4212 16244
rect 7472 16192 7524 16244
rect 9220 16192 9272 16244
rect 4436 16167 4488 16176
rect 4436 16133 4445 16167
rect 4445 16133 4479 16167
rect 4479 16133 4488 16167
rect 4436 16124 4488 16133
rect 7656 16124 7708 16176
rect 8116 16124 8168 16176
rect 10232 16124 10284 16176
rect 12992 16192 13044 16244
rect 15200 16235 15252 16244
rect 12900 16124 12952 16176
rect 15200 16201 15209 16235
rect 15209 16201 15243 16235
rect 15243 16201 15252 16235
rect 15200 16192 15252 16201
rect 1492 16099 1544 16108
rect 1492 16065 1501 16099
rect 1501 16065 1535 16099
rect 1535 16065 1544 16099
rect 1492 16056 1544 16065
rect 4344 16056 4396 16108
rect 4804 16031 4856 16040
rect 4804 15997 4813 16031
rect 4813 15997 4847 16031
rect 4847 15997 4856 16031
rect 4804 15988 4856 15997
rect 6092 15988 6144 16040
rect 7656 15988 7708 16040
rect 7932 16056 7984 16108
rect 8852 16056 8904 16108
rect 8944 16056 8996 16108
rect 11244 16056 11296 16108
rect 11428 16099 11480 16108
rect 11428 16065 11437 16099
rect 11437 16065 11471 16099
rect 11471 16065 11480 16099
rect 11428 16056 11480 16065
rect 11704 16056 11756 16108
rect 3148 15895 3200 15904
rect 3148 15861 3157 15895
rect 3157 15861 3191 15895
rect 3191 15861 3200 15895
rect 3148 15852 3200 15861
rect 3516 15895 3568 15904
rect 3516 15861 3525 15895
rect 3525 15861 3559 15895
rect 3559 15861 3568 15895
rect 3516 15852 3568 15861
rect 3700 15852 3752 15904
rect 5356 15920 5408 15972
rect 5540 15852 5592 15904
rect 9312 15988 9364 16040
rect 9680 15988 9732 16040
rect 10140 15988 10192 16040
rect 11520 15988 11572 16040
rect 11888 15988 11940 16040
rect 13820 16099 13872 16108
rect 13820 16065 13829 16099
rect 13829 16065 13863 16099
rect 13863 16065 13872 16099
rect 13820 16056 13872 16065
rect 15108 16056 15160 16108
rect 17684 16192 17736 16244
rect 20168 16192 20220 16244
rect 22376 16192 22428 16244
rect 17040 16124 17092 16176
rect 21364 16124 21416 16176
rect 20260 16099 20312 16108
rect 20260 16065 20269 16099
rect 20269 16065 20303 16099
rect 20303 16065 20312 16099
rect 20260 16056 20312 16065
rect 20812 16056 20864 16108
rect 14924 15988 14976 16040
rect 17592 15988 17644 16040
rect 17684 15988 17736 16040
rect 17868 15988 17920 16040
rect 21364 16031 21416 16040
rect 21364 15997 21373 16031
rect 21373 15997 21407 16031
rect 21407 15997 21416 16031
rect 21364 15988 21416 15997
rect 22192 15988 22244 16040
rect 7748 15895 7800 15904
rect 7748 15861 7757 15895
rect 7757 15861 7791 15895
rect 7791 15861 7800 15895
rect 7748 15852 7800 15861
rect 10416 15852 10468 15904
rect 10968 15920 11020 15972
rect 15384 15920 15436 15972
rect 15660 15920 15712 15972
rect 15844 15920 15896 15972
rect 20904 15963 20956 15972
rect 20904 15929 20913 15963
rect 20913 15929 20947 15963
rect 20947 15929 20956 15963
rect 20904 15920 20956 15929
rect 21732 15920 21784 15972
rect 11244 15895 11296 15904
rect 11244 15861 11253 15895
rect 11253 15861 11287 15895
rect 11287 15861 11296 15895
rect 11244 15852 11296 15861
rect 11796 15852 11848 15904
rect 12348 15852 12400 15904
rect 12716 15852 12768 15904
rect 12808 15895 12860 15904
rect 12808 15861 12817 15895
rect 12817 15861 12851 15895
rect 12851 15861 12860 15895
rect 12808 15852 12860 15861
rect 13268 15852 13320 15904
rect 13912 15852 13964 15904
rect 16304 15852 16356 15904
rect 16672 15852 16724 15904
rect 17500 15852 17552 15904
rect 20536 15852 20588 15904
rect 20996 15895 21048 15904
rect 20996 15861 21005 15895
rect 21005 15861 21039 15895
rect 21039 15861 21048 15895
rect 20996 15852 21048 15861
rect 22744 15895 22796 15904
rect 22744 15861 22753 15895
rect 22753 15861 22787 15895
rect 22787 15861 22796 15895
rect 22744 15852 22796 15861
rect 8379 15750 8431 15802
rect 8443 15750 8495 15802
rect 8507 15750 8559 15802
rect 8571 15750 8623 15802
rect 15776 15750 15828 15802
rect 15840 15750 15892 15802
rect 15904 15750 15956 15802
rect 15968 15750 16020 15802
rect 2872 15648 2924 15700
rect 7012 15648 7064 15700
rect 2780 15580 2832 15632
rect 4344 15580 4396 15632
rect 3976 15512 4028 15564
rect 1768 15487 1820 15496
rect 1768 15453 1777 15487
rect 1777 15453 1811 15487
rect 1811 15453 1820 15487
rect 1768 15444 1820 15453
rect 1676 15308 1728 15360
rect 4528 15444 4580 15496
rect 4344 15376 4396 15428
rect 4804 15580 4856 15632
rect 5540 15512 5592 15564
rect 6184 15580 6236 15632
rect 6552 15580 6604 15632
rect 6736 15580 6788 15632
rect 7748 15648 7800 15700
rect 9312 15648 9364 15700
rect 9496 15648 9548 15700
rect 9864 15648 9916 15700
rect 11336 15648 11388 15700
rect 6920 15512 6972 15564
rect 8944 15580 8996 15632
rect 10232 15580 10284 15632
rect 14924 15691 14976 15700
rect 14924 15657 14933 15691
rect 14933 15657 14967 15691
rect 14967 15657 14976 15691
rect 14924 15648 14976 15657
rect 15200 15648 15252 15700
rect 8116 15512 8168 15564
rect 5080 15487 5132 15496
rect 5080 15453 5089 15487
rect 5089 15453 5123 15487
rect 5123 15453 5132 15487
rect 5080 15444 5132 15453
rect 8484 15512 8536 15564
rect 10048 15555 10100 15564
rect 10048 15521 10057 15555
rect 10057 15521 10091 15555
rect 10091 15521 10100 15555
rect 10048 15512 10100 15521
rect 6736 15376 6788 15428
rect 11796 15580 11848 15632
rect 13912 15580 13964 15632
rect 16304 15648 16356 15700
rect 20996 15648 21048 15700
rect 15752 15580 15804 15632
rect 19340 15580 19392 15632
rect 19432 15580 19484 15632
rect 20720 15580 20772 15632
rect 10600 15444 10652 15496
rect 6828 15308 6880 15360
rect 8852 15308 8904 15360
rect 9680 15308 9732 15360
rect 10508 15308 10560 15360
rect 12348 15376 12400 15428
rect 11980 15308 12032 15360
rect 12808 15512 12860 15564
rect 13820 15512 13872 15564
rect 14096 15512 14148 15564
rect 14924 15512 14976 15564
rect 12716 15487 12768 15496
rect 12716 15453 12725 15487
rect 12725 15453 12759 15487
rect 12759 15453 12768 15487
rect 12716 15444 12768 15453
rect 13728 15444 13780 15496
rect 13912 15444 13964 15496
rect 17040 15512 17092 15564
rect 17500 15512 17552 15564
rect 17960 15512 18012 15564
rect 18328 15512 18380 15564
rect 20260 15512 20312 15564
rect 21364 15580 21416 15632
rect 16948 15487 17000 15496
rect 14004 15376 14056 15428
rect 15200 15376 15252 15428
rect 16948 15453 16957 15487
rect 16957 15453 16991 15487
rect 16991 15453 17000 15487
rect 16948 15444 17000 15453
rect 18052 15444 18104 15496
rect 19984 15444 20036 15496
rect 22744 15512 22796 15564
rect 20444 15376 20496 15428
rect 20628 15419 20680 15428
rect 20628 15385 20637 15419
rect 20637 15385 20671 15419
rect 20671 15385 20680 15419
rect 20628 15376 20680 15385
rect 14188 15308 14240 15360
rect 14556 15351 14608 15360
rect 14556 15317 14565 15351
rect 14565 15317 14599 15351
rect 14599 15317 14608 15351
rect 14556 15308 14608 15317
rect 15660 15308 15712 15360
rect 16948 15308 17000 15360
rect 17224 15308 17276 15360
rect 19892 15308 19944 15360
rect 20076 15308 20128 15360
rect 22376 15351 22428 15360
rect 22376 15317 22385 15351
rect 22385 15317 22419 15351
rect 22419 15317 22428 15351
rect 22376 15308 22428 15317
rect 4680 15206 4732 15258
rect 4744 15206 4796 15258
rect 4808 15206 4860 15258
rect 4872 15206 4924 15258
rect 12078 15206 12130 15258
rect 12142 15206 12194 15258
rect 12206 15206 12258 15258
rect 12270 15206 12322 15258
rect 19475 15206 19527 15258
rect 19539 15206 19591 15258
rect 19603 15206 19655 15258
rect 19667 15206 19719 15258
rect 3424 15104 3476 15156
rect 3516 15104 3568 15156
rect 5080 15104 5132 15156
rect 5540 15104 5592 15156
rect 7656 15104 7708 15156
rect 7932 15104 7984 15156
rect 5448 15036 5500 15088
rect 5724 15036 5776 15088
rect 3884 14968 3936 15020
rect 4436 14968 4488 15020
rect 8760 15036 8812 15088
rect 7840 14968 7892 15020
rect 8024 14968 8076 15020
rect 8208 14968 8260 15020
rect 9956 15104 10008 15156
rect 1400 14943 1452 14952
rect 1400 14909 1409 14943
rect 1409 14909 1443 14943
rect 1443 14909 1452 14943
rect 1400 14900 1452 14909
rect 1768 14900 1820 14952
rect 2780 14900 2832 14952
rect 3976 14943 4028 14952
rect 3976 14909 3985 14943
rect 3985 14909 4019 14943
rect 4019 14909 4028 14943
rect 3976 14900 4028 14909
rect 2504 14832 2556 14884
rect 2688 14832 2740 14884
rect 5172 14832 5224 14884
rect 6000 14900 6052 14952
rect 6828 14900 6880 14952
rect 8300 14943 8352 14952
rect 8300 14909 8309 14943
rect 8309 14909 8343 14943
rect 8343 14909 8352 14943
rect 8300 14900 8352 14909
rect 8484 14900 8536 14952
rect 8668 14900 8720 14952
rect 11888 15104 11940 15156
rect 10600 14900 10652 14952
rect 11980 14900 12032 14952
rect 12716 15104 12768 15156
rect 12808 15104 12860 15156
rect 18512 15104 18564 15156
rect 19340 15104 19392 15156
rect 13544 15036 13596 15088
rect 13728 15036 13780 15088
rect 15384 15036 15436 15088
rect 16304 15036 16356 15088
rect 15200 14968 15252 15020
rect 16212 14968 16264 15020
rect 17868 14968 17920 15020
rect 19432 14968 19484 15020
rect 4068 14807 4120 14816
rect 4068 14773 4077 14807
rect 4077 14773 4111 14807
rect 4111 14773 4120 14807
rect 4068 14764 4120 14773
rect 5080 14807 5132 14816
rect 5080 14773 5089 14807
rect 5089 14773 5123 14807
rect 5123 14773 5132 14807
rect 5080 14764 5132 14773
rect 6184 14764 6236 14816
rect 8760 14832 8812 14884
rect 9128 14875 9180 14884
rect 9128 14841 9162 14875
rect 9162 14841 9180 14875
rect 9128 14832 9180 14841
rect 12348 14832 12400 14884
rect 12992 14900 13044 14952
rect 14004 14900 14056 14952
rect 14188 14900 14240 14952
rect 15384 14900 15436 14952
rect 15752 14943 15804 14952
rect 15752 14909 15761 14943
rect 15761 14909 15795 14943
rect 15795 14909 15804 14943
rect 15752 14900 15804 14909
rect 15936 14900 15988 14952
rect 18052 14900 18104 14952
rect 13544 14832 13596 14884
rect 13912 14832 13964 14884
rect 10140 14764 10192 14816
rect 13452 14764 13504 14816
rect 13820 14807 13872 14816
rect 13820 14773 13829 14807
rect 13829 14773 13863 14807
rect 13863 14773 13872 14807
rect 13820 14764 13872 14773
rect 14188 14764 14240 14816
rect 14740 14764 14792 14816
rect 15292 14832 15344 14884
rect 16672 14832 16724 14884
rect 17224 14832 17276 14884
rect 15660 14764 15712 14816
rect 16580 14764 16632 14816
rect 16764 14764 16816 14816
rect 17500 14764 17552 14816
rect 17868 14832 17920 14884
rect 19064 14832 19116 14884
rect 19892 14832 19944 14884
rect 21732 14832 21784 14884
rect 20444 14764 20496 14816
rect 20904 14807 20956 14816
rect 20904 14773 20913 14807
rect 20913 14773 20947 14807
rect 20947 14773 20956 14807
rect 20904 14764 20956 14773
rect 21364 14807 21416 14816
rect 21364 14773 21373 14807
rect 21373 14773 21407 14807
rect 21407 14773 21416 14807
rect 21364 14764 21416 14773
rect 22284 14807 22336 14816
rect 22284 14773 22293 14807
rect 22293 14773 22327 14807
rect 22327 14773 22336 14807
rect 22284 14764 22336 14773
rect 8379 14662 8431 14714
rect 8443 14662 8495 14714
rect 8507 14662 8559 14714
rect 8571 14662 8623 14714
rect 15776 14662 15828 14714
rect 15840 14662 15892 14714
rect 15904 14662 15956 14714
rect 15968 14662 16020 14714
rect 1768 14560 1820 14612
rect 3148 14492 3200 14544
rect 4988 14560 5040 14612
rect 2044 14424 2096 14476
rect 5724 14492 5776 14544
rect 6184 14560 6236 14612
rect 8208 14560 8260 14612
rect 9128 14560 9180 14612
rect 11060 14603 11112 14612
rect 11060 14569 11069 14603
rect 11069 14569 11103 14603
rect 11103 14569 11112 14603
rect 11060 14560 11112 14569
rect 11336 14560 11388 14612
rect 12532 14560 12584 14612
rect 8668 14492 8720 14544
rect 14188 14560 14240 14612
rect 16120 14603 16172 14612
rect 16120 14569 16129 14603
rect 16129 14569 16163 14603
rect 16163 14569 16172 14603
rect 16120 14560 16172 14569
rect 17316 14560 17368 14612
rect 18512 14560 18564 14612
rect 19432 14560 19484 14612
rect 21364 14560 21416 14612
rect 21640 14560 21692 14612
rect 13084 14492 13136 14544
rect 14004 14492 14056 14544
rect 4160 14424 4212 14476
rect 5080 14424 5132 14476
rect 6000 14467 6052 14476
rect 6000 14433 6034 14467
rect 6034 14433 6052 14467
rect 6000 14424 6052 14433
rect 7748 14467 7800 14476
rect 7748 14433 7757 14467
rect 7757 14433 7791 14467
rect 7791 14433 7800 14467
rect 7748 14424 7800 14433
rect 8024 14424 8076 14476
rect 8760 14467 8812 14476
rect 8760 14433 8769 14467
rect 8769 14433 8803 14467
rect 8803 14433 8812 14467
rect 8760 14424 8812 14433
rect 2504 14288 2556 14340
rect 2136 14220 2188 14272
rect 3608 14220 3660 14272
rect 4252 14220 4304 14272
rect 5356 14356 5408 14408
rect 5264 14288 5316 14340
rect 5172 14220 5224 14272
rect 5448 14263 5500 14272
rect 5448 14229 5457 14263
rect 5457 14229 5491 14263
rect 5491 14229 5500 14263
rect 5448 14220 5500 14229
rect 8668 14356 8720 14408
rect 8024 14288 8076 14340
rect 11336 14424 11388 14476
rect 12532 14424 12584 14476
rect 13176 14424 13228 14476
rect 14832 14492 14884 14544
rect 17132 14492 17184 14544
rect 8852 14220 8904 14272
rect 9680 14399 9732 14408
rect 9680 14365 9689 14399
rect 9689 14365 9723 14399
rect 9723 14365 9732 14399
rect 9680 14356 9732 14365
rect 10968 14288 11020 14340
rect 11336 14288 11388 14340
rect 12716 14356 12768 14408
rect 14096 14399 14148 14408
rect 12808 14288 12860 14340
rect 13452 14331 13504 14340
rect 10416 14220 10468 14272
rect 11520 14220 11572 14272
rect 13452 14297 13461 14331
rect 13461 14297 13495 14331
rect 13495 14297 13504 14331
rect 13452 14288 13504 14297
rect 14096 14365 14105 14399
rect 14105 14365 14139 14399
rect 14139 14365 14148 14399
rect 14096 14356 14148 14365
rect 15016 14424 15068 14476
rect 16304 14424 16356 14476
rect 14832 14288 14884 14340
rect 14188 14220 14240 14272
rect 16580 14399 16632 14408
rect 16580 14365 16589 14399
rect 16589 14365 16623 14399
rect 16623 14365 16632 14399
rect 16580 14356 16632 14365
rect 16672 14399 16724 14408
rect 16672 14365 16681 14399
rect 16681 14365 16715 14399
rect 16715 14365 16724 14399
rect 18052 14492 18104 14544
rect 18880 14492 18932 14544
rect 19248 14424 19300 14476
rect 19432 14424 19484 14476
rect 20076 14492 20128 14544
rect 20720 14467 20772 14476
rect 20720 14433 20729 14467
rect 20729 14433 20763 14467
rect 20763 14433 20772 14467
rect 20720 14424 20772 14433
rect 16672 14356 16724 14365
rect 15108 14288 15160 14340
rect 15384 14288 15436 14340
rect 18880 14356 18932 14408
rect 19892 14356 19944 14408
rect 15660 14220 15712 14272
rect 16120 14220 16172 14272
rect 17316 14220 17368 14272
rect 20996 14288 21048 14340
rect 19064 14220 19116 14272
rect 21364 14220 21416 14272
rect 22100 14220 22152 14272
rect 22376 14492 22428 14544
rect 4680 14118 4732 14170
rect 4744 14118 4796 14170
rect 4808 14118 4860 14170
rect 4872 14118 4924 14170
rect 12078 14118 12130 14170
rect 12142 14118 12194 14170
rect 12206 14118 12258 14170
rect 12270 14118 12322 14170
rect 19475 14118 19527 14170
rect 19539 14118 19591 14170
rect 19603 14118 19655 14170
rect 19667 14118 19719 14170
rect 5080 14059 5132 14068
rect 1676 13991 1728 14000
rect 1676 13957 1685 13991
rect 1685 13957 1719 13991
rect 1719 13957 1728 13991
rect 1676 13948 1728 13957
rect 5080 14025 5089 14059
rect 5089 14025 5123 14059
rect 5123 14025 5132 14059
rect 5080 14016 5132 14025
rect 8668 14059 8720 14068
rect 5172 13948 5224 14000
rect 6184 13948 6236 14000
rect 6460 13948 6512 14000
rect 8668 14025 8677 14059
rect 8677 14025 8711 14059
rect 8711 14025 8720 14059
rect 8668 14016 8720 14025
rect 11704 14016 11756 14068
rect 12716 14016 12768 14068
rect 1676 13744 1728 13796
rect 3056 13812 3108 13864
rect 3608 13812 3660 13864
rect 6368 13880 6420 13932
rect 9312 13948 9364 14000
rect 11796 13948 11848 14000
rect 10416 13923 10468 13932
rect 3976 13855 4028 13864
rect 3976 13821 4010 13855
rect 4010 13821 4028 13855
rect 3976 13812 4028 13821
rect 5356 13812 5408 13864
rect 7564 13812 7616 13864
rect 8668 13812 8720 13864
rect 10416 13889 10425 13923
rect 10425 13889 10459 13923
rect 10459 13889 10468 13923
rect 10416 13880 10468 13889
rect 10600 13880 10652 13932
rect 11520 13880 11572 13932
rect 11244 13812 11296 13864
rect 12164 13880 12216 13932
rect 15016 14016 15068 14068
rect 16580 14016 16632 14068
rect 13452 13948 13504 14000
rect 13544 13948 13596 14000
rect 16212 13948 16264 14000
rect 16396 13991 16448 14000
rect 16396 13957 16405 13991
rect 16405 13957 16439 13991
rect 16439 13957 16448 13991
rect 16396 13948 16448 13957
rect 19340 14016 19392 14068
rect 22284 14016 22336 14068
rect 14096 13880 14148 13932
rect 14556 13880 14608 13932
rect 15108 13880 15160 13932
rect 16120 13923 16172 13932
rect 16120 13889 16129 13923
rect 16129 13889 16163 13923
rect 16163 13889 16172 13923
rect 17960 13948 18012 14000
rect 19248 13948 19300 14000
rect 16120 13880 16172 13889
rect 11888 13812 11940 13864
rect 12716 13812 12768 13864
rect 14188 13812 14240 13864
rect 16488 13812 16540 13864
rect 17132 13880 17184 13932
rect 16672 13812 16724 13864
rect 18052 13923 18104 13932
rect 18052 13889 18061 13923
rect 18061 13889 18095 13923
rect 18095 13889 18104 13923
rect 18052 13880 18104 13889
rect 20168 13880 20220 13932
rect 20720 13880 20772 13932
rect 22468 13923 22520 13932
rect 22468 13889 22477 13923
rect 22477 13889 22511 13923
rect 22511 13889 22520 13923
rect 22468 13880 22520 13889
rect 17776 13812 17828 13864
rect 18328 13855 18380 13864
rect 18328 13821 18362 13855
rect 18362 13821 18380 13855
rect 18328 13812 18380 13821
rect 20444 13812 20496 13864
rect 21272 13812 21324 13864
rect 2504 13744 2556 13796
rect 4160 13744 4212 13796
rect 10048 13744 10100 13796
rect 11152 13787 11204 13796
rect 5724 13719 5776 13728
rect 5724 13685 5733 13719
rect 5733 13685 5767 13719
rect 5767 13685 5776 13719
rect 5724 13676 5776 13685
rect 5816 13719 5868 13728
rect 5816 13685 5825 13719
rect 5825 13685 5859 13719
rect 5859 13685 5868 13719
rect 5816 13676 5868 13685
rect 7196 13676 7248 13728
rect 7564 13676 7616 13728
rect 8668 13676 8720 13728
rect 9036 13719 9088 13728
rect 9036 13685 9045 13719
rect 9045 13685 9079 13719
rect 9079 13685 9088 13719
rect 9036 13676 9088 13685
rect 10232 13719 10284 13728
rect 10232 13685 10241 13719
rect 10241 13685 10275 13719
rect 10275 13685 10284 13719
rect 10232 13676 10284 13685
rect 11152 13753 11161 13787
rect 11161 13753 11195 13787
rect 11195 13753 11204 13787
rect 11152 13744 11204 13753
rect 11244 13719 11296 13728
rect 11244 13685 11253 13719
rect 11253 13685 11287 13719
rect 11287 13685 11296 13719
rect 11244 13676 11296 13685
rect 11520 13676 11572 13728
rect 13728 13787 13780 13796
rect 13728 13753 13737 13787
rect 13737 13753 13771 13787
rect 13771 13753 13780 13787
rect 13728 13744 13780 13753
rect 13820 13744 13872 13796
rect 17132 13744 17184 13796
rect 19616 13744 19668 13796
rect 12716 13676 12768 13728
rect 13084 13676 13136 13728
rect 14280 13676 14332 13728
rect 15660 13676 15712 13728
rect 16120 13676 16172 13728
rect 16212 13676 16264 13728
rect 19340 13676 19392 13728
rect 20076 13676 20128 13728
rect 20628 13676 20680 13728
rect 21272 13676 21324 13728
rect 22376 13719 22428 13728
rect 22376 13685 22385 13719
rect 22385 13685 22419 13719
rect 22419 13685 22428 13719
rect 22376 13676 22428 13685
rect 8379 13574 8431 13626
rect 8443 13574 8495 13626
rect 8507 13574 8559 13626
rect 8571 13574 8623 13626
rect 15776 13574 15828 13626
rect 15840 13574 15892 13626
rect 15904 13574 15956 13626
rect 15968 13574 16020 13626
rect 3056 13515 3108 13524
rect 3056 13481 3065 13515
rect 3065 13481 3099 13515
rect 3099 13481 3108 13515
rect 3056 13472 3108 13481
rect 4068 13472 4120 13524
rect 6000 13472 6052 13524
rect 7748 13472 7800 13524
rect 9496 13472 9548 13524
rect 10232 13472 10284 13524
rect 2136 13404 2188 13456
rect 5448 13404 5500 13456
rect 8668 13404 8720 13456
rect 1676 13379 1728 13388
rect 1676 13345 1685 13379
rect 1685 13345 1719 13379
rect 1719 13345 1728 13379
rect 1676 13336 1728 13345
rect 3424 13379 3476 13388
rect 3424 13345 3433 13379
rect 3433 13345 3467 13379
rect 3467 13345 3476 13379
rect 3424 13336 3476 13345
rect 4160 13336 4212 13388
rect 4252 13336 4304 13388
rect 5080 13336 5132 13388
rect 7012 13336 7064 13388
rect 7932 13336 7984 13388
rect 9956 13404 10008 13456
rect 10508 13472 10560 13524
rect 11152 13472 11204 13524
rect 9220 13336 9272 13388
rect 10140 13379 10192 13388
rect 10140 13345 10149 13379
rect 10149 13345 10183 13379
rect 10183 13345 10192 13379
rect 10140 13336 10192 13345
rect 5264 13132 5316 13184
rect 5448 13132 5500 13184
rect 9680 13268 9732 13320
rect 10600 13404 10652 13456
rect 10968 13404 11020 13456
rect 12532 13472 12584 13524
rect 14096 13472 14148 13524
rect 14648 13472 14700 13524
rect 14832 13472 14884 13524
rect 16764 13472 16816 13524
rect 18512 13472 18564 13524
rect 19800 13472 19852 13524
rect 11244 13336 11296 13388
rect 16488 13404 16540 13456
rect 16580 13404 16632 13456
rect 12072 13311 12124 13320
rect 9036 13200 9088 13252
rect 10232 13200 10284 13252
rect 12072 13277 12081 13311
rect 12081 13277 12115 13311
rect 12115 13277 12124 13311
rect 12072 13268 12124 13277
rect 13544 13311 13596 13320
rect 13544 13277 13553 13311
rect 13553 13277 13587 13311
rect 13587 13277 13596 13311
rect 13544 13268 13596 13277
rect 15384 13336 15436 13388
rect 17224 13379 17276 13388
rect 17224 13345 17258 13379
rect 17258 13345 17276 13379
rect 17224 13336 17276 13345
rect 15292 13311 15344 13320
rect 15292 13277 15301 13311
rect 15301 13277 15335 13311
rect 15335 13277 15344 13311
rect 15292 13268 15344 13277
rect 16304 13268 16356 13320
rect 14556 13200 14608 13252
rect 8484 13175 8536 13184
rect 8484 13141 8493 13175
rect 8493 13141 8527 13175
rect 8527 13141 8536 13175
rect 8484 13132 8536 13141
rect 9220 13175 9272 13184
rect 9220 13141 9229 13175
rect 9229 13141 9263 13175
rect 9263 13141 9272 13175
rect 9220 13132 9272 13141
rect 9956 13132 10008 13184
rect 12440 13132 12492 13184
rect 14924 13243 14976 13252
rect 14924 13209 14933 13243
rect 14933 13209 14967 13243
rect 14967 13209 14976 13243
rect 14924 13200 14976 13209
rect 22376 13404 22428 13456
rect 18972 13336 19024 13388
rect 18052 13268 18104 13320
rect 18788 13268 18840 13320
rect 20904 13379 20956 13388
rect 18052 13132 18104 13184
rect 18512 13132 18564 13184
rect 19340 13132 19392 13184
rect 19800 13132 19852 13184
rect 20536 13175 20588 13184
rect 20536 13141 20545 13175
rect 20545 13141 20579 13175
rect 20579 13141 20588 13175
rect 20536 13132 20588 13141
rect 20904 13345 20913 13379
rect 20913 13345 20947 13379
rect 20947 13345 20956 13379
rect 20904 13336 20956 13345
rect 21364 13379 21416 13388
rect 21364 13345 21373 13379
rect 21373 13345 21407 13379
rect 21407 13345 21416 13379
rect 21364 13336 21416 13345
rect 21640 13379 21692 13388
rect 21640 13345 21674 13379
rect 21674 13345 21692 13379
rect 21640 13336 21692 13345
rect 4680 13030 4732 13082
rect 4744 13030 4796 13082
rect 4808 13030 4860 13082
rect 4872 13030 4924 13082
rect 12078 13030 12130 13082
rect 12142 13030 12194 13082
rect 12206 13030 12258 13082
rect 12270 13030 12322 13082
rect 19475 13030 19527 13082
rect 19539 13030 19591 13082
rect 19603 13030 19655 13082
rect 19667 13030 19719 13082
rect 1676 12928 1728 12980
rect 2044 12928 2096 12980
rect 3792 12928 3844 12980
rect 7656 12928 7708 12980
rect 8760 12928 8812 12980
rect 9680 12971 9732 12980
rect 9680 12937 9689 12971
rect 9689 12937 9723 12971
rect 9723 12937 9732 12971
rect 9680 12928 9732 12937
rect 11060 12928 11112 12980
rect 11244 12928 11296 12980
rect 12716 12928 12768 12980
rect 3884 12792 3936 12844
rect 4252 12792 4304 12844
rect 7012 12835 7064 12844
rect 7012 12801 7021 12835
rect 7021 12801 7055 12835
rect 7055 12801 7064 12835
rect 7012 12792 7064 12801
rect 9312 12835 9364 12844
rect 9312 12801 9321 12835
rect 9321 12801 9355 12835
rect 9355 12801 9364 12835
rect 9312 12792 9364 12801
rect 11336 12860 11388 12912
rect 19800 12928 19852 12980
rect 20168 12928 20220 12980
rect 14556 12860 14608 12912
rect 17316 12860 17368 12912
rect 18328 12860 18380 12912
rect 10140 12792 10192 12844
rect 3332 12724 3384 12776
rect 4252 12656 4304 12708
rect 3608 12631 3660 12640
rect 3608 12597 3617 12631
rect 3617 12597 3651 12631
rect 3651 12597 3660 12631
rect 3608 12588 3660 12597
rect 4068 12631 4120 12640
rect 4068 12597 4077 12631
rect 4077 12597 4111 12631
rect 4111 12597 4120 12631
rect 4068 12588 4120 12597
rect 5816 12724 5868 12776
rect 5908 12724 5960 12776
rect 8484 12724 8536 12776
rect 4436 12656 4488 12708
rect 5448 12656 5500 12708
rect 5724 12588 5776 12640
rect 8208 12588 8260 12640
rect 10039 12724 10091 12776
rect 10232 12724 10284 12776
rect 11152 12724 11204 12776
rect 11796 12724 11848 12776
rect 12624 12792 12676 12844
rect 12992 12767 13044 12776
rect 12992 12733 13001 12767
rect 13001 12733 13035 12767
rect 13035 12733 13044 12767
rect 12992 12724 13044 12733
rect 13544 12724 13596 12776
rect 14556 12724 14608 12776
rect 14924 12767 14976 12776
rect 14924 12733 14958 12767
rect 14958 12733 14976 12767
rect 14924 12724 14976 12733
rect 15292 12724 15344 12776
rect 16304 12767 16356 12776
rect 16304 12733 16313 12767
rect 16313 12733 16347 12767
rect 16347 12733 16356 12767
rect 16304 12724 16356 12733
rect 16580 12767 16632 12776
rect 16580 12733 16614 12767
rect 16614 12733 16632 12767
rect 16580 12724 16632 12733
rect 16856 12724 16908 12776
rect 17500 12792 17552 12844
rect 17868 12792 17920 12844
rect 18972 12792 19024 12844
rect 12348 12656 12400 12708
rect 12624 12699 12676 12708
rect 12624 12665 12633 12699
rect 12633 12665 12667 12699
rect 12667 12665 12676 12699
rect 12624 12656 12676 12665
rect 15660 12656 15712 12708
rect 17500 12656 17552 12708
rect 18880 12724 18932 12776
rect 19800 12792 19852 12844
rect 20996 12928 21048 12980
rect 21364 12928 21416 12980
rect 21732 12971 21784 12980
rect 21732 12937 21741 12971
rect 21741 12937 21775 12971
rect 21775 12937 21784 12971
rect 21732 12928 21784 12937
rect 22376 12835 22428 12844
rect 22376 12801 22385 12835
rect 22385 12801 22419 12835
rect 22419 12801 22428 12835
rect 22376 12792 22428 12801
rect 20168 12724 20220 12776
rect 20536 12767 20588 12776
rect 20536 12733 20559 12767
rect 20559 12733 20588 12767
rect 20536 12724 20588 12733
rect 18512 12699 18564 12708
rect 18512 12665 18521 12699
rect 18521 12665 18555 12699
rect 18555 12665 18564 12699
rect 18512 12656 18564 12665
rect 19064 12656 19116 12708
rect 9036 12631 9088 12640
rect 9036 12597 9045 12631
rect 9045 12597 9079 12631
rect 9079 12597 9088 12631
rect 9036 12588 9088 12597
rect 10692 12588 10744 12640
rect 12532 12588 12584 12640
rect 15384 12588 15436 12640
rect 16856 12588 16908 12640
rect 17684 12631 17736 12640
rect 17684 12597 17693 12631
rect 17693 12597 17727 12631
rect 17727 12597 17736 12631
rect 17684 12588 17736 12597
rect 21272 12588 21324 12640
rect 22284 12588 22336 12640
rect 8379 12486 8431 12538
rect 8443 12486 8495 12538
rect 8507 12486 8559 12538
rect 8571 12486 8623 12538
rect 15776 12486 15828 12538
rect 15840 12486 15892 12538
rect 15904 12486 15956 12538
rect 15968 12486 16020 12538
rect 2136 12384 2188 12436
rect 4528 12384 4580 12436
rect 5816 12384 5868 12436
rect 3148 12359 3200 12368
rect 3148 12325 3157 12359
rect 3157 12325 3191 12359
rect 3191 12325 3200 12359
rect 3148 12316 3200 12325
rect 3240 12316 3292 12368
rect 8208 12384 8260 12436
rect 2044 12248 2096 12300
rect 3332 12248 3384 12300
rect 9680 12384 9732 12436
rect 11520 12384 11572 12436
rect 12348 12384 12400 12436
rect 13452 12384 13504 12436
rect 15476 12384 15528 12436
rect 16212 12384 16264 12436
rect 16304 12384 16356 12436
rect 17132 12384 17184 12436
rect 17224 12384 17276 12436
rect 5816 12248 5868 12300
rect 7012 12291 7064 12300
rect 3884 12180 3936 12232
rect 4160 12180 4212 12232
rect 7012 12257 7021 12291
rect 7021 12257 7055 12291
rect 7055 12257 7064 12291
rect 7012 12248 7064 12257
rect 8852 12248 8904 12300
rect 9128 12248 9180 12300
rect 10692 12248 10744 12300
rect 11520 12248 11572 12300
rect 13636 12316 13688 12368
rect 13820 12248 13872 12300
rect 1952 12044 2004 12096
rect 3700 12044 3752 12096
rect 3884 12044 3936 12096
rect 6920 12112 6972 12164
rect 8208 12112 8260 12164
rect 12992 12112 13044 12164
rect 8300 12044 8352 12096
rect 8392 12087 8444 12096
rect 8392 12053 8401 12087
rect 8401 12053 8435 12087
rect 8435 12053 8444 12087
rect 8392 12044 8444 12053
rect 9036 12044 9088 12096
rect 10048 12044 10100 12096
rect 13268 12044 13320 12096
rect 14648 12087 14700 12096
rect 14648 12053 14657 12087
rect 14657 12053 14691 12087
rect 14691 12053 14700 12087
rect 14648 12044 14700 12053
rect 15568 12248 15620 12300
rect 16764 12316 16816 12368
rect 18052 12359 18104 12368
rect 18052 12325 18086 12359
rect 18086 12325 18104 12359
rect 18052 12316 18104 12325
rect 19064 12384 19116 12436
rect 20812 12384 20864 12436
rect 20904 12384 20956 12436
rect 21180 12384 21232 12436
rect 21272 12359 21324 12368
rect 21272 12325 21306 12359
rect 21306 12325 21324 12359
rect 21272 12316 21324 12325
rect 17592 12248 17644 12300
rect 17132 12180 17184 12232
rect 19616 12248 19668 12300
rect 19800 12291 19852 12300
rect 19800 12257 19809 12291
rect 19809 12257 19843 12291
rect 19843 12257 19852 12291
rect 19800 12248 19852 12257
rect 17408 12112 17460 12164
rect 17684 12112 17736 12164
rect 18880 12180 18932 12232
rect 20168 12248 20220 12300
rect 20996 12291 21048 12300
rect 20996 12257 21005 12291
rect 21005 12257 21039 12291
rect 21039 12257 21048 12291
rect 20996 12248 21048 12257
rect 17960 12044 18012 12096
rect 18144 12044 18196 12096
rect 20260 12044 20312 12096
rect 20996 12044 21048 12096
rect 4680 11942 4732 11994
rect 4744 11942 4796 11994
rect 4808 11942 4860 11994
rect 4872 11942 4924 11994
rect 12078 11942 12130 11994
rect 12142 11942 12194 11994
rect 12206 11942 12258 11994
rect 12270 11942 12322 11994
rect 19475 11942 19527 11994
rect 19539 11942 19591 11994
rect 19603 11942 19655 11994
rect 19667 11942 19719 11994
rect 3424 11840 3476 11892
rect 5816 11883 5868 11892
rect 3516 11772 3568 11824
rect 5816 11849 5825 11883
rect 5825 11849 5859 11883
rect 5859 11849 5868 11883
rect 5816 11840 5868 11849
rect 7472 11840 7524 11892
rect 7748 11840 7800 11892
rect 8208 11840 8260 11892
rect 8300 11840 8352 11892
rect 10968 11840 11020 11892
rect 11152 11840 11204 11892
rect 13820 11840 13872 11892
rect 1952 11747 2004 11756
rect 1952 11713 1961 11747
rect 1961 11713 1995 11747
rect 1995 11713 2004 11747
rect 1952 11704 2004 11713
rect 2136 11747 2188 11756
rect 2136 11713 2145 11747
rect 2145 11713 2179 11747
rect 2179 11713 2188 11747
rect 2136 11704 2188 11713
rect 4068 11704 4120 11756
rect 1952 11568 2004 11620
rect 4160 11636 4212 11688
rect 3332 11568 3384 11620
rect 5908 11636 5960 11688
rect 5448 11568 5500 11620
rect 8116 11772 8168 11824
rect 9956 11772 10008 11824
rect 15660 11840 15712 11892
rect 19800 11840 19852 11892
rect 20628 11840 20680 11892
rect 17684 11772 17736 11824
rect 6552 11636 6604 11688
rect 6920 11636 6972 11688
rect 9312 11704 9364 11756
rect 10048 11704 10100 11756
rect 12624 11704 12676 11756
rect 8208 11636 8260 11688
rect 9680 11679 9732 11688
rect 9680 11645 9689 11679
rect 9689 11645 9723 11679
rect 9723 11645 9732 11679
rect 10508 11679 10560 11688
rect 9680 11636 9732 11645
rect 10508 11645 10542 11679
rect 10542 11645 10560 11679
rect 10508 11636 10560 11645
rect 8392 11568 8444 11620
rect 14004 11636 14056 11688
rect 14556 11636 14608 11688
rect 14740 11679 14792 11688
rect 14740 11645 14774 11679
rect 14774 11645 14792 11679
rect 14740 11636 14792 11645
rect 3608 11500 3660 11552
rect 3792 11500 3844 11552
rect 4344 11500 4396 11552
rect 4528 11500 4580 11552
rect 7932 11500 7984 11552
rect 16764 11704 16816 11756
rect 17408 11747 17460 11756
rect 17408 11713 17417 11747
rect 17417 11713 17451 11747
rect 17451 11713 17460 11747
rect 17408 11704 17460 11713
rect 17868 11704 17920 11756
rect 19892 11704 19944 11756
rect 20352 11704 20404 11756
rect 17316 11679 17368 11688
rect 17316 11645 17325 11679
rect 17325 11645 17359 11679
rect 17359 11645 17368 11679
rect 17316 11636 17368 11645
rect 18144 11636 18196 11688
rect 19064 11636 19116 11688
rect 21916 11704 21968 11756
rect 19340 11568 19392 11620
rect 13820 11500 13872 11552
rect 14556 11500 14608 11552
rect 16212 11500 16264 11552
rect 18052 11500 18104 11552
rect 18328 11500 18380 11552
rect 18972 11500 19024 11552
rect 19616 11543 19668 11552
rect 19616 11509 19625 11543
rect 19625 11509 19659 11543
rect 19659 11509 19668 11543
rect 21272 11636 21324 11688
rect 22284 11679 22336 11688
rect 22284 11645 22293 11679
rect 22293 11645 22327 11679
rect 22327 11645 22336 11679
rect 22284 11636 22336 11645
rect 19616 11500 19668 11509
rect 20536 11500 20588 11552
rect 20812 11500 20864 11552
rect 8379 11398 8431 11450
rect 8443 11398 8495 11450
rect 8507 11398 8559 11450
rect 8571 11398 8623 11450
rect 15776 11398 15828 11450
rect 15840 11398 15892 11450
rect 15904 11398 15956 11450
rect 15968 11398 16020 11450
rect 1584 11339 1636 11348
rect 1584 11305 1593 11339
rect 1593 11305 1627 11339
rect 1627 11305 1636 11339
rect 1584 11296 1636 11305
rect 2136 11296 2188 11348
rect 3792 11296 3844 11348
rect 5448 11339 5500 11348
rect 2780 11228 2832 11280
rect 3148 11228 3200 11280
rect 4252 11228 4304 11280
rect 4160 11160 4212 11212
rect 5448 11305 5457 11339
rect 5457 11305 5491 11339
rect 5491 11305 5500 11339
rect 5448 11296 5500 11305
rect 5816 11296 5868 11348
rect 6092 11160 6144 11212
rect 9404 11296 9456 11348
rect 10508 11296 10560 11348
rect 11520 11296 11572 11348
rect 19340 11296 19392 11348
rect 9956 11228 10008 11280
rect 6920 11203 6972 11212
rect 1952 11135 2004 11144
rect 1952 11101 1961 11135
rect 1961 11101 1995 11135
rect 1995 11101 2004 11135
rect 1952 11092 2004 11101
rect 5540 11092 5592 11144
rect 6920 11169 6929 11203
rect 6929 11169 6963 11203
rect 6963 11169 6972 11203
rect 6920 11160 6972 11169
rect 8208 11160 8260 11212
rect 8760 11160 8812 11212
rect 9588 11160 9640 11212
rect 6368 11135 6420 11144
rect 6368 11101 6377 11135
rect 6377 11101 6411 11135
rect 6411 11101 6420 11135
rect 6368 11092 6420 11101
rect 9036 11135 9088 11144
rect 9036 11101 9045 11135
rect 9045 11101 9079 11135
rect 9079 11101 9088 11135
rect 9036 11092 9088 11101
rect 9312 11092 9364 11144
rect 10048 11160 10100 11212
rect 11152 11160 11204 11212
rect 11612 11203 11664 11212
rect 11612 11169 11621 11203
rect 11621 11169 11655 11203
rect 11655 11169 11664 11203
rect 11612 11160 11664 11169
rect 3332 11067 3384 11076
rect 3332 11033 3341 11067
rect 3341 11033 3375 11067
rect 3375 11033 3384 11067
rect 3332 11024 3384 11033
rect 2596 10956 2648 11008
rect 5724 10999 5776 11008
rect 5724 10965 5733 10999
rect 5733 10965 5767 10999
rect 5767 10965 5776 10999
rect 5724 10956 5776 10965
rect 8300 10999 8352 11008
rect 8300 10965 8309 10999
rect 8309 10965 8343 10999
rect 8343 10965 8352 10999
rect 8300 10956 8352 10965
rect 9864 11024 9916 11076
rect 10968 11024 11020 11076
rect 12440 11203 12492 11212
rect 12440 11169 12449 11203
rect 12449 11169 12483 11203
rect 12483 11169 12492 11203
rect 12440 11160 12492 11169
rect 12624 11160 12676 11212
rect 14280 11160 14332 11212
rect 15292 11228 15344 11280
rect 14648 11135 14700 11144
rect 14648 11101 14657 11135
rect 14657 11101 14691 11135
rect 14691 11101 14700 11135
rect 14648 11092 14700 11101
rect 15660 11160 15712 11212
rect 16488 11228 16540 11280
rect 16672 11160 16724 11212
rect 16764 11160 16816 11212
rect 18144 11228 18196 11280
rect 19616 11228 19668 11280
rect 17316 11160 17368 11212
rect 18880 11203 18932 11212
rect 18880 11169 18889 11203
rect 18889 11169 18923 11203
rect 18923 11169 18932 11203
rect 18880 11160 18932 11169
rect 20168 11296 20220 11348
rect 20444 11296 20496 11348
rect 20628 11296 20680 11348
rect 22192 11296 22244 11348
rect 17132 11092 17184 11144
rect 18328 11092 18380 11144
rect 20996 11160 21048 11212
rect 20260 11092 20312 11144
rect 20628 11092 20680 11144
rect 20904 11092 20956 11144
rect 15016 11024 15068 11076
rect 18236 11024 18288 11076
rect 19984 11024 20036 11076
rect 20444 11024 20496 11076
rect 22836 11024 22888 11076
rect 13544 10956 13596 11008
rect 13912 10999 13964 11008
rect 13912 10965 13921 10999
rect 13921 10965 13955 10999
rect 13955 10965 13964 10999
rect 13912 10956 13964 10965
rect 14188 10999 14240 11008
rect 14188 10965 14197 10999
rect 14197 10965 14231 10999
rect 14231 10965 14240 10999
rect 14188 10956 14240 10965
rect 14372 10956 14424 11008
rect 17500 10956 17552 11008
rect 18788 10956 18840 11008
rect 19064 10956 19116 11008
rect 20260 10999 20312 11008
rect 20260 10965 20269 10999
rect 20269 10965 20303 10999
rect 20303 10965 20312 10999
rect 20260 10956 20312 10965
rect 4680 10854 4732 10906
rect 4744 10854 4796 10906
rect 4808 10854 4860 10906
rect 4872 10854 4924 10906
rect 12078 10854 12130 10906
rect 12142 10854 12194 10906
rect 12206 10854 12258 10906
rect 12270 10854 12322 10906
rect 19475 10854 19527 10906
rect 19539 10854 19591 10906
rect 19603 10854 19655 10906
rect 19667 10854 19719 10906
rect 1492 10795 1544 10804
rect 1492 10761 1501 10795
rect 1501 10761 1535 10795
rect 1535 10761 1544 10795
rect 1492 10752 1544 10761
rect 1768 10795 1820 10804
rect 1768 10761 1777 10795
rect 1777 10761 1811 10795
rect 1811 10761 1820 10795
rect 1768 10752 1820 10761
rect 4252 10752 4304 10804
rect 5080 10752 5132 10804
rect 5908 10795 5960 10804
rect 5908 10761 5917 10795
rect 5917 10761 5951 10795
rect 5951 10761 5960 10795
rect 5908 10752 5960 10761
rect 4344 10684 4396 10736
rect 4620 10684 4672 10736
rect 7196 10752 7248 10804
rect 8208 10795 8260 10804
rect 8208 10761 8217 10795
rect 8217 10761 8251 10795
rect 8251 10761 8260 10795
rect 8208 10752 8260 10761
rect 7840 10684 7892 10736
rect 10876 10752 10928 10804
rect 11152 10795 11204 10804
rect 11152 10761 11161 10795
rect 11161 10761 11195 10795
rect 11195 10761 11204 10795
rect 11152 10752 11204 10761
rect 11428 10752 11480 10804
rect 9312 10684 9364 10736
rect 1492 10548 1544 10600
rect 1952 10548 2004 10600
rect 4528 10616 4580 10668
rect 5172 10591 5224 10600
rect 4068 10480 4120 10532
rect 2504 10455 2556 10464
rect 2504 10421 2513 10455
rect 2513 10421 2547 10455
rect 2547 10421 2556 10455
rect 2504 10412 2556 10421
rect 4528 10412 4580 10464
rect 5172 10557 5181 10591
rect 5181 10557 5215 10591
rect 5215 10557 5224 10591
rect 5172 10548 5224 10557
rect 5724 10548 5776 10600
rect 9220 10616 9272 10668
rect 6184 10591 6236 10600
rect 6184 10557 6193 10591
rect 6193 10557 6227 10591
rect 6227 10557 6236 10591
rect 6184 10548 6236 10557
rect 6920 10548 6972 10600
rect 7932 10548 7984 10600
rect 9772 10684 9824 10736
rect 17316 10752 17368 10804
rect 17408 10752 17460 10804
rect 18880 10752 18932 10804
rect 19248 10752 19300 10804
rect 21272 10752 21324 10804
rect 5816 10480 5868 10532
rect 8300 10480 8352 10532
rect 6184 10412 6236 10464
rect 6368 10455 6420 10464
rect 6368 10421 6377 10455
rect 6377 10421 6411 10455
rect 6411 10421 6420 10455
rect 6368 10412 6420 10421
rect 8668 10412 8720 10464
rect 8852 10455 8904 10464
rect 8852 10421 8861 10455
rect 8861 10421 8895 10455
rect 8895 10421 8904 10455
rect 8852 10412 8904 10421
rect 9864 10548 9916 10600
rect 10508 10548 10560 10600
rect 10968 10548 11020 10600
rect 11060 10480 11112 10532
rect 14280 10684 14332 10736
rect 16488 10684 16540 10736
rect 18512 10684 18564 10736
rect 12440 10591 12492 10600
rect 12440 10557 12449 10591
rect 12449 10557 12483 10591
rect 12483 10557 12492 10591
rect 12440 10548 12492 10557
rect 14372 10616 14424 10668
rect 14740 10659 14792 10668
rect 14740 10625 14749 10659
rect 14749 10625 14783 10659
rect 14783 10625 14792 10659
rect 14740 10616 14792 10625
rect 16212 10616 16264 10668
rect 17500 10659 17552 10668
rect 12532 10480 12584 10532
rect 13820 10480 13872 10532
rect 15292 10548 15344 10600
rect 15660 10480 15712 10532
rect 14096 10412 14148 10464
rect 14924 10412 14976 10464
rect 15108 10412 15160 10464
rect 16948 10548 17000 10600
rect 17500 10625 17509 10659
rect 17509 10625 17543 10659
rect 17543 10625 17552 10659
rect 17500 10616 17552 10625
rect 17592 10616 17644 10668
rect 19616 10616 19668 10668
rect 23204 10752 23256 10804
rect 21548 10616 21600 10668
rect 18052 10548 18104 10600
rect 19708 10548 19760 10600
rect 19892 10548 19944 10600
rect 16672 10480 16724 10532
rect 18144 10480 18196 10532
rect 18788 10480 18840 10532
rect 21916 10480 21968 10532
rect 16580 10412 16632 10464
rect 16856 10412 16908 10464
rect 17408 10455 17460 10464
rect 17408 10421 17417 10455
rect 17417 10421 17451 10455
rect 17451 10421 17460 10455
rect 17408 10412 17460 10421
rect 17960 10412 18012 10464
rect 19248 10412 19300 10464
rect 20444 10412 20496 10464
rect 21272 10412 21324 10464
rect 21824 10412 21876 10464
rect 22008 10455 22060 10464
rect 22008 10421 22017 10455
rect 22017 10421 22051 10455
rect 22051 10421 22060 10455
rect 22008 10412 22060 10421
rect 8379 10310 8431 10362
rect 8443 10310 8495 10362
rect 8507 10310 8559 10362
rect 8571 10310 8623 10362
rect 15776 10310 15828 10362
rect 15840 10310 15892 10362
rect 15904 10310 15956 10362
rect 15968 10310 16020 10362
rect 2596 10251 2648 10260
rect 2596 10217 2605 10251
rect 2605 10217 2639 10251
rect 2639 10217 2648 10251
rect 2596 10208 2648 10217
rect 3700 10140 3752 10192
rect 4252 10208 4304 10260
rect 4620 10208 4672 10260
rect 7840 10208 7892 10260
rect 8852 10208 8904 10260
rect 9680 10208 9732 10260
rect 11060 10251 11112 10260
rect 2688 10072 2740 10124
rect 4160 10072 4212 10124
rect 7196 10140 7248 10192
rect 8208 10140 8260 10192
rect 11060 10217 11069 10251
rect 11069 10217 11103 10251
rect 11103 10217 11112 10251
rect 11060 10208 11112 10217
rect 11980 10208 12032 10260
rect 15108 10208 15160 10260
rect 15292 10208 15344 10260
rect 17316 10208 17368 10260
rect 6368 10072 6420 10124
rect 9864 10140 9916 10192
rect 10039 10140 10091 10192
rect 11152 10140 11204 10192
rect 3608 10047 3660 10056
rect 3608 10013 3617 10047
rect 3617 10013 3651 10047
rect 3651 10013 3660 10047
rect 3608 10004 3660 10013
rect 5264 10004 5316 10056
rect 5816 10004 5868 10056
rect 9588 10072 9640 10124
rect 4252 9936 4304 9988
rect 2136 9868 2188 9920
rect 3056 9868 3108 9920
rect 5632 9868 5684 9920
rect 6092 9911 6144 9920
rect 6092 9877 6101 9911
rect 6101 9877 6135 9911
rect 6135 9877 6144 9911
rect 6092 9868 6144 9877
rect 6552 9936 6604 9988
rect 6920 10004 6972 10056
rect 9220 10004 9272 10056
rect 13544 10072 13596 10124
rect 15200 10140 15252 10192
rect 14556 10072 14608 10124
rect 15016 10072 15068 10124
rect 15660 10140 15712 10192
rect 16488 10140 16540 10192
rect 16948 10140 17000 10192
rect 19340 10208 19392 10260
rect 20444 10140 20496 10192
rect 21456 10208 21508 10260
rect 21824 10208 21876 10260
rect 22468 10208 22520 10260
rect 23020 10140 23072 10192
rect 12716 10047 12768 10056
rect 12716 10013 12725 10047
rect 12725 10013 12759 10047
rect 12759 10013 12768 10047
rect 12716 10004 12768 10013
rect 14280 10004 14332 10056
rect 7012 9936 7064 9988
rect 9588 9936 9640 9988
rect 10692 9936 10744 9988
rect 14648 10004 14700 10056
rect 15384 10072 15436 10124
rect 17132 10072 17184 10124
rect 17316 10115 17368 10124
rect 17316 10081 17350 10115
rect 17350 10081 17368 10115
rect 17316 10072 17368 10081
rect 18236 10072 18288 10124
rect 18604 10072 18656 10124
rect 18880 10072 18932 10124
rect 19432 10115 19484 10124
rect 19432 10081 19466 10115
rect 19466 10081 19484 10115
rect 11980 9868 12032 9920
rect 12440 9911 12492 9920
rect 12440 9877 12449 9911
rect 12449 9877 12483 9911
rect 12483 9877 12492 9911
rect 12440 9868 12492 9877
rect 12624 9868 12676 9920
rect 15016 9868 15068 9920
rect 18880 9936 18932 9988
rect 19064 9936 19116 9988
rect 16028 9868 16080 9920
rect 18328 9868 18380 9920
rect 18696 9868 18748 9920
rect 19432 10072 19484 10081
rect 20260 10072 20312 10124
rect 20904 10047 20956 10056
rect 20904 10013 20913 10047
rect 20913 10013 20947 10047
rect 20947 10013 20956 10047
rect 20904 10004 20956 10013
rect 22192 9936 22244 9988
rect 22928 9936 22980 9988
rect 4680 9766 4732 9818
rect 4744 9766 4796 9818
rect 4808 9766 4860 9818
rect 4872 9766 4924 9818
rect 12078 9766 12130 9818
rect 12142 9766 12194 9818
rect 12206 9766 12258 9818
rect 12270 9766 12322 9818
rect 19475 9766 19527 9818
rect 19539 9766 19591 9818
rect 19603 9766 19655 9818
rect 19667 9766 19719 9818
rect 4528 9707 4580 9716
rect 4528 9673 4537 9707
rect 4537 9673 4571 9707
rect 4571 9673 4580 9707
rect 4528 9664 4580 9673
rect 2780 9639 2832 9648
rect 2780 9605 2789 9639
rect 2789 9605 2823 9639
rect 2823 9605 2832 9639
rect 2780 9596 2832 9605
rect 7012 9664 7064 9716
rect 4252 9571 4304 9580
rect 4252 9537 4261 9571
rect 4261 9537 4295 9571
rect 4295 9537 4304 9571
rect 4252 9528 4304 9537
rect 5264 9528 5316 9580
rect 6276 9596 6328 9648
rect 9036 9596 9088 9648
rect 9772 9664 9824 9716
rect 10048 9664 10100 9716
rect 1952 9460 2004 9512
rect 2872 9460 2924 9512
rect 4896 9503 4948 9512
rect 4896 9469 4905 9503
rect 4905 9469 4939 9503
rect 4939 9469 4948 9503
rect 4896 9460 4948 9469
rect 5356 9460 5408 9512
rect 6000 9460 6052 9512
rect 7196 9503 7248 9512
rect 7196 9469 7205 9503
rect 7205 9469 7239 9503
rect 7239 9469 7248 9503
rect 7196 9460 7248 9469
rect 1492 9392 1544 9444
rect 5080 9392 5132 9444
rect 10416 9596 10468 9648
rect 8852 9460 8904 9512
rect 8944 9460 8996 9512
rect 14096 9596 14148 9648
rect 15476 9664 15528 9716
rect 17316 9664 17368 9716
rect 18236 9664 18288 9716
rect 11888 9571 11940 9580
rect 11888 9537 11897 9571
rect 11897 9537 11931 9571
rect 11931 9537 11940 9571
rect 11888 9528 11940 9537
rect 12624 9528 12676 9580
rect 14004 9571 14056 9580
rect 14004 9537 14013 9571
rect 14013 9537 14047 9571
rect 14047 9537 14056 9571
rect 14004 9528 14056 9537
rect 17408 9596 17460 9648
rect 16580 9528 16632 9580
rect 16764 9571 16816 9580
rect 16764 9537 16773 9571
rect 16773 9537 16807 9571
rect 16807 9537 16816 9571
rect 16764 9528 16816 9537
rect 18236 9528 18288 9580
rect 18788 9571 18840 9580
rect 18788 9537 18797 9571
rect 18797 9537 18831 9571
rect 18831 9537 18840 9571
rect 18788 9528 18840 9537
rect 19432 9528 19484 9580
rect 20260 9528 20312 9580
rect 20904 9528 20956 9580
rect 12808 9435 12860 9444
rect 3700 9367 3752 9376
rect 3700 9333 3709 9367
rect 3709 9333 3743 9367
rect 3743 9333 3752 9367
rect 3700 9324 3752 9333
rect 4068 9367 4120 9376
rect 4068 9333 4077 9367
rect 4077 9333 4111 9367
rect 4111 9333 4120 9367
rect 4068 9324 4120 9333
rect 5724 9367 5776 9376
rect 5724 9333 5733 9367
rect 5733 9333 5767 9367
rect 5767 9333 5776 9367
rect 5724 9324 5776 9333
rect 7472 9324 7524 9376
rect 7840 9324 7892 9376
rect 8944 9324 8996 9376
rect 12808 9401 12817 9435
rect 12817 9401 12851 9435
rect 12851 9401 12860 9435
rect 12808 9392 12860 9401
rect 13544 9460 13596 9512
rect 13636 9460 13688 9512
rect 14556 9460 14608 9512
rect 14740 9503 14792 9512
rect 14740 9469 14774 9503
rect 14774 9469 14792 9503
rect 14740 9460 14792 9469
rect 15016 9460 15068 9512
rect 12900 9367 12952 9376
rect 12900 9333 12909 9367
rect 12909 9333 12943 9367
rect 12943 9333 12952 9367
rect 12900 9324 12952 9333
rect 13820 9367 13872 9376
rect 13820 9333 13829 9367
rect 13829 9333 13863 9367
rect 13863 9333 13872 9367
rect 13820 9324 13872 9333
rect 15108 9324 15160 9376
rect 15384 9392 15436 9444
rect 17040 9460 17092 9512
rect 16580 9367 16632 9376
rect 16580 9333 16589 9367
rect 16589 9333 16623 9367
rect 16623 9333 16632 9367
rect 16580 9324 16632 9333
rect 17316 9367 17368 9376
rect 17316 9333 17325 9367
rect 17325 9333 17359 9367
rect 17359 9333 17368 9367
rect 17316 9324 17368 9333
rect 18052 9324 18104 9376
rect 19248 9460 19300 9512
rect 20444 9460 20496 9512
rect 22192 9460 22244 9512
rect 18512 9324 18564 9376
rect 18788 9324 18840 9376
rect 19892 9367 19944 9376
rect 19892 9333 19901 9367
rect 19901 9333 19935 9367
rect 19935 9333 19944 9367
rect 19892 9324 19944 9333
rect 8379 9222 8431 9274
rect 8443 9222 8495 9274
rect 8507 9222 8559 9274
rect 8571 9222 8623 9274
rect 15776 9222 15828 9274
rect 15840 9222 15892 9274
rect 15904 9222 15956 9274
rect 15968 9222 16020 9274
rect 3516 9120 3568 9172
rect 4160 9120 4212 9172
rect 5632 9120 5684 9172
rect 6552 9120 6604 9172
rect 7288 9120 7340 9172
rect 7748 9163 7800 9172
rect 7748 9129 7757 9163
rect 7757 9129 7791 9163
rect 7791 9129 7800 9163
rect 7748 9120 7800 9129
rect 8668 9120 8720 9172
rect 9680 9163 9732 9172
rect 6920 9052 6972 9104
rect 7472 9052 7524 9104
rect 3976 8984 4028 9036
rect 4436 8984 4488 9036
rect 5356 8984 5408 9036
rect 7656 8984 7708 9036
rect 8116 8984 8168 9036
rect 9312 9052 9364 9104
rect 9680 9129 9689 9163
rect 9689 9129 9723 9163
rect 9723 9129 9732 9163
rect 9680 9120 9732 9129
rect 10692 9120 10744 9172
rect 10968 9120 11020 9172
rect 12900 9120 12952 9172
rect 13728 9120 13780 9172
rect 14740 9120 14792 9172
rect 15108 9120 15160 9172
rect 15292 9163 15344 9172
rect 15292 9129 15301 9163
rect 15301 9129 15335 9163
rect 15335 9129 15344 9163
rect 15292 9120 15344 9129
rect 15384 9120 15436 9172
rect 16396 9120 16448 9172
rect 16672 9120 16724 9172
rect 19340 9120 19392 9172
rect 21916 9163 21968 9172
rect 21916 9129 21925 9163
rect 21925 9129 21959 9163
rect 21959 9129 21968 9163
rect 21916 9120 21968 9129
rect 10600 9052 10652 9104
rect 11428 9052 11480 9104
rect 11612 9052 11664 9104
rect 9042 9027 9094 9036
rect 9042 8993 9070 9027
rect 9070 8993 9094 9027
rect 9042 8984 9094 8993
rect 9864 8984 9916 9036
rect 10876 8984 10928 9036
rect 4252 8848 4304 8900
rect 7840 8916 7892 8968
rect 10508 8916 10560 8968
rect 10600 8916 10652 8968
rect 8208 8848 8260 8900
rect 9496 8848 9548 8900
rect 11152 8848 11204 8900
rect 12716 9052 12768 9104
rect 13084 8984 13136 9036
rect 14004 9052 14056 9104
rect 14464 9052 14516 9104
rect 13636 8984 13688 9036
rect 13176 8916 13228 8968
rect 14648 8984 14700 9036
rect 17592 9052 17644 9104
rect 18880 9052 18932 9104
rect 21732 9052 21784 9104
rect 15752 8959 15804 8968
rect 15752 8925 15761 8959
rect 15761 8925 15795 8959
rect 15795 8925 15804 8959
rect 15752 8916 15804 8925
rect 16488 8984 16540 9036
rect 5448 8780 5500 8832
rect 8576 8780 8628 8832
rect 10692 8780 10744 8832
rect 13452 8780 13504 8832
rect 15476 8848 15528 8900
rect 15660 8848 15712 8900
rect 16396 8916 16448 8968
rect 17960 8984 18012 9036
rect 18328 8984 18380 9036
rect 20352 8984 20404 9036
rect 18604 8916 18656 8968
rect 20628 8916 20680 8968
rect 21456 8959 21508 8968
rect 21456 8925 21465 8959
rect 21465 8925 21499 8959
rect 21499 8925 21508 8959
rect 22468 8959 22520 8968
rect 21456 8916 21508 8925
rect 22468 8925 22477 8959
rect 22477 8925 22511 8959
rect 22511 8925 22520 8959
rect 22468 8916 22520 8925
rect 16488 8848 16540 8900
rect 17960 8780 18012 8832
rect 20260 8780 20312 8832
rect 22284 8780 22336 8832
rect 4680 8678 4732 8730
rect 4744 8678 4796 8730
rect 4808 8678 4860 8730
rect 4872 8678 4924 8730
rect 12078 8678 12130 8730
rect 12142 8678 12194 8730
rect 12206 8678 12258 8730
rect 12270 8678 12322 8730
rect 19475 8678 19527 8730
rect 19539 8678 19591 8730
rect 19603 8678 19655 8730
rect 19667 8678 19719 8730
rect 4068 8576 4120 8628
rect 4712 8551 4764 8560
rect 4712 8517 4721 8551
rect 4721 8517 4755 8551
rect 4755 8517 4764 8551
rect 4712 8508 4764 8517
rect 1860 8440 1912 8492
rect 5356 8483 5408 8492
rect 5356 8449 5365 8483
rect 5365 8449 5399 8483
rect 5399 8449 5408 8483
rect 5356 8440 5408 8449
rect 1768 8415 1820 8424
rect 1768 8381 1777 8415
rect 1777 8381 1811 8415
rect 1811 8381 1820 8415
rect 1768 8372 1820 8381
rect 8392 8508 8444 8560
rect 6276 8483 6328 8492
rect 6276 8449 6285 8483
rect 6285 8449 6319 8483
rect 6319 8449 6328 8483
rect 6276 8440 6328 8449
rect 7932 8483 7984 8492
rect 7932 8449 7941 8483
rect 7941 8449 7975 8483
rect 7975 8449 7984 8483
rect 7932 8440 7984 8449
rect 11704 8576 11756 8628
rect 11796 8576 11848 8628
rect 12808 8576 12860 8628
rect 13176 8576 13228 8628
rect 15476 8619 15528 8628
rect 13452 8508 13504 8560
rect 6828 8415 6880 8424
rect 6184 8347 6236 8356
rect 6184 8313 6193 8347
rect 6193 8313 6227 8347
rect 6227 8313 6236 8347
rect 6184 8304 6236 8313
rect 6828 8381 6837 8415
rect 6837 8381 6871 8415
rect 6871 8381 6880 8415
rect 6828 8372 6880 8381
rect 12440 8483 12492 8492
rect 12440 8449 12449 8483
rect 12449 8449 12483 8483
rect 12483 8449 12492 8483
rect 12440 8440 12492 8449
rect 13636 8440 13688 8492
rect 15476 8585 15485 8619
rect 15485 8585 15519 8619
rect 15519 8585 15528 8619
rect 15476 8576 15528 8585
rect 15292 8508 15344 8560
rect 18236 8576 18288 8628
rect 18880 8619 18932 8628
rect 18880 8585 18889 8619
rect 18889 8585 18923 8619
rect 18923 8585 18932 8619
rect 18880 8576 18932 8585
rect 18144 8508 18196 8560
rect 10416 8372 10468 8424
rect 10600 8372 10652 8424
rect 7656 8304 7708 8356
rect 5264 8236 5316 8288
rect 7012 8236 7064 8288
rect 8208 8236 8260 8288
rect 10968 8347 11020 8356
rect 10968 8313 11002 8347
rect 11002 8313 11020 8347
rect 11244 8372 11296 8424
rect 15292 8372 15344 8424
rect 15476 8440 15528 8492
rect 16120 8440 16172 8492
rect 16488 8440 16540 8492
rect 16580 8483 16632 8492
rect 16580 8449 16589 8483
rect 16589 8449 16623 8483
rect 16623 8449 16632 8483
rect 16580 8440 16632 8449
rect 18420 8483 18472 8492
rect 18420 8449 18429 8483
rect 18429 8449 18463 8483
rect 18463 8449 18472 8483
rect 19156 8576 19208 8628
rect 19248 8576 19300 8628
rect 22652 8576 22704 8628
rect 22928 8576 22980 8628
rect 19892 8508 19944 8560
rect 18420 8440 18472 8449
rect 19156 8440 19208 8492
rect 19432 8483 19484 8492
rect 19432 8449 19441 8483
rect 19441 8449 19475 8483
rect 19475 8449 19484 8483
rect 19708 8483 19760 8492
rect 19432 8440 19484 8449
rect 19708 8449 19717 8483
rect 19717 8449 19751 8483
rect 19751 8449 19760 8483
rect 19708 8440 19760 8449
rect 20352 8483 20404 8492
rect 20352 8449 20364 8483
rect 20364 8449 20398 8483
rect 20398 8449 20404 8483
rect 20628 8483 20680 8492
rect 20352 8440 20404 8449
rect 20628 8449 20637 8483
rect 20637 8449 20671 8483
rect 20671 8449 20680 8483
rect 20628 8440 20680 8449
rect 22284 8440 22336 8492
rect 22652 8483 22704 8492
rect 22652 8449 22661 8483
rect 22661 8449 22695 8483
rect 22695 8449 22704 8483
rect 22652 8440 22704 8449
rect 17224 8372 17276 8424
rect 17868 8372 17920 8424
rect 10968 8304 11020 8313
rect 9588 8236 9640 8288
rect 10140 8236 10192 8288
rect 12348 8236 12400 8288
rect 12532 8304 12584 8356
rect 15752 8304 15804 8356
rect 15844 8304 15896 8356
rect 13452 8236 13504 8288
rect 15108 8236 15160 8288
rect 16304 8279 16356 8288
rect 16304 8245 16319 8279
rect 16319 8245 16353 8279
rect 16353 8245 16356 8279
rect 16304 8236 16356 8245
rect 17316 8236 17368 8288
rect 17868 8236 17920 8288
rect 18236 8372 18288 8424
rect 19800 8372 19852 8424
rect 18880 8304 18932 8356
rect 22560 8304 22612 8356
rect 18144 8236 18196 8288
rect 18420 8236 18472 8288
rect 21732 8279 21784 8288
rect 21732 8245 21741 8279
rect 21741 8245 21775 8279
rect 21775 8245 21784 8279
rect 21732 8236 21784 8245
rect 22928 8236 22980 8288
rect 8379 8134 8431 8186
rect 8443 8134 8495 8186
rect 8507 8134 8559 8186
rect 8571 8134 8623 8186
rect 15776 8134 15828 8186
rect 15840 8134 15892 8186
rect 15904 8134 15956 8186
rect 15968 8134 16020 8186
rect 4988 8032 5040 8084
rect 5080 8075 5132 8084
rect 5080 8041 5089 8075
rect 5089 8041 5123 8075
rect 5123 8041 5132 8075
rect 5080 8032 5132 8041
rect 6736 8032 6788 8084
rect 9588 8032 9640 8084
rect 12532 8075 12584 8084
rect 1768 7964 1820 8016
rect 4344 7896 4396 7948
rect 7288 7964 7340 8016
rect 6828 7939 6880 7948
rect 6828 7905 6837 7939
rect 6837 7905 6871 7939
rect 6871 7905 6880 7939
rect 6828 7896 6880 7905
rect 9956 7896 10008 7948
rect 7932 7871 7984 7880
rect 7932 7837 7941 7871
rect 7941 7837 7975 7871
rect 7975 7837 7984 7871
rect 7932 7828 7984 7837
rect 9864 7828 9916 7880
rect 10140 7871 10192 7880
rect 10140 7837 10149 7871
rect 10149 7837 10183 7871
rect 10183 7837 10192 7871
rect 10140 7828 10192 7837
rect 10968 7964 11020 8016
rect 11796 7964 11848 8016
rect 12532 8041 12541 8075
rect 12541 8041 12575 8075
rect 12575 8041 12584 8075
rect 12532 8032 12584 8041
rect 13360 8032 13412 8084
rect 14372 8032 14424 8084
rect 14832 8075 14884 8084
rect 14832 8041 14841 8075
rect 14841 8041 14875 8075
rect 14875 8041 14884 8075
rect 14832 8032 14884 8041
rect 15384 8032 15436 8084
rect 16304 8032 16356 8084
rect 16488 8032 16540 8084
rect 12992 7964 13044 8016
rect 10324 7896 10376 7948
rect 10600 7896 10652 7948
rect 11704 7896 11756 7948
rect 17316 7964 17368 8016
rect 13452 7896 13504 7948
rect 13820 7896 13872 7948
rect 15016 7939 15068 7948
rect 5632 7803 5684 7812
rect 5632 7769 5641 7803
rect 5641 7769 5675 7803
rect 5675 7769 5684 7803
rect 5632 7760 5684 7769
rect 8300 7692 8352 7744
rect 9036 7692 9088 7744
rect 9680 7760 9732 7812
rect 10324 7692 10376 7744
rect 12348 7828 12400 7880
rect 12164 7760 12216 7812
rect 12440 7692 12492 7744
rect 12624 7760 12676 7812
rect 13544 7828 13596 7880
rect 15016 7905 15025 7939
rect 15025 7905 15059 7939
rect 15059 7905 15068 7939
rect 15016 7896 15068 7905
rect 15292 7939 15344 7948
rect 15292 7905 15301 7939
rect 15301 7905 15335 7939
rect 15335 7905 15344 7939
rect 15292 7896 15344 7905
rect 17960 7896 18012 7948
rect 18144 7896 18196 7948
rect 18512 7896 18564 7948
rect 18880 7896 18932 7948
rect 20628 8032 20680 8084
rect 22468 7964 22520 8016
rect 20076 7896 20128 7948
rect 20904 7896 20956 7948
rect 14004 7760 14056 7812
rect 15752 7871 15804 7880
rect 15752 7837 15764 7871
rect 15764 7837 15798 7871
rect 15798 7837 15804 7871
rect 15752 7828 15804 7837
rect 16120 7828 16172 7880
rect 16672 7760 16724 7812
rect 17684 7760 17736 7812
rect 18328 7828 18380 7880
rect 19524 7828 19576 7880
rect 20720 7828 20772 7880
rect 20996 7828 21048 7880
rect 18512 7760 18564 7812
rect 13176 7692 13228 7744
rect 14464 7692 14516 7744
rect 14556 7692 14608 7744
rect 16948 7692 17000 7744
rect 18788 7692 18840 7744
rect 18880 7692 18932 7744
rect 21180 7760 21232 7812
rect 22376 7692 22428 7744
rect 4680 7590 4732 7642
rect 4744 7590 4796 7642
rect 4808 7590 4860 7642
rect 4872 7590 4924 7642
rect 12078 7590 12130 7642
rect 12142 7590 12194 7642
rect 12206 7590 12258 7642
rect 12270 7590 12322 7642
rect 19475 7590 19527 7642
rect 19539 7590 19591 7642
rect 19603 7590 19655 7642
rect 19667 7590 19719 7642
rect 5448 7488 5500 7540
rect 7380 7488 7432 7540
rect 8300 7488 8352 7540
rect 9956 7531 10008 7540
rect 9956 7497 9965 7531
rect 9965 7497 9999 7531
rect 9999 7497 10008 7531
rect 9956 7488 10008 7497
rect 11980 7488 12032 7540
rect 15660 7531 15712 7540
rect 5540 7284 5592 7336
rect 6920 7284 6972 7336
rect 11888 7420 11940 7472
rect 8116 7395 8168 7404
rect 8116 7361 8125 7395
rect 8125 7361 8159 7395
rect 8159 7361 8168 7395
rect 8116 7352 8168 7361
rect 9680 7352 9732 7404
rect 10232 7395 10284 7404
rect 10232 7361 10241 7395
rect 10241 7361 10275 7395
rect 10275 7361 10284 7395
rect 10232 7352 10284 7361
rect 11244 7352 11296 7404
rect 7932 7284 7984 7336
rect 6368 7216 6420 7268
rect 10140 7284 10192 7336
rect 10324 7284 10376 7336
rect 11796 7284 11848 7336
rect 13360 7284 13412 7336
rect 14280 7420 14332 7472
rect 15660 7497 15669 7531
rect 15669 7497 15703 7531
rect 15703 7497 15712 7531
rect 15660 7488 15712 7497
rect 17592 7488 17644 7540
rect 18328 7488 18380 7540
rect 22468 7488 22520 7540
rect 18052 7420 18104 7472
rect 19892 7420 19944 7472
rect 14280 7327 14332 7336
rect 14280 7293 14289 7327
rect 14289 7293 14323 7327
rect 14323 7293 14332 7327
rect 14280 7284 14332 7293
rect 14832 7284 14884 7336
rect 8760 7216 8812 7268
rect 9036 7216 9088 7268
rect 12256 7216 12308 7268
rect 15292 7216 15344 7268
rect 18144 7284 18196 7336
rect 6276 7148 6328 7200
rect 8852 7148 8904 7200
rect 8944 7148 8996 7200
rect 12440 7191 12492 7200
rect 12440 7157 12449 7191
rect 12449 7157 12483 7191
rect 12483 7157 12492 7191
rect 12808 7191 12860 7200
rect 12440 7148 12492 7157
rect 12808 7157 12817 7191
rect 12817 7157 12851 7191
rect 12851 7157 12860 7191
rect 12808 7148 12860 7157
rect 13820 7148 13872 7200
rect 17500 7216 17552 7268
rect 18604 7284 18656 7336
rect 20352 7284 20404 7336
rect 20904 7420 20956 7472
rect 20536 7352 20588 7404
rect 20904 7284 20956 7336
rect 22652 7284 22704 7336
rect 16120 7148 16172 7200
rect 21548 7216 21600 7268
rect 22376 7216 22428 7268
rect 19340 7148 19392 7200
rect 19800 7148 19852 7200
rect 21824 7148 21876 7200
rect 8379 7046 8431 7098
rect 8443 7046 8495 7098
rect 8507 7046 8559 7098
rect 8571 7046 8623 7098
rect 15776 7046 15828 7098
rect 15840 7046 15892 7098
rect 15904 7046 15956 7098
rect 15968 7046 16020 7098
rect 7564 6944 7616 6996
rect 9588 6944 9640 6996
rect 13268 6944 13320 6996
rect 6460 6851 6512 6860
rect 6460 6817 6469 6851
rect 6469 6817 6503 6851
rect 6503 6817 6512 6851
rect 6460 6808 6512 6817
rect 9036 6919 9088 6928
rect 9036 6885 9045 6919
rect 9045 6885 9079 6919
rect 9079 6885 9088 6919
rect 9036 6876 9088 6885
rect 10968 6876 11020 6928
rect 12716 6919 12768 6928
rect 8944 6851 8996 6860
rect 3700 6740 3752 6792
rect 8300 6740 8352 6792
rect 8944 6817 8953 6851
rect 8953 6817 8987 6851
rect 8987 6817 8996 6851
rect 8944 6808 8996 6817
rect 9772 6808 9824 6860
rect 9956 6851 10008 6860
rect 9956 6817 9990 6851
rect 9990 6817 10008 6851
rect 9956 6808 10008 6817
rect 11612 6808 11664 6860
rect 12716 6885 12725 6919
rect 12725 6885 12759 6919
rect 12759 6885 12768 6919
rect 12716 6876 12768 6885
rect 12900 6876 12952 6928
rect 16948 6944 17000 6996
rect 13820 6876 13872 6928
rect 16304 6876 16356 6928
rect 9496 6740 9548 6792
rect 9680 6783 9732 6792
rect 9680 6749 9689 6783
rect 9689 6749 9723 6783
rect 9723 6749 9732 6783
rect 9680 6740 9732 6749
rect 10692 6740 10744 6792
rect 11060 6740 11112 6792
rect 11152 6740 11204 6792
rect 7564 6715 7616 6724
rect 7564 6681 7573 6715
rect 7573 6681 7607 6715
rect 7607 6681 7616 6715
rect 7564 6672 7616 6681
rect 5356 6604 5408 6656
rect 6644 6647 6696 6656
rect 6644 6613 6653 6647
rect 6653 6613 6687 6647
rect 6687 6613 6696 6647
rect 6644 6604 6696 6613
rect 8484 6672 8536 6724
rect 8668 6672 8720 6724
rect 8760 6672 8812 6724
rect 8208 6604 8260 6656
rect 12256 6672 12308 6724
rect 12624 6740 12676 6792
rect 13544 6808 13596 6860
rect 14556 6851 14608 6860
rect 14556 6817 14565 6851
rect 14565 6817 14599 6851
rect 14599 6817 14608 6851
rect 14556 6808 14608 6817
rect 15568 6851 15620 6860
rect 15568 6817 15602 6851
rect 15602 6817 15620 6851
rect 15568 6808 15620 6817
rect 13084 6740 13136 6792
rect 14004 6783 14056 6792
rect 14004 6749 14013 6783
rect 14013 6749 14047 6783
rect 14047 6749 14056 6783
rect 14004 6740 14056 6749
rect 15016 6740 15068 6792
rect 16672 6876 16724 6928
rect 17408 6876 17460 6928
rect 19340 6944 19392 6996
rect 22652 6944 22704 6996
rect 20260 6876 20312 6928
rect 16764 6808 16816 6860
rect 17500 6808 17552 6860
rect 20168 6851 20220 6860
rect 18604 6740 18656 6792
rect 20168 6817 20177 6851
rect 20177 6817 20211 6851
rect 20211 6817 20220 6851
rect 20168 6808 20220 6817
rect 21456 6808 21508 6860
rect 22560 6851 22612 6860
rect 22560 6817 22569 6851
rect 22569 6817 22603 6851
rect 22603 6817 22612 6851
rect 22560 6808 22612 6817
rect 23388 6851 23440 6860
rect 23388 6817 23397 6851
rect 23397 6817 23431 6851
rect 23431 6817 23440 6851
rect 23388 6808 23440 6817
rect 20260 6783 20312 6792
rect 20260 6749 20269 6783
rect 20269 6749 20303 6783
rect 20303 6749 20312 6783
rect 20260 6740 20312 6749
rect 20904 6783 20956 6792
rect 16764 6672 16816 6724
rect 17960 6672 18012 6724
rect 11060 6647 11112 6656
rect 11060 6613 11069 6647
rect 11069 6613 11103 6647
rect 11103 6613 11112 6647
rect 11060 6604 11112 6613
rect 11336 6647 11388 6656
rect 11336 6613 11345 6647
rect 11345 6613 11379 6647
rect 11379 6613 11388 6647
rect 11336 6604 11388 6613
rect 13360 6647 13412 6656
rect 13360 6613 13369 6647
rect 13369 6613 13403 6647
rect 13403 6613 13412 6647
rect 13360 6604 13412 6613
rect 14096 6604 14148 6656
rect 17132 6604 17184 6656
rect 17592 6604 17644 6656
rect 18788 6647 18840 6656
rect 18788 6613 18797 6647
rect 18797 6613 18831 6647
rect 18831 6613 18840 6647
rect 18788 6604 18840 6613
rect 19064 6672 19116 6724
rect 20904 6749 20913 6783
rect 20913 6749 20947 6783
rect 20947 6749 20956 6783
rect 20904 6740 20956 6749
rect 20720 6604 20772 6656
rect 4680 6502 4732 6554
rect 4744 6502 4796 6554
rect 4808 6502 4860 6554
rect 4872 6502 4924 6554
rect 12078 6502 12130 6554
rect 12142 6502 12194 6554
rect 12206 6502 12258 6554
rect 12270 6502 12322 6554
rect 19475 6502 19527 6554
rect 19539 6502 19591 6554
rect 19603 6502 19655 6554
rect 19667 6502 19719 6554
rect 7104 6400 7156 6452
rect 8300 6400 8352 6452
rect 8668 6332 8720 6384
rect 9956 6400 10008 6452
rect 10600 6332 10652 6384
rect 8760 6307 8812 6316
rect 8760 6273 8769 6307
rect 8769 6273 8803 6307
rect 8803 6273 8812 6307
rect 8760 6264 8812 6273
rect 10876 6400 10928 6452
rect 10968 6307 11020 6316
rect 10968 6273 10977 6307
rect 10977 6273 11011 6307
rect 11011 6273 11020 6307
rect 10968 6264 11020 6273
rect 12348 6264 12400 6316
rect 8208 6239 8260 6248
rect 8208 6205 8217 6239
rect 8217 6205 8251 6239
rect 8251 6205 8260 6239
rect 8208 6196 8260 6205
rect 10416 6196 10468 6248
rect 11060 6196 11112 6248
rect 11520 6196 11572 6248
rect 12256 6196 12308 6248
rect 8944 6128 8996 6180
rect 13360 6128 13412 6180
rect 13728 6128 13780 6180
rect 13820 6128 13872 6180
rect 14556 6400 14608 6452
rect 15292 6400 15344 6452
rect 15660 6400 15712 6452
rect 18236 6400 18288 6452
rect 20444 6400 20496 6452
rect 21456 6400 21508 6452
rect 14372 6196 14424 6248
rect 18696 6332 18748 6384
rect 10416 6103 10468 6112
rect 10416 6069 10425 6103
rect 10425 6069 10459 6103
rect 10459 6069 10468 6103
rect 10416 6060 10468 6069
rect 11244 6060 11296 6112
rect 17408 6264 17460 6316
rect 17684 6196 17736 6248
rect 18144 6264 18196 6316
rect 19064 6307 19116 6316
rect 19064 6273 19073 6307
rect 19073 6273 19107 6307
rect 19107 6273 19116 6307
rect 19064 6264 19116 6273
rect 21824 6264 21876 6316
rect 20904 6196 20956 6248
rect 22008 6196 22060 6248
rect 19064 6128 19116 6180
rect 19248 6128 19300 6180
rect 21916 6171 21968 6180
rect 21916 6137 21925 6171
rect 21925 6137 21959 6171
rect 21959 6137 21968 6171
rect 21916 6128 21968 6137
rect 17316 6103 17368 6112
rect 17316 6069 17325 6103
rect 17325 6069 17359 6103
rect 17359 6069 17368 6103
rect 17316 6060 17368 6069
rect 17960 6060 18012 6112
rect 18420 6060 18472 6112
rect 18604 6060 18656 6112
rect 18880 6103 18932 6112
rect 18880 6069 18889 6103
rect 18889 6069 18923 6103
rect 18923 6069 18932 6103
rect 18880 6060 18932 6069
rect 20996 6060 21048 6112
rect 22008 6103 22060 6112
rect 22008 6069 22017 6103
rect 22017 6069 22051 6103
rect 22051 6069 22060 6103
rect 22008 6060 22060 6069
rect 8379 5958 8431 6010
rect 8443 5958 8495 6010
rect 8507 5958 8559 6010
rect 8571 5958 8623 6010
rect 15776 5958 15828 6010
rect 15840 5958 15892 6010
rect 15904 5958 15956 6010
rect 15968 5958 16020 6010
rect 8024 5856 8076 5908
rect 12348 5856 12400 5908
rect 13636 5856 13688 5908
rect 13728 5856 13780 5908
rect 6644 5720 6696 5772
rect 9772 5720 9824 5772
rect 11060 5720 11112 5772
rect 11612 5763 11664 5772
rect 11612 5729 11646 5763
rect 11646 5729 11664 5763
rect 11612 5720 11664 5729
rect 12532 5720 12584 5772
rect 13728 5720 13780 5772
rect 17224 5856 17276 5908
rect 17500 5899 17552 5908
rect 17500 5865 17509 5899
rect 17509 5865 17543 5899
rect 17543 5865 17552 5899
rect 17500 5856 17552 5865
rect 19248 5856 19300 5908
rect 9680 5695 9732 5704
rect 7656 5584 7708 5636
rect 9680 5661 9689 5695
rect 9689 5661 9723 5695
rect 9723 5661 9732 5695
rect 9680 5652 9732 5661
rect 11244 5652 11296 5704
rect 16120 5695 16172 5704
rect 16120 5661 16129 5695
rect 16129 5661 16163 5695
rect 16163 5661 16172 5695
rect 16120 5652 16172 5661
rect 17684 5720 17736 5772
rect 18696 5720 18748 5772
rect 19064 5763 19116 5772
rect 19064 5729 19098 5763
rect 19098 5729 19116 5763
rect 19064 5720 19116 5729
rect 20444 5788 20496 5840
rect 22560 5831 22612 5840
rect 20904 5720 20956 5772
rect 21548 5720 21600 5772
rect 22560 5797 22569 5831
rect 22569 5797 22603 5831
rect 22603 5797 22612 5831
rect 22560 5788 22612 5797
rect 17776 5652 17828 5704
rect 18328 5695 18380 5704
rect 18328 5661 18337 5695
rect 18337 5661 18371 5695
rect 18371 5661 18380 5695
rect 18328 5652 18380 5661
rect 21732 5695 21784 5704
rect 21732 5661 21741 5695
rect 21741 5661 21775 5695
rect 21775 5661 21784 5695
rect 21732 5652 21784 5661
rect 21824 5695 21876 5704
rect 21824 5661 21833 5695
rect 21833 5661 21867 5695
rect 21867 5661 21876 5695
rect 21824 5652 21876 5661
rect 11152 5584 11204 5636
rect 12624 5584 12676 5636
rect 14096 5584 14148 5636
rect 14556 5584 14608 5636
rect 16028 5584 16080 5636
rect 11980 5516 12032 5568
rect 12532 5516 12584 5568
rect 14372 5516 14424 5568
rect 18512 5516 18564 5568
rect 20444 5584 20496 5636
rect 20168 5516 20220 5568
rect 20812 5516 20864 5568
rect 4680 5414 4732 5466
rect 4744 5414 4796 5466
rect 4808 5414 4860 5466
rect 4872 5414 4924 5466
rect 12078 5414 12130 5466
rect 12142 5414 12194 5466
rect 12206 5414 12258 5466
rect 12270 5414 12322 5466
rect 19475 5414 19527 5466
rect 19539 5414 19591 5466
rect 19603 5414 19655 5466
rect 19667 5414 19719 5466
rect 11612 5312 11664 5364
rect 15108 5355 15160 5364
rect 15108 5321 15117 5355
rect 15117 5321 15151 5355
rect 15151 5321 15160 5355
rect 15108 5312 15160 5321
rect 16028 5312 16080 5364
rect 17684 5355 17736 5364
rect 13728 5244 13780 5296
rect 14372 5244 14424 5296
rect 9404 5151 9456 5160
rect 9404 5117 9413 5151
rect 9413 5117 9447 5151
rect 9447 5117 9456 5151
rect 9404 5108 9456 5117
rect 9680 5108 9732 5160
rect 11152 5108 11204 5160
rect 12256 5108 12308 5160
rect 11244 5040 11296 5092
rect 8944 5015 8996 5024
rect 8944 4981 8953 5015
rect 8953 4981 8987 5015
rect 8987 4981 8996 5015
rect 8944 4972 8996 4981
rect 12348 4972 12400 5024
rect 13912 5176 13964 5228
rect 14464 5176 14516 5228
rect 15660 5219 15712 5228
rect 15660 5185 15669 5219
rect 15669 5185 15703 5219
rect 15703 5185 15712 5219
rect 15660 5176 15712 5185
rect 16304 5219 16356 5228
rect 16304 5185 16313 5219
rect 16313 5185 16347 5219
rect 16347 5185 16356 5219
rect 16304 5176 16356 5185
rect 17684 5321 17693 5355
rect 17693 5321 17727 5355
rect 17727 5321 17736 5355
rect 17684 5312 17736 5321
rect 18052 5355 18104 5364
rect 18052 5321 18061 5355
rect 18061 5321 18095 5355
rect 18095 5321 18104 5355
rect 18052 5312 18104 5321
rect 18144 5312 18196 5364
rect 19800 5312 19852 5364
rect 20904 5312 20956 5364
rect 17592 5244 17644 5296
rect 18328 5176 18380 5228
rect 18512 5219 18564 5228
rect 18512 5185 18521 5219
rect 18521 5185 18555 5219
rect 18555 5185 18564 5219
rect 18512 5176 18564 5185
rect 12716 5151 12768 5160
rect 12716 5117 12750 5151
rect 12750 5117 12768 5151
rect 12716 5108 12768 5117
rect 13820 5108 13872 5160
rect 16396 5108 16448 5160
rect 17500 5108 17552 5160
rect 17868 5108 17920 5160
rect 19616 5176 19668 5228
rect 20812 5219 20864 5228
rect 20812 5185 20821 5219
rect 20821 5185 20855 5219
rect 20855 5185 20864 5219
rect 20812 5176 20864 5185
rect 20904 5219 20956 5228
rect 20904 5185 20913 5219
rect 20913 5185 20947 5219
rect 20947 5185 20956 5219
rect 20904 5176 20956 5185
rect 18696 5108 18748 5160
rect 20628 5108 20680 5160
rect 20996 5108 21048 5160
rect 21180 5108 21232 5160
rect 13084 5040 13136 5092
rect 14188 5040 14240 5092
rect 15660 5040 15712 5092
rect 18880 5040 18932 5092
rect 19064 5040 19116 5092
rect 12532 4972 12584 5024
rect 13820 4972 13872 5024
rect 14464 5015 14516 5024
rect 14464 4981 14473 5015
rect 14473 4981 14507 5015
rect 14507 4981 14516 5015
rect 14464 4972 14516 4981
rect 14556 4972 14608 5024
rect 18420 5015 18472 5024
rect 18420 4981 18429 5015
rect 18429 4981 18463 5015
rect 18463 4981 18472 5015
rect 18420 4972 18472 4981
rect 19616 5015 19668 5024
rect 19616 4981 19625 5015
rect 19625 4981 19659 5015
rect 19659 4981 19668 5015
rect 19616 4972 19668 4981
rect 19800 4972 19852 5024
rect 20904 5040 20956 5092
rect 21640 5083 21692 5092
rect 21640 5049 21652 5083
rect 21652 5049 21692 5083
rect 21640 5040 21692 5049
rect 8379 4870 8431 4922
rect 8443 4870 8495 4922
rect 8507 4870 8559 4922
rect 8571 4870 8623 4922
rect 15776 4870 15828 4922
rect 15840 4870 15892 4922
rect 15904 4870 15956 4922
rect 15968 4870 16020 4922
rect 9404 4768 9456 4820
rect 10416 4768 10468 4820
rect 11520 4768 11572 4820
rect 12716 4811 12768 4820
rect 12716 4777 12725 4811
rect 12725 4777 12759 4811
rect 12759 4777 12768 4811
rect 12716 4768 12768 4777
rect 12808 4768 12860 4820
rect 13360 4811 13412 4820
rect 13360 4777 13369 4811
rect 13369 4777 13403 4811
rect 13403 4777 13412 4811
rect 13360 4768 13412 4777
rect 13728 4768 13780 4820
rect 14372 4811 14424 4820
rect 14372 4777 14381 4811
rect 14381 4777 14415 4811
rect 14415 4777 14424 4811
rect 14372 4768 14424 4777
rect 15660 4768 15712 4820
rect 11336 4700 11388 4752
rect 12624 4700 12676 4752
rect 17224 4768 17276 4820
rect 18420 4768 18472 4820
rect 19616 4768 19668 4820
rect 21640 4768 21692 4820
rect 17684 4700 17736 4752
rect 18328 4700 18380 4752
rect 18972 4700 19024 4752
rect 15292 4675 15344 4684
rect 11244 4564 11296 4616
rect 12348 4564 12400 4616
rect 13452 4564 13504 4616
rect 13544 4607 13596 4616
rect 13544 4573 13553 4607
rect 13553 4573 13587 4607
rect 13587 4573 13596 4607
rect 15292 4641 15301 4675
rect 15301 4641 15335 4675
rect 15335 4641 15344 4675
rect 15292 4632 15344 4641
rect 13544 4564 13596 4573
rect 14648 4607 14700 4616
rect 14648 4573 14657 4607
rect 14657 4573 14691 4607
rect 14691 4573 14700 4607
rect 14648 4564 14700 4573
rect 15660 4564 15712 4616
rect 15936 4632 15988 4684
rect 17132 4632 17184 4684
rect 18144 4632 18196 4684
rect 13176 4496 13228 4548
rect 8944 4428 8996 4480
rect 13360 4428 13412 4480
rect 16580 4428 16632 4480
rect 18328 4564 18380 4616
rect 20720 4700 20772 4752
rect 20812 4632 20864 4684
rect 21916 4632 21968 4684
rect 20168 4607 20220 4616
rect 17408 4496 17460 4548
rect 20168 4573 20177 4607
rect 20177 4573 20211 4607
rect 20211 4573 20220 4607
rect 20168 4564 20220 4573
rect 20996 4564 21048 4616
rect 21180 4564 21232 4616
rect 20352 4496 20404 4548
rect 17960 4428 18012 4480
rect 18696 4428 18748 4480
rect 20628 4428 20680 4480
rect 4680 4326 4732 4378
rect 4744 4326 4796 4378
rect 4808 4326 4860 4378
rect 4872 4326 4924 4378
rect 12078 4326 12130 4378
rect 12142 4326 12194 4378
rect 12206 4326 12258 4378
rect 12270 4326 12322 4378
rect 19475 4326 19527 4378
rect 19539 4326 19591 4378
rect 19603 4326 19655 4378
rect 19667 4326 19719 4378
rect 8116 4224 8168 4276
rect 11428 4156 11480 4208
rect 6920 4088 6972 4140
rect 13360 4224 13412 4276
rect 17132 4267 17184 4276
rect 13452 4156 13504 4208
rect 17132 4233 17141 4267
rect 17141 4233 17175 4267
rect 17175 4233 17184 4267
rect 17132 4224 17184 4233
rect 17224 4224 17276 4276
rect 19064 4224 19116 4276
rect 19800 4224 19852 4276
rect 10784 4063 10836 4072
rect 10784 4029 10793 4063
rect 10793 4029 10827 4063
rect 10827 4029 10836 4063
rect 10784 4020 10836 4029
rect 11704 4063 11756 4072
rect 11704 4029 11713 4063
rect 11713 4029 11747 4063
rect 11747 4029 11756 4063
rect 11704 4020 11756 4029
rect 14280 4131 14332 4140
rect 14280 4097 14289 4131
rect 14289 4097 14323 4131
rect 14323 4097 14332 4131
rect 14280 4088 14332 4097
rect 15016 4088 15068 4140
rect 17868 4156 17920 4208
rect 20352 4156 20404 4208
rect 13176 4063 13228 4072
rect 7288 3952 7340 4004
rect 5172 3884 5224 3936
rect 11612 3952 11664 4004
rect 13176 4029 13185 4063
rect 13185 4029 13219 4063
rect 13219 4029 13228 4063
rect 13176 4020 13228 4029
rect 14740 4020 14792 4072
rect 15200 4020 15252 4072
rect 15660 4020 15712 4072
rect 16580 4020 16632 4072
rect 17500 4020 17552 4072
rect 17776 4020 17828 4072
rect 12808 3952 12860 4004
rect 14556 3952 14608 4004
rect 13176 3884 13228 3936
rect 15292 3952 15344 4004
rect 17960 3952 18012 4004
rect 17316 3884 17368 3936
rect 18604 4020 18656 4072
rect 19248 4020 19300 4072
rect 18880 3952 18932 4004
rect 20536 4020 20588 4072
rect 20904 4063 20956 4072
rect 20904 4029 20913 4063
rect 20913 4029 20947 4063
rect 20947 4029 20956 4063
rect 20904 4020 20956 4029
rect 20996 4020 21048 4072
rect 22008 4020 22060 4072
rect 21824 3952 21876 4004
rect 19064 3884 19116 3936
rect 19432 3927 19484 3936
rect 19432 3893 19441 3927
rect 19441 3893 19475 3927
rect 19475 3893 19484 3927
rect 19432 3884 19484 3893
rect 20444 3884 20496 3936
rect 21916 3884 21968 3936
rect 8379 3782 8431 3834
rect 8443 3782 8495 3834
rect 8507 3782 8559 3834
rect 8571 3782 8623 3834
rect 15776 3782 15828 3834
rect 15840 3782 15892 3834
rect 15904 3782 15956 3834
rect 15968 3782 16020 3834
rect 10324 3680 10376 3732
rect 12808 3723 12860 3732
rect 12808 3689 12817 3723
rect 12817 3689 12851 3723
rect 12851 3689 12860 3723
rect 12808 3680 12860 3689
rect 3884 3612 3936 3664
rect 1768 3476 1820 3528
rect 12440 3544 12492 3596
rect 13636 3612 13688 3664
rect 13544 3587 13596 3596
rect 13544 3553 13553 3587
rect 13553 3553 13587 3587
rect 13587 3553 13596 3587
rect 13544 3544 13596 3553
rect 12072 3476 12124 3528
rect 13636 3519 13688 3528
rect 12808 3408 12860 3460
rect 2504 3340 2556 3392
rect 11612 3340 11664 3392
rect 11980 3340 12032 3392
rect 13636 3485 13645 3519
rect 13645 3485 13679 3519
rect 13679 3485 13688 3519
rect 13636 3476 13688 3485
rect 16948 3680 17000 3732
rect 18880 3723 18932 3732
rect 18880 3689 18889 3723
rect 18889 3689 18923 3723
rect 18923 3689 18932 3723
rect 18880 3680 18932 3689
rect 21548 3680 21600 3732
rect 14924 3612 14976 3664
rect 17132 3612 17184 3664
rect 19432 3655 19484 3664
rect 19432 3621 19466 3655
rect 19466 3621 19484 3655
rect 19432 3612 19484 3621
rect 21732 3612 21784 3664
rect 14832 3544 14884 3596
rect 17592 3544 17644 3596
rect 17776 3587 17828 3596
rect 17776 3553 17810 3587
rect 17810 3553 17828 3587
rect 17776 3544 17828 3553
rect 19064 3544 19116 3596
rect 14280 3476 14332 3528
rect 15568 3476 15620 3528
rect 15660 3476 15712 3528
rect 17500 3519 17552 3528
rect 17500 3485 17509 3519
rect 17509 3485 17543 3519
rect 17543 3485 17552 3519
rect 17500 3476 17552 3485
rect 20904 3519 20956 3528
rect 20904 3485 20913 3519
rect 20913 3485 20947 3519
rect 20947 3485 20956 3519
rect 20904 3476 20956 3485
rect 12992 3408 13044 3460
rect 17408 3408 17460 3460
rect 14372 3340 14424 3392
rect 20260 3340 20312 3392
rect 20444 3340 20496 3392
rect 4680 3238 4732 3290
rect 4744 3238 4796 3290
rect 4808 3238 4860 3290
rect 4872 3238 4924 3290
rect 12078 3238 12130 3290
rect 12142 3238 12194 3290
rect 12206 3238 12258 3290
rect 12270 3238 12322 3290
rect 19475 3238 19527 3290
rect 19539 3238 19591 3290
rect 19603 3238 19655 3290
rect 19667 3238 19719 3290
rect 13084 3179 13136 3188
rect 13084 3145 13093 3179
rect 13093 3145 13127 3179
rect 13127 3145 13136 3179
rect 13084 3136 13136 3145
rect 13636 3136 13688 3188
rect 2596 3068 2648 3120
rect 1952 3043 2004 3052
rect 1952 3009 1961 3043
rect 1961 3009 1995 3043
rect 1995 3009 2004 3043
rect 1952 3000 2004 3009
rect 15476 3000 15528 3052
rect 15568 3043 15620 3052
rect 15568 3009 15577 3043
rect 15577 3009 15611 3043
rect 15611 3009 15620 3043
rect 16396 3136 16448 3188
rect 18144 3136 18196 3188
rect 20168 3136 20220 3188
rect 21732 3136 21784 3188
rect 17500 3068 17552 3120
rect 18052 3068 18104 3120
rect 15568 3000 15620 3009
rect 1768 2975 1820 2984
rect 1768 2941 1777 2975
rect 1777 2941 1811 2975
rect 1811 2941 1820 2975
rect 1768 2932 1820 2941
rect 2504 2975 2556 2984
rect 2504 2941 2513 2975
rect 2513 2941 2547 2975
rect 2547 2941 2556 2975
rect 2504 2932 2556 2941
rect 5080 2975 5132 2984
rect 5080 2941 5089 2975
rect 5089 2941 5123 2975
rect 5123 2941 5132 2975
rect 5080 2932 5132 2941
rect 11888 2932 11940 2984
rect 13912 2932 13964 2984
rect 16120 2932 16172 2984
rect 17408 2932 17460 2984
rect 18788 2932 18840 2984
rect 2136 2864 2188 2916
rect 17040 2864 17092 2916
rect 20444 2932 20496 2984
rect 20812 2975 20864 2984
rect 20812 2941 20846 2975
rect 20846 2941 20864 2975
rect 19064 2864 19116 2916
rect 20812 2932 20864 2941
rect 22100 2932 22152 2984
rect 20904 2864 20956 2916
rect 22560 2864 22612 2916
rect 1676 2796 1728 2848
rect 7012 2796 7064 2848
rect 12992 2796 13044 2848
rect 14188 2796 14240 2848
rect 14464 2839 14516 2848
rect 14464 2805 14473 2839
rect 14473 2805 14507 2839
rect 14507 2805 14516 2839
rect 14464 2796 14516 2805
rect 17684 2796 17736 2848
rect 22744 2796 22796 2848
rect 8379 2694 8431 2746
rect 8443 2694 8495 2746
rect 8507 2694 8559 2746
rect 8571 2694 8623 2746
rect 15776 2694 15828 2746
rect 15840 2694 15892 2746
rect 15904 2694 15956 2746
rect 15968 2694 16020 2746
rect 14372 2592 14424 2644
rect 14464 2524 14516 2576
rect 15568 2524 15620 2576
rect 3056 2456 3108 2508
rect 15936 2499 15988 2508
rect 15936 2465 15945 2499
rect 15945 2465 15979 2499
rect 15979 2465 15988 2499
rect 15936 2456 15988 2465
rect 14832 2431 14884 2440
rect 14832 2397 14841 2431
rect 14841 2397 14875 2431
rect 14875 2397 14884 2431
rect 14832 2388 14884 2397
rect 15016 2431 15068 2440
rect 15016 2397 15025 2431
rect 15025 2397 15059 2431
rect 15059 2397 15068 2431
rect 15016 2388 15068 2397
rect 16396 2456 16448 2508
rect 17776 2592 17828 2644
rect 18144 2524 18196 2576
rect 18880 2592 18932 2644
rect 20168 2524 20220 2576
rect 20812 2592 20864 2644
rect 21824 2592 21876 2644
rect 21088 2524 21140 2576
rect 21640 2524 21692 2576
rect 19064 2456 19116 2508
rect 20904 2456 20956 2508
rect 18972 2431 19024 2440
rect 18972 2397 18981 2431
rect 18981 2397 19015 2431
rect 19015 2397 19024 2431
rect 18972 2388 19024 2397
rect 6184 2320 6236 2372
rect 9864 2252 9916 2304
rect 15200 2252 15252 2304
rect 4680 2150 4732 2202
rect 4744 2150 4796 2202
rect 4808 2150 4860 2202
rect 4872 2150 4924 2202
rect 12078 2150 12130 2202
rect 12142 2150 12194 2202
rect 12206 2150 12258 2202
rect 12270 2150 12322 2202
rect 19475 2150 19527 2202
rect 19539 2150 19591 2202
rect 19603 2150 19655 2202
rect 19667 2150 19719 2202
rect 14832 2048 14884 2100
rect 19984 2048 20036 2100
rect 15016 1980 15068 2032
rect 21456 1980 21508 2032
rect 16856 1912 16908 1964
rect 19892 1912 19944 1964
<< metal2 >>
rect 294 23600 350 24400
rect 846 23600 902 24400
rect 1490 23600 1546 24400
rect 2134 23600 2190 24400
rect 2778 23600 2834 24400
rect 3422 23600 3478 24400
rect 4066 23600 4122 24400
rect 4710 23600 4766 24400
rect 5354 23600 5410 24400
rect 5998 23600 6054 24400
rect 6642 23600 6698 24400
rect 7286 23600 7342 24400
rect 7930 23600 7986 24400
rect 8574 23600 8630 24400
rect 9218 23600 9274 24400
rect 9862 23600 9918 24400
rect 10506 23600 10562 24400
rect 11150 23600 11206 24400
rect 11794 23600 11850 24400
rect 12438 23610 12494 24400
rect 13082 23610 13138 24400
rect 12438 23600 12664 23610
rect 13082 23600 13676 23610
rect 13726 23600 13782 24400
rect 14370 23610 14426 24400
rect 14370 23600 14596 23610
rect 15014 23600 15070 24400
rect 15658 23600 15714 24400
rect 16302 23600 16358 24400
rect 16946 23600 17002 24400
rect 17590 23600 17646 24400
rect 18234 23600 18290 24400
rect 18878 23600 18934 24400
rect 19430 24032 19486 24041
rect 19430 23967 19486 23976
rect 308 21146 336 23600
rect 296 21140 348 21146
rect 296 21082 348 21088
rect 860 20602 888 23600
rect 1400 21344 1452 21350
rect 1400 21286 1452 21292
rect 848 20596 900 20602
rect 848 20538 900 20544
rect 1412 14958 1440 21286
rect 1504 19446 1532 23600
rect 2044 21956 2096 21962
rect 2044 21898 2096 21904
rect 1584 21412 1636 21418
rect 1584 21354 1636 21360
rect 1492 19440 1544 19446
rect 1492 19382 1544 19388
rect 1596 19174 1624 21354
rect 2056 21010 2084 21898
rect 2044 21004 2096 21010
rect 2044 20946 2096 20952
rect 2148 20262 2176 23600
rect 2792 22250 2820 23600
rect 2792 22222 2912 22250
rect 2884 21486 2912 22222
rect 3056 21548 3108 21554
rect 3056 21490 3108 21496
rect 2872 21480 2924 21486
rect 2872 21422 2924 21428
rect 2228 21344 2280 21350
rect 2228 21286 2280 21292
rect 2136 20256 2188 20262
rect 2136 20198 2188 20204
rect 1860 19984 1912 19990
rect 1860 19926 1912 19932
rect 1676 19916 1728 19922
rect 1676 19858 1728 19864
rect 1584 19168 1636 19174
rect 1584 19110 1636 19116
rect 1688 18834 1716 19858
rect 1872 19825 1900 19926
rect 1858 19816 1914 19825
rect 1858 19751 1914 19760
rect 2240 19310 2268 21286
rect 2780 20800 2832 20806
rect 2780 20742 2832 20748
rect 3068 20754 3096 21490
rect 3148 21344 3200 21350
rect 3148 21286 3200 21292
rect 3240 21344 3292 21350
rect 3240 21286 3292 21292
rect 3160 21146 3188 21286
rect 3148 21140 3200 21146
rect 3148 21082 3200 21088
rect 3252 21010 3280 21286
rect 3240 21004 3292 21010
rect 3240 20946 3292 20952
rect 2792 20398 2820 20742
rect 3068 20726 3188 20754
rect 3056 20596 3108 20602
rect 3056 20538 3108 20544
rect 2780 20392 2832 20398
rect 2780 20334 2832 20340
rect 2964 20324 3016 20330
rect 2964 20266 3016 20272
rect 2976 20058 3004 20266
rect 3068 20058 3096 20538
rect 2964 20052 3016 20058
rect 2964 19994 3016 20000
rect 3056 20052 3108 20058
rect 3056 19994 3108 20000
rect 2778 19816 2834 19825
rect 2778 19751 2834 19760
rect 2228 19304 2280 19310
rect 2228 19246 2280 19252
rect 1952 19168 2004 19174
rect 1952 19110 2004 19116
rect 1964 18902 1992 19110
rect 2792 18970 2820 19751
rect 3056 19440 3108 19446
rect 3056 19382 3108 19388
rect 2872 19168 2924 19174
rect 2872 19110 2924 19116
rect 2780 18964 2832 18970
rect 2780 18906 2832 18912
rect 1952 18896 2004 18902
rect 1952 18838 2004 18844
rect 1676 18828 1728 18834
rect 1676 18770 1728 18776
rect 1688 18204 1716 18770
rect 1768 18216 1820 18222
rect 1688 18176 1768 18204
rect 1820 18176 1900 18204
rect 1768 18158 1820 18164
rect 1872 17746 1900 18176
rect 1860 17740 1912 17746
rect 1860 17682 1912 17688
rect 1768 17536 1820 17542
rect 1768 17478 1820 17484
rect 1780 16794 1808 17478
rect 1872 17134 1900 17682
rect 1860 17128 1912 17134
rect 1860 17070 1912 17076
rect 2136 16992 2188 16998
rect 2136 16934 2188 16940
rect 1768 16788 1820 16794
rect 1768 16730 1820 16736
rect 2148 16590 2176 16934
rect 1492 16584 1544 16590
rect 1492 16526 1544 16532
rect 2136 16584 2188 16590
rect 2136 16526 2188 16532
rect 1504 16114 1532 16526
rect 2780 16244 2832 16250
rect 2780 16186 2832 16192
rect 1492 16108 1544 16114
rect 1492 16050 1544 16056
rect 2792 15638 2820 16186
rect 2884 15706 2912 19110
rect 3068 18970 3096 19382
rect 3160 19378 3188 20726
rect 3252 20602 3280 20946
rect 3332 20936 3384 20942
rect 3332 20878 3384 20884
rect 3240 20596 3292 20602
rect 3240 20538 3292 20544
rect 3344 20398 3372 20878
rect 3332 20392 3384 20398
rect 3332 20334 3384 20340
rect 3238 20224 3294 20233
rect 3238 20159 3294 20168
rect 3148 19372 3200 19378
rect 3148 19314 3200 19320
rect 3148 19236 3200 19242
rect 3148 19178 3200 19184
rect 3056 18964 3108 18970
rect 3056 18906 3108 18912
rect 3056 18828 3108 18834
rect 3056 18770 3108 18776
rect 3068 18426 3096 18770
rect 3056 18420 3108 18426
rect 3056 18362 3108 18368
rect 3160 18154 3188 19178
rect 3148 18148 3200 18154
rect 3148 18090 3200 18096
rect 3160 17882 3188 18090
rect 3148 17876 3200 17882
rect 3148 17818 3200 17824
rect 3148 15904 3200 15910
rect 3148 15846 3200 15852
rect 2872 15700 2924 15706
rect 2872 15642 2924 15648
rect 2780 15632 2832 15638
rect 2780 15574 2832 15580
rect 1768 15496 1820 15502
rect 1490 15464 1546 15473
rect 1768 15438 1820 15444
rect 1490 15399 1546 15408
rect 1400 14952 1452 14958
rect 1400 14894 1452 14900
rect 1504 10810 1532 15399
rect 1676 15360 1728 15366
rect 1676 15302 1728 15308
rect 1688 14498 1716 15302
rect 1780 14958 1808 15438
rect 1858 15192 1914 15201
rect 1858 15127 1914 15136
rect 1768 14952 1820 14958
rect 1768 14894 1820 14900
rect 1780 14618 1808 14894
rect 1768 14612 1820 14618
rect 1768 14554 1820 14560
rect 1688 14470 1808 14498
rect 1674 14376 1730 14385
rect 1674 14311 1730 14320
rect 1688 14006 1716 14311
rect 1676 14000 1728 14006
rect 1676 13942 1728 13948
rect 1676 13796 1728 13802
rect 1676 13738 1728 13744
rect 1688 13394 1716 13738
rect 1676 13388 1728 13394
rect 1676 13330 1728 13336
rect 1688 12986 1716 13330
rect 1676 12980 1728 12986
rect 1676 12922 1728 12928
rect 1582 12336 1638 12345
rect 1582 12271 1638 12280
rect 1596 11354 1624 12271
rect 1584 11348 1636 11354
rect 1584 11290 1636 11296
rect 1780 10810 1808 14470
rect 1492 10804 1544 10810
rect 1492 10746 1544 10752
rect 1768 10804 1820 10810
rect 1768 10746 1820 10752
rect 1504 10606 1532 10746
rect 1492 10600 1544 10606
rect 1492 10542 1544 10548
rect 1492 9444 1544 9450
rect 1492 9386 1544 9392
rect 1504 9081 1532 9386
rect 1490 9072 1546 9081
rect 1490 9007 1546 9016
rect 1872 8498 1900 15127
rect 2884 15042 2912 15642
rect 2792 15014 2912 15042
rect 2792 14958 2820 15014
rect 2780 14952 2832 14958
rect 2780 14894 2832 14900
rect 2504 14884 2556 14890
rect 2504 14826 2556 14832
rect 2688 14884 2740 14890
rect 2688 14826 2740 14832
rect 2044 14476 2096 14482
rect 2044 14418 2096 14424
rect 2056 12986 2084 14418
rect 2516 14346 2544 14826
rect 2504 14340 2556 14346
rect 2504 14282 2556 14288
rect 2136 14272 2188 14278
rect 2136 14214 2188 14220
rect 2148 13462 2176 14214
rect 2516 13802 2544 14282
rect 2504 13796 2556 13802
rect 2504 13738 2556 13744
rect 2136 13456 2188 13462
rect 2136 13398 2188 13404
rect 2044 12980 2096 12986
rect 2044 12922 2096 12928
rect 2056 12306 2084 12922
rect 2148 12442 2176 13398
rect 2136 12436 2188 12442
rect 2136 12378 2188 12384
rect 2044 12300 2096 12306
rect 2044 12242 2096 12248
rect 1952 12096 2004 12102
rect 1952 12038 2004 12044
rect 1964 11762 1992 12038
rect 1952 11756 2004 11762
rect 1952 11698 2004 11704
rect 2136 11756 2188 11762
rect 2136 11698 2188 11704
rect 1952 11620 2004 11626
rect 1952 11562 2004 11568
rect 1964 11150 1992 11562
rect 2148 11354 2176 11698
rect 2136 11348 2188 11354
rect 2136 11290 2188 11296
rect 1952 11144 2004 11150
rect 1952 11086 2004 11092
rect 1964 10606 1992 11086
rect 2596 11008 2648 11014
rect 2596 10950 2648 10956
rect 1952 10600 2004 10606
rect 1952 10542 2004 10548
rect 1964 9518 1992 10542
rect 2504 10464 2556 10470
rect 2504 10406 2556 10412
rect 2136 9920 2188 9926
rect 2136 9862 2188 9868
rect 1952 9512 2004 9518
rect 1952 9454 2004 9460
rect 1860 8492 1912 8498
rect 1860 8434 1912 8440
rect 1768 8424 1820 8430
rect 1768 8366 1820 8372
rect 1780 8022 1808 8366
rect 1768 8016 1820 8022
rect 1768 7958 1820 7964
rect 1768 3528 1820 3534
rect 1768 3470 1820 3476
rect 1780 2990 1808 3470
rect 1950 3088 2006 3097
rect 1950 3023 1952 3032
rect 2004 3023 2006 3032
rect 1952 2994 2004 3000
rect 1768 2984 1820 2990
rect 1768 2926 1820 2932
rect 2148 2922 2176 9862
rect 2516 4978 2544 10406
rect 2608 10266 2636 10950
rect 2596 10260 2648 10266
rect 2596 10202 2648 10208
rect 2700 10130 2728 14826
rect 3160 14550 3188 15846
rect 3148 14544 3200 14550
rect 3148 14486 3200 14492
rect 3056 13864 3108 13870
rect 2870 13832 2926 13841
rect 3056 13806 3108 13812
rect 2870 13767 2926 13776
rect 2780 11280 2832 11286
rect 2780 11222 2832 11228
rect 2688 10124 2740 10130
rect 2688 10066 2740 10072
rect 2792 9654 2820 11222
rect 2780 9648 2832 9654
rect 2780 9590 2832 9596
rect 2884 9518 2912 13767
rect 3068 13530 3096 13806
rect 3056 13524 3108 13530
rect 3056 13466 3108 13472
rect 3252 12374 3280 20159
rect 3344 19378 3372 20334
rect 3436 19922 3464 23600
rect 3516 21140 3568 21146
rect 3516 21082 3568 21088
rect 3528 20398 3556 21082
rect 3516 20392 3568 20398
rect 3516 20334 3568 20340
rect 3976 20392 4028 20398
rect 3976 20334 4028 20340
rect 3608 20256 3660 20262
rect 3608 20198 3660 20204
rect 3424 19916 3476 19922
rect 3424 19858 3476 19864
rect 3332 19372 3384 19378
rect 3332 19314 3384 19320
rect 3344 18222 3372 19314
rect 3516 19168 3568 19174
rect 3516 19110 3568 19116
rect 3528 18970 3556 19110
rect 3516 18964 3568 18970
rect 3516 18906 3568 18912
rect 3516 18828 3568 18834
rect 3516 18770 3568 18776
rect 3424 18760 3476 18766
rect 3424 18702 3476 18708
rect 3332 18216 3384 18222
rect 3332 18158 3384 18164
rect 3344 17678 3372 18158
rect 3332 17672 3384 17678
rect 3332 17614 3384 17620
rect 3344 16998 3372 17614
rect 3332 16992 3384 16998
rect 3332 16934 3384 16940
rect 3436 16726 3464 18702
rect 3528 17134 3556 18770
rect 3620 17882 3648 20198
rect 3790 19952 3846 19961
rect 3790 19887 3846 19896
rect 3700 18964 3752 18970
rect 3700 18906 3752 18912
rect 3608 17876 3660 17882
rect 3608 17818 3660 17824
rect 3516 17128 3568 17134
rect 3516 17070 3568 17076
rect 3528 16794 3556 17070
rect 3516 16788 3568 16794
rect 3516 16730 3568 16736
rect 3424 16720 3476 16726
rect 3330 16688 3386 16697
rect 3424 16662 3476 16668
rect 3330 16623 3386 16632
rect 3344 12782 3372 16623
rect 3436 15162 3464 16662
rect 3712 16250 3740 18906
rect 3804 17746 3832 19887
rect 3884 19848 3936 19854
rect 3884 19790 3936 19796
rect 3896 19446 3924 19790
rect 3884 19440 3936 19446
rect 3884 19382 3936 19388
rect 3884 19236 3936 19242
rect 3884 19178 3936 19184
rect 3896 18086 3924 19178
rect 3884 18080 3936 18086
rect 3884 18022 3936 18028
rect 3896 17814 3924 18022
rect 3884 17808 3936 17814
rect 3884 17750 3936 17756
rect 3792 17740 3844 17746
rect 3792 17682 3844 17688
rect 3700 16244 3752 16250
rect 3700 16186 3752 16192
rect 3516 15904 3568 15910
rect 3516 15846 3568 15852
rect 3700 15904 3752 15910
rect 3700 15846 3752 15852
rect 3528 15162 3556 15846
rect 3424 15156 3476 15162
rect 3424 15098 3476 15104
rect 3516 15156 3568 15162
rect 3516 15098 3568 15104
rect 3608 14272 3660 14278
rect 3608 14214 3660 14220
rect 3620 13870 3648 14214
rect 3608 13864 3660 13870
rect 3608 13806 3660 13812
rect 3424 13388 3476 13394
rect 3424 13330 3476 13336
rect 3332 12776 3384 12782
rect 3332 12718 3384 12724
rect 3148 12368 3200 12374
rect 3148 12310 3200 12316
rect 3240 12368 3292 12374
rect 3240 12310 3292 12316
rect 3160 11286 3188 12310
rect 3332 12300 3384 12306
rect 3332 12242 3384 12248
rect 3344 11626 3372 12242
rect 3436 11898 3464 13330
rect 3608 12640 3660 12646
rect 3608 12582 3660 12588
rect 3424 11892 3476 11898
rect 3424 11834 3476 11840
rect 3516 11824 3568 11830
rect 3516 11766 3568 11772
rect 3332 11620 3384 11626
rect 3332 11562 3384 11568
rect 3148 11280 3200 11286
rect 3148 11222 3200 11228
rect 3344 11082 3372 11562
rect 3332 11076 3384 11082
rect 3332 11018 3384 11024
rect 3056 9920 3108 9926
rect 3056 9862 3108 9868
rect 2872 9512 2924 9518
rect 2872 9454 2924 9460
rect 2516 4950 2636 4978
rect 2504 3392 2556 3398
rect 2504 3334 2556 3340
rect 2516 2990 2544 3334
rect 2608 3126 2636 4950
rect 2596 3120 2648 3126
rect 2596 3062 2648 3068
rect 2504 2984 2556 2990
rect 2504 2926 2556 2932
rect 2136 2916 2188 2922
rect 2136 2858 2188 2864
rect 1676 2848 1728 2854
rect 1676 2790 1728 2796
rect 1688 800 1716 2790
rect 3068 2514 3096 9862
rect 3528 9178 3556 11766
rect 3620 11558 3648 12582
rect 3712 12102 3740 15846
rect 3988 15570 4016 20334
rect 4080 19786 4108 23600
rect 4724 22930 4752 23600
rect 4724 22902 5028 22930
rect 4654 21788 4950 21808
rect 4710 21786 4734 21788
rect 4790 21786 4814 21788
rect 4870 21786 4894 21788
rect 4732 21734 4734 21786
rect 4796 21734 4808 21786
rect 4870 21734 4872 21786
rect 4710 21732 4734 21734
rect 4790 21732 4814 21734
rect 4870 21732 4894 21734
rect 4654 21712 4950 21732
rect 4342 21448 4398 21457
rect 4342 21383 4398 21392
rect 4356 21350 4384 21383
rect 4344 21344 4396 21350
rect 4344 21286 4396 21292
rect 4528 21344 4580 21350
rect 4528 21286 4580 21292
rect 4344 21004 4396 21010
rect 4344 20946 4396 20952
rect 4356 20602 4384 20946
rect 4436 20800 4488 20806
rect 4436 20742 4488 20748
rect 4344 20596 4396 20602
rect 4344 20538 4396 20544
rect 4160 20324 4212 20330
rect 4160 20266 4212 20272
rect 4068 19780 4120 19786
rect 4068 19722 4120 19728
rect 4172 19514 4200 20266
rect 4344 20256 4396 20262
rect 4344 20198 4396 20204
rect 4252 19916 4304 19922
rect 4252 19858 4304 19864
rect 4160 19508 4212 19514
rect 4160 19450 4212 19456
rect 4068 19168 4120 19174
rect 4068 19110 4120 19116
rect 4080 18222 4108 19110
rect 4068 18216 4120 18222
rect 4068 18158 4120 18164
rect 4080 17270 4108 18158
rect 4264 17882 4292 19858
rect 4252 17876 4304 17882
rect 4252 17818 4304 17824
rect 4068 17264 4120 17270
rect 4068 17206 4120 17212
rect 4252 17264 4304 17270
rect 4252 17206 4304 17212
rect 4160 17128 4212 17134
rect 4160 17070 4212 17076
rect 4172 16250 4200 17070
rect 4160 16244 4212 16250
rect 4160 16186 4212 16192
rect 3976 15564 4028 15570
rect 3976 15506 4028 15512
rect 3790 15056 3846 15065
rect 3790 14991 3846 15000
rect 3884 15020 3936 15026
rect 3804 12986 3832 14991
rect 3884 14962 3936 14968
rect 3792 12980 3844 12986
rect 3792 12922 3844 12928
rect 3896 12850 3924 14962
rect 3976 14952 4028 14958
rect 3976 14894 4028 14900
rect 3988 13870 4016 14894
rect 4068 14816 4120 14822
rect 4068 14758 4120 14764
rect 3976 13864 4028 13870
rect 3976 13806 4028 13812
rect 4080 13530 4108 14758
rect 4172 14482 4200 16186
rect 4160 14476 4212 14482
rect 4160 14418 4212 14424
rect 4264 14278 4292 17206
rect 4356 16726 4384 20198
rect 4344 16720 4396 16726
rect 4344 16662 4396 16668
rect 4448 16658 4476 20742
rect 4540 20058 4568 21286
rect 4654 20700 4950 20720
rect 4710 20698 4734 20700
rect 4790 20698 4814 20700
rect 4870 20698 4894 20700
rect 4732 20646 4734 20698
rect 4796 20646 4808 20698
rect 4870 20646 4872 20698
rect 4710 20644 4734 20646
rect 4790 20644 4814 20646
rect 4870 20644 4894 20646
rect 4654 20624 4950 20644
rect 4528 20052 4580 20058
rect 4528 19994 4580 20000
rect 4620 19984 4672 19990
rect 4540 19932 4620 19938
rect 4540 19926 4672 19932
rect 4540 19910 4660 19926
rect 4804 19916 4856 19922
rect 4540 19378 4568 19910
rect 4804 19858 4856 19864
rect 4816 19825 4844 19858
rect 4802 19816 4858 19825
rect 4802 19751 4858 19760
rect 4654 19612 4950 19632
rect 4710 19610 4734 19612
rect 4790 19610 4814 19612
rect 4870 19610 4894 19612
rect 4732 19558 4734 19610
rect 4796 19558 4808 19610
rect 4870 19558 4872 19610
rect 4710 19556 4734 19558
rect 4790 19556 4814 19558
rect 4870 19556 4894 19558
rect 4654 19536 4950 19556
rect 5000 19514 5028 22902
rect 5264 21548 5316 21554
rect 5264 21490 5316 21496
rect 5172 21072 5224 21078
rect 5172 21014 5224 21020
rect 5080 20936 5132 20942
rect 5080 20878 5132 20884
rect 4988 19508 5040 19514
rect 4988 19450 5040 19456
rect 4620 19440 4672 19446
rect 4620 19382 4672 19388
rect 4528 19372 4580 19378
rect 4528 19314 4580 19320
rect 4632 18766 4660 19382
rect 4620 18760 4672 18766
rect 4620 18702 4672 18708
rect 4654 18524 4950 18544
rect 4710 18522 4734 18524
rect 4790 18522 4814 18524
rect 4870 18522 4894 18524
rect 4732 18470 4734 18522
rect 4796 18470 4808 18522
rect 4870 18470 4872 18522
rect 4710 18468 4734 18470
rect 4790 18468 4814 18470
rect 4870 18468 4894 18470
rect 4654 18448 4950 18468
rect 4988 18352 5040 18358
rect 4988 18294 5040 18300
rect 4528 18216 4580 18222
rect 4528 18158 4580 18164
rect 4540 16998 4568 18158
rect 4896 17740 4948 17746
rect 4896 17682 4948 17688
rect 4908 17649 4936 17682
rect 4894 17640 4950 17649
rect 4894 17575 4950 17584
rect 4654 17436 4950 17456
rect 4710 17434 4734 17436
rect 4790 17434 4814 17436
rect 4870 17434 4894 17436
rect 4732 17382 4734 17434
rect 4796 17382 4808 17434
rect 4870 17382 4872 17434
rect 4710 17380 4734 17382
rect 4790 17380 4814 17382
rect 4870 17380 4894 17382
rect 4654 17360 4950 17380
rect 4802 17232 4858 17241
rect 4802 17167 4858 17176
rect 4528 16992 4580 16998
rect 4528 16934 4580 16940
rect 4436 16652 4488 16658
rect 4436 16594 4488 16600
rect 4816 16590 4844 17167
rect 5000 17134 5028 18294
rect 4988 17128 5040 17134
rect 4988 17070 5040 17076
rect 4804 16584 4856 16590
rect 4804 16526 4856 16532
rect 4528 16448 4580 16454
rect 4528 16390 4580 16396
rect 4436 16176 4488 16182
rect 4436 16118 4488 16124
rect 4344 16108 4396 16114
rect 4344 16050 4396 16056
rect 4356 15638 4384 16050
rect 4344 15632 4396 15638
rect 4344 15574 4396 15580
rect 4356 15434 4384 15574
rect 4344 15428 4396 15434
rect 4344 15370 4396 15376
rect 4252 14272 4304 14278
rect 4252 14214 4304 14220
rect 4160 13796 4212 13802
rect 4160 13738 4212 13744
rect 4068 13524 4120 13530
rect 4068 13466 4120 13472
rect 4172 13394 4200 13738
rect 4264 13394 4292 14214
rect 4160 13388 4212 13394
rect 4160 13330 4212 13336
rect 4252 13388 4304 13394
rect 4252 13330 4304 13336
rect 3974 13288 4030 13297
rect 3974 13223 4030 13232
rect 3884 12844 3936 12850
rect 3884 12786 3936 12792
rect 3896 12481 3924 12786
rect 3882 12472 3938 12481
rect 3882 12407 3938 12416
rect 3896 12238 3924 12407
rect 3884 12232 3936 12238
rect 3884 12174 3936 12180
rect 3700 12096 3752 12102
rect 3700 12038 3752 12044
rect 3884 12096 3936 12102
rect 3884 12038 3936 12044
rect 3608 11552 3660 11558
rect 3608 11494 3660 11500
rect 3792 11552 3844 11558
rect 3792 11494 3844 11500
rect 3804 11354 3832 11494
rect 3792 11348 3844 11354
rect 3792 11290 3844 11296
rect 3700 10192 3752 10198
rect 3700 10134 3752 10140
rect 3608 10056 3660 10062
rect 3606 10024 3608 10033
rect 3660 10024 3662 10033
rect 3606 9959 3662 9968
rect 3712 9382 3740 10134
rect 3700 9376 3752 9382
rect 3700 9318 3752 9324
rect 3516 9172 3568 9178
rect 3516 9114 3568 9120
rect 3712 6798 3740 9318
rect 3700 6792 3752 6798
rect 3700 6734 3752 6740
rect 3896 3670 3924 12038
rect 3988 9042 4016 13223
rect 4264 12850 4292 13330
rect 4252 12844 4304 12850
rect 4252 12786 4304 12792
rect 4252 12708 4304 12714
rect 4252 12650 4304 12656
rect 4068 12640 4120 12646
rect 4068 12582 4120 12588
rect 4080 11762 4108 12582
rect 4160 12232 4212 12238
rect 4160 12174 4212 12180
rect 4068 11756 4120 11762
rect 4068 11698 4120 11704
rect 4080 10538 4108 11698
rect 4172 11694 4200 12174
rect 4160 11688 4212 11694
rect 4160 11630 4212 11636
rect 4172 11218 4200 11630
rect 4264 11286 4292 12650
rect 4356 11558 4384 15370
rect 4448 15026 4476 16118
rect 4540 15502 4568 16390
rect 4654 16348 4950 16368
rect 4710 16346 4734 16348
rect 4790 16346 4814 16348
rect 4870 16346 4894 16348
rect 4732 16294 4734 16346
rect 4796 16294 4808 16346
rect 4870 16294 4872 16346
rect 4710 16292 4734 16294
rect 4790 16292 4814 16294
rect 4870 16292 4894 16294
rect 4654 16272 4950 16292
rect 4804 16040 4856 16046
rect 4804 15982 4856 15988
rect 4816 15638 4844 15982
rect 5092 15892 5120 20878
rect 5184 19310 5212 21014
rect 5276 20874 5304 21490
rect 5264 20868 5316 20874
rect 5264 20810 5316 20816
rect 5264 20596 5316 20602
rect 5264 20538 5316 20544
rect 5172 19304 5224 19310
rect 5172 19246 5224 19252
rect 5276 18902 5304 20538
rect 5264 18896 5316 18902
rect 5264 18838 5316 18844
rect 5172 18148 5224 18154
rect 5172 18090 5224 18096
rect 5184 17134 5212 18090
rect 5264 17876 5316 17882
rect 5264 17818 5316 17824
rect 5276 17542 5304 17818
rect 5264 17536 5316 17542
rect 5264 17478 5316 17484
rect 5172 17128 5224 17134
rect 5172 17070 5224 17076
rect 5262 16960 5318 16969
rect 5262 16895 5318 16904
rect 5000 15864 5120 15892
rect 4804 15632 4856 15638
rect 4804 15574 4856 15580
rect 4528 15496 4580 15502
rect 4528 15438 4580 15444
rect 4654 15260 4950 15280
rect 4710 15258 4734 15260
rect 4790 15258 4814 15260
rect 4870 15258 4894 15260
rect 4732 15206 4734 15258
rect 4796 15206 4808 15258
rect 4870 15206 4872 15258
rect 4710 15204 4734 15206
rect 4790 15204 4814 15206
rect 4870 15204 4894 15206
rect 4654 15184 4950 15204
rect 5000 15042 5028 15864
rect 5080 15496 5132 15502
rect 5080 15438 5132 15444
rect 5092 15162 5120 15438
rect 5080 15156 5132 15162
rect 5080 15098 5132 15104
rect 4436 15020 4488 15026
rect 4436 14962 4488 14968
rect 4540 15014 5028 15042
rect 4436 12708 4488 12714
rect 4436 12650 4488 12656
rect 4344 11552 4396 11558
rect 4344 11494 4396 11500
rect 4252 11280 4304 11286
rect 4252 11222 4304 11228
rect 4160 11212 4212 11218
rect 4160 11154 4212 11160
rect 4264 10810 4292 11222
rect 4252 10804 4304 10810
rect 4252 10746 4304 10752
rect 4344 10736 4396 10742
rect 4344 10678 4396 10684
rect 4068 10532 4120 10538
rect 4068 10474 4120 10480
rect 4252 10260 4304 10266
rect 4252 10202 4304 10208
rect 4160 10124 4212 10130
rect 4160 10066 4212 10072
rect 4068 9376 4120 9382
rect 4068 9318 4120 9324
rect 3976 9036 4028 9042
rect 3976 8978 4028 8984
rect 4080 8634 4108 9318
rect 4172 9178 4200 10066
rect 4264 9994 4292 10202
rect 4252 9988 4304 9994
rect 4252 9930 4304 9936
rect 4252 9580 4304 9586
rect 4252 9522 4304 9528
rect 4160 9172 4212 9178
rect 4160 9114 4212 9120
rect 4264 8906 4292 9522
rect 4252 8900 4304 8906
rect 4252 8842 4304 8848
rect 4068 8628 4120 8634
rect 4068 8570 4120 8576
rect 4356 7954 4384 10678
rect 4448 9042 4476 12650
rect 4540 12442 4568 15014
rect 5172 14884 5224 14890
rect 5172 14826 5224 14832
rect 5080 14816 5132 14822
rect 5080 14758 5132 14764
rect 4988 14612 5040 14618
rect 4988 14554 5040 14560
rect 4654 14172 4950 14192
rect 4710 14170 4734 14172
rect 4790 14170 4814 14172
rect 4870 14170 4894 14172
rect 4732 14118 4734 14170
rect 4796 14118 4808 14170
rect 4870 14118 4872 14170
rect 4710 14116 4734 14118
rect 4790 14116 4814 14118
rect 4870 14116 4894 14118
rect 4654 14096 4950 14116
rect 4654 13084 4950 13104
rect 4710 13082 4734 13084
rect 4790 13082 4814 13084
rect 4870 13082 4894 13084
rect 4732 13030 4734 13082
rect 4796 13030 4808 13082
rect 4870 13030 4872 13082
rect 4710 13028 4734 13030
rect 4790 13028 4814 13030
rect 4870 13028 4894 13030
rect 4654 13008 4950 13028
rect 4528 12436 4580 12442
rect 4528 12378 4580 12384
rect 4654 11996 4950 12016
rect 4710 11994 4734 11996
rect 4790 11994 4814 11996
rect 4870 11994 4894 11996
rect 4732 11942 4734 11994
rect 4796 11942 4808 11994
rect 4870 11942 4872 11994
rect 4710 11940 4734 11942
rect 4790 11940 4814 11942
rect 4870 11940 4894 11942
rect 4654 11920 4950 11940
rect 4528 11552 4580 11558
rect 4528 11494 4580 11500
rect 4540 10674 4568 11494
rect 4654 10908 4950 10928
rect 4710 10906 4734 10908
rect 4790 10906 4814 10908
rect 4870 10906 4894 10908
rect 4732 10854 4734 10906
rect 4796 10854 4808 10906
rect 4870 10854 4872 10906
rect 4710 10852 4734 10854
rect 4790 10852 4814 10854
rect 4870 10852 4894 10854
rect 4654 10832 4950 10852
rect 4620 10736 4672 10742
rect 4620 10678 4672 10684
rect 4528 10668 4580 10674
rect 4528 10610 4580 10616
rect 4528 10464 4580 10470
rect 4528 10406 4580 10412
rect 4540 9722 4568 10406
rect 4632 10266 4660 10678
rect 4620 10260 4672 10266
rect 4620 10202 4672 10208
rect 4654 9820 4950 9840
rect 4710 9818 4734 9820
rect 4790 9818 4814 9820
rect 4870 9818 4894 9820
rect 4732 9766 4734 9818
rect 4796 9766 4808 9818
rect 4870 9766 4872 9818
rect 4710 9764 4734 9766
rect 4790 9764 4814 9766
rect 4870 9764 4894 9766
rect 4654 9744 4950 9764
rect 4528 9716 4580 9722
rect 4528 9658 4580 9664
rect 4894 9616 4950 9625
rect 4894 9551 4950 9560
rect 4908 9518 4936 9551
rect 4896 9512 4948 9518
rect 4896 9454 4948 9460
rect 4436 9036 4488 9042
rect 4436 8978 4488 8984
rect 4654 8732 4950 8752
rect 4710 8730 4734 8732
rect 4790 8730 4814 8732
rect 4870 8730 4894 8732
rect 4732 8678 4734 8730
rect 4796 8678 4808 8730
rect 4870 8678 4872 8730
rect 4710 8676 4734 8678
rect 4790 8676 4814 8678
rect 4870 8676 4894 8678
rect 4654 8656 4950 8676
rect 4712 8560 4764 8566
rect 4712 8502 4764 8508
rect 4724 8401 4752 8502
rect 4710 8392 4766 8401
rect 4710 8327 4766 8336
rect 5000 8090 5028 14554
rect 5092 14482 5120 14758
rect 5080 14476 5132 14482
rect 5080 14418 5132 14424
rect 5092 14074 5120 14418
rect 5184 14278 5212 14826
rect 5276 14498 5304 16895
rect 5368 15978 5396 23600
rect 5632 21616 5684 21622
rect 5632 21558 5684 21564
rect 5540 21344 5592 21350
rect 5540 21286 5592 21292
rect 5552 21146 5580 21286
rect 5540 21140 5592 21146
rect 5540 21082 5592 21088
rect 5448 20868 5500 20874
rect 5448 20810 5500 20816
rect 5460 20346 5488 20810
rect 5644 20448 5672 21558
rect 5816 20800 5868 20806
rect 5816 20742 5868 20748
rect 5724 20460 5776 20466
rect 5644 20420 5724 20448
rect 5724 20402 5776 20408
rect 5460 20318 5580 20346
rect 5448 20256 5500 20262
rect 5448 20198 5500 20204
rect 5460 18970 5488 20198
rect 5448 18964 5500 18970
rect 5448 18906 5500 18912
rect 5552 18850 5580 20318
rect 5632 20256 5684 20262
rect 5630 20224 5632 20233
rect 5684 20224 5686 20233
rect 5630 20159 5686 20168
rect 5736 19825 5764 20402
rect 5828 19990 5856 20742
rect 6012 20534 6040 23600
rect 6182 21992 6238 22001
rect 6182 21927 6238 21936
rect 6090 21584 6146 21593
rect 6090 21519 6146 21528
rect 6104 21486 6132 21519
rect 6092 21480 6144 21486
rect 6092 21422 6144 21428
rect 6000 20528 6052 20534
rect 6000 20470 6052 20476
rect 5816 19984 5868 19990
rect 5816 19926 5868 19932
rect 5722 19816 5778 19825
rect 5722 19751 5778 19760
rect 5828 19174 5856 19926
rect 5816 19168 5868 19174
rect 5816 19110 5868 19116
rect 5632 18964 5684 18970
rect 5632 18906 5684 18912
rect 5460 18822 5580 18850
rect 5356 15972 5408 15978
rect 5356 15914 5408 15920
rect 5460 15094 5488 18822
rect 5644 18714 5672 18906
rect 6092 18828 6144 18834
rect 6092 18770 6144 18776
rect 5552 18686 5672 18714
rect 5816 18760 5868 18766
rect 5816 18702 5868 18708
rect 5552 15910 5580 18686
rect 5828 18290 5856 18702
rect 5816 18284 5868 18290
rect 5816 18226 5868 18232
rect 5724 18148 5776 18154
rect 5724 18090 5776 18096
rect 5632 18080 5684 18086
rect 5632 18022 5684 18028
rect 5644 16726 5672 18022
rect 5736 17542 5764 18090
rect 5724 17536 5776 17542
rect 5724 17478 5776 17484
rect 5908 17196 5960 17202
rect 5908 17138 5960 17144
rect 5920 16794 5948 17138
rect 6104 16794 6132 18770
rect 5908 16788 5960 16794
rect 5908 16730 5960 16736
rect 6092 16788 6144 16794
rect 6092 16730 6144 16736
rect 5632 16720 5684 16726
rect 5632 16662 5684 16668
rect 6104 16046 6132 16730
rect 6092 16040 6144 16046
rect 6092 15982 6144 15988
rect 5540 15904 5592 15910
rect 5540 15846 5592 15852
rect 6196 15722 6224 21927
rect 6656 21894 6684 23600
rect 6644 21888 6696 21894
rect 6644 21830 6696 21836
rect 6644 21548 6696 21554
rect 6644 21490 6696 21496
rect 6736 21548 6788 21554
rect 6736 21490 6788 21496
rect 6276 21480 6328 21486
rect 6276 21422 6328 21428
rect 6288 19310 6316 21422
rect 6552 21004 6604 21010
rect 6552 20946 6604 20952
rect 6460 20936 6512 20942
rect 6460 20878 6512 20884
rect 6472 20398 6500 20878
rect 6460 20392 6512 20398
rect 6460 20334 6512 20340
rect 6472 20058 6500 20334
rect 6460 20052 6512 20058
rect 6460 19994 6512 20000
rect 6368 19916 6420 19922
rect 6368 19858 6420 19864
rect 6276 19304 6328 19310
rect 6276 19246 6328 19252
rect 6380 18630 6408 19858
rect 6472 18834 6500 19994
rect 6460 18828 6512 18834
rect 6460 18770 6512 18776
rect 6368 18624 6420 18630
rect 6564 18601 6592 20946
rect 6656 19553 6684 21490
rect 6748 21078 6776 21490
rect 6920 21344 6972 21350
rect 6920 21286 6972 21292
rect 6736 21072 6788 21078
rect 6736 21014 6788 21020
rect 6642 19544 6698 19553
rect 6642 19479 6698 19488
rect 6734 19272 6790 19281
rect 6734 19207 6790 19216
rect 6368 18566 6420 18572
rect 6550 18592 6606 18601
rect 6550 18527 6606 18536
rect 6564 18358 6592 18527
rect 6552 18352 6604 18358
rect 6552 18294 6604 18300
rect 6458 17776 6514 17785
rect 6458 17711 6514 17720
rect 6276 16992 6328 16998
rect 6276 16934 6328 16940
rect 6288 16726 6316 16934
rect 6276 16720 6328 16726
rect 6276 16662 6328 16668
rect 6196 15694 6316 15722
rect 6184 15632 6236 15638
rect 6184 15574 6236 15580
rect 5540 15564 5592 15570
rect 5540 15506 5592 15512
rect 5552 15162 5580 15506
rect 5540 15156 5592 15162
rect 5540 15098 5592 15104
rect 5448 15088 5500 15094
rect 5448 15030 5500 15036
rect 5724 15088 5776 15094
rect 5724 15030 5776 15036
rect 5736 14550 5764 15030
rect 6000 14952 6052 14958
rect 6000 14894 6052 14900
rect 5724 14544 5776 14550
rect 5276 14470 5580 14498
rect 5724 14486 5776 14492
rect 6012 14482 6040 14894
rect 6196 14822 6224 15574
rect 6184 14816 6236 14822
rect 6184 14758 6236 14764
rect 6196 14618 6224 14758
rect 6184 14612 6236 14618
rect 6184 14554 6236 14560
rect 5356 14408 5408 14414
rect 5356 14350 5408 14356
rect 5264 14340 5316 14346
rect 5264 14282 5316 14288
rect 5172 14272 5224 14278
rect 5172 14214 5224 14220
rect 5080 14068 5132 14074
rect 5080 14010 5132 14016
rect 5172 14000 5224 14006
rect 5172 13942 5224 13948
rect 5080 13388 5132 13394
rect 5080 13330 5132 13336
rect 5092 10810 5120 13330
rect 5080 10804 5132 10810
rect 5080 10746 5132 10752
rect 5184 10606 5212 13942
rect 5276 13190 5304 14282
rect 5368 13870 5396 14350
rect 5448 14272 5500 14278
rect 5448 14214 5500 14220
rect 5356 13864 5408 13870
rect 5356 13806 5408 13812
rect 5460 13462 5488 14214
rect 5448 13456 5500 13462
rect 5448 13398 5500 13404
rect 5552 13274 5580 14470
rect 6000 14476 6052 14482
rect 6000 14418 6052 14424
rect 5724 13728 5776 13734
rect 5724 13670 5776 13676
rect 5816 13728 5868 13734
rect 5816 13670 5868 13676
rect 5368 13246 5580 13274
rect 5264 13184 5316 13190
rect 5264 13126 5316 13132
rect 5172 10600 5224 10606
rect 5172 10542 5224 10548
rect 5264 10056 5316 10062
rect 5170 10024 5226 10033
rect 5264 9998 5316 10004
rect 5170 9959 5226 9968
rect 5080 9444 5132 9450
rect 5080 9386 5132 9392
rect 5092 8090 5120 9386
rect 4988 8084 5040 8090
rect 4988 8026 5040 8032
rect 5080 8084 5132 8090
rect 5080 8026 5132 8032
rect 4344 7948 4396 7954
rect 4344 7890 4396 7896
rect 4654 7644 4950 7664
rect 4710 7642 4734 7644
rect 4790 7642 4814 7644
rect 4870 7642 4894 7644
rect 4732 7590 4734 7642
rect 4796 7590 4808 7642
rect 4870 7590 4872 7642
rect 4710 7588 4734 7590
rect 4790 7588 4814 7590
rect 4870 7588 4894 7590
rect 4654 7568 4950 7588
rect 4654 6556 4950 6576
rect 4710 6554 4734 6556
rect 4790 6554 4814 6556
rect 4870 6554 4894 6556
rect 4732 6502 4734 6554
rect 4796 6502 4808 6554
rect 4870 6502 4872 6554
rect 4710 6500 4734 6502
rect 4790 6500 4814 6502
rect 4870 6500 4894 6502
rect 4654 6480 4950 6500
rect 4654 5468 4950 5488
rect 4710 5466 4734 5468
rect 4790 5466 4814 5468
rect 4870 5466 4894 5468
rect 4732 5414 4734 5466
rect 4796 5414 4808 5466
rect 4870 5414 4872 5466
rect 4710 5412 4734 5414
rect 4790 5412 4814 5414
rect 4870 5412 4894 5414
rect 4654 5392 4950 5412
rect 4654 4380 4950 4400
rect 4710 4378 4734 4380
rect 4790 4378 4814 4380
rect 4870 4378 4894 4380
rect 4732 4326 4734 4378
rect 4796 4326 4808 4378
rect 4870 4326 4872 4378
rect 4710 4324 4734 4326
rect 4790 4324 4814 4326
rect 4870 4324 4894 4326
rect 4654 4304 4950 4324
rect 5184 3942 5212 9959
rect 5276 9586 5304 9998
rect 5264 9580 5316 9586
rect 5264 9522 5316 9528
rect 5276 8378 5304 9522
rect 5368 9518 5396 13246
rect 5448 13184 5500 13190
rect 5448 13126 5500 13132
rect 5460 12714 5488 13126
rect 5448 12708 5500 12714
rect 5448 12650 5500 12656
rect 5736 12646 5764 13670
rect 5828 12782 5856 13670
rect 6012 13530 6040 14418
rect 6184 14000 6236 14006
rect 6184 13942 6236 13948
rect 6000 13524 6052 13530
rect 6000 13466 6052 13472
rect 5998 13424 6054 13433
rect 5998 13359 6054 13368
rect 5816 12776 5868 12782
rect 5816 12718 5868 12724
rect 5908 12776 5960 12782
rect 5908 12718 5960 12724
rect 5724 12640 5776 12646
rect 5724 12582 5776 12588
rect 5828 12442 5856 12718
rect 5816 12436 5868 12442
rect 5816 12378 5868 12384
rect 5816 12300 5868 12306
rect 5816 12242 5868 12248
rect 5828 11898 5856 12242
rect 5816 11892 5868 11898
rect 5816 11834 5868 11840
rect 5448 11620 5500 11626
rect 5448 11562 5500 11568
rect 5460 11354 5488 11562
rect 5828 11354 5856 11834
rect 5920 11694 5948 12718
rect 5908 11688 5960 11694
rect 5908 11630 5960 11636
rect 5448 11348 5500 11354
rect 5448 11290 5500 11296
rect 5816 11348 5868 11354
rect 5816 11290 5868 11296
rect 5540 11144 5592 11150
rect 5540 11086 5592 11092
rect 5356 9512 5408 9518
rect 5356 9454 5408 9460
rect 5356 9036 5408 9042
rect 5356 8978 5408 8984
rect 5368 8616 5396 8978
rect 5448 8832 5500 8838
rect 5446 8800 5448 8809
rect 5500 8800 5502 8809
rect 5446 8735 5502 8744
rect 5368 8588 5488 8616
rect 5354 8528 5410 8537
rect 5354 8463 5356 8472
rect 5408 8463 5410 8472
rect 5356 8434 5408 8440
rect 5276 8350 5396 8378
rect 5264 8288 5316 8294
rect 5264 8230 5316 8236
rect 5276 4729 5304 8230
rect 5368 6662 5396 8350
rect 5460 7546 5488 8588
rect 5448 7540 5500 7546
rect 5448 7482 5500 7488
rect 5552 7342 5580 11086
rect 5724 11008 5776 11014
rect 5724 10950 5776 10956
rect 5736 10606 5764 10950
rect 5920 10810 5948 11630
rect 5908 10804 5960 10810
rect 5908 10746 5960 10752
rect 5724 10600 5776 10606
rect 5724 10542 5776 10548
rect 5816 10532 5868 10538
rect 5816 10474 5868 10480
rect 5828 10062 5856 10474
rect 5816 10056 5868 10062
rect 5816 9998 5868 10004
rect 5632 9920 5684 9926
rect 5632 9862 5684 9868
rect 5644 9178 5672 9862
rect 6012 9518 6040 13359
rect 6092 11212 6144 11218
rect 6092 11154 6144 11160
rect 6104 9926 6132 11154
rect 6196 10606 6224 13942
rect 6184 10600 6236 10606
rect 6184 10542 6236 10548
rect 6184 10464 6236 10470
rect 6184 10406 6236 10412
rect 6092 9920 6144 9926
rect 6092 9862 6144 9868
rect 6000 9512 6052 9518
rect 6000 9454 6052 9460
rect 5724 9376 5776 9382
rect 5724 9318 5776 9324
rect 5632 9172 5684 9178
rect 5632 9114 5684 9120
rect 5736 9081 5764 9318
rect 5722 9072 5778 9081
rect 5722 9007 5778 9016
rect 6196 8480 6224 10406
rect 6288 9654 6316 15694
rect 6472 14006 6500 17711
rect 6644 17672 6696 17678
rect 6644 17614 6696 17620
rect 6656 17241 6684 17614
rect 6642 17232 6698 17241
rect 6642 17167 6698 17176
rect 6748 15722 6776 19207
rect 6932 18222 6960 21286
rect 7196 21072 7248 21078
rect 7196 21014 7248 21020
rect 7010 20360 7066 20369
rect 7010 20295 7066 20304
rect 7104 20324 7156 20330
rect 7024 19922 7052 20295
rect 7104 20266 7156 20272
rect 7012 19916 7064 19922
rect 7012 19858 7064 19864
rect 7116 19718 7144 20266
rect 7104 19712 7156 19718
rect 7104 19654 7156 19660
rect 7104 19168 7156 19174
rect 7104 19110 7156 19116
rect 7116 18290 7144 19110
rect 7104 18284 7156 18290
rect 7104 18226 7156 18232
rect 6920 18216 6972 18222
rect 6920 18158 6972 18164
rect 7104 18080 7156 18086
rect 7104 18022 7156 18028
rect 7010 17232 7066 17241
rect 7010 17167 7066 17176
rect 7024 17134 7052 17167
rect 7012 17128 7064 17134
rect 7012 17070 7064 17076
rect 7116 16998 7144 18022
rect 7208 17202 7236 21014
rect 7196 17196 7248 17202
rect 7196 17138 7248 17144
rect 7194 17096 7250 17105
rect 7194 17031 7250 17040
rect 7104 16992 7156 16998
rect 7104 16934 7156 16940
rect 7012 16652 7064 16658
rect 7012 16594 7064 16600
rect 6920 16584 6972 16590
rect 6920 16526 6972 16532
rect 6656 15694 6776 15722
rect 6552 15632 6604 15638
rect 6552 15574 6604 15580
rect 6460 14000 6512 14006
rect 6460 13942 6512 13948
rect 6368 13932 6420 13938
rect 6368 13874 6420 13880
rect 6380 12481 6408 13874
rect 6458 12880 6514 12889
rect 6458 12815 6514 12824
rect 6366 12472 6422 12481
rect 6366 12407 6422 12416
rect 6380 11150 6408 12407
rect 6368 11144 6420 11150
rect 6368 11086 6420 11092
rect 6366 10568 6422 10577
rect 6366 10503 6422 10512
rect 6380 10470 6408 10503
rect 6368 10464 6420 10470
rect 6368 10406 6420 10412
rect 6368 10124 6420 10130
rect 6368 10066 6420 10072
rect 6276 9648 6328 9654
rect 6276 9590 6328 9596
rect 6276 8492 6328 8498
rect 6196 8452 6276 8480
rect 6276 8434 6328 8440
rect 6184 8356 6236 8362
rect 6184 8298 6236 8304
rect 5630 7848 5686 7857
rect 5630 7783 5632 7792
rect 5684 7783 5686 7792
rect 5632 7754 5684 7760
rect 5540 7336 5592 7342
rect 5540 7278 5592 7284
rect 5356 6656 5408 6662
rect 5356 6598 5408 6604
rect 5262 4720 5318 4729
rect 5262 4655 5318 4664
rect 5172 3936 5224 3942
rect 5172 3878 5224 3884
rect 3884 3664 3936 3670
rect 3884 3606 3936 3612
rect 4654 3292 4950 3312
rect 4710 3290 4734 3292
rect 4790 3290 4814 3292
rect 4870 3290 4894 3292
rect 4732 3238 4734 3290
rect 4796 3238 4808 3290
rect 4870 3238 4872 3290
rect 4710 3236 4734 3238
rect 4790 3236 4814 3238
rect 4870 3236 4894 3238
rect 4654 3216 4950 3236
rect 5080 2984 5132 2990
rect 5080 2926 5132 2932
rect 3056 2508 3108 2514
rect 3056 2450 3108 2456
rect 4654 2204 4950 2224
rect 4710 2202 4734 2204
rect 4790 2202 4814 2204
rect 4870 2202 4894 2204
rect 4732 2150 4734 2202
rect 4796 2150 4808 2202
rect 4870 2150 4872 2202
rect 4710 2148 4734 2150
rect 4790 2148 4814 2150
rect 4870 2148 4894 2150
rect 4654 2128 4950 2148
rect 5092 800 5120 2926
rect 6196 2378 6224 8298
rect 6288 7206 6316 8434
rect 6380 7274 6408 10066
rect 6368 7268 6420 7274
rect 6368 7210 6420 7216
rect 6276 7200 6328 7206
rect 6276 7142 6328 7148
rect 6472 6866 6500 12815
rect 6564 11694 6592 15574
rect 6552 11688 6604 11694
rect 6552 11630 6604 11636
rect 6550 11520 6606 11529
rect 6550 11455 6606 11464
rect 6564 9994 6592 11455
rect 6552 9988 6604 9994
rect 6552 9930 6604 9936
rect 6656 9874 6684 15694
rect 6736 15632 6788 15638
rect 6736 15574 6788 15580
rect 6748 15434 6776 15574
rect 6932 15570 6960 16526
rect 7024 15706 7052 16594
rect 7012 15700 7064 15706
rect 7012 15642 7064 15648
rect 7102 15600 7158 15609
rect 6920 15564 6972 15570
rect 7102 15535 7158 15544
rect 6920 15506 6972 15512
rect 6736 15428 6788 15434
rect 6736 15370 6788 15376
rect 6828 15360 6880 15366
rect 6828 15302 6880 15308
rect 6840 14958 6868 15302
rect 6828 14952 6880 14958
rect 6828 14894 6880 14900
rect 6826 14240 6882 14249
rect 6826 14175 6882 14184
rect 6840 13988 6868 14175
rect 6564 9846 6684 9874
rect 6748 13960 6868 13988
rect 6564 9178 6592 9846
rect 6552 9172 6604 9178
rect 6552 9114 6604 9120
rect 6748 8090 6776 13960
rect 7012 13388 7064 13394
rect 7012 13330 7064 13336
rect 7024 12850 7052 13330
rect 7012 12844 7064 12850
rect 7012 12786 7064 12792
rect 6826 12744 6882 12753
rect 6826 12679 6882 12688
rect 6840 8430 6868 12679
rect 7024 12306 7052 12786
rect 7012 12300 7064 12306
rect 7012 12242 7064 12248
rect 6918 12200 6974 12209
rect 6918 12135 6920 12144
rect 6972 12135 6974 12144
rect 6920 12106 6972 12112
rect 6920 11688 6972 11694
rect 7024 11676 7052 12242
rect 6972 11648 7052 11676
rect 6920 11630 6972 11636
rect 6932 11218 6960 11630
rect 6920 11212 6972 11218
rect 6920 11154 6972 11160
rect 6932 10606 6960 11154
rect 6920 10600 6972 10606
rect 6920 10542 6972 10548
rect 6932 10062 6960 10542
rect 6920 10056 6972 10062
rect 6920 9998 6972 10004
rect 7010 10024 7066 10033
rect 7010 9959 7012 9968
rect 7064 9959 7066 9968
rect 7012 9930 7064 9936
rect 7024 9722 7052 9930
rect 7012 9716 7064 9722
rect 7012 9658 7064 9664
rect 6920 9104 6972 9110
rect 6920 9046 6972 9052
rect 6828 8424 6880 8430
rect 6828 8366 6880 8372
rect 6736 8084 6788 8090
rect 6736 8026 6788 8032
rect 6828 7948 6880 7954
rect 6828 7890 6880 7896
rect 6460 6860 6512 6866
rect 6460 6802 6512 6808
rect 6644 6656 6696 6662
rect 6644 6598 6696 6604
rect 6656 5778 6684 6598
rect 6840 6497 6868 7890
rect 6932 7449 6960 9046
rect 7012 8288 7064 8294
rect 7012 8230 7064 8236
rect 6918 7440 6974 7449
rect 6918 7375 6974 7384
rect 6920 7336 6972 7342
rect 6920 7278 6972 7284
rect 6826 6488 6882 6497
rect 6826 6423 6882 6432
rect 6644 5772 6696 5778
rect 6644 5714 6696 5720
rect 6932 4146 6960 7278
rect 6920 4140 6972 4146
rect 6920 4082 6972 4088
rect 7024 2854 7052 8230
rect 7116 6458 7144 15535
rect 7208 13734 7236 17031
rect 7300 16794 7328 23600
rect 7944 22098 7972 23600
rect 8588 22914 8616 23600
rect 8576 22908 8628 22914
rect 8576 22850 8628 22856
rect 9232 22166 9260 23600
rect 9496 22908 9548 22914
rect 9496 22850 9548 22856
rect 9220 22160 9272 22166
rect 9220 22102 9272 22108
rect 7932 22092 7984 22098
rect 7932 22034 7984 22040
rect 9404 22092 9456 22098
rect 9404 22034 9456 22040
rect 8760 22024 8812 22030
rect 8760 21966 8812 21972
rect 7748 21888 7800 21894
rect 7748 21830 7800 21836
rect 8208 21888 8260 21894
rect 8208 21830 8260 21836
rect 7656 21548 7708 21554
rect 7656 21490 7708 21496
rect 7380 21344 7432 21350
rect 7380 21286 7432 21292
rect 7392 21078 7420 21286
rect 7380 21072 7432 21078
rect 7380 21014 7432 21020
rect 7472 21072 7524 21078
rect 7472 21014 7524 21020
rect 7484 19990 7512 21014
rect 7472 19984 7524 19990
rect 7472 19926 7524 19932
rect 7668 19417 7696 21490
rect 7760 19990 7788 21830
rect 8220 21570 8248 21830
rect 8036 21542 8248 21570
rect 8392 21616 8444 21622
rect 8392 21558 8444 21564
rect 7840 21140 7892 21146
rect 7840 21082 7892 21088
rect 7852 20942 7880 21082
rect 8036 21010 8064 21542
rect 8404 21486 8432 21558
rect 8668 21548 8720 21554
rect 8668 21490 8720 21496
rect 8392 21480 8444 21486
rect 8392 21422 8444 21428
rect 8353 21244 8649 21264
rect 8409 21242 8433 21244
rect 8489 21242 8513 21244
rect 8569 21242 8593 21244
rect 8431 21190 8433 21242
rect 8495 21190 8507 21242
rect 8569 21190 8571 21242
rect 8409 21188 8433 21190
rect 8489 21188 8513 21190
rect 8569 21188 8593 21190
rect 8353 21168 8649 21188
rect 8024 21004 8076 21010
rect 8024 20946 8076 20952
rect 7840 20936 7892 20942
rect 7840 20878 7892 20884
rect 8036 20618 8064 20946
rect 8680 20874 8708 21490
rect 8668 20868 8720 20874
rect 8668 20810 8720 20816
rect 8576 20800 8628 20806
rect 8576 20742 8628 20748
rect 8036 20602 8156 20618
rect 8588 20602 8616 20742
rect 8036 20596 8168 20602
rect 8036 20590 8116 20596
rect 8116 20538 8168 20544
rect 8576 20596 8628 20602
rect 8576 20538 8628 20544
rect 8588 20380 8616 20538
rect 8588 20352 8708 20380
rect 8353 20156 8649 20176
rect 8409 20154 8433 20156
rect 8489 20154 8513 20156
rect 8569 20154 8593 20156
rect 8431 20102 8433 20154
rect 8495 20102 8507 20154
rect 8569 20102 8571 20154
rect 8409 20100 8433 20102
rect 8489 20100 8513 20102
rect 8569 20100 8593 20102
rect 8353 20080 8649 20100
rect 8680 20058 8708 20352
rect 8668 20052 8720 20058
rect 8668 19994 8720 20000
rect 7748 19984 7800 19990
rect 7748 19926 7800 19932
rect 7840 19916 7892 19922
rect 7840 19858 7892 19864
rect 7654 19408 7710 19417
rect 7654 19343 7710 19352
rect 7748 19372 7800 19378
rect 7748 19314 7800 19320
rect 7656 19304 7708 19310
rect 7656 19246 7708 19252
rect 7668 18902 7696 19246
rect 7656 18896 7708 18902
rect 7656 18838 7708 18844
rect 7380 18828 7432 18834
rect 7380 18770 7432 18776
rect 7472 18828 7524 18834
rect 7472 18770 7524 18776
rect 7392 18737 7420 18770
rect 7378 18728 7434 18737
rect 7378 18663 7434 18672
rect 7484 17882 7512 18770
rect 7760 18442 7788 19314
rect 7668 18414 7788 18442
rect 7668 18290 7696 18414
rect 7656 18284 7708 18290
rect 7656 18226 7708 18232
rect 7472 17876 7524 17882
rect 7472 17818 7524 17824
rect 7564 17876 7616 17882
rect 7564 17818 7616 17824
rect 7472 16992 7524 16998
rect 7472 16934 7524 16940
rect 7288 16788 7340 16794
rect 7288 16730 7340 16736
rect 7378 16552 7434 16561
rect 7378 16487 7434 16496
rect 7286 13968 7342 13977
rect 7286 13903 7342 13912
rect 7196 13728 7248 13734
rect 7196 13670 7248 13676
rect 7300 10826 7328 13903
rect 7208 10810 7328 10826
rect 7196 10804 7328 10810
rect 7248 10798 7328 10804
rect 7196 10746 7248 10752
rect 7196 10192 7248 10198
rect 7286 10160 7342 10169
rect 7248 10140 7286 10146
rect 7196 10134 7286 10140
rect 7208 10118 7286 10134
rect 7286 10095 7342 10104
rect 7196 9512 7248 9518
rect 7196 9454 7248 9460
rect 7208 8945 7236 9454
rect 7300 9178 7328 10095
rect 7288 9172 7340 9178
rect 7288 9114 7340 9120
rect 7194 8936 7250 8945
rect 7194 8871 7250 8880
rect 7288 8016 7340 8022
rect 7288 7958 7340 7964
rect 7104 6452 7156 6458
rect 7104 6394 7156 6400
rect 7300 4010 7328 7958
rect 7392 7546 7420 16487
rect 7484 16250 7512 16934
rect 7472 16244 7524 16250
rect 7472 16186 7524 16192
rect 7576 16130 7604 17818
rect 7748 17672 7800 17678
rect 7748 17614 7800 17620
rect 7760 17270 7788 17614
rect 7748 17264 7800 17270
rect 7748 17206 7800 17212
rect 7656 16176 7708 16182
rect 7576 16124 7656 16130
rect 7576 16118 7708 16124
rect 7576 16102 7696 16118
rect 7470 14512 7526 14521
rect 7470 14447 7526 14456
rect 7484 11898 7512 14447
rect 7576 13870 7604 16102
rect 7656 16040 7708 16046
rect 7656 15982 7708 15988
rect 7668 15162 7696 15982
rect 7748 15904 7800 15910
rect 7748 15846 7800 15852
rect 7760 15706 7788 15846
rect 7748 15700 7800 15706
rect 7748 15642 7800 15648
rect 7656 15156 7708 15162
rect 7656 15098 7708 15104
rect 7852 15026 7880 19858
rect 8772 19718 8800 21966
rect 9034 21584 9090 21593
rect 9034 21519 9090 21528
rect 9048 21486 9076 21519
rect 8944 21480 8996 21486
rect 8942 21448 8944 21457
rect 9036 21480 9088 21486
rect 8996 21448 8998 21457
rect 9036 21422 9088 21428
rect 8942 21383 8998 21392
rect 9036 20936 9088 20942
rect 9036 20878 9088 20884
rect 8852 20800 8904 20806
rect 8852 20742 8904 20748
rect 8864 20398 8892 20742
rect 8852 20392 8904 20398
rect 8850 20360 8852 20369
rect 8904 20360 8906 20369
rect 8850 20295 8906 20304
rect 8942 19816 8998 19825
rect 8942 19751 8998 19760
rect 8116 19712 8168 19718
rect 8116 19654 8168 19660
rect 8300 19712 8352 19718
rect 8300 19654 8352 19660
rect 8760 19712 8812 19718
rect 8760 19654 8812 19660
rect 7930 19408 7986 19417
rect 7930 19343 7932 19352
rect 7984 19343 7986 19352
rect 7932 19314 7984 19320
rect 8024 18896 8076 18902
rect 8024 18838 8076 18844
rect 7932 18760 7984 18766
rect 7932 18702 7984 18708
rect 7944 17066 7972 18702
rect 8036 18222 8064 18838
rect 8128 18222 8156 19654
rect 8208 19304 8260 19310
rect 8312 19292 8340 19654
rect 8260 19264 8340 19292
rect 8208 19246 8260 19252
rect 8353 19068 8649 19088
rect 8409 19066 8433 19068
rect 8489 19066 8513 19068
rect 8569 19066 8593 19068
rect 8431 19014 8433 19066
rect 8495 19014 8507 19066
rect 8569 19014 8571 19066
rect 8409 19012 8433 19014
rect 8489 19012 8513 19014
rect 8569 19012 8593 19014
rect 8353 18992 8649 19012
rect 8760 18692 8812 18698
rect 8760 18634 8812 18640
rect 8208 18624 8260 18630
rect 8484 18624 8536 18630
rect 8208 18566 8260 18572
rect 8482 18592 8484 18601
rect 8536 18592 8538 18601
rect 8024 18216 8076 18222
rect 8024 18158 8076 18164
rect 8116 18216 8168 18222
rect 8116 18158 8168 18164
rect 8220 17864 8248 18566
rect 8482 18527 8538 18536
rect 8353 17980 8649 18000
rect 8409 17978 8433 17980
rect 8489 17978 8513 17980
rect 8569 17978 8593 17980
rect 8431 17926 8433 17978
rect 8495 17926 8507 17978
rect 8569 17926 8571 17978
rect 8409 17924 8433 17926
rect 8489 17924 8513 17926
rect 8569 17924 8593 17926
rect 8353 17904 8649 17924
rect 8128 17836 8248 17864
rect 8128 17746 8156 17836
rect 8772 17814 8800 18634
rect 8852 18420 8904 18426
rect 8852 18362 8904 18368
rect 8864 17882 8892 18362
rect 8852 17876 8904 17882
rect 8852 17818 8904 17824
rect 8760 17808 8812 17814
rect 8760 17750 8812 17756
rect 8116 17740 8168 17746
rect 8116 17682 8168 17688
rect 7932 17060 7984 17066
rect 7932 17002 7984 17008
rect 8128 16998 8156 17682
rect 8956 17678 8984 19751
rect 9048 19242 9076 20878
rect 9312 20324 9364 20330
rect 9312 20266 9364 20272
rect 9126 20088 9182 20097
rect 9126 20023 9182 20032
rect 9140 19446 9168 20023
rect 9220 19916 9272 19922
rect 9220 19858 9272 19864
rect 9128 19440 9180 19446
rect 9128 19382 9180 19388
rect 9128 19304 9180 19310
rect 9128 19246 9180 19252
rect 9036 19236 9088 19242
rect 9036 19178 9088 19184
rect 9140 18426 9168 19246
rect 9128 18420 9180 18426
rect 9128 18362 9180 18368
rect 9128 17740 9180 17746
rect 9128 17682 9180 17688
rect 8944 17672 8996 17678
rect 9140 17649 9168 17682
rect 8944 17614 8996 17620
rect 9126 17640 9182 17649
rect 9126 17575 9182 17584
rect 8392 17536 8444 17542
rect 8392 17478 8444 17484
rect 8404 17338 8432 17478
rect 8392 17332 8444 17338
rect 8392 17274 8444 17280
rect 8300 17128 8352 17134
rect 8220 17088 8300 17116
rect 8116 16992 8168 16998
rect 8116 16934 8168 16940
rect 8220 16794 8248 17088
rect 8300 17070 8352 17076
rect 8353 16892 8649 16912
rect 8409 16890 8433 16892
rect 8489 16890 8513 16892
rect 8569 16890 8593 16892
rect 8431 16838 8433 16890
rect 8495 16838 8507 16890
rect 8569 16838 8571 16890
rect 8409 16836 8433 16838
rect 8489 16836 8513 16838
rect 8569 16836 8593 16838
rect 8353 16816 8649 16836
rect 8208 16788 8260 16794
rect 8208 16730 8260 16736
rect 7932 16652 7984 16658
rect 7932 16594 7984 16600
rect 8208 16652 8260 16658
rect 8208 16594 8260 16600
rect 8760 16652 8812 16658
rect 8760 16594 8812 16600
rect 7944 16114 7972 16594
rect 8116 16176 8168 16182
rect 8116 16118 8168 16124
rect 7932 16108 7984 16114
rect 7932 16050 7984 16056
rect 8128 15570 8156 16118
rect 8116 15564 8168 15570
rect 8116 15506 8168 15512
rect 7932 15156 7984 15162
rect 7932 15098 7984 15104
rect 7840 15020 7892 15026
rect 7840 14962 7892 14968
rect 7748 14476 7800 14482
rect 7748 14418 7800 14424
rect 7564 13864 7616 13870
rect 7564 13806 7616 13812
rect 7564 13728 7616 13734
rect 7564 13670 7616 13676
rect 7472 11892 7524 11898
rect 7472 11834 7524 11840
rect 7470 9480 7526 9489
rect 7470 9415 7526 9424
rect 7484 9382 7512 9415
rect 7472 9376 7524 9382
rect 7472 9318 7524 9324
rect 7472 9104 7524 9110
rect 7472 9046 7524 9052
rect 7484 8673 7512 9046
rect 7470 8664 7526 8673
rect 7470 8599 7526 8608
rect 7380 7540 7432 7546
rect 7380 7482 7432 7488
rect 7576 7002 7604 13670
rect 7760 13530 7788 14418
rect 7748 13524 7800 13530
rect 7748 13466 7800 13472
rect 7944 13394 7972 15098
rect 8220 15026 8248 16594
rect 8353 15804 8649 15824
rect 8409 15802 8433 15804
rect 8489 15802 8513 15804
rect 8569 15802 8593 15804
rect 8431 15750 8433 15802
rect 8495 15750 8507 15802
rect 8569 15750 8571 15802
rect 8409 15748 8433 15750
rect 8489 15748 8513 15750
rect 8569 15748 8593 15750
rect 8353 15728 8649 15748
rect 8484 15564 8536 15570
rect 8484 15506 8536 15512
rect 8024 15020 8076 15026
rect 8024 14962 8076 14968
rect 8208 15020 8260 15026
rect 8208 14962 8260 14968
rect 8036 14482 8064 14962
rect 8496 14958 8524 15506
rect 8772 15094 8800 16594
rect 9232 16454 9260 19858
rect 9324 19825 9352 20266
rect 9416 20233 9444 22034
rect 9508 20330 9536 22850
rect 9680 22092 9732 22098
rect 9680 22034 9732 22040
rect 9692 22001 9720 22034
rect 9678 21992 9734 22001
rect 9678 21927 9734 21936
rect 9772 21344 9824 21350
rect 9772 21286 9824 21292
rect 9588 20868 9640 20874
rect 9588 20810 9640 20816
rect 9496 20324 9548 20330
rect 9496 20266 9548 20272
rect 9402 20224 9458 20233
rect 9600 20210 9628 20810
rect 9402 20159 9458 20168
rect 9508 20182 9628 20210
rect 9508 19938 9536 20182
rect 9586 20088 9642 20097
rect 9642 20058 9720 20074
rect 9642 20052 9732 20058
rect 9642 20046 9680 20052
rect 9586 20023 9642 20032
rect 9680 19994 9732 20000
rect 9508 19922 9720 19938
rect 9508 19916 9732 19922
rect 9508 19910 9680 19916
rect 9680 19858 9732 19864
rect 9310 19816 9366 19825
rect 9310 19751 9366 19760
rect 9402 19680 9458 19689
rect 9402 19615 9458 19624
rect 9416 19446 9444 19615
rect 9494 19544 9550 19553
rect 9494 19479 9550 19488
rect 9404 19440 9456 19446
rect 9404 19382 9456 19388
rect 9312 17672 9364 17678
rect 9310 17640 9312 17649
rect 9364 17640 9366 17649
rect 9310 17575 9366 17584
rect 9416 17338 9444 19382
rect 9508 18766 9536 19479
rect 9680 19304 9732 19310
rect 9586 19272 9642 19281
rect 9680 19246 9732 19252
rect 9586 19207 9642 19216
rect 9600 19174 9628 19207
rect 9588 19168 9640 19174
rect 9588 19110 9640 19116
rect 9496 18760 9548 18766
rect 9496 18702 9548 18708
rect 9508 18057 9536 18702
rect 9494 18048 9550 18057
rect 9494 17983 9550 17992
rect 9496 17672 9548 17678
rect 9496 17614 9548 17620
rect 9404 17332 9456 17338
rect 9404 17274 9456 17280
rect 9508 17134 9536 17614
rect 9496 17128 9548 17134
rect 9496 17070 9548 17076
rect 9496 16652 9548 16658
rect 9496 16594 9548 16600
rect 9220 16448 9272 16454
rect 9048 16396 9220 16402
rect 9048 16390 9272 16396
rect 9048 16374 9260 16390
rect 8942 16144 8998 16153
rect 8852 16108 8904 16114
rect 8942 16079 8944 16088
rect 8852 16050 8904 16056
rect 8996 16079 8998 16088
rect 8944 16050 8996 16056
rect 8864 15366 8892 16050
rect 8944 15632 8996 15638
rect 8944 15574 8996 15580
rect 8852 15360 8904 15366
rect 8852 15302 8904 15308
rect 8760 15088 8812 15094
rect 8760 15030 8812 15036
rect 8300 14952 8352 14958
rect 8220 14900 8300 14906
rect 8220 14894 8352 14900
rect 8484 14952 8536 14958
rect 8484 14894 8536 14900
rect 8668 14952 8720 14958
rect 8668 14894 8720 14900
rect 8220 14878 8340 14894
rect 8220 14618 8248 14878
rect 8353 14716 8649 14736
rect 8409 14714 8433 14716
rect 8489 14714 8513 14716
rect 8569 14714 8593 14716
rect 8431 14662 8433 14714
rect 8495 14662 8507 14714
rect 8569 14662 8571 14714
rect 8409 14660 8433 14662
rect 8489 14660 8513 14662
rect 8569 14660 8593 14662
rect 8353 14640 8649 14660
rect 8208 14612 8260 14618
rect 8208 14554 8260 14560
rect 8680 14550 8708 14894
rect 8772 14890 8800 15030
rect 8760 14884 8812 14890
rect 8760 14826 8812 14832
rect 8668 14544 8720 14550
rect 8668 14486 8720 14492
rect 8024 14476 8076 14482
rect 8024 14418 8076 14424
rect 8760 14476 8812 14482
rect 8760 14418 8812 14424
rect 8668 14408 8720 14414
rect 8668 14350 8720 14356
rect 8024 14340 8076 14346
rect 8024 14282 8076 14288
rect 7932 13388 7984 13394
rect 7932 13330 7984 13336
rect 7656 12980 7708 12986
rect 7656 12922 7708 12928
rect 7668 9042 7696 12922
rect 7748 11892 7800 11898
rect 7748 11834 7800 11840
rect 7760 9178 7788 11834
rect 7932 11552 7984 11558
rect 7932 11494 7984 11500
rect 7840 10736 7892 10742
rect 7840 10678 7892 10684
rect 7852 10266 7880 10678
rect 7944 10606 7972 11494
rect 7932 10600 7984 10606
rect 7932 10542 7984 10548
rect 7840 10260 7892 10266
rect 7840 10202 7892 10208
rect 7930 9480 7986 9489
rect 7930 9415 7986 9424
rect 7840 9376 7892 9382
rect 7840 9318 7892 9324
rect 7748 9172 7800 9178
rect 7748 9114 7800 9120
rect 7656 9036 7708 9042
rect 7656 8978 7708 8984
rect 7852 8974 7880 9318
rect 7840 8968 7892 8974
rect 7840 8910 7892 8916
rect 7944 8498 7972 9415
rect 7932 8492 7984 8498
rect 7932 8434 7984 8440
rect 7656 8356 7708 8362
rect 7656 8298 7708 8304
rect 7564 6996 7616 7002
rect 7564 6938 7616 6944
rect 7562 6760 7618 6769
rect 7562 6695 7564 6704
rect 7616 6695 7618 6704
rect 7564 6666 7616 6672
rect 7668 5642 7696 8298
rect 7932 7880 7984 7886
rect 7932 7822 7984 7828
rect 7944 7342 7972 7822
rect 7932 7336 7984 7342
rect 7932 7278 7984 7284
rect 8036 5914 8064 14282
rect 8680 14074 8708 14350
rect 8668 14068 8720 14074
rect 8668 14010 8720 14016
rect 8668 13864 8720 13870
rect 8668 13806 8720 13812
rect 8680 13734 8708 13806
rect 8668 13728 8720 13734
rect 8668 13670 8720 13676
rect 8353 13628 8649 13648
rect 8409 13626 8433 13628
rect 8489 13626 8513 13628
rect 8569 13626 8593 13628
rect 8431 13574 8433 13626
rect 8495 13574 8507 13626
rect 8569 13574 8571 13626
rect 8409 13572 8433 13574
rect 8489 13572 8513 13574
rect 8569 13572 8593 13574
rect 8353 13552 8649 13572
rect 8680 13462 8708 13670
rect 8668 13456 8720 13462
rect 8668 13398 8720 13404
rect 8484 13184 8536 13190
rect 8484 13126 8536 13132
rect 8496 12782 8524 13126
rect 8772 12986 8800 14418
rect 8852 14272 8904 14278
rect 8852 14214 8904 14220
rect 8760 12980 8812 12986
rect 8760 12922 8812 12928
rect 8484 12776 8536 12782
rect 8484 12718 8536 12724
rect 8208 12640 8260 12646
rect 8208 12582 8260 12588
rect 8220 12442 8248 12582
rect 8353 12540 8649 12560
rect 8409 12538 8433 12540
rect 8489 12538 8513 12540
rect 8569 12538 8593 12540
rect 8431 12486 8433 12538
rect 8495 12486 8507 12538
rect 8569 12486 8571 12538
rect 8409 12484 8433 12486
rect 8489 12484 8513 12486
rect 8569 12484 8593 12486
rect 8353 12464 8649 12484
rect 8208 12436 8260 12442
rect 8208 12378 8260 12384
rect 8864 12306 8892 14214
rect 8956 12345 8984 15574
rect 9048 14498 9076 16374
rect 9220 16244 9272 16250
rect 9220 16186 9272 16192
rect 9128 14884 9180 14890
rect 9128 14826 9180 14832
rect 9140 14618 9168 14826
rect 9128 14612 9180 14618
rect 9128 14554 9180 14560
rect 9048 14470 9168 14498
rect 9036 13728 9088 13734
rect 9036 13670 9088 13676
rect 9048 13258 9076 13670
rect 9036 13252 9088 13258
rect 9036 13194 9088 13200
rect 9036 12640 9088 12646
rect 9036 12582 9088 12588
rect 8942 12336 8998 12345
rect 8852 12300 8904 12306
rect 8942 12271 8998 12280
rect 8852 12242 8904 12248
rect 8208 12164 8260 12170
rect 8208 12106 8260 12112
rect 8220 11898 8248 12106
rect 9048 12102 9076 12582
rect 9140 12306 9168 14470
rect 9232 13394 9260 16186
rect 9312 16040 9364 16046
rect 9312 15982 9364 15988
rect 9324 15706 9352 15982
rect 9402 15872 9458 15881
rect 9402 15807 9458 15816
rect 9312 15700 9364 15706
rect 9312 15642 9364 15648
rect 9312 14000 9364 14006
rect 9312 13942 9364 13948
rect 9220 13388 9272 13394
rect 9220 13330 9272 13336
rect 9220 13184 9272 13190
rect 9218 13152 9220 13161
rect 9272 13152 9274 13161
rect 9218 13087 9274 13096
rect 9324 12850 9352 13942
rect 9312 12844 9364 12850
rect 9312 12786 9364 12792
rect 9128 12300 9180 12306
rect 9128 12242 9180 12248
rect 8300 12096 8352 12102
rect 8300 12038 8352 12044
rect 8392 12096 8444 12102
rect 8392 12038 8444 12044
rect 9036 12096 9088 12102
rect 9036 12038 9088 12044
rect 8312 11898 8340 12038
rect 8208 11892 8260 11898
rect 8208 11834 8260 11840
rect 8300 11892 8352 11898
rect 8300 11834 8352 11840
rect 8116 11824 8168 11830
rect 8116 11766 8168 11772
rect 8128 9042 8156 11766
rect 8208 11688 8260 11694
rect 8208 11630 8260 11636
rect 8220 11218 8248 11630
rect 8404 11626 8432 12038
rect 9324 11762 9352 12786
rect 9312 11756 9364 11762
rect 9312 11698 9364 11704
rect 8392 11620 8444 11626
rect 8392 11562 8444 11568
rect 8353 11452 8649 11472
rect 8409 11450 8433 11452
rect 8489 11450 8513 11452
rect 8569 11450 8593 11452
rect 8431 11398 8433 11450
rect 8495 11398 8507 11450
rect 8569 11398 8571 11450
rect 8409 11396 8433 11398
rect 8489 11396 8513 11398
rect 8569 11396 8593 11398
rect 8353 11376 8649 11396
rect 8208 11212 8260 11218
rect 8208 11154 8260 11160
rect 8760 11212 8812 11218
rect 8760 11154 8812 11160
rect 8220 10810 8248 11154
rect 8300 11008 8352 11014
rect 8300 10950 8352 10956
rect 8208 10804 8260 10810
rect 8208 10746 8260 10752
rect 8312 10538 8340 10950
rect 8300 10532 8352 10538
rect 8220 10492 8300 10520
rect 8220 10198 8248 10492
rect 8300 10474 8352 10480
rect 8312 10409 8340 10474
rect 8668 10464 8720 10470
rect 8668 10406 8720 10412
rect 8353 10364 8649 10384
rect 8409 10362 8433 10364
rect 8489 10362 8513 10364
rect 8569 10362 8593 10364
rect 8431 10310 8433 10362
rect 8495 10310 8507 10362
rect 8569 10310 8571 10362
rect 8409 10308 8433 10310
rect 8489 10308 8513 10310
rect 8569 10308 8593 10310
rect 8353 10288 8649 10308
rect 8208 10192 8260 10198
rect 8208 10134 8260 10140
rect 8353 9276 8649 9296
rect 8409 9274 8433 9276
rect 8489 9274 8513 9276
rect 8569 9274 8593 9276
rect 8431 9222 8433 9274
rect 8495 9222 8507 9274
rect 8569 9222 8571 9274
rect 8409 9220 8433 9222
rect 8489 9220 8513 9222
rect 8569 9220 8593 9222
rect 8353 9200 8649 9220
rect 8680 9178 8708 10406
rect 8668 9172 8720 9178
rect 8668 9114 8720 9120
rect 8772 9058 8800 11154
rect 9324 11150 9352 11698
rect 9416 11354 9444 15807
rect 9508 15706 9536 16594
rect 9600 16028 9628 19110
rect 9692 18834 9720 19246
rect 9680 18828 9732 18834
rect 9680 18770 9732 18776
rect 9784 18222 9812 21286
rect 9876 20262 9904 23600
rect 10048 21956 10100 21962
rect 10048 21898 10100 21904
rect 10060 21690 10088 21898
rect 10048 21684 10100 21690
rect 10048 21626 10100 21632
rect 10232 21004 10284 21010
rect 10232 20946 10284 20952
rect 9956 20800 10008 20806
rect 9956 20742 10008 20748
rect 9968 20466 9996 20742
rect 10244 20602 10272 20946
rect 10520 20913 10548 23600
rect 10968 22160 11020 22166
rect 10968 22102 11020 22108
rect 10506 20904 10562 20913
rect 10506 20839 10562 20848
rect 10232 20596 10284 20602
rect 10232 20538 10284 20544
rect 10414 20496 10470 20505
rect 9956 20460 10008 20466
rect 9956 20402 10008 20408
rect 10232 20460 10284 20466
rect 10414 20431 10470 20440
rect 10232 20402 10284 20408
rect 9864 20256 9916 20262
rect 9864 20198 9916 20204
rect 9862 20088 9918 20097
rect 9862 20023 9864 20032
rect 9916 20023 9918 20032
rect 9864 19994 9916 20000
rect 10244 19718 10272 20402
rect 10428 20398 10456 20431
rect 10416 20392 10468 20398
rect 10416 20334 10468 20340
rect 10600 20052 10652 20058
rect 10600 19994 10652 20000
rect 10416 19780 10468 19786
rect 10416 19722 10468 19728
rect 10232 19712 10284 19718
rect 10232 19654 10284 19660
rect 10046 19408 10102 19417
rect 10046 19343 10102 19352
rect 9864 19168 9916 19174
rect 10060 19145 10088 19343
rect 10244 19292 10272 19654
rect 10324 19304 10376 19310
rect 10244 19264 10324 19292
rect 10324 19246 10376 19252
rect 9864 19110 9916 19116
rect 10046 19136 10102 19145
rect 9680 18216 9732 18222
rect 9680 18158 9732 18164
rect 9772 18216 9824 18222
rect 9772 18158 9824 18164
rect 9692 16266 9720 18158
rect 9784 17354 9812 18158
rect 9876 17814 9904 19110
rect 10046 19071 10102 19080
rect 10060 18766 10088 19071
rect 10324 18828 10376 18834
rect 10428 18816 10456 19722
rect 10508 19304 10560 19310
rect 10508 19246 10560 19252
rect 10376 18788 10456 18816
rect 10324 18770 10376 18776
rect 10048 18760 10100 18766
rect 10048 18702 10100 18708
rect 10140 18760 10192 18766
rect 10140 18702 10192 18708
rect 10060 18154 10088 18702
rect 10048 18148 10100 18154
rect 10048 18090 10100 18096
rect 9864 17808 9916 17814
rect 9864 17750 9916 17756
rect 9784 17338 9904 17354
rect 9784 17332 9916 17338
rect 9784 17326 9864 17332
rect 9864 17274 9916 17280
rect 9956 17060 10008 17066
rect 9956 17002 10008 17008
rect 9968 16289 9996 17002
rect 10060 16726 10088 18090
rect 10048 16720 10100 16726
rect 10048 16662 10100 16668
rect 10152 16658 10180 18702
rect 10140 16652 10192 16658
rect 10140 16594 10192 16600
rect 10324 16652 10376 16658
rect 10324 16594 10376 16600
rect 9954 16280 10010 16289
rect 9692 16238 9904 16266
rect 9680 16040 9732 16046
rect 9600 16000 9680 16028
rect 9680 15982 9732 15988
rect 9876 15706 9904 16238
rect 9954 16215 10010 16224
rect 9496 15700 9548 15706
rect 9496 15642 9548 15648
rect 9864 15700 9916 15706
rect 9864 15642 9916 15648
rect 9508 13530 9536 15642
rect 9680 15360 9732 15366
rect 9680 15302 9732 15308
rect 9692 14414 9720 15302
rect 9968 15162 9996 16215
rect 10232 16176 10284 16182
rect 10336 16153 10364 16594
rect 10428 16590 10456 18788
rect 10520 18222 10548 19246
rect 10612 19145 10640 19994
rect 10598 19136 10654 19145
rect 10598 19071 10654 19080
rect 10980 18714 11008 22102
rect 11060 20800 11112 20806
rect 11060 20742 11112 20748
rect 11072 20330 11100 20742
rect 11060 20324 11112 20330
rect 11060 20266 11112 20272
rect 11164 20262 11192 23600
rect 11612 21888 11664 21894
rect 11612 21830 11664 21836
rect 11336 21616 11388 21622
rect 11336 21558 11388 21564
rect 11428 21616 11480 21622
rect 11428 21558 11480 21564
rect 11244 21344 11296 21350
rect 11244 21286 11296 21292
rect 11256 20806 11284 21286
rect 11244 20800 11296 20806
rect 11244 20742 11296 20748
rect 11152 20256 11204 20262
rect 11058 20224 11114 20233
rect 11152 20198 11204 20204
rect 11058 20159 11114 20168
rect 11072 19836 11100 20159
rect 11256 20074 11284 20742
rect 11164 20046 11284 20074
rect 11164 19961 11192 20046
rect 11150 19952 11206 19961
rect 11150 19887 11206 19896
rect 11072 19808 11192 19836
rect 11060 19712 11112 19718
rect 11060 19654 11112 19660
rect 11072 19242 11100 19654
rect 11060 19236 11112 19242
rect 11060 19178 11112 19184
rect 11072 18834 11100 19178
rect 11164 18834 11192 19808
rect 11348 19242 11376 21558
rect 11440 21350 11468 21558
rect 11624 21554 11652 21830
rect 11520 21548 11572 21554
rect 11520 21490 11572 21496
rect 11612 21548 11664 21554
rect 11612 21490 11664 21496
rect 11428 21344 11480 21350
rect 11428 21286 11480 21292
rect 11532 21078 11560 21490
rect 11612 21344 11664 21350
rect 11612 21286 11664 21292
rect 11520 21072 11572 21078
rect 11520 21014 11572 21020
rect 11532 20602 11560 21014
rect 11520 20596 11572 20602
rect 11520 20538 11572 20544
rect 11624 20346 11652 21286
rect 11532 20318 11652 20346
rect 11704 20324 11756 20330
rect 11428 19848 11480 19854
rect 11428 19790 11480 19796
rect 11336 19236 11388 19242
rect 11336 19178 11388 19184
rect 11060 18828 11112 18834
rect 11060 18770 11112 18776
rect 11152 18828 11204 18834
rect 11152 18770 11204 18776
rect 10980 18686 11376 18714
rect 11058 18320 11114 18329
rect 11058 18255 11114 18264
rect 10508 18216 10560 18222
rect 10508 18158 10560 18164
rect 10520 17882 10548 18158
rect 10508 17876 10560 17882
rect 10508 17818 10560 17824
rect 10600 17876 10652 17882
rect 11072 17864 11100 18255
rect 11244 18148 11296 18154
rect 11244 18090 11296 18096
rect 10600 17818 10652 17824
rect 10980 17836 11100 17864
rect 10612 17785 10640 17818
rect 10598 17776 10654 17785
rect 10598 17711 10654 17720
rect 10980 17218 11008 17836
rect 11152 17808 11204 17814
rect 11152 17750 11204 17756
rect 11060 17740 11112 17746
rect 11060 17682 11112 17688
rect 11072 17338 11100 17682
rect 11164 17338 11192 17750
rect 11256 17542 11284 18090
rect 11348 17762 11376 18686
rect 11440 17882 11468 19790
rect 11532 18426 11560 20318
rect 11704 20266 11756 20272
rect 11612 20256 11664 20262
rect 11612 20198 11664 20204
rect 11520 18420 11572 18426
rect 11520 18362 11572 18368
rect 11428 17876 11480 17882
rect 11428 17818 11480 17824
rect 11348 17734 11560 17762
rect 11244 17536 11296 17542
rect 11244 17478 11296 17484
rect 11060 17332 11112 17338
rect 11060 17274 11112 17280
rect 11152 17332 11204 17338
rect 11152 17274 11204 17280
rect 10980 17190 11192 17218
rect 10416 16584 10468 16590
rect 10692 16584 10744 16590
rect 10468 16532 10548 16538
rect 10416 16526 10548 16532
rect 10692 16526 10744 16532
rect 10968 16584 11020 16590
rect 10968 16526 11020 16532
rect 10428 16510 10548 16526
rect 10232 16118 10284 16124
rect 10322 16144 10378 16153
rect 10140 16040 10192 16046
rect 10140 15982 10192 15988
rect 10048 15564 10100 15570
rect 10048 15506 10100 15512
rect 9956 15156 10008 15162
rect 9956 15098 10008 15104
rect 9680 14408 9732 14414
rect 9680 14350 9732 14356
rect 9496 13524 9548 13530
rect 9496 13466 9548 13472
rect 9692 13410 9720 14350
rect 9954 13832 10010 13841
rect 10060 13802 10088 15506
rect 10152 14822 10180 15982
rect 10244 15638 10272 16118
rect 10322 16079 10378 16088
rect 10232 15632 10284 15638
rect 10232 15574 10284 15580
rect 10140 14816 10192 14822
rect 10140 14758 10192 14764
rect 9954 13767 10010 13776
rect 10048 13796 10100 13802
rect 9968 13462 9996 13767
rect 10048 13738 10100 13744
rect 10152 13682 10180 14758
rect 10060 13654 10180 13682
rect 10232 13728 10284 13734
rect 10232 13670 10284 13676
rect 9600 13382 9720 13410
rect 9956 13456 10008 13462
rect 9956 13398 10008 13404
rect 9600 12730 9628 13382
rect 9680 13320 9732 13326
rect 9680 13262 9732 13268
rect 9692 12986 9720 13262
rect 9956 13184 10008 13190
rect 9956 13126 10008 13132
rect 9680 12980 9732 12986
rect 9680 12922 9732 12928
rect 9692 12832 9720 12922
rect 9692 12804 9812 12832
rect 9600 12702 9720 12730
rect 9692 12442 9720 12702
rect 9680 12436 9732 12442
rect 9680 12378 9732 12384
rect 9680 11688 9732 11694
rect 9586 11656 9642 11665
rect 9680 11630 9732 11636
rect 9586 11591 9642 11600
rect 9404 11348 9456 11354
rect 9404 11290 9456 11296
rect 9600 11218 9628 11591
rect 9588 11212 9640 11218
rect 9588 11154 9640 11160
rect 9036 11144 9088 11150
rect 9312 11144 9364 11150
rect 9036 11086 9088 11092
rect 9232 11104 9312 11132
rect 8852 10464 8904 10470
rect 8852 10406 8904 10412
rect 8864 10266 8892 10406
rect 8852 10260 8904 10266
rect 8852 10202 8904 10208
rect 8864 9518 8892 10202
rect 9048 9654 9076 11086
rect 9232 10674 9260 11104
rect 9312 11086 9364 11092
rect 9312 10736 9364 10742
rect 9692 10713 9720 11630
rect 9784 10742 9812 12804
rect 9968 11830 9996 13126
rect 10060 12782 10088 13654
rect 10244 13530 10272 13670
rect 10232 13524 10284 13530
rect 10232 13466 10284 13472
rect 10140 13388 10192 13394
rect 10140 13330 10192 13336
rect 10152 12850 10180 13330
rect 10232 13252 10284 13258
rect 10232 13194 10284 13200
rect 10140 12844 10192 12850
rect 10140 12786 10192 12792
rect 10244 12782 10272 13194
rect 10039 12776 10091 12782
rect 10039 12718 10091 12724
rect 10232 12776 10284 12782
rect 10232 12718 10284 12724
rect 10244 12594 10272 12718
rect 10060 12566 10272 12594
rect 10060 12102 10088 12566
rect 10336 12458 10364 16079
rect 10416 15904 10468 15910
rect 10520 15892 10548 16510
rect 10468 15864 10548 15892
rect 10416 15846 10468 15852
rect 10520 15366 10548 15864
rect 10600 15496 10652 15502
rect 10600 15438 10652 15444
rect 10508 15360 10560 15366
rect 10508 15302 10560 15308
rect 10612 14958 10640 15438
rect 10600 14952 10652 14958
rect 10598 14920 10600 14929
rect 10652 14920 10654 14929
rect 10598 14855 10654 14864
rect 10416 14272 10468 14278
rect 10416 14214 10468 14220
rect 10428 13938 10456 14214
rect 10416 13932 10468 13938
rect 10416 13874 10468 13880
rect 10600 13932 10652 13938
rect 10600 13874 10652 13880
rect 10244 12430 10364 12458
rect 10048 12096 10100 12102
rect 10048 12038 10100 12044
rect 9956 11824 10008 11830
rect 9956 11766 10008 11772
rect 10060 11762 10088 12038
rect 10048 11756 10100 11762
rect 10048 11698 10100 11704
rect 9956 11280 10008 11286
rect 9956 11222 10008 11228
rect 9864 11076 9916 11082
rect 9864 11018 9916 11024
rect 9876 10985 9904 11018
rect 9862 10976 9918 10985
rect 9862 10911 9918 10920
rect 9772 10736 9824 10742
rect 9312 10678 9364 10684
rect 9678 10704 9734 10713
rect 9220 10668 9272 10674
rect 9220 10610 9272 10616
rect 9232 10062 9260 10610
rect 9220 10056 9272 10062
rect 9220 9998 9272 10004
rect 9036 9648 9088 9654
rect 9036 9590 9088 9596
rect 8852 9512 8904 9518
rect 8852 9454 8904 9460
rect 8944 9512 8996 9518
rect 8944 9454 8996 9460
rect 8956 9382 8984 9454
rect 8944 9376 8996 9382
rect 8944 9318 8996 9324
rect 9324 9110 9352 10678
rect 9772 10678 9824 10684
rect 9862 10704 9918 10713
rect 9678 10639 9734 10648
rect 9862 10639 9918 10648
rect 9876 10606 9904 10639
rect 9864 10600 9916 10606
rect 9864 10542 9916 10548
rect 9658 10296 9714 10305
rect 9876 10282 9904 10542
rect 9714 10266 9720 10282
rect 9714 10260 9732 10266
rect 9658 10231 9680 10240
rect 9680 10202 9732 10208
rect 9784 10254 9904 10282
rect 9784 10146 9812 10254
rect 9600 10130 9812 10146
rect 9864 10192 9916 10198
rect 9968 10180 9996 11222
rect 10060 11218 10088 11698
rect 10048 11212 10100 11218
rect 10048 11154 10100 11160
rect 10060 10713 10088 11154
rect 10046 10704 10102 10713
rect 10046 10639 10102 10648
rect 10046 10432 10102 10441
rect 10046 10367 10102 10376
rect 10060 10198 10088 10367
rect 9916 10152 9996 10180
rect 9864 10134 9916 10140
rect 9588 10124 9812 10130
rect 9640 10118 9812 10124
rect 9588 10066 9640 10072
rect 9588 9988 9640 9994
rect 9588 9930 9640 9936
rect 9312 9104 9364 9110
rect 8116 9036 8168 9042
rect 8116 8978 8168 8984
rect 8404 9030 8800 9058
rect 9218 9072 9274 9081
rect 9042 9036 9094 9042
rect 8208 8900 8260 8906
rect 8404 8888 8432 9030
rect 8956 8996 9042 9024
rect 8260 8860 8432 8888
rect 8496 8894 8708 8922
rect 8208 8842 8260 8848
rect 8392 8560 8444 8566
rect 8496 8548 8524 8894
rect 8576 8832 8628 8838
rect 8576 8774 8628 8780
rect 8444 8520 8524 8548
rect 8588 8548 8616 8774
rect 8680 8650 8708 8894
rect 8956 8650 8984 8996
rect 9312 9046 9364 9052
rect 9600 9058 9628 9930
rect 9672 9908 9700 10118
rect 9672 9880 9812 9908
rect 9678 9752 9734 9761
rect 9784 9722 9812 9880
rect 9862 9888 9918 9897
rect 9862 9823 9918 9832
rect 9678 9687 9734 9696
rect 9772 9716 9824 9722
rect 9692 9178 9720 9687
rect 9772 9658 9824 9664
rect 9680 9172 9732 9178
rect 9680 9114 9732 9120
rect 9600 9030 9720 9058
rect 9876 9042 9904 9823
rect 9968 9704 9996 10152
rect 10039 10192 10091 10198
rect 10039 10134 10091 10140
rect 10048 9716 10100 9722
rect 9968 9676 10048 9704
rect 10048 9658 10100 9664
rect 9218 9007 9274 9016
rect 9042 8978 9094 8984
rect 9232 8809 9260 9007
rect 9496 8900 9548 8906
rect 9496 8842 9548 8848
rect 9218 8800 9274 8809
rect 9218 8735 9274 8744
rect 8680 8622 8984 8650
rect 9508 8548 9536 8842
rect 8588 8520 9536 8548
rect 8392 8502 8444 8508
rect 8208 8288 8260 8294
rect 8208 8230 8260 8236
rect 9588 8288 9640 8294
rect 9588 8230 9640 8236
rect 8220 8072 8248 8230
rect 8353 8188 8649 8208
rect 8409 8186 8433 8188
rect 8489 8186 8513 8188
rect 8569 8186 8593 8188
rect 8431 8134 8433 8186
rect 8495 8134 8507 8186
rect 8569 8134 8571 8186
rect 8409 8132 8433 8134
rect 8489 8132 8513 8134
rect 8569 8132 8593 8134
rect 8353 8112 8649 8132
rect 9600 8090 9628 8230
rect 9588 8084 9640 8090
rect 8220 8044 8708 8072
rect 8300 7744 8352 7750
rect 8300 7686 8352 7692
rect 8312 7546 8340 7686
rect 8300 7540 8352 7546
rect 8300 7482 8352 7488
rect 8116 7404 8168 7410
rect 8116 7346 8168 7352
rect 8024 5908 8076 5914
rect 8024 5850 8076 5856
rect 7656 5636 7708 5642
rect 7656 5578 7708 5584
rect 8128 4282 8156 7346
rect 8353 7100 8649 7120
rect 8409 7098 8433 7100
rect 8489 7098 8513 7100
rect 8569 7098 8593 7100
rect 8431 7046 8433 7098
rect 8495 7046 8507 7098
rect 8569 7046 8571 7098
rect 8409 7044 8433 7046
rect 8489 7044 8513 7046
rect 8569 7044 8593 7046
rect 8353 7024 8649 7044
rect 8300 6792 8352 6798
rect 8300 6734 8352 6740
rect 8208 6656 8260 6662
rect 8208 6598 8260 6604
rect 8220 6254 8248 6598
rect 8312 6458 8340 6734
rect 8680 6730 8708 8044
rect 9588 8026 9640 8032
rect 9692 7818 9720 9030
rect 9864 9036 9916 9042
rect 9864 8978 9916 8984
rect 10244 8412 10272 12430
rect 10428 10588 10456 13874
rect 10508 13524 10560 13530
rect 10508 13466 10560 13472
rect 10520 11694 10548 13466
rect 10612 13462 10640 13874
rect 10600 13456 10652 13462
rect 10600 13398 10652 13404
rect 10704 12646 10732 16526
rect 10782 16144 10838 16153
rect 10782 16079 10838 16088
rect 10692 12640 10744 12646
rect 10692 12582 10744 12588
rect 10692 12300 10744 12306
rect 10692 12242 10744 12248
rect 10508 11688 10560 11694
rect 10508 11630 10560 11636
rect 10520 11354 10548 11630
rect 10508 11348 10560 11354
rect 10508 11290 10560 11296
rect 10704 11132 10732 12242
rect 10612 11104 10732 11132
rect 10508 10600 10560 10606
rect 10428 10560 10508 10588
rect 10508 10542 10560 10548
rect 10416 9648 10468 9654
rect 10416 9590 10468 9596
rect 10428 8430 10456 9590
rect 10520 8974 10548 10542
rect 10612 9110 10640 11104
rect 10692 9988 10744 9994
rect 10692 9930 10744 9936
rect 10704 9178 10732 9930
rect 10692 9172 10744 9178
rect 10692 9114 10744 9120
rect 10600 9104 10652 9110
rect 10600 9046 10652 9052
rect 10508 8968 10560 8974
rect 10508 8910 10560 8916
rect 10600 8968 10652 8974
rect 10600 8910 10652 8916
rect 10612 8430 10640 8910
rect 10692 8832 10744 8838
rect 10692 8774 10744 8780
rect 9876 8384 10272 8412
rect 9876 7886 9904 8384
rect 10140 8288 10192 8294
rect 10140 8230 10192 8236
rect 9956 7948 10008 7954
rect 9956 7890 10008 7896
rect 9864 7880 9916 7886
rect 9864 7822 9916 7828
rect 9680 7812 9732 7818
rect 9680 7754 9732 7760
rect 9036 7744 9088 7750
rect 9036 7686 9088 7692
rect 9048 7274 9076 7686
rect 9692 7562 9720 7754
rect 9508 7534 9720 7562
rect 9968 7546 9996 7890
rect 10152 7886 10180 8230
rect 10244 8129 10272 8384
rect 10416 8424 10468 8430
rect 10416 8366 10468 8372
rect 10600 8424 10652 8430
rect 10600 8366 10652 8372
rect 10230 8120 10286 8129
rect 10230 8055 10286 8064
rect 10612 7954 10640 8366
rect 10704 8265 10732 8774
rect 10690 8256 10746 8265
rect 10690 8191 10746 8200
rect 10324 7948 10376 7954
rect 10244 7908 10324 7936
rect 10140 7880 10192 7886
rect 10140 7822 10192 7828
rect 9956 7540 10008 7546
rect 8760 7268 8812 7274
rect 8760 7210 8812 7216
rect 9036 7268 9088 7274
rect 9036 7210 9088 7216
rect 8772 6730 8800 7210
rect 8852 7200 8904 7206
rect 8852 7142 8904 7148
rect 8944 7200 8996 7206
rect 8944 7142 8996 7148
rect 8864 7041 8892 7142
rect 8850 7032 8906 7041
rect 8850 6967 8906 6976
rect 8956 6866 8984 7142
rect 9048 6934 9076 7210
rect 9036 6928 9088 6934
rect 9036 6870 9088 6876
rect 8944 6860 8996 6866
rect 8944 6802 8996 6808
rect 8484 6724 8536 6730
rect 8484 6666 8536 6672
rect 8668 6724 8720 6730
rect 8668 6666 8720 6672
rect 8760 6724 8812 6730
rect 8760 6666 8812 6672
rect 8300 6452 8352 6458
rect 8300 6394 8352 6400
rect 8496 6361 8524 6666
rect 8668 6384 8720 6390
rect 8482 6352 8538 6361
rect 8668 6326 8720 6332
rect 8482 6287 8538 6296
rect 8208 6248 8260 6254
rect 8208 6190 8260 6196
rect 8353 6012 8649 6032
rect 8409 6010 8433 6012
rect 8489 6010 8513 6012
rect 8569 6010 8593 6012
rect 8431 5958 8433 6010
rect 8495 5958 8507 6010
rect 8569 5958 8571 6010
rect 8409 5956 8433 5958
rect 8489 5956 8513 5958
rect 8569 5956 8593 5958
rect 8353 5936 8649 5956
rect 8680 5273 8708 6326
rect 8772 6322 8800 6666
rect 8760 6316 8812 6322
rect 8760 6258 8812 6264
rect 8956 6186 8984 6802
rect 9508 6798 9536 7534
rect 9956 7482 10008 7488
rect 9680 7404 9732 7410
rect 9680 7346 9732 7352
rect 9586 7032 9642 7041
rect 9586 6967 9588 6976
rect 9640 6967 9642 6976
rect 9588 6938 9640 6944
rect 9692 6798 9720 7346
rect 10152 7342 10180 7822
rect 10244 7410 10272 7908
rect 10324 7890 10376 7896
rect 10600 7948 10652 7954
rect 10600 7890 10652 7896
rect 10324 7744 10376 7750
rect 10324 7686 10376 7692
rect 10232 7404 10284 7410
rect 10232 7346 10284 7352
rect 10336 7342 10364 7686
rect 10140 7336 10192 7342
rect 10140 7278 10192 7284
rect 10324 7336 10376 7342
rect 10324 7278 10376 7284
rect 10414 6896 10470 6905
rect 9772 6860 9824 6866
rect 9956 6860 10008 6866
rect 9824 6820 9904 6848
rect 9772 6802 9824 6808
rect 9496 6792 9548 6798
rect 9496 6734 9548 6740
rect 9680 6792 9732 6798
rect 9680 6734 9732 6740
rect 8944 6180 8996 6186
rect 8944 6122 8996 6128
rect 9692 5710 9720 6734
rect 9770 5808 9826 5817
rect 9770 5743 9772 5752
rect 9824 5743 9826 5752
rect 9772 5714 9824 5720
rect 9680 5704 9732 5710
rect 9680 5646 9732 5652
rect 8666 5264 8722 5273
rect 8666 5199 8722 5208
rect 9692 5166 9720 5646
rect 9404 5160 9456 5166
rect 9404 5102 9456 5108
rect 9680 5160 9732 5166
rect 9680 5102 9732 5108
rect 8944 5024 8996 5030
rect 8944 4966 8996 4972
rect 8353 4924 8649 4944
rect 8409 4922 8433 4924
rect 8489 4922 8513 4924
rect 8569 4922 8593 4924
rect 8431 4870 8433 4922
rect 8495 4870 8507 4922
rect 8569 4870 8571 4922
rect 8409 4868 8433 4870
rect 8489 4868 8513 4870
rect 8569 4868 8593 4870
rect 8353 4848 8649 4868
rect 8956 4486 8984 4966
rect 9416 4826 9444 5102
rect 9404 4820 9456 4826
rect 9404 4762 9456 4768
rect 8944 4480 8996 4486
rect 8944 4422 8996 4428
rect 8116 4276 8168 4282
rect 8116 4218 8168 4224
rect 7288 4004 7340 4010
rect 7288 3946 7340 3952
rect 8353 3836 8649 3856
rect 8409 3834 8433 3836
rect 8489 3834 8513 3836
rect 8569 3834 8593 3836
rect 8431 3782 8433 3834
rect 8495 3782 8507 3834
rect 8569 3782 8571 3834
rect 8409 3780 8433 3782
rect 8489 3780 8513 3782
rect 8569 3780 8593 3782
rect 8353 3760 8649 3780
rect 7012 2848 7064 2854
rect 7012 2790 7064 2796
rect 8353 2748 8649 2768
rect 8409 2746 8433 2748
rect 8489 2746 8513 2748
rect 8569 2746 8593 2748
rect 8431 2694 8433 2746
rect 8495 2694 8507 2746
rect 8569 2694 8571 2746
rect 8409 2692 8433 2694
rect 8489 2692 8513 2694
rect 8569 2692 8593 2694
rect 8353 2672 8649 2692
rect 6184 2372 6236 2378
rect 6184 2314 6236 2320
rect 9876 2310 9904 6820
rect 10414 6831 10470 6840
rect 9956 6802 10008 6808
rect 9968 6458 9996 6802
rect 9956 6452 10008 6458
rect 9956 6394 10008 6400
rect 10428 6254 10456 6831
rect 10692 6792 10744 6798
rect 10692 6734 10744 6740
rect 10704 6474 10732 6734
rect 10612 6446 10732 6474
rect 10612 6390 10640 6446
rect 10600 6384 10652 6390
rect 10600 6326 10652 6332
rect 10416 6248 10468 6254
rect 10416 6190 10468 6196
rect 10416 6112 10468 6118
rect 10416 6054 10468 6060
rect 10428 4826 10456 6054
rect 10416 4820 10468 4826
rect 10416 4762 10468 4768
rect 10796 4078 10824 16079
rect 10980 15978 11008 16526
rect 10968 15972 11020 15978
rect 10968 15914 11020 15920
rect 10966 14920 11022 14929
rect 10966 14855 11022 14864
rect 10980 14346 11008 14855
rect 11060 14612 11112 14618
rect 11060 14554 11112 14560
rect 11072 14521 11100 14554
rect 11058 14512 11114 14521
rect 11058 14447 11114 14456
rect 10968 14340 11020 14346
rect 10968 14282 11020 14288
rect 11164 14249 11192 17190
rect 11256 16658 11284 17478
rect 11336 16992 11388 16998
rect 11336 16934 11388 16940
rect 11244 16652 11296 16658
rect 11244 16594 11296 16600
rect 11244 16108 11296 16114
rect 11244 16050 11296 16056
rect 11256 16017 11284 16050
rect 11242 16008 11298 16017
rect 11242 15943 11298 15952
rect 11244 15904 11296 15910
rect 11244 15846 11296 15852
rect 11150 14240 11206 14249
rect 11150 14175 11206 14184
rect 11256 13870 11284 15846
rect 11348 15706 11376 16934
rect 11428 16108 11480 16114
rect 11428 16050 11480 16056
rect 11336 15700 11388 15706
rect 11336 15642 11388 15648
rect 11336 14612 11388 14618
rect 11336 14554 11388 14560
rect 11348 14482 11376 14554
rect 11336 14476 11388 14482
rect 11336 14418 11388 14424
rect 11336 14340 11388 14346
rect 11336 14282 11388 14288
rect 11244 13864 11296 13870
rect 11244 13806 11296 13812
rect 11152 13796 11204 13802
rect 11152 13738 11204 13744
rect 11164 13530 11192 13738
rect 11244 13728 11296 13734
rect 11244 13670 11296 13676
rect 11152 13524 11204 13530
rect 11152 13466 11204 13472
rect 10968 13456 11020 13462
rect 10968 13398 11020 13404
rect 10980 11898 11008 13398
rect 11256 13394 11284 13670
rect 11348 13569 11376 14282
rect 11334 13560 11390 13569
rect 11334 13495 11390 13504
rect 11244 13388 11296 13394
rect 11244 13330 11296 13336
rect 11256 12986 11284 13330
rect 11060 12980 11112 12986
rect 11060 12922 11112 12928
rect 11244 12980 11296 12986
rect 11244 12922 11296 12928
rect 11072 12617 11100 12922
rect 11336 12912 11388 12918
rect 11336 12854 11388 12860
rect 11152 12776 11204 12782
rect 11152 12718 11204 12724
rect 11058 12608 11114 12617
rect 11058 12543 11114 12552
rect 11164 11898 11192 12718
rect 11348 12696 11376 12854
rect 11256 12668 11376 12696
rect 10968 11892 11020 11898
rect 10968 11834 11020 11840
rect 11152 11892 11204 11898
rect 11152 11834 11204 11840
rect 11152 11212 11204 11218
rect 11152 11154 11204 11160
rect 10968 11076 11020 11082
rect 10968 11018 11020 11024
rect 10876 10804 10928 10810
rect 10876 10746 10928 10752
rect 10888 10713 10916 10746
rect 10874 10704 10930 10713
rect 10874 10639 10930 10648
rect 10980 10606 11008 11018
rect 11164 10810 11192 11154
rect 11152 10804 11204 10810
rect 11152 10746 11204 10752
rect 10968 10600 11020 10606
rect 10968 10542 11020 10548
rect 11060 10532 11112 10538
rect 11060 10474 11112 10480
rect 11072 10266 11100 10474
rect 11060 10260 11112 10266
rect 11060 10202 11112 10208
rect 11164 10198 11192 10746
rect 11152 10192 11204 10198
rect 11152 10134 11204 10140
rect 10968 9172 11020 9178
rect 10968 9114 11020 9120
rect 10876 9036 10928 9042
rect 10876 8978 10928 8984
rect 10888 7041 10916 8978
rect 10980 8362 11008 9114
rect 11152 8900 11204 8906
rect 11152 8842 11204 8848
rect 11164 8412 11192 8842
rect 11256 8650 11284 12668
rect 11440 10810 11468 16050
rect 11532 16046 11560 17734
rect 11520 16040 11572 16046
rect 11520 15982 11572 15988
rect 11520 14272 11572 14278
rect 11520 14214 11572 14220
rect 11532 13938 11560 14214
rect 11520 13932 11572 13938
rect 11520 13874 11572 13880
rect 11520 13728 11572 13734
rect 11520 13670 11572 13676
rect 11532 12442 11560 13670
rect 11520 12436 11572 12442
rect 11520 12378 11572 12384
rect 11520 12300 11572 12306
rect 11520 12242 11572 12248
rect 11532 12209 11560 12242
rect 11518 12200 11574 12209
rect 11518 12135 11574 12144
rect 11520 11348 11572 11354
rect 11520 11290 11572 11296
rect 11428 10804 11480 10810
rect 11428 10746 11480 10752
rect 11532 10305 11560 11290
rect 11624 11218 11652 20198
rect 11716 19378 11744 20266
rect 11808 19446 11836 23600
rect 12452 23582 12664 23600
rect 13096 23582 13676 23600
rect 12052 21788 12348 21808
rect 12108 21786 12132 21788
rect 12188 21786 12212 21788
rect 12268 21786 12292 21788
rect 12130 21734 12132 21786
rect 12194 21734 12206 21786
rect 12268 21734 12270 21786
rect 12108 21732 12132 21734
rect 12188 21732 12212 21734
rect 12268 21732 12292 21734
rect 12052 21712 12348 21732
rect 11888 21616 11940 21622
rect 11888 21558 11940 21564
rect 11796 19440 11848 19446
rect 11796 19382 11848 19388
rect 11704 19372 11756 19378
rect 11704 19314 11756 19320
rect 11704 19168 11756 19174
rect 11704 19110 11756 19116
rect 11716 18902 11744 19110
rect 11704 18896 11756 18902
rect 11704 18838 11756 18844
rect 11794 18728 11850 18737
rect 11704 18692 11756 18698
rect 11794 18663 11850 18672
rect 11704 18634 11756 18640
rect 11716 17066 11744 18634
rect 11808 18630 11836 18663
rect 11796 18624 11848 18630
rect 11796 18566 11848 18572
rect 11900 18086 11928 21558
rect 11980 21548 12032 21554
rect 11980 21490 12032 21496
rect 11992 21010 12020 21490
rect 12532 21412 12584 21418
rect 12532 21354 12584 21360
rect 12072 21344 12124 21350
rect 12072 21286 12124 21292
rect 12084 21146 12112 21286
rect 12072 21140 12124 21146
rect 12072 21082 12124 21088
rect 12544 21078 12572 21354
rect 12532 21072 12584 21078
rect 12532 21014 12584 21020
rect 11980 21004 12032 21010
rect 11980 20946 12032 20952
rect 12440 20868 12492 20874
rect 12440 20810 12492 20816
rect 11980 20800 12032 20806
rect 11980 20742 12032 20748
rect 11992 20330 12020 20742
rect 12052 20700 12348 20720
rect 12108 20698 12132 20700
rect 12188 20698 12212 20700
rect 12268 20698 12292 20700
rect 12130 20646 12132 20698
rect 12194 20646 12206 20698
rect 12268 20646 12270 20698
rect 12108 20644 12132 20646
rect 12188 20644 12212 20646
rect 12268 20644 12292 20646
rect 12052 20624 12348 20644
rect 12452 20534 12480 20810
rect 12532 20800 12584 20806
rect 12532 20742 12584 20748
rect 12440 20528 12492 20534
rect 12440 20470 12492 20476
rect 12440 20392 12492 20398
rect 12440 20334 12492 20340
rect 11980 20324 12032 20330
rect 11980 20266 12032 20272
rect 12052 19612 12348 19632
rect 12108 19610 12132 19612
rect 12188 19610 12212 19612
rect 12268 19610 12292 19612
rect 12130 19558 12132 19610
rect 12194 19558 12206 19610
rect 12268 19558 12270 19610
rect 12108 19556 12132 19558
rect 12188 19556 12212 19558
rect 12268 19556 12292 19558
rect 12052 19536 12348 19556
rect 11980 19168 12032 19174
rect 12452 19156 12480 20334
rect 12544 19310 12572 20742
rect 12532 19304 12584 19310
rect 12532 19246 12584 19252
rect 12452 19128 12572 19156
rect 11980 19110 12032 19116
rect 11888 18080 11940 18086
rect 11794 18048 11850 18057
rect 11888 18022 11940 18028
rect 11794 17983 11850 17992
rect 11704 17060 11756 17066
rect 11704 17002 11756 17008
rect 11702 16280 11758 16289
rect 11702 16215 11758 16224
rect 11716 16114 11744 16215
rect 11704 16108 11756 16114
rect 11704 16050 11756 16056
rect 11808 15910 11836 17983
rect 11992 17678 12020 19110
rect 12070 18728 12126 18737
rect 12070 18663 12072 18672
rect 12124 18663 12126 18672
rect 12072 18634 12124 18640
rect 12052 18524 12348 18544
rect 12108 18522 12132 18524
rect 12188 18522 12212 18524
rect 12268 18522 12292 18524
rect 12130 18470 12132 18522
rect 12194 18470 12206 18522
rect 12268 18470 12270 18522
rect 12108 18468 12132 18470
rect 12188 18468 12212 18470
rect 12268 18468 12292 18470
rect 12052 18448 12348 18468
rect 12440 18080 12492 18086
rect 12440 18022 12492 18028
rect 12452 17882 12480 18022
rect 12440 17876 12492 17882
rect 12440 17818 12492 17824
rect 12544 17746 12572 19128
rect 12532 17740 12584 17746
rect 12532 17682 12584 17688
rect 11980 17672 12032 17678
rect 11980 17614 12032 17620
rect 12530 17640 12586 17649
rect 12530 17575 12532 17584
rect 12584 17575 12586 17584
rect 12532 17546 12584 17552
rect 12052 17436 12348 17456
rect 12108 17434 12132 17436
rect 12188 17434 12212 17436
rect 12268 17434 12292 17436
rect 12130 17382 12132 17434
rect 12194 17382 12206 17434
rect 12268 17382 12270 17434
rect 12108 17380 12132 17382
rect 12188 17380 12212 17382
rect 12268 17380 12292 17382
rect 12052 17360 12348 17380
rect 12438 17368 12494 17377
rect 12438 17303 12494 17312
rect 12452 17218 12480 17303
rect 12268 17190 12480 17218
rect 11980 17128 12032 17134
rect 11978 17096 11980 17105
rect 12032 17096 12034 17105
rect 11978 17031 12034 17040
rect 12268 16522 12296 17190
rect 12440 17128 12492 17134
rect 12438 17096 12440 17105
rect 12492 17096 12494 17105
rect 12438 17031 12494 17040
rect 12348 16992 12400 16998
rect 12348 16934 12400 16940
rect 12360 16590 12388 16934
rect 12348 16584 12400 16590
rect 12348 16526 12400 16532
rect 12256 16516 12308 16522
rect 12256 16458 12308 16464
rect 11888 16448 11940 16454
rect 11888 16390 11940 16396
rect 12438 16416 12494 16425
rect 11900 16046 11928 16390
rect 12052 16348 12348 16368
rect 12438 16351 12494 16360
rect 12108 16346 12132 16348
rect 12188 16346 12212 16348
rect 12268 16346 12292 16348
rect 12130 16294 12132 16346
rect 12194 16294 12206 16346
rect 12268 16294 12270 16346
rect 12108 16292 12132 16294
rect 12188 16292 12212 16294
rect 12268 16292 12292 16294
rect 12052 16272 12348 16292
rect 11888 16040 11940 16046
rect 11888 15982 11940 15988
rect 11796 15904 11848 15910
rect 11796 15846 11848 15852
rect 12348 15904 12400 15910
rect 12348 15846 12400 15852
rect 11796 15632 11848 15638
rect 11796 15574 11848 15580
rect 11808 15065 11836 15574
rect 12360 15434 12388 15846
rect 12348 15428 12400 15434
rect 12348 15370 12400 15376
rect 11980 15360 12032 15366
rect 11980 15302 12032 15308
rect 11888 15156 11940 15162
rect 11888 15098 11940 15104
rect 11794 15056 11850 15065
rect 11794 14991 11850 15000
rect 11702 14920 11758 14929
rect 11702 14855 11758 14864
rect 11716 14074 11744 14855
rect 11900 14396 11928 15098
rect 11992 14958 12020 15302
rect 12052 15260 12348 15280
rect 12108 15258 12132 15260
rect 12188 15258 12212 15260
rect 12268 15258 12292 15260
rect 12130 15206 12132 15258
rect 12194 15206 12206 15258
rect 12268 15206 12270 15258
rect 12108 15204 12132 15206
rect 12188 15204 12212 15206
rect 12268 15204 12292 15206
rect 12052 15184 12348 15204
rect 12346 15056 12402 15065
rect 12346 14991 12402 15000
rect 11980 14952 12032 14958
rect 11980 14894 12032 14900
rect 11992 14793 12020 14894
rect 12360 14890 12388 14991
rect 12348 14884 12400 14890
rect 12348 14826 12400 14832
rect 11978 14784 12034 14793
rect 11978 14719 12034 14728
rect 11900 14368 12020 14396
rect 11704 14068 11756 14074
rect 11704 14010 11756 14016
rect 11796 14000 11848 14006
rect 11796 13942 11848 13948
rect 11992 13954 12020 14368
rect 12052 14172 12348 14192
rect 12108 14170 12132 14172
rect 12188 14170 12212 14172
rect 12268 14170 12292 14172
rect 12130 14118 12132 14170
rect 12194 14118 12206 14170
rect 12268 14118 12270 14170
rect 12108 14116 12132 14118
rect 12188 14116 12212 14118
rect 12268 14116 12292 14118
rect 12052 14096 12348 14116
rect 11808 12782 11836 13942
rect 11992 13938 12204 13954
rect 11992 13932 12216 13938
rect 11992 13926 12164 13932
rect 12164 13874 12216 13880
rect 11888 13864 11940 13870
rect 11888 13806 11940 13812
rect 11900 13161 11928 13806
rect 12070 13560 12126 13569
rect 12070 13495 12126 13504
rect 12084 13326 12112 13495
rect 12072 13320 12124 13326
rect 12072 13262 12124 13268
rect 12452 13190 12480 16351
rect 12530 15192 12586 15201
rect 12530 15127 12586 15136
rect 12544 14618 12572 15127
rect 12532 14612 12584 14618
rect 12532 14554 12584 14560
rect 12532 14476 12584 14482
rect 12532 14418 12584 14424
rect 12544 13530 12572 14418
rect 12532 13524 12584 13530
rect 12532 13466 12584 13472
rect 12440 13184 12492 13190
rect 11886 13152 11942 13161
rect 12440 13126 12492 13132
rect 11886 13087 11942 13096
rect 12052 13084 12348 13104
rect 12108 13082 12132 13084
rect 12188 13082 12212 13084
rect 12268 13082 12292 13084
rect 12130 13030 12132 13082
rect 12194 13030 12206 13082
rect 12268 13030 12270 13082
rect 12108 13028 12132 13030
rect 12188 13028 12212 13030
rect 12268 13028 12292 13030
rect 12052 13008 12348 13028
rect 11796 12776 11848 12782
rect 11796 12718 11848 12724
rect 12544 12730 12572 13466
rect 12636 12850 12664 23582
rect 12716 22024 12768 22030
rect 12716 21966 12768 21972
rect 12728 19990 12756 21966
rect 13452 21956 13504 21962
rect 13452 21898 13504 21904
rect 12992 21344 13044 21350
rect 12992 21286 13044 21292
rect 13084 21344 13136 21350
rect 13084 21286 13136 21292
rect 12900 20868 12952 20874
rect 12900 20810 12952 20816
rect 12912 19990 12940 20810
rect 13004 20097 13032 21286
rect 12990 20088 13046 20097
rect 12990 20023 13046 20032
rect 12716 19984 12768 19990
rect 12716 19926 12768 19932
rect 12900 19984 12952 19990
rect 12900 19926 12952 19932
rect 12716 19168 12768 19174
rect 12716 19110 12768 19116
rect 12728 18834 12756 19110
rect 12716 18828 12768 18834
rect 12716 18770 12768 18776
rect 12912 18630 12940 19926
rect 13096 19281 13124 21286
rect 13360 21140 13412 21146
rect 13360 21082 13412 21088
rect 13176 19984 13228 19990
rect 13176 19926 13228 19932
rect 13188 19514 13216 19926
rect 13176 19508 13228 19514
rect 13176 19450 13228 19456
rect 13082 19272 13138 19281
rect 13082 19207 13138 19216
rect 12992 19168 13044 19174
rect 12992 19110 13044 19116
rect 13084 19168 13136 19174
rect 13084 19110 13136 19116
rect 13004 18737 13032 19110
rect 12990 18728 13046 18737
rect 12990 18663 13046 18672
rect 12900 18624 12952 18630
rect 12820 18584 12900 18612
rect 12820 18222 12848 18584
rect 12900 18566 12952 18572
rect 12900 18352 12952 18358
rect 12952 18312 13032 18340
rect 12900 18294 12952 18300
rect 12808 18216 12860 18222
rect 12860 18176 12940 18204
rect 12808 18158 12860 18164
rect 12808 18080 12860 18086
rect 12808 18022 12860 18028
rect 12716 17604 12768 17610
rect 12716 17546 12768 17552
rect 12728 16998 12756 17546
rect 12716 16992 12768 16998
rect 12716 16934 12768 16940
rect 12714 16552 12770 16561
rect 12714 16487 12770 16496
rect 12728 16454 12756 16487
rect 12716 16448 12768 16454
rect 12716 16390 12768 16396
rect 12820 15994 12848 18022
rect 12912 17610 12940 18176
rect 12900 17604 12952 17610
rect 12900 17546 12952 17552
rect 12900 17332 12952 17338
rect 12900 17274 12952 17280
rect 12912 17241 12940 17274
rect 12898 17232 12954 17241
rect 12898 17167 12954 17176
rect 12900 16992 12952 16998
rect 12900 16934 12952 16940
rect 12912 16182 12940 16934
rect 13004 16658 13032 18312
rect 13096 17746 13124 19110
rect 13174 18048 13230 18057
rect 13174 17983 13230 17992
rect 13084 17740 13136 17746
rect 13084 17682 13136 17688
rect 12992 16652 13044 16658
rect 12992 16594 13044 16600
rect 12990 16280 13046 16289
rect 12990 16215 12992 16224
rect 13044 16215 13046 16224
rect 12992 16186 13044 16192
rect 12900 16176 12952 16182
rect 12900 16118 12952 16124
rect 12728 15966 12848 15994
rect 12898 16008 12954 16017
rect 12728 15910 12756 15966
rect 12898 15943 12954 15952
rect 12716 15904 12768 15910
rect 12716 15846 12768 15852
rect 12808 15904 12860 15910
rect 12808 15846 12860 15852
rect 12820 15745 12848 15846
rect 12806 15736 12862 15745
rect 12806 15671 12862 15680
rect 12808 15564 12860 15570
rect 12808 15506 12860 15512
rect 12716 15496 12768 15502
rect 12716 15438 12768 15444
rect 12728 15162 12756 15438
rect 12820 15337 12848 15506
rect 12806 15328 12862 15337
rect 12806 15263 12862 15272
rect 12716 15156 12768 15162
rect 12716 15098 12768 15104
rect 12808 15156 12860 15162
rect 12808 15098 12860 15104
rect 12820 14929 12848 15098
rect 12806 14920 12862 14929
rect 12806 14855 12862 14864
rect 12716 14408 12768 14414
rect 12716 14350 12768 14356
rect 12728 14074 12756 14350
rect 12808 14340 12860 14346
rect 12808 14282 12860 14288
rect 12716 14068 12768 14074
rect 12716 14010 12768 14016
rect 12716 13864 12768 13870
rect 12820 13852 12848 14282
rect 12912 14249 12940 15943
rect 12992 14952 13044 14958
rect 12992 14894 13044 14900
rect 12898 14240 12954 14249
rect 12898 14175 12954 14184
rect 12768 13824 12848 13852
rect 12716 13806 12768 13812
rect 12716 13728 12768 13734
rect 12716 13670 12768 13676
rect 12728 12986 12756 13670
rect 12716 12980 12768 12986
rect 12716 12922 12768 12928
rect 12624 12844 12676 12850
rect 12624 12786 12676 12792
rect 13004 12782 13032 14894
rect 13084 14544 13136 14550
rect 13084 14486 13136 14492
rect 13096 13734 13124 14486
rect 13188 14482 13216 17983
rect 13372 17513 13400 21082
rect 13358 17504 13414 17513
rect 13358 17439 13414 17448
rect 13268 17128 13320 17134
rect 13268 17070 13320 17076
rect 13280 15910 13308 17070
rect 13360 17060 13412 17066
rect 13360 17002 13412 17008
rect 13268 15904 13320 15910
rect 13268 15846 13320 15852
rect 13176 14476 13228 14482
rect 13176 14418 13228 14424
rect 13084 13728 13136 13734
rect 13084 13670 13136 13676
rect 13082 13560 13138 13569
rect 13082 13495 13138 13504
rect 12992 12776 13044 12782
rect 12544 12714 12664 12730
rect 12992 12718 13044 12724
rect 12348 12708 12400 12714
rect 12544 12708 12676 12714
rect 12544 12702 12624 12708
rect 12348 12650 12400 12656
rect 12624 12650 12676 12656
rect 12360 12442 12388 12650
rect 12532 12640 12584 12646
rect 12532 12582 12584 12588
rect 12348 12436 12400 12442
rect 12400 12396 12480 12424
rect 12348 12378 12400 12384
rect 12052 11996 12348 12016
rect 12108 11994 12132 11996
rect 12188 11994 12212 11996
rect 12268 11994 12292 11996
rect 12130 11942 12132 11994
rect 12194 11942 12206 11994
rect 12268 11942 12270 11994
rect 12108 11940 12132 11942
rect 12188 11940 12212 11942
rect 12268 11940 12292 11942
rect 12052 11920 12348 11940
rect 12452 11218 12480 12396
rect 11612 11212 11664 11218
rect 11612 11154 11664 11160
rect 12440 11212 12492 11218
rect 12440 11154 12492 11160
rect 12052 10908 12348 10928
rect 12108 10906 12132 10908
rect 12188 10906 12212 10908
rect 12268 10906 12292 10908
rect 12130 10854 12132 10906
rect 12194 10854 12206 10906
rect 12268 10854 12270 10906
rect 12108 10852 12132 10854
rect 12188 10852 12212 10854
rect 12268 10852 12292 10854
rect 12052 10832 12348 10852
rect 12440 10600 12492 10606
rect 12440 10542 12492 10548
rect 11518 10296 11574 10305
rect 11518 10231 11574 10240
rect 11980 10260 12032 10266
rect 11980 10202 12032 10208
rect 11992 9926 12020 10202
rect 12452 9926 12480 10542
rect 12544 10538 12572 12582
rect 13004 12170 13032 12718
rect 12992 12164 13044 12170
rect 12992 12106 13044 12112
rect 12624 11756 12676 11762
rect 12624 11698 12676 11704
rect 12636 11218 12664 11698
rect 12624 11212 12676 11218
rect 12624 11154 12676 11160
rect 12532 10532 12584 10538
rect 12532 10474 12584 10480
rect 12636 9926 12664 11154
rect 12990 10840 13046 10849
rect 12990 10775 13046 10784
rect 12716 10056 12768 10062
rect 12716 9998 12768 10004
rect 11980 9920 12032 9926
rect 11980 9862 12032 9868
rect 12440 9920 12492 9926
rect 12440 9862 12492 9868
rect 12624 9920 12676 9926
rect 12728 9874 12756 9998
rect 12676 9868 12756 9874
rect 12624 9862 12756 9868
rect 12052 9820 12348 9840
rect 12108 9818 12132 9820
rect 12188 9818 12212 9820
rect 12268 9818 12292 9820
rect 12130 9766 12132 9818
rect 12194 9766 12206 9818
rect 12268 9766 12270 9818
rect 12108 9764 12132 9766
rect 12188 9764 12212 9766
rect 12268 9764 12292 9766
rect 12052 9744 12348 9764
rect 11888 9580 11940 9586
rect 11888 9522 11940 9528
rect 11900 9489 11928 9522
rect 11886 9480 11942 9489
rect 11886 9415 11942 9424
rect 11428 9104 11480 9110
rect 11612 9104 11664 9110
rect 11480 9064 11560 9092
rect 11428 9046 11480 9052
rect 11256 8622 11468 8650
rect 11244 8424 11296 8430
rect 11164 8384 11244 8412
rect 11244 8366 11296 8372
rect 10968 8356 11020 8362
rect 10968 8298 11020 8304
rect 10968 8016 11020 8022
rect 10968 7958 11020 7964
rect 11058 7984 11114 7993
rect 10874 7032 10930 7041
rect 10874 6967 10930 6976
rect 10980 6934 11008 7958
rect 11058 7919 11114 7928
rect 10968 6928 11020 6934
rect 10968 6870 11020 6876
rect 10874 6488 10930 6497
rect 10874 6423 10876 6432
rect 10928 6423 10930 6432
rect 10876 6394 10928 6400
rect 10980 6322 11008 6870
rect 11072 6798 11100 7919
rect 11244 7404 11296 7410
rect 11244 7346 11296 7352
rect 11060 6792 11112 6798
rect 11060 6734 11112 6740
rect 11152 6792 11204 6798
rect 11152 6734 11204 6740
rect 11060 6656 11112 6662
rect 11060 6598 11112 6604
rect 10968 6316 11020 6322
rect 10968 6258 11020 6264
rect 11072 6254 11100 6598
rect 11060 6248 11112 6254
rect 11060 6190 11112 6196
rect 11072 5778 11100 6190
rect 11060 5772 11112 5778
rect 11060 5714 11112 5720
rect 11164 5642 11192 6734
rect 11256 6225 11284 7346
rect 11336 6656 11388 6662
rect 11336 6598 11388 6604
rect 11242 6216 11298 6225
rect 11242 6151 11298 6160
rect 11244 6112 11296 6118
rect 11244 6054 11296 6060
rect 11256 5710 11284 6054
rect 11244 5704 11296 5710
rect 11244 5646 11296 5652
rect 11152 5636 11204 5642
rect 11152 5578 11204 5584
rect 11164 5166 11192 5578
rect 11152 5160 11204 5166
rect 11152 5102 11204 5108
rect 11256 5098 11284 5646
rect 11244 5092 11296 5098
rect 11244 5034 11296 5040
rect 11256 4622 11284 5034
rect 11348 4758 11376 6598
rect 11336 4752 11388 4758
rect 11336 4694 11388 4700
rect 11244 4616 11296 4622
rect 11244 4558 11296 4564
rect 11440 4214 11468 8622
rect 11532 6254 11560 9064
rect 11612 9046 11664 9052
rect 11624 8673 11652 9046
rect 11610 8664 11666 8673
rect 11610 8599 11666 8608
rect 11704 8628 11756 8634
rect 11704 8570 11756 8576
rect 11796 8628 11848 8634
rect 11796 8570 11848 8576
rect 11716 7954 11744 8570
rect 11808 8022 11836 8570
rect 11796 8016 11848 8022
rect 11796 7958 11848 7964
rect 11704 7948 11756 7954
rect 11704 7890 11756 7896
rect 11900 7478 11928 9415
rect 12052 8732 12348 8752
rect 12108 8730 12132 8732
rect 12188 8730 12212 8732
rect 12268 8730 12292 8732
rect 12130 8678 12132 8730
rect 12194 8678 12206 8730
rect 12268 8678 12270 8730
rect 12108 8676 12132 8678
rect 12188 8676 12212 8678
rect 12268 8676 12292 8678
rect 12052 8656 12348 8676
rect 12452 8498 12480 9862
rect 12636 9846 12756 9862
rect 12624 9580 12676 9586
rect 12624 9522 12676 9528
rect 12440 8492 12492 8498
rect 12440 8434 12492 8440
rect 12532 8356 12584 8362
rect 12532 8298 12584 8304
rect 12348 8288 12400 8294
rect 12348 8230 12400 8236
rect 12360 7886 12388 8230
rect 12544 8090 12572 8298
rect 12532 8084 12584 8090
rect 12532 8026 12584 8032
rect 12348 7880 12400 7886
rect 12348 7822 12400 7828
rect 12636 7818 12664 9522
rect 12728 9110 12756 9846
rect 12808 9444 12860 9450
rect 12808 9386 12860 9392
rect 12716 9104 12768 9110
rect 12716 9046 12768 9052
rect 12820 8634 12848 9386
rect 12900 9376 12952 9382
rect 12900 9318 12952 9324
rect 12912 9178 12940 9318
rect 12900 9172 12952 9178
rect 12900 9114 12952 9120
rect 13004 9058 13032 10775
rect 12912 9030 13032 9058
rect 13096 9042 13124 13495
rect 13280 12102 13308 15846
rect 13268 12096 13320 12102
rect 13268 12038 13320 12044
rect 13372 9058 13400 17002
rect 13464 15314 13492 21898
rect 13544 19168 13596 19174
rect 13544 19110 13596 19116
rect 13556 18902 13584 19110
rect 13544 18896 13596 18902
rect 13544 18838 13596 18844
rect 13464 15286 13584 15314
rect 13556 15094 13584 15286
rect 13544 15088 13596 15094
rect 13544 15030 13596 15036
rect 13544 14884 13596 14890
rect 13544 14826 13596 14832
rect 13452 14816 13504 14822
rect 13452 14758 13504 14764
rect 13464 14346 13492 14758
rect 13452 14340 13504 14346
rect 13452 14282 13504 14288
rect 13556 14006 13584 14826
rect 13452 14000 13504 14006
rect 13452 13942 13504 13948
rect 13544 14000 13596 14006
rect 13544 13942 13596 13948
rect 13464 12442 13492 13942
rect 13544 13320 13596 13326
rect 13544 13262 13596 13268
rect 13556 12782 13584 13262
rect 13544 12776 13596 12782
rect 13544 12718 13596 12724
rect 13452 12436 13504 12442
rect 13452 12378 13504 12384
rect 13648 12374 13676 23582
rect 13740 19446 13768 23600
rect 14384 23582 14596 23600
rect 14188 21888 14240 21894
rect 14188 21830 14240 21836
rect 14200 21554 14228 21830
rect 14188 21548 14240 21554
rect 14188 21490 14240 21496
rect 14464 21412 14516 21418
rect 14464 21354 14516 21360
rect 13820 21344 13872 21350
rect 13820 21286 13872 21292
rect 14004 21344 14056 21350
rect 14004 21286 14056 21292
rect 13832 20641 13860 21286
rect 13818 20632 13874 20641
rect 13818 20567 13874 20576
rect 14016 20505 14044 21286
rect 14476 21146 14504 21354
rect 14464 21140 14516 21146
rect 14464 21082 14516 21088
rect 14096 21004 14148 21010
rect 14096 20946 14148 20952
rect 14108 20602 14136 20946
rect 14372 20936 14424 20942
rect 14372 20878 14424 20884
rect 14384 20806 14412 20878
rect 14372 20800 14424 20806
rect 14372 20742 14424 20748
rect 14096 20596 14148 20602
rect 14096 20538 14148 20544
rect 14002 20496 14058 20505
rect 14384 20466 14412 20742
rect 14002 20431 14058 20440
rect 14372 20460 14424 20466
rect 14372 20402 14424 20408
rect 14476 20398 14504 21082
rect 13912 20392 13964 20398
rect 13912 20334 13964 20340
rect 14464 20392 14516 20398
rect 14464 20334 14516 20340
rect 13924 19938 13952 20334
rect 14004 20324 14056 20330
rect 14004 20266 14056 20272
rect 14016 20058 14044 20266
rect 14004 20052 14056 20058
rect 14004 19994 14056 20000
rect 13924 19910 14228 19938
rect 14004 19848 14056 19854
rect 14004 19790 14056 19796
rect 13728 19440 13780 19446
rect 13728 19382 13780 19388
rect 14016 18970 14044 19790
rect 14200 19514 14228 19910
rect 14464 19712 14516 19718
rect 14278 19680 14334 19689
rect 14464 19654 14516 19660
rect 14278 19615 14334 19624
rect 14096 19508 14148 19514
rect 14096 19450 14148 19456
rect 14188 19508 14240 19514
rect 14188 19450 14240 19456
rect 14004 18964 14056 18970
rect 14004 18906 14056 18912
rect 13820 17740 13872 17746
rect 13820 17682 13872 17688
rect 13728 17536 13780 17542
rect 13728 17478 13780 17484
rect 13740 16998 13768 17478
rect 13832 17270 13860 17682
rect 13820 17264 13872 17270
rect 13820 17206 13872 17212
rect 14004 17060 14056 17066
rect 14004 17002 14056 17008
rect 13728 16992 13780 16998
rect 13780 16952 13860 16980
rect 13728 16934 13780 16940
rect 13728 16448 13780 16454
rect 13728 16390 13780 16396
rect 13740 15502 13768 16390
rect 13832 16114 13860 16952
rect 14016 16522 14044 17002
rect 14004 16516 14056 16522
rect 14004 16458 14056 16464
rect 13820 16108 13872 16114
rect 13820 16050 13872 16056
rect 13912 15904 13964 15910
rect 13912 15846 13964 15852
rect 13924 15638 13952 15846
rect 13912 15632 13964 15638
rect 13912 15574 13964 15580
rect 14108 15570 14136 19450
rect 14292 19394 14320 19615
rect 14200 19366 14320 19394
rect 14200 18034 14228 19366
rect 14278 19272 14334 19281
rect 14278 19207 14334 19216
rect 14292 18902 14320 19207
rect 14372 18964 14424 18970
rect 14372 18906 14424 18912
rect 14280 18896 14332 18902
rect 14280 18838 14332 18844
rect 14384 18222 14412 18906
rect 14372 18216 14424 18222
rect 14372 18158 14424 18164
rect 14200 18006 14320 18034
rect 14188 17876 14240 17882
rect 14188 17818 14240 17824
rect 14200 17785 14228 17818
rect 14186 17776 14242 17785
rect 14186 17711 14242 17720
rect 14188 16720 14240 16726
rect 14188 16662 14240 16668
rect 14200 16522 14228 16662
rect 14188 16516 14240 16522
rect 14188 16458 14240 16464
rect 13820 15564 13872 15570
rect 13820 15506 13872 15512
rect 14096 15564 14148 15570
rect 14096 15506 14148 15512
rect 13728 15496 13780 15502
rect 13728 15438 13780 15444
rect 13728 15088 13780 15094
rect 13728 15030 13780 15036
rect 13740 13802 13768 15030
rect 13832 14822 13860 15506
rect 13912 15496 13964 15502
rect 14292 15450 14320 18006
rect 14384 17882 14412 18158
rect 14372 17876 14424 17882
rect 14372 17818 14424 17824
rect 14476 16096 14504 19654
rect 14568 19553 14596 23582
rect 14648 21480 14700 21486
rect 14648 21422 14700 21428
rect 14660 21146 14688 21422
rect 14648 21140 14700 21146
rect 14648 21082 14700 21088
rect 14924 20392 14976 20398
rect 14924 20334 14976 20340
rect 14936 20074 14964 20334
rect 14660 20046 14964 20074
rect 14660 19990 14688 20046
rect 14648 19984 14700 19990
rect 14648 19926 14700 19932
rect 15028 19922 15056 23600
rect 15384 22908 15436 22914
rect 15384 22850 15436 22856
rect 15108 21480 15160 21486
rect 15108 21422 15160 21428
rect 15120 20602 15148 21422
rect 15200 21140 15252 21146
rect 15200 21082 15252 21088
rect 15108 20596 15160 20602
rect 15108 20538 15160 20544
rect 15016 19916 15068 19922
rect 15016 19858 15068 19864
rect 14554 19544 14610 19553
rect 15212 19496 15240 21082
rect 14554 19479 14610 19488
rect 15028 19468 15332 19496
rect 14556 19440 14608 19446
rect 14556 19382 14608 19388
rect 13912 15438 13964 15444
rect 13924 14890 13952 15438
rect 14004 15428 14056 15434
rect 14004 15370 14056 15376
rect 14108 15422 14320 15450
rect 14384 16068 14504 16096
rect 14016 14958 14044 15370
rect 14004 14952 14056 14958
rect 14004 14894 14056 14900
rect 13912 14884 13964 14890
rect 13912 14826 13964 14832
rect 13820 14816 13872 14822
rect 13820 14758 13872 14764
rect 13832 13802 13860 14758
rect 14108 14634 14136 15422
rect 14188 15360 14240 15366
rect 14188 15302 14240 15308
rect 14278 15328 14334 15337
rect 14200 14958 14228 15302
rect 14278 15263 14334 15272
rect 14188 14952 14240 14958
rect 14188 14894 14240 14900
rect 14188 14816 14240 14822
rect 14188 14758 14240 14764
rect 13924 14606 14136 14634
rect 14200 14618 14228 14758
rect 14188 14612 14240 14618
rect 13728 13796 13780 13802
rect 13728 13738 13780 13744
rect 13820 13796 13872 13802
rect 13820 13738 13872 13744
rect 13924 13682 13952 14606
rect 14188 14554 14240 14560
rect 14004 14544 14056 14550
rect 14004 14486 14056 14492
rect 14186 14512 14242 14521
rect 13740 13654 13952 13682
rect 13636 12368 13688 12374
rect 13636 12310 13688 12316
rect 13544 11008 13596 11014
rect 13544 10950 13596 10956
rect 13556 10130 13584 10950
rect 13544 10124 13596 10130
rect 13544 10066 13596 10072
rect 13544 9512 13596 9518
rect 13544 9454 13596 9460
rect 13636 9512 13688 9518
rect 13636 9454 13688 9460
rect 13084 9036 13136 9042
rect 12808 8628 12860 8634
rect 12808 8570 12860 8576
rect 12164 7812 12216 7818
rect 11992 7772 12164 7800
rect 11992 7546 12020 7772
rect 12164 7754 12216 7760
rect 12624 7812 12676 7818
rect 12624 7754 12676 7760
rect 12440 7744 12492 7750
rect 12912 7698 12940 9030
rect 13084 8978 13136 8984
rect 13280 9030 13400 9058
rect 13176 8968 13228 8974
rect 13176 8910 13228 8916
rect 13188 8634 13216 8910
rect 13176 8628 13228 8634
rect 13176 8570 13228 8576
rect 12992 8016 13044 8022
rect 12992 7958 13044 7964
rect 13004 7857 13032 7958
rect 12990 7848 13046 7857
rect 12990 7783 13046 7792
rect 12440 7686 12492 7692
rect 12052 7644 12348 7664
rect 12108 7642 12132 7644
rect 12188 7642 12212 7644
rect 12268 7642 12292 7644
rect 12130 7590 12132 7642
rect 12194 7590 12206 7642
rect 12268 7590 12270 7642
rect 12108 7588 12132 7590
rect 12188 7588 12212 7590
rect 12268 7588 12292 7590
rect 12052 7568 12348 7588
rect 12452 7585 12480 7686
rect 12544 7670 12940 7698
rect 13176 7744 13228 7750
rect 13176 7686 13228 7692
rect 12438 7576 12494 7585
rect 11980 7540 12032 7546
rect 12438 7511 12494 7520
rect 11980 7482 12032 7488
rect 11888 7472 11940 7478
rect 11888 7414 11940 7420
rect 11796 7336 11848 7342
rect 11796 7278 11848 7284
rect 11612 6860 11664 6866
rect 11612 6802 11664 6808
rect 11520 6248 11572 6254
rect 11520 6190 11572 6196
rect 11518 6080 11574 6089
rect 11518 6015 11574 6024
rect 11532 4826 11560 6015
rect 11624 5778 11652 6802
rect 11702 6352 11758 6361
rect 11702 6287 11758 6296
rect 11612 5772 11664 5778
rect 11612 5714 11664 5720
rect 11624 5370 11652 5714
rect 11612 5364 11664 5370
rect 11612 5306 11664 5312
rect 11520 4820 11572 4826
rect 11520 4762 11572 4768
rect 11610 4584 11666 4593
rect 11610 4519 11666 4528
rect 11428 4208 11480 4214
rect 11428 4150 11480 4156
rect 10784 4072 10836 4078
rect 10784 4014 10836 4020
rect 11624 4010 11652 4519
rect 11716 4078 11744 6287
rect 11704 4072 11756 4078
rect 11704 4014 11756 4020
rect 11808 4026 11836 7278
rect 12256 7268 12308 7274
rect 12256 7210 12308 7216
rect 12268 6730 12296 7210
rect 12440 7200 12492 7206
rect 12440 7142 12492 7148
rect 12256 6724 12308 6730
rect 12256 6666 12308 6672
rect 12052 6556 12348 6576
rect 12108 6554 12132 6556
rect 12188 6554 12212 6556
rect 12268 6554 12292 6556
rect 12130 6502 12132 6554
rect 12194 6502 12206 6554
rect 12268 6502 12270 6554
rect 12108 6500 12132 6502
rect 12188 6500 12212 6502
rect 12268 6500 12292 6502
rect 12052 6480 12348 6500
rect 12348 6316 12400 6322
rect 12348 6258 12400 6264
rect 12256 6248 12308 6254
rect 12256 6190 12308 6196
rect 12268 5681 12296 6190
rect 12360 5914 12388 6258
rect 12348 5908 12400 5914
rect 12348 5850 12400 5856
rect 12254 5672 12310 5681
rect 12254 5607 12310 5616
rect 11980 5568 12032 5574
rect 11980 5510 12032 5516
rect 11612 4004 11664 4010
rect 11808 3998 11928 4026
rect 11612 3946 11664 3952
rect 10324 3732 10376 3738
rect 10324 3674 10376 3680
rect 10336 3641 10364 3674
rect 10322 3632 10378 3641
rect 10322 3567 10378 3576
rect 11624 3398 11652 3946
rect 11612 3392 11664 3398
rect 11612 3334 11664 3340
rect 11900 2990 11928 3998
rect 11992 3618 12020 5510
rect 12052 5468 12348 5488
rect 12108 5466 12132 5468
rect 12188 5466 12212 5468
rect 12268 5466 12292 5468
rect 12130 5414 12132 5466
rect 12194 5414 12206 5466
rect 12268 5414 12270 5466
rect 12108 5412 12132 5414
rect 12188 5412 12212 5414
rect 12268 5412 12292 5414
rect 12052 5392 12348 5412
rect 12256 5160 12308 5166
rect 12254 5128 12256 5137
rect 12308 5128 12310 5137
rect 12254 5063 12310 5072
rect 12348 5024 12400 5030
rect 12348 4966 12400 4972
rect 12360 4622 12388 4966
rect 12348 4616 12400 4622
rect 12348 4558 12400 4564
rect 12052 4380 12348 4400
rect 12108 4378 12132 4380
rect 12188 4378 12212 4380
rect 12268 4378 12292 4380
rect 12130 4326 12132 4378
rect 12194 4326 12206 4378
rect 12268 4326 12270 4378
rect 12108 4324 12132 4326
rect 12188 4324 12212 4326
rect 12268 4324 12292 4326
rect 12052 4304 12348 4324
rect 11992 3590 12112 3618
rect 12452 3602 12480 7142
rect 12544 5778 12572 7670
rect 12990 7440 13046 7449
rect 12990 7375 13046 7384
rect 12808 7200 12860 7206
rect 12808 7142 12860 7148
rect 12716 6928 12768 6934
rect 12716 6870 12768 6876
rect 12624 6792 12676 6798
rect 12624 6734 12676 6740
rect 12532 5772 12584 5778
rect 12532 5714 12584 5720
rect 12636 5642 12664 6734
rect 12624 5636 12676 5642
rect 12624 5578 12676 5584
rect 12532 5568 12584 5574
rect 12532 5510 12584 5516
rect 12544 5030 12572 5510
rect 12532 5024 12584 5030
rect 12532 4966 12584 4972
rect 12636 4758 12664 5578
rect 12728 5166 12756 6870
rect 12716 5160 12768 5166
rect 12716 5102 12768 5108
rect 12728 4826 12756 5102
rect 12820 4826 12848 7142
rect 12900 6928 12952 6934
rect 12900 6870 12952 6876
rect 12716 4820 12768 4826
rect 12716 4762 12768 4768
rect 12808 4820 12860 4826
rect 12808 4762 12860 4768
rect 12624 4752 12676 4758
rect 12624 4694 12676 4700
rect 12808 4004 12860 4010
rect 12808 3946 12860 3952
rect 12820 3738 12848 3946
rect 12808 3732 12860 3738
rect 12808 3674 12860 3680
rect 12084 3534 12112 3590
rect 12440 3596 12492 3602
rect 12440 3538 12492 3544
rect 12072 3528 12124 3534
rect 12912 3482 12940 6870
rect 13004 4978 13032 7375
rect 13084 6792 13136 6798
rect 13084 6734 13136 6740
rect 13096 5098 13124 6734
rect 13084 5092 13136 5098
rect 13084 5034 13136 5040
rect 13004 4950 13124 4978
rect 12072 3470 12124 3476
rect 12820 3466 12940 3482
rect 12808 3460 12940 3466
rect 12860 3454 12940 3460
rect 12992 3460 13044 3466
rect 12808 3402 12860 3408
rect 12992 3402 13044 3408
rect 11980 3392 12032 3398
rect 11980 3334 12032 3340
rect 11888 2984 11940 2990
rect 11888 2926 11940 2932
rect 9864 2304 9916 2310
rect 9864 2246 9916 2252
rect 11992 2088 12020 3334
rect 12052 3292 12348 3312
rect 12108 3290 12132 3292
rect 12188 3290 12212 3292
rect 12268 3290 12292 3292
rect 12130 3238 12132 3290
rect 12194 3238 12206 3290
rect 12268 3238 12270 3290
rect 12108 3236 12132 3238
rect 12188 3236 12212 3238
rect 12268 3236 12292 3238
rect 12052 3216 12348 3236
rect 13004 2854 13032 3402
rect 13096 3194 13124 4950
rect 13188 4554 13216 7686
rect 13280 7154 13308 9030
rect 13452 8832 13504 8838
rect 13450 8800 13452 8809
rect 13504 8800 13506 8809
rect 13450 8735 13506 8744
rect 13452 8560 13504 8566
rect 13452 8502 13504 8508
rect 13464 8294 13492 8502
rect 13452 8288 13504 8294
rect 13358 8256 13414 8265
rect 13452 8230 13504 8236
rect 13358 8191 13414 8200
rect 13372 8090 13400 8191
rect 13360 8084 13412 8090
rect 13360 8026 13412 8032
rect 13464 7954 13492 8230
rect 13452 7948 13504 7954
rect 13452 7890 13504 7896
rect 13556 7886 13584 9454
rect 13648 9042 13676 9454
rect 13740 9178 13768 13654
rect 13820 12300 13872 12306
rect 13820 12242 13872 12248
rect 13832 11898 13860 12242
rect 13820 11892 13872 11898
rect 13820 11834 13872 11840
rect 14016 11694 14044 14486
rect 14186 14447 14242 14456
rect 14096 14408 14148 14414
rect 14096 14350 14148 14356
rect 14108 13938 14136 14350
rect 14200 14278 14228 14447
rect 14188 14272 14240 14278
rect 14188 14214 14240 14220
rect 14096 13932 14148 13938
rect 14096 13874 14148 13880
rect 14188 13864 14240 13870
rect 14188 13806 14240 13812
rect 14200 13705 14228 13806
rect 14292 13734 14320 15263
rect 14280 13728 14332 13734
rect 14186 13696 14242 13705
rect 14280 13670 14332 13676
rect 14186 13631 14242 13640
rect 14096 13524 14148 13530
rect 14096 13466 14148 13472
rect 14004 11688 14056 11694
rect 14004 11630 14056 11636
rect 13820 11552 13872 11558
rect 13820 11494 13872 11500
rect 13832 10538 13860 11494
rect 13912 11008 13964 11014
rect 13910 10976 13912 10985
rect 13964 10976 13966 10985
rect 13910 10911 13966 10920
rect 14108 10826 14136 13466
rect 14278 12336 14334 12345
rect 14278 12271 14334 12280
rect 14292 11218 14320 12271
rect 14384 11937 14412 16068
rect 14568 15994 14596 19382
rect 14832 19168 14884 19174
rect 14832 19110 14884 19116
rect 14844 17746 14872 19110
rect 14924 18284 14976 18290
rect 14924 18226 14976 18232
rect 14936 17814 14964 18226
rect 14924 17808 14976 17814
rect 14924 17750 14976 17756
rect 14648 17740 14700 17746
rect 14648 17682 14700 17688
rect 14832 17740 14884 17746
rect 14832 17682 14884 17688
rect 14476 15966 14596 15994
rect 14370 11928 14426 11937
rect 14370 11863 14426 11872
rect 14280 11212 14332 11218
rect 14280 11154 14332 11160
rect 14188 11008 14240 11014
rect 14188 10950 14240 10956
rect 13924 10798 14136 10826
rect 13820 10532 13872 10538
rect 13820 10474 13872 10480
rect 13820 9376 13872 9382
rect 13820 9318 13872 9324
rect 13728 9172 13780 9178
rect 13728 9114 13780 9120
rect 13636 9036 13688 9042
rect 13636 8978 13688 8984
rect 13648 8498 13676 8978
rect 13636 8492 13688 8498
rect 13636 8434 13688 8440
rect 13726 8256 13782 8265
rect 13726 8191 13782 8200
rect 13544 7880 13596 7886
rect 13544 7822 13596 7828
rect 13358 7440 13414 7449
rect 13358 7375 13414 7384
rect 13372 7342 13400 7375
rect 13360 7336 13412 7342
rect 13360 7278 13412 7284
rect 13280 7126 13492 7154
rect 13358 7032 13414 7041
rect 13268 6996 13320 7002
rect 13358 6967 13414 6976
rect 13268 6938 13320 6944
rect 13176 4548 13228 4554
rect 13176 4490 13228 4496
rect 13280 4264 13308 6938
rect 13372 6662 13400 6967
rect 13360 6656 13412 6662
rect 13360 6598 13412 6604
rect 13360 6180 13412 6186
rect 13360 6122 13412 6128
rect 13372 4826 13400 6122
rect 13360 4820 13412 4826
rect 13360 4762 13412 4768
rect 13464 4706 13492 7126
rect 13556 6866 13584 7822
rect 13544 6860 13596 6866
rect 13544 6802 13596 6808
rect 13372 4678 13492 4706
rect 13372 4486 13400 4678
rect 13556 4622 13584 6802
rect 13634 6624 13690 6633
rect 13634 6559 13690 6568
rect 13648 5914 13676 6559
rect 13740 6304 13768 8191
rect 13832 7954 13860 9318
rect 13820 7948 13872 7954
rect 13820 7890 13872 7896
rect 13820 7200 13872 7206
rect 13820 7142 13872 7148
rect 13832 6934 13860 7142
rect 13820 6928 13872 6934
rect 13820 6870 13872 6876
rect 13924 6769 13952 10798
rect 14096 10464 14148 10470
rect 14200 10441 14228 10950
rect 14292 10742 14320 11154
rect 14372 11008 14424 11014
rect 14372 10950 14424 10956
rect 14280 10736 14332 10742
rect 14280 10678 14332 10684
rect 14384 10674 14412 10950
rect 14372 10668 14424 10674
rect 14372 10610 14424 10616
rect 14096 10406 14148 10412
rect 14186 10432 14242 10441
rect 14108 9654 14136 10406
rect 14186 10367 14242 10376
rect 14280 10056 14332 10062
rect 14280 9998 14332 10004
rect 14370 10024 14426 10033
rect 14186 9888 14242 9897
rect 14186 9823 14242 9832
rect 14096 9648 14148 9654
rect 14096 9590 14148 9596
rect 14004 9580 14056 9586
rect 14004 9522 14056 9528
rect 14016 9110 14044 9522
rect 14004 9104 14056 9110
rect 14004 9046 14056 9052
rect 14004 7812 14056 7818
rect 14004 7754 14056 7760
rect 14016 6798 14044 7754
rect 14004 6792 14056 6798
rect 13910 6760 13966 6769
rect 14004 6734 14056 6740
rect 13910 6695 13966 6704
rect 14096 6656 14148 6662
rect 14096 6598 14148 6604
rect 13740 6276 13860 6304
rect 13832 6186 13860 6276
rect 13728 6180 13780 6186
rect 13728 6122 13780 6128
rect 13820 6180 13872 6186
rect 13820 6122 13872 6128
rect 13740 5914 13768 6122
rect 13636 5908 13688 5914
rect 13636 5850 13688 5856
rect 13728 5908 13780 5914
rect 13728 5850 13780 5856
rect 13728 5772 13780 5778
rect 13728 5714 13780 5720
rect 13740 5302 13768 5714
rect 14108 5642 14136 6598
rect 14200 5817 14228 9823
rect 14292 8106 14320 9998
rect 14370 9959 14426 9968
rect 14384 8922 14412 9959
rect 14476 9110 14504 15966
rect 14556 15360 14608 15366
rect 14556 15302 14608 15308
rect 14568 13938 14596 15302
rect 14556 13932 14608 13938
rect 14556 13874 14608 13880
rect 14660 13530 14688 17682
rect 15028 17270 15056 19468
rect 15304 19417 15332 19468
rect 15290 19408 15346 19417
rect 15200 19372 15252 19378
rect 15290 19343 15346 19352
rect 15200 19314 15252 19320
rect 15108 18828 15160 18834
rect 15108 18770 15160 18776
rect 15120 18601 15148 18770
rect 15106 18592 15162 18601
rect 15106 18527 15162 18536
rect 15212 18290 15240 19314
rect 15292 19168 15344 19174
rect 15292 19110 15344 19116
rect 15200 18284 15252 18290
rect 15200 18226 15252 18232
rect 15304 17814 15332 19110
rect 15396 17882 15424 22850
rect 15476 21344 15528 21350
rect 15476 21286 15528 21292
rect 15488 21146 15516 21286
rect 15476 21140 15528 21146
rect 15476 21082 15528 21088
rect 15568 21072 15620 21078
rect 15568 21014 15620 21020
rect 15476 20800 15528 20806
rect 15476 20742 15528 20748
rect 15384 17876 15436 17882
rect 15384 17818 15436 17824
rect 15200 17808 15252 17814
rect 15200 17750 15252 17756
rect 15292 17808 15344 17814
rect 15292 17750 15344 17756
rect 15108 17672 15160 17678
rect 15108 17614 15160 17620
rect 15016 17264 15068 17270
rect 14922 17232 14978 17241
rect 14832 17196 14884 17202
rect 15016 17206 15068 17212
rect 14922 17167 14978 17176
rect 14832 17138 14884 17144
rect 14844 16658 14872 17138
rect 14936 16794 14964 17167
rect 15120 16998 15148 17614
rect 15108 16992 15160 16998
rect 15108 16934 15160 16940
rect 14924 16788 14976 16794
rect 14924 16730 14976 16736
rect 15120 16658 15148 16934
rect 14832 16652 14884 16658
rect 14832 16594 14884 16600
rect 15108 16652 15160 16658
rect 15108 16594 15160 16600
rect 14740 16584 14792 16590
rect 14740 16526 14792 16532
rect 14752 15881 14780 16526
rect 15120 16114 15148 16594
rect 15212 16250 15240 17750
rect 15304 16998 15332 17750
rect 15292 16992 15344 16998
rect 15292 16934 15344 16940
rect 15488 16810 15516 20742
rect 15580 20262 15608 21014
rect 15568 20256 15620 20262
rect 15568 20198 15620 20204
rect 15580 19990 15608 20198
rect 15568 19984 15620 19990
rect 15568 19926 15620 19932
rect 15672 19446 15700 23600
rect 16960 22030 16988 23600
rect 16948 22024 17000 22030
rect 16948 21966 17000 21972
rect 17604 21690 17632 23600
rect 17684 22636 17736 22642
rect 17684 22578 17736 22584
rect 17592 21684 17644 21690
rect 17592 21626 17644 21632
rect 16212 21548 16264 21554
rect 16212 21490 16264 21496
rect 16776 21542 16988 21570
rect 15750 21244 16046 21264
rect 15806 21242 15830 21244
rect 15886 21242 15910 21244
rect 15966 21242 15990 21244
rect 15828 21190 15830 21242
rect 15892 21190 15904 21242
rect 15966 21190 15968 21242
rect 15806 21188 15830 21190
rect 15886 21188 15910 21190
rect 15966 21188 15990 21190
rect 15750 21168 16046 21188
rect 16120 20392 16172 20398
rect 16120 20334 16172 20340
rect 15750 20156 16046 20176
rect 15806 20154 15830 20156
rect 15886 20154 15910 20156
rect 15966 20154 15990 20156
rect 15828 20102 15830 20154
rect 15892 20102 15904 20154
rect 15966 20102 15968 20154
rect 15806 20100 15830 20102
rect 15886 20100 15910 20102
rect 15966 20100 15990 20102
rect 15750 20080 16046 20100
rect 16028 19916 16080 19922
rect 16028 19858 16080 19864
rect 16040 19689 16068 19858
rect 16132 19854 16160 20334
rect 16120 19848 16172 19854
rect 16120 19790 16172 19796
rect 16026 19680 16082 19689
rect 16026 19615 16082 19624
rect 15660 19440 15712 19446
rect 15660 19382 15712 19388
rect 16132 19258 16160 19790
rect 16224 19786 16252 21490
rect 16776 21486 16804 21542
rect 16764 21480 16816 21486
rect 16764 21422 16816 21428
rect 16856 21480 16908 21486
rect 16856 21422 16908 21428
rect 16488 21344 16540 21350
rect 16488 21286 16540 21292
rect 16500 20806 16528 21286
rect 16488 20800 16540 20806
rect 16488 20742 16540 20748
rect 16580 20800 16632 20806
rect 16580 20742 16632 20748
rect 16592 20330 16620 20742
rect 16580 20324 16632 20330
rect 16580 20266 16632 20272
rect 16212 19780 16264 19786
rect 16212 19722 16264 19728
rect 16224 19378 16252 19722
rect 16592 19514 16620 20266
rect 16764 20256 16816 20262
rect 16764 20198 16816 20204
rect 16776 19990 16804 20198
rect 16764 19984 16816 19990
rect 16764 19926 16816 19932
rect 16762 19544 16818 19553
rect 16580 19508 16632 19514
rect 16762 19479 16818 19488
rect 16580 19450 16632 19456
rect 16212 19372 16264 19378
rect 16264 19332 16436 19360
rect 16212 19314 16264 19320
rect 16132 19230 16344 19258
rect 15568 19168 15620 19174
rect 15568 19110 15620 19116
rect 16120 19168 16172 19174
rect 16120 19110 16172 19116
rect 16212 19168 16264 19174
rect 16212 19110 16264 19116
rect 15580 18902 15608 19110
rect 15750 19068 16046 19088
rect 15806 19066 15830 19068
rect 15886 19066 15910 19068
rect 15966 19066 15990 19068
rect 15828 19014 15830 19066
rect 15892 19014 15904 19066
rect 15966 19014 15968 19066
rect 15806 19012 15830 19014
rect 15886 19012 15910 19014
rect 15966 19012 15990 19014
rect 15750 18992 16046 19012
rect 16132 18970 16160 19110
rect 16120 18964 16172 18970
rect 16120 18906 16172 18912
rect 15568 18896 15620 18902
rect 15568 18838 15620 18844
rect 16026 18864 16082 18873
rect 15580 18426 15608 18838
rect 16026 18799 16082 18808
rect 15752 18760 15804 18766
rect 15750 18728 15752 18737
rect 15804 18728 15806 18737
rect 15750 18663 15806 18672
rect 15568 18420 15620 18426
rect 15568 18362 15620 18368
rect 16040 18290 16068 18799
rect 16028 18284 16080 18290
rect 16028 18226 16080 18232
rect 15568 18148 15620 18154
rect 15568 18090 15620 18096
rect 15580 18034 15608 18090
rect 15580 18006 15700 18034
rect 15488 16782 15608 16810
rect 15200 16244 15252 16250
rect 15200 16186 15252 16192
rect 15108 16108 15160 16114
rect 15108 16050 15160 16056
rect 14924 16040 14976 16046
rect 14924 15982 14976 15988
rect 14738 15872 14794 15881
rect 14738 15807 14794 15816
rect 14936 15706 14964 15982
rect 15106 15736 15162 15745
rect 14924 15700 14976 15706
rect 15212 15706 15240 16186
rect 15384 15972 15436 15978
rect 15384 15914 15436 15920
rect 15106 15671 15162 15680
rect 15200 15700 15252 15706
rect 14924 15642 14976 15648
rect 14924 15564 14976 15570
rect 14924 15506 14976 15512
rect 14830 15192 14886 15201
rect 14830 15127 14886 15136
rect 14740 14816 14792 14822
rect 14740 14758 14792 14764
rect 14752 14464 14780 14758
rect 14844 14550 14872 15127
rect 14832 14544 14884 14550
rect 14832 14486 14884 14492
rect 14743 14436 14780 14464
rect 14743 14328 14771 14436
rect 14832 14340 14884 14346
rect 14743 14300 14832 14328
rect 14832 14282 14884 14288
rect 14936 13682 14964 15506
rect 15016 14476 15068 14482
rect 15016 14418 15068 14424
rect 15028 14074 15056 14418
rect 15120 14346 15148 15671
rect 15200 15642 15252 15648
rect 15200 15428 15252 15434
rect 15200 15370 15252 15376
rect 15212 15201 15240 15370
rect 15198 15192 15254 15201
rect 15198 15127 15254 15136
rect 15396 15094 15424 15914
rect 15384 15088 15436 15094
rect 15384 15030 15436 15036
rect 15200 15020 15252 15026
rect 15200 14962 15252 14968
rect 15108 14340 15160 14346
rect 15108 14282 15160 14288
rect 15016 14068 15068 14074
rect 15016 14010 15068 14016
rect 15120 13938 15148 14282
rect 15108 13932 15160 13938
rect 15108 13874 15160 13880
rect 14936 13654 15056 13682
rect 14648 13524 14700 13530
rect 14648 13466 14700 13472
rect 14832 13524 14884 13530
rect 14832 13466 14884 13472
rect 14556 13252 14608 13258
rect 14556 13194 14608 13200
rect 14568 12918 14596 13194
rect 14556 12912 14608 12918
rect 14556 12854 14608 12860
rect 14556 12776 14608 12782
rect 14556 12718 14608 12724
rect 14568 11694 14596 12718
rect 14844 12617 14872 13466
rect 14924 13252 14976 13258
rect 14924 13194 14976 13200
rect 14936 13161 14964 13194
rect 14922 13152 14978 13161
rect 14922 13087 14978 13096
rect 14936 12782 14964 13087
rect 14924 12776 14976 12782
rect 14924 12718 14976 12724
rect 14830 12608 14886 12617
rect 14830 12543 14886 12552
rect 14648 12096 14700 12102
rect 14646 12064 14648 12073
rect 14700 12064 14702 12073
rect 14646 11999 14702 12008
rect 14556 11688 14608 11694
rect 14660 11676 14688 11999
rect 14740 11688 14792 11694
rect 14660 11648 14740 11676
rect 14556 11630 14608 11636
rect 14740 11630 14792 11636
rect 14556 11552 14608 11558
rect 14556 11494 14608 11500
rect 14568 10130 14596 11494
rect 14648 11144 14700 11150
rect 14648 11086 14700 11092
rect 14830 11112 14886 11121
rect 14660 10305 14688 11086
rect 15028 11082 15056 13654
rect 14830 11047 14886 11056
rect 15016 11076 15068 11082
rect 14740 10668 14792 10674
rect 14740 10610 14792 10616
rect 14646 10296 14702 10305
rect 14646 10231 14702 10240
rect 14556 10124 14608 10130
rect 14556 10066 14608 10072
rect 14648 10056 14700 10062
rect 14648 9998 14700 10004
rect 14556 9512 14608 9518
rect 14660 9500 14688 9998
rect 14752 9518 14780 10610
rect 14608 9472 14688 9500
rect 14740 9512 14792 9518
rect 14556 9454 14608 9460
rect 14740 9454 14792 9460
rect 14646 9208 14702 9217
rect 14752 9178 14780 9454
rect 14646 9143 14702 9152
rect 14740 9172 14792 9178
rect 14464 9104 14516 9110
rect 14464 9046 14516 9052
rect 14660 9042 14688 9143
rect 14740 9114 14792 9120
rect 14648 9036 14700 9042
rect 14648 8978 14700 8984
rect 14384 8894 14596 8922
rect 14568 8786 14596 8894
rect 14568 8758 14688 8786
rect 14292 8090 14412 8106
rect 14292 8084 14424 8090
rect 14292 8078 14372 8084
rect 14372 8026 14424 8032
rect 14292 7806 14596 7834
rect 14292 7478 14320 7806
rect 14568 7750 14596 7806
rect 14464 7744 14516 7750
rect 14464 7686 14516 7692
rect 14556 7744 14608 7750
rect 14556 7686 14608 7692
rect 14280 7472 14332 7478
rect 14280 7414 14332 7420
rect 14280 7336 14332 7342
rect 14280 7278 14332 7284
rect 14292 6474 14320 7278
rect 14370 6488 14426 6497
rect 14292 6446 14370 6474
rect 14370 6423 14426 6432
rect 14384 6254 14412 6423
rect 14372 6248 14424 6254
rect 14372 6190 14424 6196
rect 14186 5808 14242 5817
rect 14186 5743 14242 5752
rect 14096 5636 14148 5642
rect 14096 5578 14148 5584
rect 13728 5296 13780 5302
rect 13728 5238 13780 5244
rect 14200 5250 14228 5743
rect 14384 5574 14412 6190
rect 14372 5568 14424 5574
rect 14372 5510 14424 5516
rect 14372 5296 14424 5302
rect 14370 5264 14372 5273
rect 14424 5264 14426 5273
rect 13740 4826 13768 5238
rect 13912 5228 13964 5234
rect 14200 5222 14320 5250
rect 13912 5170 13964 5176
rect 13820 5160 13872 5166
rect 13818 5128 13820 5137
rect 13872 5128 13874 5137
rect 13818 5063 13874 5072
rect 13820 5024 13872 5030
rect 13820 4966 13872 4972
rect 13728 4820 13780 4826
rect 13728 4762 13780 4768
rect 13452 4616 13504 4622
rect 13452 4558 13504 4564
rect 13544 4616 13596 4622
rect 13544 4558 13596 4564
rect 13360 4480 13412 4486
rect 13360 4422 13412 4428
rect 13360 4276 13412 4282
rect 13280 4236 13360 4264
rect 13360 4218 13412 4224
rect 13464 4214 13492 4558
rect 13452 4208 13504 4214
rect 13452 4150 13504 4156
rect 13176 4072 13228 4078
rect 13174 4040 13176 4049
rect 13228 4040 13230 4049
rect 13174 3975 13230 3984
rect 13176 3936 13228 3942
rect 13174 3904 13176 3913
rect 13228 3904 13230 3913
rect 13174 3839 13230 3848
rect 13832 3754 13860 4966
rect 13648 3726 13860 3754
rect 13648 3670 13676 3726
rect 13636 3664 13688 3670
rect 13636 3606 13688 3612
rect 13544 3596 13596 3602
rect 13544 3538 13596 3544
rect 13556 3233 13584 3538
rect 13636 3528 13688 3534
rect 13636 3470 13688 3476
rect 13542 3224 13598 3233
rect 13084 3188 13136 3194
rect 13648 3194 13676 3470
rect 13542 3159 13598 3168
rect 13636 3188 13688 3194
rect 13084 3130 13136 3136
rect 13636 3130 13688 3136
rect 13924 2990 13952 5170
rect 14188 5092 14240 5098
rect 14188 5034 14240 5040
rect 13912 2984 13964 2990
rect 13912 2926 13964 2932
rect 14200 2854 14228 5034
rect 14292 4146 14320 5222
rect 14476 5234 14504 7686
rect 14556 6860 14608 6866
rect 14556 6802 14608 6808
rect 14568 6458 14596 6802
rect 14556 6452 14608 6458
rect 14556 6394 14608 6400
rect 14556 5636 14608 5642
rect 14556 5578 14608 5584
rect 14370 5199 14426 5208
rect 14464 5228 14516 5234
rect 14464 5170 14516 5176
rect 14370 5128 14426 5137
rect 14568 5114 14596 5578
rect 14370 5063 14426 5072
rect 14476 5086 14596 5114
rect 14384 4826 14412 5063
rect 14476 5030 14504 5086
rect 14464 5024 14516 5030
rect 14464 4966 14516 4972
rect 14556 5024 14608 5030
rect 14556 4966 14608 4972
rect 14372 4820 14424 4826
rect 14372 4762 14424 4768
rect 14280 4140 14332 4146
rect 14280 4082 14332 4088
rect 14292 3534 14320 4082
rect 14568 4010 14596 4966
rect 14660 4622 14688 8758
rect 14844 8242 14872 11047
rect 15016 11018 15068 11024
rect 14924 10464 14976 10470
rect 14924 10406 14976 10412
rect 14752 8214 14872 8242
rect 14648 4616 14700 4622
rect 14648 4558 14700 4564
rect 14752 4078 14780 8214
rect 14832 8084 14884 8090
rect 14832 8026 14884 8032
rect 14844 7342 14872 8026
rect 14832 7336 14884 7342
rect 14936 7313 14964 10406
rect 15028 10130 15056 11018
rect 15108 10464 15160 10470
rect 15108 10406 15160 10412
rect 15120 10266 15148 10406
rect 15108 10260 15160 10266
rect 15108 10202 15160 10208
rect 15212 10198 15240 14962
rect 15384 14952 15436 14958
rect 15384 14894 15436 14900
rect 15292 14884 15344 14890
rect 15292 14826 15344 14832
rect 15304 14793 15332 14826
rect 15290 14784 15346 14793
rect 15290 14719 15346 14728
rect 15396 14346 15424 14894
rect 15474 14784 15530 14793
rect 15474 14719 15530 14728
rect 15384 14340 15436 14346
rect 15384 14282 15436 14288
rect 15384 13388 15436 13394
rect 15384 13330 15436 13336
rect 15292 13320 15344 13326
rect 15292 13262 15344 13268
rect 15304 12782 15332 13262
rect 15292 12776 15344 12782
rect 15292 12718 15344 12724
rect 15396 12646 15424 13330
rect 15384 12640 15436 12646
rect 15384 12582 15436 12588
rect 15488 12442 15516 14719
rect 15476 12436 15528 12442
rect 15476 12378 15528 12384
rect 15580 12306 15608 16782
rect 15672 15978 15700 18006
rect 15750 17980 16046 18000
rect 15806 17978 15830 17980
rect 15886 17978 15910 17980
rect 15966 17978 15990 17980
rect 15828 17926 15830 17978
rect 15892 17926 15904 17978
rect 15966 17926 15968 17978
rect 15806 17924 15830 17926
rect 15886 17924 15910 17926
rect 15966 17924 15990 17926
rect 15750 17904 16046 17924
rect 15750 16892 16046 16912
rect 15806 16890 15830 16892
rect 15886 16890 15910 16892
rect 15966 16890 15990 16892
rect 15828 16838 15830 16890
rect 15892 16838 15904 16890
rect 15966 16838 15968 16890
rect 15806 16836 15830 16838
rect 15886 16836 15910 16838
rect 15966 16836 15990 16838
rect 15750 16816 16046 16836
rect 16028 16720 16080 16726
rect 16028 16662 16080 16668
rect 15842 16280 15898 16289
rect 15842 16215 15898 16224
rect 15856 15978 15884 16215
rect 16040 16017 16068 16662
rect 16118 16552 16174 16561
rect 16118 16487 16174 16496
rect 16026 16008 16082 16017
rect 15660 15972 15712 15978
rect 15660 15914 15712 15920
rect 15844 15972 15896 15978
rect 16026 15943 16082 15952
rect 15844 15914 15896 15920
rect 15672 15366 15700 15914
rect 15750 15804 16046 15824
rect 15806 15802 15830 15804
rect 15886 15802 15910 15804
rect 15966 15802 15990 15804
rect 15828 15750 15830 15802
rect 15892 15750 15904 15802
rect 15966 15750 15968 15802
rect 15806 15748 15830 15750
rect 15886 15748 15910 15750
rect 15966 15748 15990 15750
rect 15750 15728 16046 15748
rect 15752 15632 15804 15638
rect 15752 15574 15804 15580
rect 15764 15473 15792 15574
rect 15750 15464 15806 15473
rect 15750 15399 15806 15408
rect 15660 15360 15712 15366
rect 15660 15302 15712 15308
rect 15750 15328 15806 15337
rect 15750 15263 15806 15272
rect 15764 14958 15792 15263
rect 15934 15192 15990 15201
rect 15934 15127 15990 15136
rect 15948 14958 15976 15127
rect 15752 14952 15804 14958
rect 15752 14894 15804 14900
rect 15936 14952 15988 14958
rect 15936 14894 15988 14900
rect 16026 14920 16082 14929
rect 16132 14906 16160 16487
rect 16224 15026 16252 19110
rect 16316 18737 16344 19230
rect 16302 18728 16358 18737
rect 16302 18663 16358 18672
rect 16408 17762 16436 19332
rect 16486 19000 16542 19009
rect 16486 18935 16542 18944
rect 16500 18834 16528 18935
rect 16488 18828 16540 18834
rect 16488 18770 16540 18776
rect 16580 18828 16632 18834
rect 16580 18770 16632 18776
rect 16592 18465 16620 18770
rect 16578 18456 16634 18465
rect 16578 18391 16634 18400
rect 16488 18216 16540 18222
rect 16488 18158 16540 18164
rect 16316 17734 16436 17762
rect 16316 17202 16344 17734
rect 16396 17672 16448 17678
rect 16396 17614 16448 17620
rect 16304 17196 16356 17202
rect 16304 17138 16356 17144
rect 16304 16992 16356 16998
rect 16304 16934 16356 16940
rect 16316 16425 16344 16934
rect 16302 16416 16358 16425
rect 16302 16351 16358 16360
rect 16304 15904 16356 15910
rect 16304 15846 16356 15852
rect 16316 15706 16344 15846
rect 16304 15700 16356 15706
rect 16304 15642 16356 15648
rect 16304 15088 16356 15094
rect 16304 15030 16356 15036
rect 16212 15020 16264 15026
rect 16212 14962 16264 14968
rect 16082 14878 16160 14906
rect 16026 14855 16082 14864
rect 15660 14816 15712 14822
rect 15660 14758 15712 14764
rect 15672 14278 15700 14758
rect 15750 14716 16046 14736
rect 15806 14714 15830 14716
rect 15886 14714 15910 14716
rect 15966 14714 15990 14716
rect 15828 14662 15830 14714
rect 15892 14662 15904 14714
rect 15966 14662 15968 14714
rect 15806 14660 15830 14662
rect 15886 14660 15910 14662
rect 15966 14660 15990 14662
rect 15750 14640 16046 14660
rect 16120 14612 16172 14618
rect 16120 14554 16172 14560
rect 16132 14362 16160 14554
rect 16316 14482 16344 15030
rect 16304 14476 16356 14482
rect 16304 14418 16356 14424
rect 16040 14334 16160 14362
rect 15660 14272 15712 14278
rect 16040 14249 16068 14334
rect 16120 14272 16172 14278
rect 15660 14214 15712 14220
rect 16026 14240 16082 14249
rect 16120 14214 16172 14220
rect 16026 14175 16082 14184
rect 16026 14104 16082 14113
rect 16026 14039 16082 14048
rect 15660 13728 15712 13734
rect 16040 13716 16068 14039
rect 16132 13938 16160 14214
rect 16302 14104 16358 14113
rect 16302 14039 16358 14048
rect 16212 14000 16264 14006
rect 16212 13942 16264 13948
rect 16120 13932 16172 13938
rect 16120 13874 16172 13880
rect 16224 13734 16252 13942
rect 16120 13728 16172 13734
rect 16040 13688 16120 13716
rect 15660 13670 15712 13676
rect 16120 13670 16172 13676
rect 16212 13728 16264 13734
rect 16212 13670 16264 13676
rect 15672 13025 15700 13670
rect 15750 13628 16046 13648
rect 15806 13626 15830 13628
rect 15886 13626 15910 13628
rect 15966 13626 15990 13628
rect 15828 13574 15830 13626
rect 15892 13574 15904 13626
rect 15966 13574 15968 13626
rect 15806 13572 15830 13574
rect 15886 13572 15910 13574
rect 15966 13572 15990 13574
rect 15750 13552 16046 13572
rect 16210 13560 16266 13569
rect 16132 13518 16210 13546
rect 15658 13016 15714 13025
rect 15658 12951 15714 12960
rect 15660 12708 15712 12714
rect 15660 12650 15712 12656
rect 15568 12300 15620 12306
rect 15568 12242 15620 12248
rect 15672 11898 15700 12650
rect 15750 12540 16046 12560
rect 15806 12538 15830 12540
rect 15886 12538 15910 12540
rect 15966 12538 15990 12540
rect 15828 12486 15830 12538
rect 15892 12486 15904 12538
rect 15966 12486 15968 12538
rect 15806 12484 15830 12486
rect 15886 12484 15910 12486
rect 15966 12484 15990 12486
rect 15750 12464 16046 12484
rect 15660 11892 15712 11898
rect 15660 11834 15712 11840
rect 15750 11452 16046 11472
rect 15806 11450 15830 11452
rect 15886 11450 15910 11452
rect 15966 11450 15990 11452
rect 15828 11398 15830 11450
rect 15892 11398 15904 11450
rect 15966 11398 15968 11450
rect 15806 11396 15830 11398
rect 15886 11396 15910 11398
rect 15966 11396 15990 11398
rect 15750 11376 16046 11396
rect 15292 11280 15344 11286
rect 15292 11222 15344 11228
rect 15658 11248 15714 11257
rect 15304 10606 15332 11222
rect 15658 11183 15660 11192
rect 15712 11183 15714 11192
rect 15660 11154 15712 11160
rect 15292 10600 15344 10606
rect 15292 10542 15344 10548
rect 15304 10266 15332 10542
rect 15660 10532 15712 10538
rect 15660 10474 15712 10480
rect 15382 10296 15438 10305
rect 15292 10260 15344 10266
rect 15382 10231 15438 10240
rect 15292 10202 15344 10208
rect 15200 10192 15252 10198
rect 15200 10134 15252 10140
rect 15396 10130 15424 10231
rect 15672 10198 15700 10474
rect 15750 10364 16046 10384
rect 15806 10362 15830 10364
rect 15886 10362 15910 10364
rect 15966 10362 15990 10364
rect 15828 10310 15830 10362
rect 15892 10310 15904 10362
rect 15966 10310 15968 10362
rect 15806 10308 15830 10310
rect 15886 10308 15910 10310
rect 15966 10308 15990 10310
rect 15750 10288 16046 10308
rect 15660 10192 15712 10198
rect 15660 10134 15712 10140
rect 15016 10124 15068 10130
rect 15016 10066 15068 10072
rect 15384 10124 15436 10130
rect 15384 10066 15436 10072
rect 15016 9920 15068 9926
rect 15016 9862 15068 9868
rect 15198 9888 15254 9897
rect 15028 9518 15056 9862
rect 15198 9823 15254 9832
rect 15016 9512 15068 9518
rect 15016 9454 15068 9460
rect 15028 7954 15056 9454
rect 15108 9376 15160 9382
rect 15108 9318 15160 9324
rect 15120 9178 15148 9318
rect 15108 9172 15160 9178
rect 15108 9114 15160 9120
rect 15108 8288 15160 8294
rect 15108 8230 15160 8236
rect 15016 7948 15068 7954
rect 15016 7890 15068 7896
rect 14832 7278 14884 7284
rect 14922 7304 14978 7313
rect 14922 7239 14978 7248
rect 15016 6792 15068 6798
rect 15016 6734 15068 6740
rect 15028 6497 15056 6734
rect 15014 6488 15070 6497
rect 15014 6423 15070 6432
rect 15120 5370 15148 8230
rect 15108 5364 15160 5370
rect 15108 5306 15160 5312
rect 14830 5264 14886 5273
rect 14830 5199 14886 5208
rect 14740 4072 14792 4078
rect 14740 4014 14792 4020
rect 14556 4004 14608 4010
rect 14556 3946 14608 3952
rect 14844 3602 14872 5199
rect 14922 4448 14978 4457
rect 14922 4383 14978 4392
rect 14936 3670 14964 4383
rect 15212 4162 15240 9823
rect 15396 9704 15424 10066
rect 16028 9920 16080 9926
rect 16132 9908 16160 13518
rect 16210 13495 16266 13504
rect 16316 13326 16344 14039
rect 16408 14006 16436 17614
rect 16500 17241 16528 18158
rect 16486 17232 16542 17241
rect 16486 17167 16542 17176
rect 16488 16992 16540 16998
rect 16488 16934 16540 16940
rect 16500 16794 16528 16934
rect 16488 16788 16540 16794
rect 16488 16730 16540 16736
rect 16488 16652 16540 16658
rect 16488 16594 16540 16600
rect 16396 14000 16448 14006
rect 16396 13942 16448 13948
rect 16500 13870 16528 16594
rect 16592 15337 16620 18391
rect 16776 17898 16804 19479
rect 16868 18834 16896 21422
rect 16856 18828 16908 18834
rect 16856 18770 16908 18776
rect 16776 17870 16896 17898
rect 16764 17808 16816 17814
rect 16762 17776 16764 17785
rect 16816 17776 16818 17785
rect 16868 17746 16896 17870
rect 16762 17711 16818 17720
rect 16856 17740 16908 17746
rect 16856 17682 16908 17688
rect 16764 17196 16816 17202
rect 16764 17138 16816 17144
rect 16672 17128 16724 17134
rect 16672 17070 16724 17076
rect 16684 16522 16712 17070
rect 16776 16658 16804 17138
rect 16960 17082 16988 21542
rect 17408 21480 17460 21486
rect 17144 21440 17408 21468
rect 17144 18737 17172 21440
rect 17408 21422 17460 21428
rect 17408 20936 17460 20942
rect 17408 20878 17460 20884
rect 17592 20936 17644 20942
rect 17592 20878 17644 20884
rect 17222 20496 17278 20505
rect 17222 20431 17278 20440
rect 17130 18728 17186 18737
rect 17130 18663 17186 18672
rect 17040 18624 17092 18630
rect 17040 18566 17092 18572
rect 17132 18624 17184 18630
rect 17132 18566 17184 18572
rect 17052 17882 17080 18566
rect 17040 17876 17092 17882
rect 17040 17818 17092 17824
rect 17040 17740 17092 17746
rect 17040 17682 17092 17688
rect 17052 17116 17080 17682
rect 17144 17241 17172 18566
rect 17130 17232 17186 17241
rect 17130 17167 17186 17176
rect 17236 17134 17264 20431
rect 17420 19718 17448 20878
rect 17500 19780 17552 19786
rect 17500 19722 17552 19728
rect 17408 19712 17460 19718
rect 17408 19654 17460 19660
rect 17512 19446 17540 19722
rect 17500 19440 17552 19446
rect 17500 19382 17552 19388
rect 17604 19378 17632 20878
rect 17592 19372 17644 19378
rect 17592 19314 17644 19320
rect 17500 18828 17552 18834
rect 17500 18770 17552 18776
rect 17408 18624 17460 18630
rect 17408 18566 17460 18572
rect 17420 18154 17448 18566
rect 17408 18148 17460 18154
rect 17408 18090 17460 18096
rect 17316 17740 17368 17746
rect 17316 17682 17368 17688
rect 17224 17128 17276 17134
rect 17052 17088 17172 17116
rect 16868 17054 16988 17082
rect 16764 16652 16816 16658
rect 16764 16594 16816 16600
rect 16672 16516 16724 16522
rect 16672 16458 16724 16464
rect 16764 16516 16816 16522
rect 16764 16458 16816 16464
rect 16776 16425 16804 16458
rect 16762 16416 16818 16425
rect 16762 16351 16818 16360
rect 16670 16008 16726 16017
rect 16670 15943 16726 15952
rect 16684 15910 16712 15943
rect 16672 15904 16724 15910
rect 16672 15846 16724 15852
rect 16578 15328 16634 15337
rect 16578 15263 16634 15272
rect 16578 15192 16634 15201
rect 16578 15127 16634 15136
rect 16592 14822 16620 15127
rect 16672 14884 16724 14890
rect 16672 14826 16724 14832
rect 16580 14816 16632 14822
rect 16580 14758 16632 14764
rect 16684 14414 16712 14826
rect 16764 14816 16816 14822
rect 16764 14758 16816 14764
rect 16580 14408 16632 14414
rect 16580 14350 16632 14356
rect 16672 14408 16724 14414
rect 16672 14350 16724 14356
rect 16592 14074 16620 14350
rect 16580 14068 16632 14074
rect 16580 14010 16632 14016
rect 16776 13977 16804 14758
rect 16762 13968 16818 13977
rect 16762 13903 16818 13912
rect 16488 13864 16540 13870
rect 16488 13806 16540 13812
rect 16672 13864 16724 13870
rect 16672 13806 16724 13812
rect 16394 13696 16450 13705
rect 16394 13631 16450 13640
rect 16304 13320 16356 13326
rect 16304 13262 16356 13268
rect 16316 12782 16344 13262
rect 16304 12776 16356 12782
rect 16304 12718 16356 12724
rect 16210 12608 16266 12617
rect 16210 12543 16266 12552
rect 16224 12442 16252 12543
rect 16316 12442 16344 12718
rect 16212 12436 16264 12442
rect 16212 12378 16264 12384
rect 16304 12436 16356 12442
rect 16304 12378 16356 12384
rect 16302 12064 16358 12073
rect 16302 11999 16358 12008
rect 16212 11552 16264 11558
rect 16316 11529 16344 11999
rect 16212 11494 16264 11500
rect 16302 11520 16358 11529
rect 16224 10792 16252 11494
rect 16302 11455 16358 11464
rect 16224 10764 16344 10792
rect 16212 10668 16264 10674
rect 16212 10610 16264 10616
rect 16080 9880 16160 9908
rect 16028 9862 16080 9868
rect 15566 9752 15622 9761
rect 15476 9716 15528 9722
rect 15396 9676 15476 9704
rect 15566 9687 15622 9696
rect 15476 9658 15528 9664
rect 15384 9444 15436 9450
rect 15384 9386 15436 9392
rect 15396 9330 15424 9386
rect 15304 9302 15424 9330
rect 15304 9178 15332 9302
rect 15580 9194 15608 9687
rect 16118 9616 16174 9625
rect 16118 9551 16174 9560
rect 15750 9276 16046 9296
rect 15806 9274 15830 9276
rect 15886 9274 15910 9276
rect 15966 9274 15990 9276
rect 15828 9222 15830 9274
rect 15892 9222 15904 9274
rect 15966 9222 15968 9274
rect 15806 9220 15830 9222
rect 15886 9220 15910 9222
rect 15966 9220 15990 9222
rect 15750 9200 16046 9220
rect 15292 9172 15344 9178
rect 15292 9114 15344 9120
rect 15384 9172 15436 9178
rect 15384 9114 15436 9120
rect 15571 9166 15608 9194
rect 15292 8560 15344 8566
rect 15292 8502 15344 8508
rect 15304 8430 15332 8502
rect 15292 8424 15344 8430
rect 15292 8366 15344 8372
rect 15396 8265 15424 9114
rect 15571 9092 15599 9166
rect 15571 9064 15608 9092
rect 16132 9081 16160 9551
rect 15476 8900 15528 8906
rect 15476 8842 15528 8848
rect 15488 8634 15516 8842
rect 15476 8628 15528 8634
rect 15476 8570 15528 8576
rect 15476 8492 15528 8498
rect 15476 8434 15528 8440
rect 15382 8256 15438 8265
rect 15382 8191 15438 8200
rect 15382 8120 15438 8129
rect 15382 8055 15384 8064
rect 15436 8055 15438 8064
rect 15384 8026 15436 8032
rect 15488 7970 15516 8434
rect 15304 7954 15516 7970
rect 15292 7948 15516 7954
rect 15344 7942 15516 7948
rect 15292 7890 15344 7896
rect 15292 7268 15344 7274
rect 15292 7210 15344 7216
rect 15304 6458 15332 7210
rect 15580 6984 15608 9064
rect 16118 9072 16174 9081
rect 16118 9007 16174 9016
rect 15752 8968 15804 8974
rect 15804 8928 15884 8956
rect 15752 8910 15804 8916
rect 15660 8900 15712 8906
rect 15660 8842 15712 8848
rect 15672 7546 15700 8842
rect 15750 8664 15806 8673
rect 15750 8599 15806 8608
rect 15764 8362 15792 8599
rect 15856 8362 15884 8928
rect 16120 8492 16172 8498
rect 16120 8434 16172 8440
rect 15752 8356 15804 8362
rect 15752 8298 15804 8304
rect 15844 8356 15896 8362
rect 15844 8298 15896 8304
rect 15750 8188 16046 8208
rect 15806 8186 15830 8188
rect 15886 8186 15910 8188
rect 15966 8186 15990 8188
rect 15828 8134 15830 8186
rect 15892 8134 15904 8186
rect 15966 8134 15968 8186
rect 15806 8132 15830 8134
rect 15886 8132 15910 8134
rect 15966 8132 15990 8134
rect 15750 8112 16046 8132
rect 16132 7886 16160 8434
rect 15752 7880 15804 7886
rect 15752 7822 15804 7828
rect 16120 7880 16172 7886
rect 16120 7822 16172 7828
rect 15660 7540 15712 7546
rect 15660 7482 15712 7488
rect 15488 6956 15608 6984
rect 15292 6452 15344 6458
rect 15292 6394 15344 6400
rect 15292 4684 15344 4690
rect 15292 4626 15344 4632
rect 15028 4146 15240 4162
rect 15016 4140 15240 4146
rect 15068 4134 15240 4140
rect 15016 4082 15068 4088
rect 15200 4072 15252 4078
rect 15200 4014 15252 4020
rect 14924 3664 14976 3670
rect 14924 3606 14976 3612
rect 14832 3596 14884 3602
rect 14832 3538 14884 3544
rect 14280 3528 14332 3534
rect 14280 3470 14332 3476
rect 14372 3392 14424 3398
rect 14372 3334 14424 3340
rect 12992 2848 13044 2854
rect 12992 2790 13044 2796
rect 14188 2848 14240 2854
rect 14188 2790 14240 2796
rect 14384 2650 14412 3334
rect 14464 2848 14516 2854
rect 14464 2790 14516 2796
rect 14372 2644 14424 2650
rect 14372 2586 14424 2592
rect 14476 2582 14504 2790
rect 14464 2576 14516 2582
rect 14464 2518 14516 2524
rect 14832 2440 14884 2446
rect 14832 2382 14884 2388
rect 15016 2440 15068 2446
rect 15016 2382 15068 2388
rect 12052 2204 12348 2224
rect 12108 2202 12132 2204
rect 12188 2202 12212 2204
rect 12268 2202 12292 2204
rect 12130 2150 12132 2202
rect 12194 2150 12206 2202
rect 12268 2150 12270 2202
rect 12108 2148 12132 2150
rect 12188 2148 12212 2150
rect 12268 2148 12292 2150
rect 12052 2128 12348 2148
rect 14844 2106 14872 2382
rect 14832 2100 14884 2106
rect 11992 2060 12112 2088
rect 12084 800 12112 2060
rect 14832 2042 14884 2048
rect 15028 2038 15056 2382
rect 15212 2310 15240 4014
rect 15304 4010 15332 4626
rect 15292 4004 15344 4010
rect 15292 3946 15344 3952
rect 15488 3058 15516 6956
rect 15568 6860 15620 6866
rect 15672 6848 15700 7482
rect 15764 7313 15792 7822
rect 16224 7449 16252 10610
rect 16316 8480 16344 10764
rect 16408 9178 16436 13631
rect 16500 13462 16528 13806
rect 16488 13456 16540 13462
rect 16488 13398 16540 13404
rect 16580 13456 16632 13462
rect 16684 13444 16712 13806
rect 16764 13524 16816 13530
rect 16764 13466 16816 13472
rect 16632 13416 16712 13444
rect 16580 13398 16632 13404
rect 16776 13240 16804 13466
rect 16592 13212 16804 13240
rect 16592 12782 16620 13212
rect 16868 13172 16896 17054
rect 16948 16992 17000 16998
rect 16948 16934 17000 16940
rect 17040 16992 17092 16998
rect 17040 16934 17092 16940
rect 16960 16726 16988 16934
rect 16948 16720 17000 16726
rect 16948 16662 17000 16668
rect 16948 16584 17000 16590
rect 16948 16526 17000 16532
rect 16960 15502 16988 16526
rect 17052 16425 17080 16934
rect 17038 16416 17094 16425
rect 17038 16351 17094 16360
rect 17040 16176 17092 16182
rect 17040 16118 17092 16124
rect 17052 15570 17080 16118
rect 17040 15564 17092 15570
rect 17040 15506 17092 15512
rect 16948 15496 17000 15502
rect 16948 15438 17000 15444
rect 16948 15360 17000 15366
rect 17144 15314 17172 17088
rect 17224 17070 17276 17076
rect 17224 16652 17276 16658
rect 17224 16594 17276 16600
rect 17236 15366 17264 16594
rect 16948 15302 17000 15308
rect 16684 13144 16896 13172
rect 16580 12776 16632 12782
rect 16580 12718 16632 12724
rect 16684 12152 16712 13144
rect 16856 12776 16908 12782
rect 16856 12718 16908 12724
rect 16868 12646 16896 12718
rect 16856 12640 16908 12646
rect 16856 12582 16908 12588
rect 16854 12472 16910 12481
rect 16854 12407 16910 12416
rect 16764 12368 16816 12374
rect 16764 12310 16816 12316
rect 16592 12124 16712 12152
rect 16488 11280 16540 11286
rect 16488 11222 16540 11228
rect 16500 10742 16528 11222
rect 16488 10736 16540 10742
rect 16488 10678 16540 10684
rect 16592 10470 16620 12124
rect 16670 12064 16726 12073
rect 16670 11999 16726 12008
rect 16684 11218 16712 11999
rect 16776 11762 16804 12310
rect 16764 11756 16816 11762
rect 16764 11698 16816 11704
rect 16762 11248 16818 11257
rect 16672 11212 16724 11218
rect 16762 11183 16764 11192
rect 16672 11154 16724 11160
rect 16816 11183 16818 11192
rect 16764 11154 16816 11160
rect 16868 10713 16896 12407
rect 16670 10704 16726 10713
rect 16670 10639 16726 10648
rect 16854 10704 16910 10713
rect 16854 10639 16910 10648
rect 16684 10538 16712 10639
rect 16960 10606 16988 15302
rect 17052 15286 17172 15314
rect 17224 15360 17276 15366
rect 17224 15302 17276 15308
rect 16948 10600 17000 10606
rect 16948 10542 17000 10548
rect 16672 10532 16724 10538
rect 16672 10474 16724 10480
rect 16580 10464 16632 10470
rect 16580 10406 16632 10412
rect 16856 10464 16908 10470
rect 16856 10406 16908 10412
rect 16488 10192 16540 10198
rect 16488 10134 16540 10140
rect 16396 9172 16448 9178
rect 16396 9114 16448 9120
rect 16394 9072 16450 9081
rect 16500 9042 16528 10134
rect 16580 9580 16632 9586
rect 16764 9580 16816 9586
rect 16632 9540 16712 9568
rect 16580 9522 16632 9528
rect 16580 9376 16632 9382
rect 16580 9318 16632 9324
rect 16394 9007 16450 9016
rect 16488 9036 16540 9042
rect 16408 8974 16436 9007
rect 16488 8978 16540 8984
rect 16396 8968 16448 8974
rect 16396 8910 16448 8916
rect 16488 8900 16540 8906
rect 16488 8842 16540 8848
rect 16500 8809 16528 8842
rect 16486 8800 16542 8809
rect 16486 8735 16542 8744
rect 16500 8498 16528 8735
rect 16592 8498 16620 9318
rect 16684 9178 16712 9540
rect 16764 9522 16816 9528
rect 16672 9172 16724 9178
rect 16672 9114 16724 9120
rect 16488 8492 16540 8498
rect 16316 8452 16436 8480
rect 16304 8288 16356 8294
rect 16304 8230 16356 8236
rect 16316 8090 16344 8230
rect 16304 8084 16356 8090
rect 16304 8026 16356 8032
rect 16408 7970 16436 8452
rect 16488 8434 16540 8440
rect 16580 8492 16632 8498
rect 16580 8434 16632 8440
rect 16488 8084 16540 8090
rect 16592 8072 16620 8434
rect 16540 8044 16620 8072
rect 16488 8026 16540 8032
rect 16408 7942 16528 7970
rect 16210 7440 16266 7449
rect 16210 7375 16266 7384
rect 15750 7304 15806 7313
rect 15750 7239 15806 7248
rect 16120 7200 16172 7206
rect 16120 7142 16172 7148
rect 15750 7100 16046 7120
rect 15806 7098 15830 7100
rect 15886 7098 15910 7100
rect 15966 7098 15990 7100
rect 15828 7046 15830 7098
rect 15892 7046 15904 7098
rect 15966 7046 15968 7098
rect 15806 7044 15830 7046
rect 15886 7044 15910 7046
rect 15966 7044 15990 7046
rect 15750 7024 16046 7044
rect 15620 6820 15700 6848
rect 15568 6802 15620 6808
rect 16132 6497 16160 7142
rect 16304 6928 16356 6934
rect 16500 6905 16528 7942
rect 16672 7812 16724 7818
rect 16672 7754 16724 7760
rect 16684 7585 16712 7754
rect 16670 7576 16726 7585
rect 16670 7511 16726 7520
rect 16672 6928 16724 6934
rect 16304 6870 16356 6876
rect 16486 6896 16542 6905
rect 16118 6488 16174 6497
rect 15660 6452 15712 6458
rect 16118 6423 16174 6432
rect 15660 6394 15712 6400
rect 15672 5234 15700 6394
rect 15750 6012 16046 6032
rect 15806 6010 15830 6012
rect 15886 6010 15910 6012
rect 15966 6010 15990 6012
rect 15828 5958 15830 6010
rect 15892 5958 15904 6010
rect 15966 5958 15968 6010
rect 15806 5956 15830 5958
rect 15886 5956 15910 5958
rect 15966 5956 15990 5958
rect 15750 5936 16046 5956
rect 16132 5710 16160 6423
rect 16316 5817 16344 6870
rect 16672 6870 16724 6876
rect 16486 6831 16542 6840
rect 16302 5808 16358 5817
rect 16302 5743 16358 5752
rect 16120 5704 16172 5710
rect 16120 5646 16172 5652
rect 16028 5636 16080 5642
rect 16028 5578 16080 5584
rect 16040 5370 16068 5578
rect 16028 5364 16080 5370
rect 16028 5306 16080 5312
rect 15660 5228 15712 5234
rect 15660 5170 15712 5176
rect 15660 5092 15712 5098
rect 15660 5034 15712 5040
rect 15672 4826 15700 5034
rect 15750 4924 16046 4944
rect 15806 4922 15830 4924
rect 15886 4922 15910 4924
rect 15966 4922 15990 4924
rect 15828 4870 15830 4922
rect 15892 4870 15904 4922
rect 15966 4870 15968 4922
rect 15806 4868 15830 4870
rect 15886 4868 15910 4870
rect 15966 4868 15990 4870
rect 15750 4848 16046 4868
rect 15660 4820 15712 4826
rect 15660 4762 15712 4768
rect 15936 4684 15988 4690
rect 16132 4672 16160 5646
rect 16316 5234 16344 5743
rect 16304 5228 16356 5234
rect 16304 5170 16356 5176
rect 16396 5160 16448 5166
rect 16684 5148 16712 6870
rect 16776 6866 16804 9522
rect 16764 6860 16816 6866
rect 16764 6802 16816 6808
rect 16776 6730 16804 6802
rect 16764 6724 16816 6730
rect 16764 6666 16816 6672
rect 16448 5120 16712 5148
rect 16396 5102 16448 5108
rect 15988 4644 16160 4672
rect 15936 4626 15988 4632
rect 15660 4616 15712 4622
rect 15660 4558 15712 4564
rect 15672 4078 15700 4558
rect 16580 4480 16632 4486
rect 16580 4422 16632 4428
rect 16118 4176 16174 4185
rect 16118 4111 16174 4120
rect 15660 4072 15712 4078
rect 15660 4014 15712 4020
rect 15672 3534 15700 4014
rect 15750 3836 16046 3856
rect 15806 3834 15830 3836
rect 15886 3834 15910 3836
rect 15966 3834 15990 3836
rect 15828 3782 15830 3834
rect 15892 3782 15904 3834
rect 15966 3782 15968 3834
rect 15806 3780 15830 3782
rect 15886 3780 15910 3782
rect 15966 3780 15990 3782
rect 15750 3760 16046 3780
rect 15568 3528 15620 3534
rect 15568 3470 15620 3476
rect 15660 3528 15712 3534
rect 15660 3470 15712 3476
rect 15580 3058 15608 3470
rect 15476 3052 15528 3058
rect 15476 2994 15528 3000
rect 15568 3052 15620 3058
rect 15568 2994 15620 3000
rect 15580 2582 15608 2994
rect 16132 2990 16160 4111
rect 16592 4078 16620 4422
rect 16580 4072 16632 4078
rect 16580 4014 16632 4020
rect 16396 3188 16448 3194
rect 16396 3130 16448 3136
rect 16120 2984 16172 2990
rect 16120 2926 16172 2932
rect 15750 2748 16046 2768
rect 15806 2746 15830 2748
rect 15886 2746 15910 2748
rect 15966 2746 15990 2748
rect 15828 2694 15830 2746
rect 15892 2694 15904 2746
rect 15966 2694 15968 2746
rect 15806 2692 15830 2694
rect 15886 2692 15910 2694
rect 15966 2692 15990 2694
rect 15750 2672 16046 2692
rect 15568 2576 15620 2582
rect 15568 2518 15620 2524
rect 15934 2544 15990 2553
rect 16408 2514 16436 3130
rect 15934 2479 15936 2488
rect 15988 2479 15990 2488
rect 16396 2508 16448 2514
rect 15936 2450 15988 2456
rect 16396 2450 16448 2456
rect 15200 2304 15252 2310
rect 15200 2246 15252 2252
rect 15016 2032 15068 2038
rect 15016 1974 15068 1980
rect 16868 1970 16896 10406
rect 16948 10192 17000 10198
rect 16948 10134 17000 10140
rect 16960 7750 16988 10134
rect 17052 9518 17080 15286
rect 17224 14884 17276 14890
rect 17224 14826 17276 14832
rect 17132 14544 17184 14550
rect 17132 14486 17184 14492
rect 17144 13938 17172 14486
rect 17132 13932 17184 13938
rect 17132 13874 17184 13880
rect 17132 13796 17184 13802
rect 17132 13738 17184 13744
rect 17144 13161 17172 13738
rect 17236 13394 17264 14826
rect 17328 14618 17356 17682
rect 17408 17536 17460 17542
rect 17408 17478 17460 17484
rect 17316 14612 17368 14618
rect 17316 14554 17368 14560
rect 17314 14512 17370 14521
rect 17314 14447 17370 14456
rect 17328 14278 17356 14447
rect 17316 14272 17368 14278
rect 17316 14214 17368 14220
rect 17314 13696 17370 13705
rect 17314 13631 17370 13640
rect 17224 13388 17276 13394
rect 17224 13330 17276 13336
rect 17130 13152 17186 13161
rect 17130 13087 17186 13096
rect 17236 12442 17264 13330
rect 17328 13297 17356 13631
rect 17314 13288 17370 13297
rect 17314 13223 17370 13232
rect 17316 12912 17368 12918
rect 17316 12854 17368 12860
rect 17132 12436 17184 12442
rect 17132 12378 17184 12384
rect 17224 12436 17276 12442
rect 17224 12378 17276 12384
rect 17144 12238 17172 12378
rect 17132 12232 17184 12238
rect 17132 12174 17184 12180
rect 17222 12200 17278 12209
rect 17222 12135 17278 12144
rect 17132 11144 17184 11150
rect 17132 11086 17184 11092
rect 17144 10130 17172 11086
rect 17132 10124 17184 10130
rect 17132 10066 17184 10072
rect 17130 10024 17186 10033
rect 17130 9959 17186 9968
rect 17040 9512 17092 9518
rect 17040 9454 17092 9460
rect 17038 8936 17094 8945
rect 17144 8922 17172 9959
rect 17094 8894 17172 8922
rect 17038 8871 17094 8880
rect 17236 8616 17264 12135
rect 17328 11801 17356 12854
rect 17420 12170 17448 17478
rect 17512 15910 17540 18770
rect 17604 17678 17632 19314
rect 17592 17672 17644 17678
rect 17592 17614 17644 17620
rect 17604 16130 17632 17614
rect 17696 16250 17724 22578
rect 18248 21486 18276 23600
rect 18328 22364 18380 22370
rect 18328 22306 18380 22312
rect 18236 21480 18288 21486
rect 18236 21422 18288 21428
rect 17776 21344 17828 21350
rect 17776 21286 17828 21292
rect 18052 21344 18104 21350
rect 18052 21286 18104 21292
rect 17788 19718 17816 21286
rect 17960 20936 18012 20942
rect 17960 20878 18012 20884
rect 17972 20398 18000 20878
rect 17960 20392 18012 20398
rect 17960 20334 18012 20340
rect 17972 19990 18000 20334
rect 17960 19984 18012 19990
rect 17960 19926 18012 19932
rect 17776 19712 17828 19718
rect 17776 19654 17828 19660
rect 17684 16244 17736 16250
rect 17684 16186 17736 16192
rect 17604 16102 17724 16130
rect 17696 16046 17724 16102
rect 17592 16040 17644 16046
rect 17592 15982 17644 15988
rect 17684 16040 17736 16046
rect 17684 15982 17736 15988
rect 17500 15904 17552 15910
rect 17500 15846 17552 15852
rect 17500 15564 17552 15570
rect 17500 15506 17552 15512
rect 17512 14822 17540 15506
rect 17500 14816 17552 14822
rect 17500 14758 17552 14764
rect 17498 12880 17554 12889
rect 17498 12815 17500 12824
rect 17552 12815 17554 12824
rect 17500 12786 17552 12792
rect 17500 12708 17552 12714
rect 17500 12650 17552 12656
rect 17408 12164 17460 12170
rect 17408 12106 17460 12112
rect 17314 11792 17370 11801
rect 17314 11727 17370 11736
rect 17408 11756 17460 11762
rect 17408 11698 17460 11704
rect 17316 11688 17368 11694
rect 17316 11630 17368 11636
rect 17328 11393 17356 11630
rect 17314 11384 17370 11393
rect 17314 11319 17370 11328
rect 17316 11212 17368 11218
rect 17316 11154 17368 11160
rect 17328 10810 17356 11154
rect 17420 10810 17448 11698
rect 17512 11014 17540 12650
rect 17604 12481 17632 15982
rect 17696 15337 17724 15982
rect 17682 15328 17738 15337
rect 17682 15263 17738 15272
rect 17788 13870 17816 19654
rect 18064 19496 18092 21286
rect 18234 20632 18290 20641
rect 18234 20567 18290 20576
rect 18144 20392 18196 20398
rect 18144 20334 18196 20340
rect 18156 20058 18184 20334
rect 18248 20058 18276 20567
rect 18144 20052 18196 20058
rect 18144 19994 18196 20000
rect 18236 20052 18288 20058
rect 18236 19994 18288 20000
rect 18236 19848 18288 19854
rect 18142 19816 18198 19825
rect 18236 19790 18288 19796
rect 18142 19751 18198 19760
rect 17880 19468 18092 19496
rect 17880 19156 17908 19468
rect 17960 19304 18012 19310
rect 18156 19292 18184 19751
rect 18012 19264 18184 19292
rect 17960 19246 18012 19252
rect 18144 19168 18196 19174
rect 17880 19128 18092 19156
rect 17960 18828 18012 18834
rect 17960 18770 18012 18776
rect 17868 18284 17920 18290
rect 17868 18226 17920 18232
rect 17880 16998 17908 18226
rect 17972 17105 18000 18770
rect 18064 18290 18092 19128
rect 18144 19110 18196 19116
rect 18156 18970 18184 19110
rect 18144 18964 18196 18970
rect 18144 18906 18196 18912
rect 18052 18284 18104 18290
rect 18052 18226 18104 18232
rect 18052 18148 18104 18154
rect 18052 18090 18104 18096
rect 18064 17678 18092 18090
rect 18052 17672 18104 17678
rect 18052 17614 18104 17620
rect 18064 17134 18092 17614
rect 18052 17128 18104 17134
rect 17958 17096 18014 17105
rect 18052 17070 18104 17076
rect 17958 17031 18014 17040
rect 17868 16992 17920 16998
rect 17868 16934 17920 16940
rect 18064 16658 18092 17070
rect 18144 17060 18196 17066
rect 18144 17002 18196 17008
rect 18156 16969 18184 17002
rect 18142 16960 18198 16969
rect 18142 16895 18198 16904
rect 18156 16726 18184 16895
rect 18144 16720 18196 16726
rect 18144 16662 18196 16668
rect 18052 16652 18104 16658
rect 18052 16594 18104 16600
rect 17868 16448 17920 16454
rect 17868 16390 17920 16396
rect 18144 16448 18196 16454
rect 18144 16390 18196 16396
rect 17880 16046 17908 16390
rect 17868 16040 17920 16046
rect 17868 15982 17920 15988
rect 17866 15736 17922 15745
rect 17866 15671 17922 15680
rect 17880 15026 17908 15671
rect 17960 15564 18012 15570
rect 17960 15506 18012 15512
rect 17868 15020 17920 15026
rect 17868 14962 17920 14968
rect 17868 14884 17920 14890
rect 17868 14826 17920 14832
rect 17776 13864 17828 13870
rect 17776 13806 17828 13812
rect 17880 13274 17908 14826
rect 17972 14006 18000 15506
rect 18052 15496 18104 15502
rect 18052 15438 18104 15444
rect 18064 14958 18092 15438
rect 18052 14952 18104 14958
rect 18052 14894 18104 14900
rect 18064 14550 18092 14894
rect 18052 14544 18104 14550
rect 18052 14486 18104 14492
rect 18064 14113 18092 14486
rect 18050 14104 18106 14113
rect 18050 14039 18106 14048
rect 17960 14000 18012 14006
rect 17960 13942 18012 13948
rect 18064 13938 18092 14039
rect 18052 13932 18104 13938
rect 18052 13874 18104 13880
rect 18064 13326 18092 13874
rect 18052 13320 18104 13326
rect 17696 13246 17908 13274
rect 17958 13288 18014 13297
rect 17696 12646 17724 13246
rect 18052 13262 18104 13268
rect 17958 13223 18014 13232
rect 17774 13152 17830 13161
rect 17774 13087 17830 13096
rect 17684 12640 17736 12646
rect 17684 12582 17736 12588
rect 17590 12472 17646 12481
rect 17590 12407 17646 12416
rect 17592 12300 17644 12306
rect 17696 12288 17724 12582
rect 17644 12260 17724 12288
rect 17592 12242 17644 12248
rect 17684 12164 17736 12170
rect 17684 12106 17736 12112
rect 17696 11830 17724 12106
rect 17684 11824 17736 11830
rect 17684 11766 17736 11772
rect 17682 11384 17738 11393
rect 17682 11319 17738 11328
rect 17500 11008 17552 11014
rect 17500 10950 17552 10956
rect 17316 10804 17368 10810
rect 17316 10746 17368 10752
rect 17408 10804 17460 10810
rect 17408 10746 17460 10752
rect 17328 10266 17356 10746
rect 17500 10668 17552 10674
rect 17500 10610 17552 10616
rect 17592 10668 17644 10674
rect 17592 10610 17644 10616
rect 17408 10464 17460 10470
rect 17408 10406 17460 10412
rect 17316 10260 17368 10266
rect 17316 10202 17368 10208
rect 17316 10124 17368 10130
rect 17316 10066 17368 10072
rect 17328 9722 17356 10066
rect 17316 9716 17368 9722
rect 17316 9658 17368 9664
rect 17420 9654 17448 10406
rect 17408 9648 17460 9654
rect 17408 9590 17460 9596
rect 17316 9376 17368 9382
rect 17316 9318 17368 9324
rect 17406 9344 17462 9353
rect 17328 9217 17356 9318
rect 17406 9279 17462 9288
rect 17314 9208 17370 9217
rect 17314 9143 17370 9152
rect 17144 8588 17264 8616
rect 17038 8120 17094 8129
rect 17038 8055 17094 8064
rect 16948 7744 17000 7750
rect 16948 7686 17000 7692
rect 16948 6996 17000 7002
rect 16948 6938 17000 6944
rect 16960 6361 16988 6938
rect 16946 6352 17002 6361
rect 16946 6287 17002 6296
rect 16946 4992 17002 5001
rect 16946 4927 17002 4936
rect 16960 3738 16988 4927
rect 16948 3732 17000 3738
rect 16948 3674 17000 3680
rect 17052 2922 17080 8055
rect 17144 6662 17172 8588
rect 17224 8424 17276 8430
rect 17224 8366 17276 8372
rect 17132 6656 17184 6662
rect 17132 6598 17184 6604
rect 17236 5914 17264 8366
rect 17316 8288 17368 8294
rect 17316 8230 17368 8236
rect 17328 8022 17356 8230
rect 17316 8016 17368 8022
rect 17316 7958 17368 7964
rect 17420 6934 17448 9279
rect 17512 7274 17540 10610
rect 17604 9110 17632 10610
rect 17592 9104 17644 9110
rect 17592 9046 17644 9052
rect 17604 7546 17632 9046
rect 17696 7818 17724 11319
rect 17684 7812 17736 7818
rect 17684 7754 17736 7760
rect 17592 7540 17644 7546
rect 17592 7482 17644 7488
rect 17500 7268 17552 7274
rect 17552 7228 17632 7256
rect 17500 7210 17552 7216
rect 17408 6928 17460 6934
rect 17408 6870 17460 6876
rect 17500 6860 17552 6866
rect 17500 6802 17552 6808
rect 17408 6316 17460 6322
rect 17512 6304 17540 6802
rect 17604 6662 17632 7228
rect 17592 6656 17644 6662
rect 17592 6598 17644 6604
rect 17460 6276 17540 6304
rect 17408 6258 17460 6264
rect 17684 6248 17736 6254
rect 17684 6190 17736 6196
rect 17316 6112 17368 6118
rect 17696 6089 17724 6190
rect 17316 6054 17368 6060
rect 17682 6080 17738 6089
rect 17224 5908 17276 5914
rect 17224 5850 17276 5856
rect 17224 4820 17276 4826
rect 17224 4762 17276 4768
rect 17132 4684 17184 4690
rect 17132 4626 17184 4632
rect 17144 4282 17172 4626
rect 17236 4282 17264 4762
rect 17132 4276 17184 4282
rect 17132 4218 17184 4224
rect 17224 4276 17276 4282
rect 17224 4218 17276 4224
rect 17144 3670 17172 4218
rect 17328 3942 17356 6054
rect 17682 6015 17738 6024
rect 17500 5908 17552 5914
rect 17500 5850 17552 5856
rect 17512 5166 17540 5850
rect 17684 5772 17736 5778
rect 17684 5714 17736 5720
rect 17696 5370 17724 5714
rect 17788 5710 17816 13087
rect 17868 12844 17920 12850
rect 17868 12786 17920 12792
rect 17880 12073 17908 12786
rect 17972 12209 18000 13223
rect 18052 13184 18104 13190
rect 18052 13126 18104 13132
rect 18064 12374 18092 13126
rect 18052 12368 18104 12374
rect 18052 12310 18104 12316
rect 17958 12200 18014 12209
rect 17958 12135 18014 12144
rect 17960 12096 18012 12102
rect 17866 12064 17922 12073
rect 17960 12038 18012 12044
rect 17866 11999 17922 12008
rect 17868 11756 17920 11762
rect 17868 11698 17920 11704
rect 17880 8786 17908 11698
rect 17972 11121 18000 12038
rect 18064 11558 18092 12310
rect 18156 12102 18184 16390
rect 18248 13569 18276 19790
rect 18340 19009 18368 22306
rect 18788 21072 18840 21078
rect 18788 21014 18840 21020
rect 18510 20088 18566 20097
rect 18510 20023 18566 20032
rect 18420 19712 18472 19718
rect 18420 19654 18472 19660
rect 18326 19000 18382 19009
rect 18326 18935 18382 18944
rect 18328 18828 18380 18834
rect 18328 18770 18380 18776
rect 18340 15570 18368 18770
rect 18328 15564 18380 15570
rect 18328 15506 18380 15512
rect 18328 13864 18380 13870
rect 18328 13806 18380 13812
rect 18234 13560 18290 13569
rect 18234 13495 18290 13504
rect 18340 13444 18368 13806
rect 18248 13416 18368 13444
rect 18144 12096 18196 12102
rect 18144 12038 18196 12044
rect 18144 11688 18196 11694
rect 18248 11665 18276 13416
rect 18328 12912 18380 12918
rect 18328 12854 18380 12860
rect 18144 11630 18196 11636
rect 18234 11656 18290 11665
rect 18052 11552 18104 11558
rect 18052 11494 18104 11500
rect 18156 11286 18184 11630
rect 18234 11591 18290 11600
rect 18144 11280 18196 11286
rect 18144 11222 18196 11228
rect 17958 11112 18014 11121
rect 18248 11082 18276 11591
rect 18340 11558 18368 12854
rect 18328 11552 18380 11558
rect 18328 11494 18380 11500
rect 18328 11144 18380 11150
rect 18328 11086 18380 11092
rect 17958 11047 18014 11056
rect 18236 11076 18288 11082
rect 18236 11018 18288 11024
rect 18052 10600 18104 10606
rect 18052 10542 18104 10548
rect 17960 10464 18012 10470
rect 17960 10406 18012 10412
rect 17972 9042 18000 10406
rect 18064 9382 18092 10542
rect 18144 10532 18196 10538
rect 18144 10474 18196 10480
rect 18052 9376 18104 9382
rect 18052 9318 18104 9324
rect 17960 9036 18012 9042
rect 17960 8978 18012 8984
rect 17960 8832 18012 8838
rect 17880 8780 17960 8786
rect 17880 8774 18012 8780
rect 17880 8758 18000 8774
rect 17880 8673 17908 8758
rect 17866 8664 17922 8673
rect 17866 8599 17922 8608
rect 17866 8528 17922 8537
rect 17866 8463 17922 8472
rect 17880 8430 17908 8463
rect 17868 8424 17920 8430
rect 17868 8366 17920 8372
rect 17868 8288 17920 8294
rect 17866 8256 17868 8265
rect 17920 8256 17922 8265
rect 17866 8191 17922 8200
rect 17960 7948 18012 7954
rect 17960 7890 18012 7896
rect 17972 7313 18000 7890
rect 18064 7478 18092 9318
rect 18156 8566 18184 10474
rect 18236 10124 18288 10130
rect 18236 10066 18288 10072
rect 18248 9722 18276 10066
rect 18340 10033 18368 11086
rect 18326 10024 18382 10033
rect 18326 9959 18382 9968
rect 18328 9920 18380 9926
rect 18328 9862 18380 9868
rect 18236 9716 18288 9722
rect 18236 9658 18288 9664
rect 18236 9580 18288 9586
rect 18236 9522 18288 9528
rect 18248 8634 18276 9522
rect 18340 9217 18368 9862
rect 18326 9208 18382 9217
rect 18326 9143 18382 9152
rect 18328 9036 18380 9042
rect 18328 8978 18380 8984
rect 18236 8628 18288 8634
rect 18236 8570 18288 8576
rect 18144 8560 18196 8566
rect 18144 8502 18196 8508
rect 18236 8424 18288 8430
rect 18236 8366 18288 8372
rect 18144 8288 18196 8294
rect 18144 8230 18196 8236
rect 18156 7954 18184 8230
rect 18144 7948 18196 7954
rect 18144 7890 18196 7896
rect 18052 7472 18104 7478
rect 18052 7414 18104 7420
rect 18144 7336 18196 7342
rect 17958 7304 18014 7313
rect 18144 7278 18196 7284
rect 17958 7239 18014 7248
rect 17960 6724 18012 6730
rect 17960 6666 18012 6672
rect 17972 6633 18000 6666
rect 17958 6624 18014 6633
rect 17958 6559 18014 6568
rect 18156 6322 18184 7278
rect 18248 6458 18276 8366
rect 18340 7886 18368 8978
rect 18432 8498 18460 19654
rect 18524 19378 18552 20023
rect 18604 19984 18656 19990
rect 18604 19926 18656 19932
rect 18512 19372 18564 19378
rect 18512 19314 18564 19320
rect 18524 18834 18552 19314
rect 18512 18828 18564 18834
rect 18512 18770 18564 18776
rect 18616 18714 18644 19926
rect 18696 19848 18748 19854
rect 18696 19790 18748 19796
rect 18524 18686 18644 18714
rect 18708 18698 18736 19790
rect 18800 19378 18828 21014
rect 18892 19718 18920 23600
rect 19338 23352 19394 23361
rect 19338 23287 19394 23296
rect 19352 22642 19380 23287
rect 19444 22914 19472 23967
rect 19522 23600 19578 24400
rect 20166 23600 20222 24400
rect 20810 23600 20866 24400
rect 21454 23600 21510 24400
rect 22098 23600 22154 24400
rect 22742 23600 22798 24400
rect 23386 23600 23442 24400
rect 24030 23600 24086 24400
rect 19432 22908 19484 22914
rect 19432 22850 19484 22856
rect 19340 22636 19392 22642
rect 19340 22578 19392 22584
rect 19536 22114 19564 23600
rect 19798 22672 19854 22681
rect 19798 22607 19854 22616
rect 19812 22370 19840 22607
rect 19800 22364 19852 22370
rect 19800 22306 19852 22312
rect 19536 22086 19656 22114
rect 19628 21962 19656 22086
rect 19156 21956 19208 21962
rect 19156 21898 19208 21904
rect 19616 21956 19668 21962
rect 19616 21898 19668 21904
rect 18972 21684 19024 21690
rect 18972 21626 19024 21632
rect 18880 19712 18932 19718
rect 18880 19654 18932 19660
rect 18788 19372 18840 19378
rect 18840 19332 18920 19360
rect 18788 19314 18840 19320
rect 18788 19168 18840 19174
rect 18788 19110 18840 19116
rect 18800 19009 18828 19110
rect 18786 19000 18842 19009
rect 18786 18935 18842 18944
rect 18892 18884 18920 19332
rect 18800 18856 18920 18884
rect 18800 18850 18828 18856
rect 18791 18822 18828 18850
rect 18791 18714 18819 18822
rect 18696 18692 18748 18698
rect 18524 18222 18552 18686
rect 18791 18686 18828 18714
rect 18696 18634 18748 18640
rect 18604 18624 18656 18630
rect 18604 18566 18656 18572
rect 18512 18216 18564 18222
rect 18512 18158 18564 18164
rect 18616 17814 18644 18566
rect 18604 17808 18656 17814
rect 18604 17750 18656 17756
rect 18512 16992 18564 16998
rect 18512 16934 18564 16940
rect 18524 16153 18552 16934
rect 18510 16144 18566 16153
rect 18510 16079 18566 16088
rect 18512 15156 18564 15162
rect 18512 15098 18564 15104
rect 18524 14618 18552 15098
rect 18512 14612 18564 14618
rect 18512 14554 18564 14560
rect 18510 14512 18566 14521
rect 18510 14447 18566 14456
rect 18524 13530 18552 14447
rect 18512 13524 18564 13530
rect 18512 13466 18564 13472
rect 18512 13184 18564 13190
rect 18512 13126 18564 13132
rect 18524 12889 18552 13126
rect 18510 12880 18566 12889
rect 18510 12815 18566 12824
rect 18512 12708 18564 12714
rect 18512 12650 18564 12656
rect 18524 10742 18552 12650
rect 18512 10736 18564 10742
rect 18512 10678 18564 10684
rect 18616 10282 18644 17750
rect 18524 10254 18644 10282
rect 18524 9489 18552 10254
rect 18604 10124 18656 10130
rect 18604 10066 18656 10072
rect 18510 9480 18566 9489
rect 18510 9415 18566 9424
rect 18512 9376 18564 9382
rect 18512 9318 18564 9324
rect 18420 8492 18472 8498
rect 18420 8434 18472 8440
rect 18420 8288 18472 8294
rect 18420 8230 18472 8236
rect 18328 7880 18380 7886
rect 18328 7822 18380 7828
rect 18340 7546 18368 7822
rect 18328 7540 18380 7546
rect 18328 7482 18380 7488
rect 18236 6452 18288 6458
rect 18236 6394 18288 6400
rect 18144 6316 18196 6322
rect 18144 6258 18196 6264
rect 18432 6118 18460 8230
rect 18524 7954 18552 9318
rect 18616 8974 18644 10066
rect 18708 9926 18736 18634
rect 18800 18426 18828 18686
rect 18788 18420 18840 18426
rect 18788 18362 18840 18368
rect 18880 18420 18932 18426
rect 18880 18362 18932 18368
rect 18788 17808 18840 17814
rect 18788 17750 18840 17756
rect 18800 15201 18828 17750
rect 18892 16561 18920 18362
rect 18984 16810 19012 21626
rect 19168 21418 19196 21898
rect 19800 21888 19852 21894
rect 19800 21830 19852 21836
rect 19449 21788 19745 21808
rect 19505 21786 19529 21788
rect 19585 21786 19609 21788
rect 19665 21786 19689 21788
rect 19527 21734 19529 21786
rect 19591 21734 19603 21786
rect 19665 21734 19667 21786
rect 19505 21732 19529 21734
rect 19585 21732 19609 21734
rect 19665 21732 19689 21734
rect 19449 21712 19745 21732
rect 19340 21548 19392 21554
rect 19340 21490 19392 21496
rect 19156 21412 19208 21418
rect 19156 21354 19208 21360
rect 19352 21321 19380 21490
rect 19812 21350 19840 21830
rect 19892 21548 19944 21554
rect 19892 21490 19944 21496
rect 19432 21344 19484 21350
rect 19338 21312 19394 21321
rect 19432 21286 19484 21292
rect 19800 21344 19852 21350
rect 19800 21286 19852 21292
rect 19338 21247 19394 21256
rect 19444 21162 19472 21286
rect 19352 21134 19472 21162
rect 19156 20868 19208 20874
rect 19156 20810 19208 20816
rect 19168 20398 19196 20810
rect 19352 20602 19380 21134
rect 19904 21010 19932 21490
rect 20076 21344 20128 21350
rect 20076 21286 20128 21292
rect 20088 21146 20116 21286
rect 20076 21140 20128 21146
rect 20076 21082 20128 21088
rect 19892 21004 19944 21010
rect 19892 20946 19944 20952
rect 19800 20800 19852 20806
rect 19800 20742 19852 20748
rect 19449 20700 19745 20720
rect 19505 20698 19529 20700
rect 19585 20698 19609 20700
rect 19665 20698 19689 20700
rect 19527 20646 19529 20698
rect 19591 20646 19603 20698
rect 19665 20646 19667 20698
rect 19505 20644 19529 20646
rect 19585 20644 19609 20646
rect 19665 20644 19689 20646
rect 19449 20624 19745 20644
rect 19340 20596 19392 20602
rect 19340 20538 19392 20544
rect 19812 20398 19840 20742
rect 19904 20602 19932 20946
rect 19892 20596 19944 20602
rect 19892 20538 19944 20544
rect 19156 20392 19208 20398
rect 19156 20334 19208 20340
rect 19708 20392 19760 20398
rect 19708 20334 19760 20340
rect 19800 20392 19852 20398
rect 20180 20369 20208 23600
rect 20442 21992 20498 22001
rect 20442 21927 20498 21936
rect 20352 21480 20404 21486
rect 20352 21422 20404 21428
rect 20364 21078 20392 21422
rect 20260 21072 20312 21078
rect 20260 21014 20312 21020
rect 20352 21072 20404 21078
rect 20352 21014 20404 21020
rect 20272 20618 20300 21014
rect 20272 20602 20392 20618
rect 20272 20596 20404 20602
rect 20272 20590 20352 20596
rect 19800 20334 19852 20340
rect 19890 20360 19946 20369
rect 19720 19700 19748 20334
rect 20166 20360 20222 20369
rect 19890 20295 19892 20304
rect 19944 20295 19946 20304
rect 20076 20324 20128 20330
rect 19892 20266 19944 20272
rect 20166 20295 20222 20304
rect 20076 20266 20128 20272
rect 19800 19712 19852 19718
rect 19720 19672 19800 19700
rect 19800 19654 19852 19660
rect 19449 19612 19745 19632
rect 19505 19610 19529 19612
rect 19585 19610 19609 19612
rect 19665 19610 19689 19612
rect 19527 19558 19529 19610
rect 19591 19558 19603 19610
rect 19665 19558 19667 19610
rect 19505 19556 19529 19558
rect 19585 19556 19609 19558
rect 19665 19556 19689 19558
rect 19449 19536 19745 19556
rect 19812 19378 19840 19654
rect 20088 19514 20116 20266
rect 20166 19816 20222 19825
rect 20166 19751 20222 19760
rect 20076 19508 20128 19514
rect 20076 19450 20128 19456
rect 19800 19372 19852 19378
rect 19800 19314 19852 19320
rect 20088 19174 20116 19205
rect 19064 19168 19116 19174
rect 19064 19110 19116 19116
rect 20076 19168 20128 19174
rect 20180 19122 20208 19751
rect 20128 19116 20208 19122
rect 20076 19110 20208 19116
rect 19076 17814 19104 19110
rect 20088 19094 20208 19110
rect 19984 18964 20036 18970
rect 19984 18906 20036 18912
rect 19800 18828 19852 18834
rect 19800 18770 19852 18776
rect 19892 18828 19944 18834
rect 19892 18770 19944 18776
rect 19248 18760 19300 18766
rect 19248 18702 19300 18708
rect 19156 18624 19208 18630
rect 19156 18566 19208 18572
rect 19168 18465 19196 18566
rect 19154 18456 19210 18465
rect 19260 18426 19288 18702
rect 19449 18524 19745 18544
rect 19505 18522 19529 18524
rect 19585 18522 19609 18524
rect 19665 18522 19689 18524
rect 19527 18470 19529 18522
rect 19591 18470 19603 18522
rect 19665 18470 19667 18522
rect 19505 18468 19529 18470
rect 19585 18468 19609 18470
rect 19665 18468 19689 18470
rect 19449 18448 19745 18468
rect 19154 18391 19210 18400
rect 19248 18420 19300 18426
rect 19248 18362 19300 18368
rect 19524 18352 19576 18358
rect 19524 18294 19576 18300
rect 19156 18148 19208 18154
rect 19156 18090 19208 18096
rect 19064 17808 19116 17814
rect 19064 17750 19116 17756
rect 19168 17542 19196 18090
rect 19248 18080 19300 18086
rect 19248 18022 19300 18028
rect 19260 17678 19288 18022
rect 19340 17876 19392 17882
rect 19340 17818 19392 17824
rect 19248 17672 19300 17678
rect 19248 17614 19300 17620
rect 19156 17536 19208 17542
rect 19156 17478 19208 17484
rect 19064 17264 19116 17270
rect 19064 17206 19116 17212
rect 19076 16998 19104 17206
rect 19064 16992 19116 16998
rect 19064 16934 19116 16940
rect 18984 16782 19104 16810
rect 18972 16652 19024 16658
rect 18972 16594 19024 16600
rect 18878 16552 18934 16561
rect 18878 16487 18934 16496
rect 18786 15192 18842 15201
rect 18786 15127 18842 15136
rect 18880 14544 18932 14550
rect 18880 14486 18932 14492
rect 18892 14414 18920 14486
rect 18880 14408 18932 14414
rect 18880 14350 18932 14356
rect 18984 13394 19012 16594
rect 19076 14890 19104 16782
rect 19064 14884 19116 14890
rect 19064 14826 19116 14832
rect 19076 14278 19104 14826
rect 19064 14272 19116 14278
rect 19064 14214 19116 14220
rect 18972 13388 19024 13394
rect 18972 13330 19024 13336
rect 18788 13320 18840 13326
rect 18788 13262 18840 13268
rect 18800 11014 18828 13262
rect 18970 13016 19026 13025
rect 18970 12951 19026 12960
rect 18984 12850 19012 12951
rect 19062 12880 19118 12889
rect 18972 12844 19024 12850
rect 19062 12815 19118 12824
rect 18972 12786 19024 12792
rect 18880 12776 18932 12782
rect 18880 12718 18932 12724
rect 18892 12594 18920 12718
rect 19076 12714 19104 12815
rect 19064 12708 19116 12714
rect 19064 12650 19116 12656
rect 18892 12566 19012 12594
rect 18880 12232 18932 12238
rect 18880 12174 18932 12180
rect 18892 12073 18920 12174
rect 18878 12064 18934 12073
rect 18878 11999 18934 12008
rect 18984 11642 19012 12566
rect 19064 12436 19116 12442
rect 19064 12378 19116 12384
rect 19076 11694 19104 12378
rect 18892 11614 19012 11642
rect 19064 11688 19116 11694
rect 19064 11630 19116 11636
rect 18892 11393 18920 11614
rect 18972 11552 19024 11558
rect 18972 11494 19024 11500
rect 18878 11384 18934 11393
rect 18878 11319 18934 11328
rect 18880 11212 18932 11218
rect 18880 11154 18932 11160
rect 18788 11008 18840 11014
rect 18788 10950 18840 10956
rect 18892 10810 18920 11154
rect 18880 10804 18932 10810
rect 18880 10746 18932 10752
rect 18788 10532 18840 10538
rect 18788 10474 18840 10480
rect 18696 9920 18748 9926
rect 18696 9862 18748 9868
rect 18800 9586 18828 10474
rect 18892 10130 18920 10746
rect 18880 10124 18932 10130
rect 18880 10066 18932 10072
rect 18880 9988 18932 9994
rect 18880 9930 18932 9936
rect 18788 9580 18840 9586
rect 18788 9522 18840 9528
rect 18892 9466 18920 9930
rect 18708 9438 18920 9466
rect 18604 8968 18656 8974
rect 18604 8910 18656 8916
rect 18512 7948 18564 7954
rect 18512 7890 18564 7896
rect 18524 7818 18552 7890
rect 18512 7812 18564 7818
rect 18512 7754 18564 7760
rect 18524 7721 18552 7754
rect 18510 7712 18566 7721
rect 18510 7647 18566 7656
rect 18616 7342 18644 8910
rect 18708 7993 18736 9438
rect 18788 9376 18840 9382
rect 18788 9318 18840 9324
rect 18694 7984 18750 7993
rect 18694 7919 18750 7928
rect 18800 7750 18828 9318
rect 18880 9104 18932 9110
rect 18880 9046 18932 9052
rect 18892 8634 18920 9046
rect 18880 8628 18932 8634
rect 18880 8570 18932 8576
rect 18892 8362 18920 8570
rect 18880 8356 18932 8362
rect 18880 8298 18932 8304
rect 18878 7984 18934 7993
rect 18878 7919 18880 7928
rect 18932 7919 18934 7928
rect 18880 7890 18932 7896
rect 18878 7848 18934 7857
rect 18878 7783 18934 7792
rect 18892 7750 18920 7783
rect 18788 7744 18840 7750
rect 18788 7686 18840 7692
rect 18880 7744 18932 7750
rect 18880 7686 18932 7692
rect 18604 7336 18656 7342
rect 18604 7278 18656 7284
rect 18604 6792 18656 6798
rect 18604 6734 18656 6740
rect 18616 6118 18644 6734
rect 18788 6656 18840 6662
rect 18788 6598 18840 6604
rect 18696 6384 18748 6390
rect 18696 6326 18748 6332
rect 17960 6112 18012 6118
rect 18420 6112 18472 6118
rect 17960 6054 18012 6060
rect 18050 6080 18106 6089
rect 17866 5808 17922 5817
rect 17866 5743 17922 5752
rect 17776 5704 17828 5710
rect 17776 5646 17828 5652
rect 17684 5364 17736 5370
rect 17684 5306 17736 5312
rect 17592 5296 17644 5302
rect 17592 5238 17644 5244
rect 17500 5160 17552 5166
rect 17500 5102 17552 5108
rect 17408 4548 17460 4554
rect 17408 4490 17460 4496
rect 17316 3936 17368 3942
rect 17316 3878 17368 3884
rect 17132 3664 17184 3670
rect 17132 3606 17184 3612
rect 17420 3466 17448 4490
rect 17500 4072 17552 4078
rect 17500 4014 17552 4020
rect 17512 3534 17540 4014
rect 17604 3602 17632 5238
rect 17696 4758 17724 5306
rect 17880 5250 17908 5743
rect 17788 5222 17908 5250
rect 17684 4752 17736 4758
rect 17684 4694 17736 4700
rect 17788 4078 17816 5222
rect 17868 5160 17920 5166
rect 17868 5102 17920 5108
rect 17880 4214 17908 5102
rect 17972 4570 18000 6054
rect 18420 6054 18472 6060
rect 18604 6112 18656 6118
rect 18604 6054 18656 6060
rect 18050 6015 18106 6024
rect 18064 5370 18092 6015
rect 18328 5704 18380 5710
rect 18328 5646 18380 5652
rect 18052 5364 18104 5370
rect 18052 5306 18104 5312
rect 18144 5364 18196 5370
rect 18144 5306 18196 5312
rect 18156 5273 18184 5306
rect 18142 5264 18198 5273
rect 18340 5234 18368 5646
rect 18512 5568 18564 5574
rect 18512 5510 18564 5516
rect 18524 5234 18552 5510
rect 18142 5199 18198 5208
rect 18328 5228 18380 5234
rect 18328 5170 18380 5176
rect 18512 5228 18564 5234
rect 18512 5170 18564 5176
rect 18340 4758 18368 5170
rect 18420 5024 18472 5030
rect 18420 4966 18472 4972
rect 18432 4826 18460 4966
rect 18420 4820 18472 4826
rect 18420 4762 18472 4768
rect 18328 4752 18380 4758
rect 18328 4694 18380 4700
rect 18144 4684 18196 4690
rect 18144 4626 18196 4632
rect 17972 4542 18092 4570
rect 17960 4480 18012 4486
rect 17960 4422 18012 4428
rect 17868 4208 17920 4214
rect 17868 4150 17920 4156
rect 17776 4072 17828 4078
rect 17776 4014 17828 4020
rect 17972 4010 18000 4422
rect 17960 4004 18012 4010
rect 17960 3946 18012 3952
rect 17592 3596 17644 3602
rect 17592 3538 17644 3544
rect 17776 3596 17828 3602
rect 17776 3538 17828 3544
rect 17500 3528 17552 3534
rect 17500 3470 17552 3476
rect 17408 3460 17460 3466
rect 17408 3402 17460 3408
rect 17420 2990 17448 3402
rect 17512 3126 17540 3470
rect 17682 3224 17738 3233
rect 17682 3159 17738 3168
rect 17500 3120 17552 3126
rect 17500 3062 17552 3068
rect 17408 2984 17460 2990
rect 17408 2926 17460 2932
rect 17040 2916 17092 2922
rect 17040 2858 17092 2864
rect 17696 2854 17724 3159
rect 17684 2848 17736 2854
rect 17684 2790 17736 2796
rect 17788 2650 17816 3538
rect 18064 3126 18092 4542
rect 18156 3194 18184 4626
rect 18340 4622 18368 4694
rect 18328 4616 18380 4622
rect 18328 4558 18380 4564
rect 18616 4078 18644 6054
rect 18708 5817 18736 6326
rect 18694 5808 18750 5817
rect 18694 5743 18696 5752
rect 18748 5743 18750 5752
rect 18696 5714 18748 5720
rect 18696 5160 18748 5166
rect 18694 5128 18696 5137
rect 18748 5128 18750 5137
rect 18694 5063 18750 5072
rect 18696 4480 18748 4486
rect 18694 4448 18696 4457
rect 18748 4448 18750 4457
rect 18694 4383 18750 4392
rect 18604 4072 18656 4078
rect 18604 4014 18656 4020
rect 18144 3188 18196 3194
rect 18144 3130 18196 3136
rect 18052 3120 18104 3126
rect 18052 3062 18104 3068
rect 17776 2644 17828 2650
rect 17776 2586 17828 2592
rect 18156 2582 18184 3130
rect 18800 2990 18828 6598
rect 18880 6112 18932 6118
rect 18880 6054 18932 6060
rect 18892 5098 18920 6054
rect 18880 5092 18932 5098
rect 18880 5034 18932 5040
rect 18984 4842 19012 11494
rect 19064 11008 19116 11014
rect 19064 10950 19116 10956
rect 19076 9994 19104 10950
rect 19064 9988 19116 9994
rect 19064 9930 19116 9936
rect 19168 9738 19196 17478
rect 19352 17202 19380 17818
rect 19536 17649 19564 18294
rect 19522 17640 19578 17649
rect 19522 17575 19578 17584
rect 19449 17436 19745 17456
rect 19505 17434 19529 17436
rect 19585 17434 19609 17436
rect 19665 17434 19689 17436
rect 19527 17382 19529 17434
rect 19591 17382 19603 17434
rect 19665 17382 19667 17434
rect 19505 17380 19529 17382
rect 19585 17380 19609 17382
rect 19665 17380 19689 17382
rect 19449 17360 19745 17380
rect 19340 17196 19392 17202
rect 19340 17138 19392 17144
rect 19246 17096 19302 17105
rect 19246 17031 19302 17040
rect 19260 16998 19288 17031
rect 19248 16992 19300 16998
rect 19248 16934 19300 16940
rect 19449 16348 19745 16368
rect 19505 16346 19529 16348
rect 19585 16346 19609 16348
rect 19665 16346 19689 16348
rect 19527 16294 19529 16346
rect 19591 16294 19603 16346
rect 19665 16294 19667 16346
rect 19505 16292 19529 16294
rect 19585 16292 19609 16294
rect 19665 16292 19689 16294
rect 19246 16280 19302 16289
rect 19449 16272 19745 16292
rect 19246 16215 19302 16224
rect 19260 14482 19288 16215
rect 19340 15632 19392 15638
rect 19340 15574 19392 15580
rect 19432 15632 19484 15638
rect 19432 15574 19484 15580
rect 19352 15473 19380 15574
rect 19338 15464 19394 15473
rect 19338 15399 19394 15408
rect 19444 15348 19472 15574
rect 19352 15320 19472 15348
rect 19352 15162 19380 15320
rect 19449 15260 19745 15280
rect 19505 15258 19529 15260
rect 19585 15258 19609 15260
rect 19665 15258 19689 15260
rect 19527 15206 19529 15258
rect 19591 15206 19603 15258
rect 19665 15206 19667 15258
rect 19505 15204 19529 15206
rect 19585 15204 19609 15206
rect 19665 15204 19689 15206
rect 19449 15184 19745 15204
rect 19340 15156 19392 15162
rect 19340 15098 19392 15104
rect 19432 15020 19484 15026
rect 19432 14962 19484 14968
rect 19338 14784 19394 14793
rect 19338 14719 19394 14728
rect 19248 14476 19300 14482
rect 19248 14418 19300 14424
rect 19260 14006 19288 14418
rect 19352 14074 19380 14719
rect 19444 14618 19472 14962
rect 19432 14612 19484 14618
rect 19432 14554 19484 14560
rect 19430 14512 19486 14521
rect 19430 14447 19432 14456
rect 19484 14447 19486 14456
rect 19432 14418 19484 14424
rect 19449 14172 19745 14192
rect 19505 14170 19529 14172
rect 19585 14170 19609 14172
rect 19665 14170 19689 14172
rect 19527 14118 19529 14170
rect 19591 14118 19603 14170
rect 19665 14118 19667 14170
rect 19505 14116 19529 14118
rect 19585 14116 19609 14118
rect 19665 14116 19689 14118
rect 19449 14096 19745 14116
rect 19340 14068 19392 14074
rect 19340 14010 19392 14016
rect 19248 14000 19300 14006
rect 19248 13942 19300 13948
rect 19616 13796 19668 13802
rect 19616 13738 19668 13744
rect 19340 13728 19392 13734
rect 19340 13670 19392 13676
rect 19352 13190 19380 13670
rect 19628 13569 19656 13738
rect 19614 13560 19670 13569
rect 19812 13530 19840 18770
rect 19904 17785 19932 18770
rect 19996 18136 20024 18906
rect 20088 18465 20116 19094
rect 20168 18964 20220 18970
rect 20168 18906 20220 18912
rect 20180 18737 20208 18906
rect 20166 18728 20222 18737
rect 20166 18663 20222 18672
rect 20168 18624 20220 18630
rect 20168 18566 20220 18572
rect 20074 18456 20130 18465
rect 20074 18391 20130 18400
rect 20180 18329 20208 18566
rect 20166 18320 20222 18329
rect 20166 18255 20222 18264
rect 20076 18216 20128 18222
rect 20076 18158 20128 18164
rect 19987 18108 20024 18136
rect 19987 18068 20015 18108
rect 19987 18040 20024 18068
rect 19890 17776 19946 17785
rect 19890 17711 19946 17720
rect 19890 17368 19946 17377
rect 19890 17303 19946 17312
rect 19904 17134 19932 17303
rect 19892 17128 19944 17134
rect 19892 17070 19944 17076
rect 19892 16992 19944 16998
rect 19892 16934 19944 16940
rect 19904 15745 19932 16934
rect 19890 15736 19946 15745
rect 19890 15671 19946 15680
rect 19904 15366 19932 15671
rect 19996 15586 20024 18040
rect 20088 16726 20116 18158
rect 20272 17882 20300 20590
rect 20352 20538 20404 20544
rect 20352 19168 20404 19174
rect 20352 19110 20404 19116
rect 20364 18426 20392 19110
rect 20352 18420 20404 18426
rect 20352 18362 20404 18368
rect 20352 18148 20404 18154
rect 20352 18090 20404 18096
rect 20260 17876 20312 17882
rect 20260 17818 20312 17824
rect 20168 17536 20220 17542
rect 20168 17478 20220 17484
rect 20180 17202 20208 17478
rect 20258 17232 20314 17241
rect 20168 17196 20220 17202
rect 20258 17167 20260 17176
rect 20168 17138 20220 17144
rect 20312 17167 20314 17176
rect 20260 17138 20312 17144
rect 20076 16720 20128 16726
rect 20076 16662 20128 16668
rect 20168 16584 20220 16590
rect 20168 16526 20220 16532
rect 20180 16250 20208 16526
rect 20260 16516 20312 16522
rect 20260 16458 20312 16464
rect 20168 16244 20220 16250
rect 20168 16186 20220 16192
rect 20272 16114 20300 16458
rect 20260 16108 20312 16114
rect 20260 16050 20312 16056
rect 19996 15558 20208 15586
rect 19984 15496 20036 15502
rect 19984 15438 20036 15444
rect 19892 15360 19944 15366
rect 19892 15302 19944 15308
rect 19892 14884 19944 14890
rect 19892 14826 19944 14832
rect 19904 14414 19932 14826
rect 19892 14408 19944 14414
rect 19892 14350 19944 14356
rect 19614 13495 19670 13504
rect 19800 13524 19852 13530
rect 19800 13466 19852 13472
rect 19340 13184 19392 13190
rect 19340 13126 19392 13132
rect 19800 13184 19852 13190
rect 19904 13161 19932 14350
rect 19800 13126 19852 13132
rect 19890 13152 19946 13161
rect 19449 13084 19745 13104
rect 19505 13082 19529 13084
rect 19585 13082 19609 13084
rect 19665 13082 19689 13084
rect 19527 13030 19529 13082
rect 19591 13030 19603 13082
rect 19665 13030 19667 13082
rect 19505 13028 19529 13030
rect 19585 13028 19609 13030
rect 19665 13028 19689 13030
rect 19449 13008 19745 13028
rect 19812 12986 19840 13126
rect 19890 13087 19946 13096
rect 19800 12980 19852 12986
rect 19800 12922 19852 12928
rect 19800 12844 19852 12850
rect 19904 12832 19932 13087
rect 19852 12804 19932 12832
rect 19800 12786 19852 12792
rect 19996 12730 20024 15438
rect 20076 15360 20128 15366
rect 20076 15302 20128 15308
rect 20088 14929 20116 15302
rect 20074 14920 20130 14929
rect 20074 14855 20130 14864
rect 20076 14544 20128 14550
rect 20076 14486 20128 14492
rect 20088 13734 20116 14486
rect 20180 13938 20208 15558
rect 20260 15564 20312 15570
rect 20260 15506 20312 15512
rect 20168 13932 20220 13938
rect 20168 13874 20220 13880
rect 20076 13728 20128 13734
rect 20076 13670 20128 13676
rect 20180 12986 20208 13874
rect 20168 12980 20220 12986
rect 19260 12702 19380 12730
rect 19260 11665 19288 12702
rect 19352 12481 19380 12702
rect 19720 12702 20024 12730
rect 20088 12940 20168 12968
rect 19338 12472 19394 12481
rect 19338 12407 19394 12416
rect 19338 12336 19394 12345
rect 19338 12271 19394 12280
rect 19616 12300 19668 12306
rect 19246 11656 19302 11665
rect 19352 11626 19380 12271
rect 19720 12288 19748 12702
rect 20088 12594 20116 12940
rect 20168 12922 20220 12928
rect 20168 12776 20220 12782
rect 20168 12718 20220 12724
rect 19904 12566 20116 12594
rect 19668 12260 19748 12288
rect 19800 12300 19852 12306
rect 19616 12242 19668 12248
rect 19800 12242 19852 12248
rect 19628 12209 19656 12242
rect 19614 12200 19670 12209
rect 19614 12135 19670 12144
rect 19449 11996 19745 12016
rect 19505 11994 19529 11996
rect 19585 11994 19609 11996
rect 19665 11994 19689 11996
rect 19527 11942 19529 11994
rect 19591 11942 19603 11994
rect 19665 11942 19667 11994
rect 19505 11940 19529 11942
rect 19585 11940 19609 11942
rect 19665 11940 19689 11942
rect 19449 11920 19745 11940
rect 19812 11898 19840 12242
rect 19800 11892 19852 11898
rect 19800 11834 19852 11840
rect 19904 11762 19932 12566
rect 20074 12472 20130 12481
rect 20074 12407 20130 12416
rect 19892 11756 19944 11762
rect 19812 11716 19892 11744
rect 19246 11591 19302 11600
rect 19340 11620 19392 11626
rect 19340 11562 19392 11568
rect 19616 11552 19668 11558
rect 19338 11520 19394 11529
rect 19616 11494 19668 11500
rect 19338 11455 19394 11464
rect 19352 11354 19380 11455
rect 19340 11348 19392 11354
rect 19340 11290 19392 11296
rect 19628 11286 19656 11494
rect 19616 11280 19668 11286
rect 19616 11222 19668 11228
rect 19449 10908 19745 10928
rect 19505 10906 19529 10908
rect 19585 10906 19609 10908
rect 19665 10906 19689 10908
rect 19527 10854 19529 10906
rect 19591 10854 19603 10906
rect 19665 10854 19667 10906
rect 19505 10852 19529 10854
rect 19585 10852 19609 10854
rect 19665 10852 19689 10854
rect 19246 10840 19302 10849
rect 19449 10832 19745 10852
rect 19246 10775 19248 10784
rect 19300 10775 19302 10784
rect 19248 10746 19300 10752
rect 19616 10668 19668 10674
rect 19616 10610 19668 10616
rect 19628 10577 19656 10610
rect 19708 10600 19760 10606
rect 19614 10568 19670 10577
rect 19812 10588 19840 11716
rect 19892 11698 19944 11704
rect 19984 11076 20036 11082
rect 19984 11018 20036 11024
rect 19760 10560 19840 10588
rect 19708 10542 19760 10548
rect 19614 10503 19670 10512
rect 19248 10464 19300 10470
rect 19248 10406 19300 10412
rect 19076 9710 19196 9738
rect 19076 8129 19104 9710
rect 19260 9518 19288 10406
rect 19340 10260 19392 10266
rect 19340 10202 19392 10208
rect 19352 10169 19380 10202
rect 19338 10160 19394 10169
rect 19338 10095 19394 10104
rect 19432 10124 19484 10130
rect 19432 10066 19484 10072
rect 19444 10010 19472 10066
rect 19435 9982 19472 10010
rect 19435 9976 19463 9982
rect 19352 9948 19463 9976
rect 19248 9512 19300 9518
rect 19248 9454 19300 9460
rect 19260 8634 19288 9454
rect 19352 9178 19380 9948
rect 19449 9820 19745 9840
rect 19505 9818 19529 9820
rect 19585 9818 19609 9820
rect 19665 9818 19689 9820
rect 19527 9766 19529 9818
rect 19591 9766 19603 9818
rect 19665 9766 19667 9818
rect 19505 9764 19529 9766
rect 19585 9764 19609 9766
rect 19665 9764 19689 9766
rect 19449 9744 19745 9764
rect 19432 9580 19484 9586
rect 19432 9522 19484 9528
rect 19340 9172 19392 9178
rect 19340 9114 19392 9120
rect 19444 8820 19472 9522
rect 19352 8792 19472 8820
rect 19156 8628 19208 8634
rect 19156 8570 19208 8576
rect 19248 8628 19300 8634
rect 19352 8616 19380 8792
rect 19449 8732 19745 8752
rect 19505 8730 19529 8732
rect 19585 8730 19609 8732
rect 19665 8730 19689 8732
rect 19527 8678 19529 8730
rect 19591 8678 19603 8730
rect 19665 8678 19667 8730
rect 19505 8676 19529 8678
rect 19585 8676 19609 8678
rect 19665 8676 19689 8678
rect 19449 8656 19745 8676
rect 19352 8588 19656 8616
rect 19248 8570 19300 8576
rect 19168 8498 19196 8570
rect 19156 8492 19208 8498
rect 19432 8492 19484 8498
rect 19156 8434 19208 8440
rect 19260 8452 19432 8480
rect 19062 8120 19118 8129
rect 19062 8055 19118 8064
rect 19064 6724 19116 6730
rect 19064 6666 19116 6672
rect 19076 6322 19104 6666
rect 19064 6316 19116 6322
rect 19064 6258 19116 6264
rect 19260 6186 19288 8452
rect 19432 8434 19484 8440
rect 19338 8392 19394 8401
rect 19522 8392 19578 8401
rect 19338 8327 19394 8336
rect 19444 8350 19522 8378
rect 19352 8129 19380 8327
rect 19338 8120 19394 8129
rect 19338 8055 19394 8064
rect 19444 7834 19472 8350
rect 19522 8327 19578 8336
rect 19352 7806 19472 7834
rect 19524 7880 19576 7886
rect 19628 7868 19656 8588
rect 19708 8492 19760 8498
rect 19708 8434 19760 8440
rect 19720 7993 19748 8434
rect 19812 8430 19840 10560
rect 19892 10600 19944 10606
rect 19892 10542 19944 10548
rect 19904 9382 19932 10542
rect 19892 9376 19944 9382
rect 19892 9318 19944 9324
rect 19904 8566 19932 9318
rect 19892 8560 19944 8566
rect 19892 8502 19944 8508
rect 19800 8424 19852 8430
rect 19800 8366 19852 8372
rect 19706 7984 19762 7993
rect 19706 7919 19762 7928
rect 19576 7840 19656 7868
rect 19812 7857 19840 8366
rect 19890 8256 19946 8265
rect 19890 8191 19946 8200
rect 19798 7848 19854 7857
rect 19524 7822 19576 7828
rect 19352 7290 19380 7806
rect 19798 7783 19854 7792
rect 19449 7644 19745 7664
rect 19505 7642 19529 7644
rect 19585 7642 19609 7644
rect 19665 7642 19689 7644
rect 19527 7590 19529 7642
rect 19591 7590 19603 7642
rect 19665 7590 19667 7642
rect 19505 7588 19529 7590
rect 19585 7588 19609 7590
rect 19665 7588 19689 7590
rect 19449 7568 19745 7588
rect 19904 7478 19932 8191
rect 19892 7472 19944 7478
rect 19892 7414 19944 7420
rect 19352 7262 19472 7290
rect 19340 7200 19392 7206
rect 19340 7142 19392 7148
rect 19352 7002 19380 7142
rect 19340 6996 19392 7002
rect 19340 6938 19392 6944
rect 19444 6746 19472 7262
rect 19800 7200 19852 7206
rect 19800 7142 19852 7148
rect 19352 6718 19472 6746
rect 19064 6180 19116 6186
rect 19064 6122 19116 6128
rect 19248 6180 19300 6186
rect 19248 6122 19300 6128
rect 19076 5778 19104 6122
rect 19260 5914 19288 6122
rect 19248 5908 19300 5914
rect 19248 5850 19300 5856
rect 19064 5772 19116 5778
rect 19064 5714 19116 5720
rect 19076 5098 19104 5714
rect 19246 5672 19302 5681
rect 19246 5607 19302 5616
rect 19064 5092 19116 5098
rect 19064 5034 19116 5040
rect 18984 4814 19104 4842
rect 18972 4752 19024 4758
rect 18972 4694 19024 4700
rect 18880 4004 18932 4010
rect 18880 3946 18932 3952
rect 18892 3738 18920 3946
rect 18880 3732 18932 3738
rect 18880 3674 18932 3680
rect 18788 2984 18840 2990
rect 18788 2926 18840 2932
rect 18892 2650 18920 3674
rect 18880 2644 18932 2650
rect 18880 2586 18932 2592
rect 18144 2576 18196 2582
rect 18144 2518 18196 2524
rect 18984 2446 19012 4694
rect 19076 4282 19104 4814
rect 19064 4276 19116 4282
rect 19064 4218 19116 4224
rect 19260 4078 19288 5607
rect 19352 4185 19380 6718
rect 19449 6556 19745 6576
rect 19505 6554 19529 6556
rect 19585 6554 19609 6556
rect 19665 6554 19689 6556
rect 19527 6502 19529 6554
rect 19591 6502 19603 6554
rect 19665 6502 19667 6554
rect 19505 6500 19529 6502
rect 19585 6500 19609 6502
rect 19665 6500 19689 6502
rect 19449 6480 19745 6500
rect 19449 5468 19745 5488
rect 19505 5466 19529 5468
rect 19585 5466 19609 5468
rect 19665 5466 19689 5468
rect 19527 5414 19529 5466
rect 19591 5414 19603 5466
rect 19665 5414 19667 5466
rect 19505 5412 19529 5414
rect 19585 5412 19609 5414
rect 19665 5412 19689 5414
rect 19449 5392 19745 5412
rect 19812 5370 19840 7142
rect 19904 6361 19932 7414
rect 19890 6352 19946 6361
rect 19890 6287 19946 6296
rect 19800 5364 19852 5370
rect 19800 5306 19852 5312
rect 19614 5264 19670 5273
rect 19614 5199 19616 5208
rect 19668 5199 19670 5208
rect 19616 5170 19668 5176
rect 19616 5024 19668 5030
rect 19616 4966 19668 4972
rect 19800 5024 19852 5030
rect 19800 4966 19852 4972
rect 19628 4826 19656 4966
rect 19616 4820 19668 4826
rect 19616 4762 19668 4768
rect 19449 4380 19745 4400
rect 19505 4378 19529 4380
rect 19585 4378 19609 4380
rect 19665 4378 19689 4380
rect 19527 4326 19529 4378
rect 19591 4326 19603 4378
rect 19665 4326 19667 4378
rect 19505 4324 19529 4326
rect 19585 4324 19609 4326
rect 19665 4324 19689 4326
rect 19449 4304 19745 4324
rect 19812 4282 19840 4966
rect 19800 4276 19852 4282
rect 19800 4218 19852 4224
rect 19338 4176 19394 4185
rect 19338 4111 19394 4120
rect 19248 4072 19300 4078
rect 19248 4014 19300 4020
rect 19064 3936 19116 3942
rect 19064 3878 19116 3884
rect 19432 3936 19484 3942
rect 19432 3878 19484 3884
rect 19076 3602 19104 3878
rect 19444 3670 19472 3878
rect 19432 3664 19484 3670
rect 19432 3606 19484 3612
rect 19064 3596 19116 3602
rect 19064 3538 19116 3544
rect 19076 2922 19104 3538
rect 19449 3292 19745 3312
rect 19505 3290 19529 3292
rect 19585 3290 19609 3292
rect 19665 3290 19689 3292
rect 19527 3238 19529 3290
rect 19591 3238 19603 3290
rect 19665 3238 19667 3290
rect 19505 3236 19529 3238
rect 19585 3236 19609 3238
rect 19665 3236 19689 3238
rect 19449 3216 19745 3236
rect 19064 2916 19116 2922
rect 19064 2858 19116 2864
rect 19076 2514 19104 2858
rect 19064 2508 19116 2514
rect 19064 2450 19116 2456
rect 18972 2440 19024 2446
rect 18972 2382 19024 2388
rect 19890 2272 19946 2281
rect 19449 2204 19745 2224
rect 19890 2207 19946 2216
rect 19505 2202 19529 2204
rect 19585 2202 19609 2204
rect 19665 2202 19689 2204
rect 19527 2150 19529 2202
rect 19591 2150 19603 2202
rect 19665 2150 19667 2202
rect 19505 2148 19529 2150
rect 19585 2148 19609 2150
rect 19665 2148 19689 2150
rect 19449 2128 19745 2148
rect 19904 1970 19932 2207
rect 19996 2106 20024 11018
rect 20088 7954 20116 12407
rect 20180 12306 20208 12718
rect 20272 12617 20300 15506
rect 20258 12608 20314 12617
rect 20258 12543 20314 12552
rect 20168 12300 20220 12306
rect 20168 12242 20220 12248
rect 20166 12200 20222 12209
rect 20166 12135 20222 12144
rect 20180 11354 20208 12135
rect 20260 12096 20312 12102
rect 20260 12038 20312 12044
rect 20168 11348 20220 11354
rect 20168 11290 20220 11296
rect 20272 11150 20300 12038
rect 20364 11937 20392 18090
rect 20456 15434 20484 21927
rect 20628 21888 20680 21894
rect 20628 21830 20680 21836
rect 20640 21622 20668 21830
rect 20536 21616 20588 21622
rect 20536 21558 20588 21564
rect 20628 21616 20680 21622
rect 20628 21558 20680 21564
rect 20548 19961 20576 21558
rect 20628 21344 20680 21350
rect 20628 21286 20680 21292
rect 20640 21146 20668 21286
rect 20628 21140 20680 21146
rect 20628 21082 20680 21088
rect 20626 20632 20682 20641
rect 20626 20567 20682 20576
rect 20534 19952 20590 19961
rect 20534 19887 20590 19896
rect 20536 19848 20588 19854
rect 20536 19790 20588 19796
rect 20548 18902 20576 19790
rect 20536 18896 20588 18902
rect 20536 18838 20588 18844
rect 20548 17678 20576 18838
rect 20536 17672 20588 17678
rect 20536 17614 20588 17620
rect 20536 15904 20588 15910
rect 20536 15846 20588 15852
rect 20444 15428 20496 15434
rect 20444 15370 20496 15376
rect 20548 15178 20576 15846
rect 20640 15434 20668 20567
rect 20720 20460 20772 20466
rect 20720 20402 20772 20408
rect 20732 20262 20760 20402
rect 20720 20256 20772 20262
rect 20720 20198 20772 20204
rect 20824 20058 20852 23600
rect 21272 21480 21324 21486
rect 21272 21422 21324 21428
rect 21180 21344 21232 21350
rect 21180 21286 21232 21292
rect 21192 20913 21220 21286
rect 21178 20904 21234 20913
rect 21088 20868 21140 20874
rect 21178 20839 21234 20848
rect 21088 20810 21140 20816
rect 20904 20800 20956 20806
rect 20904 20742 20956 20748
rect 20916 20534 20944 20742
rect 20904 20528 20956 20534
rect 20904 20470 20956 20476
rect 20812 20052 20864 20058
rect 20812 19994 20864 20000
rect 20916 19281 20944 20470
rect 21100 20262 21128 20810
rect 21180 20800 21232 20806
rect 21180 20742 21232 20748
rect 21088 20256 21140 20262
rect 21088 20198 21140 20204
rect 21100 19990 21128 20198
rect 21088 19984 21140 19990
rect 21088 19926 21140 19932
rect 20996 19848 21048 19854
rect 20996 19790 21048 19796
rect 20902 19272 20958 19281
rect 20902 19207 20958 19216
rect 20904 19168 20956 19174
rect 21008 19156 21036 19790
rect 20956 19128 21036 19156
rect 20904 19110 20956 19116
rect 20812 18760 20864 18766
rect 20718 18728 20774 18737
rect 20812 18702 20864 18708
rect 20718 18663 20774 18672
rect 20732 17134 20760 18663
rect 20720 17128 20772 17134
rect 20720 17070 20772 17076
rect 20824 16232 20852 18702
rect 20916 18222 20944 19110
rect 21192 18970 21220 20742
rect 21180 18964 21232 18970
rect 21180 18906 21232 18912
rect 21180 18828 21232 18834
rect 21180 18770 21232 18776
rect 20996 18692 21048 18698
rect 20996 18634 21048 18640
rect 20904 18216 20956 18222
rect 20904 18158 20956 18164
rect 20916 17678 20944 18158
rect 21008 18057 21036 18634
rect 20994 18048 21050 18057
rect 20994 17983 21050 17992
rect 20996 17808 21048 17814
rect 20996 17750 21048 17756
rect 21088 17808 21140 17814
rect 21088 17750 21140 17756
rect 20904 17672 20956 17678
rect 20904 17614 20956 17620
rect 20916 17202 20944 17614
rect 20904 17196 20956 17202
rect 20904 17138 20956 17144
rect 21008 16794 21036 17750
rect 20904 16788 20956 16794
rect 20904 16730 20956 16736
rect 20996 16788 21048 16794
rect 20996 16730 21048 16736
rect 20916 16697 20944 16730
rect 20902 16688 20958 16697
rect 20902 16623 20958 16632
rect 20732 16204 20852 16232
rect 20732 15638 20760 16204
rect 20812 16108 20864 16114
rect 20812 16050 20864 16056
rect 20720 15632 20772 15638
rect 20720 15574 20772 15580
rect 20628 15428 20680 15434
rect 20628 15370 20680 15376
rect 20548 15150 20760 15178
rect 20626 15056 20682 15065
rect 20626 14991 20682 15000
rect 20444 14816 20496 14822
rect 20444 14758 20496 14764
rect 20456 14657 20484 14758
rect 20442 14648 20498 14657
rect 20442 14583 20498 14592
rect 20640 14113 20668 14991
rect 20732 14482 20760 15150
rect 20720 14476 20772 14482
rect 20720 14418 20772 14424
rect 20626 14104 20682 14113
rect 20626 14039 20682 14048
rect 20720 13932 20772 13938
rect 20720 13874 20772 13880
rect 20444 13864 20496 13870
rect 20444 13806 20496 13812
rect 20350 11928 20406 11937
rect 20350 11863 20406 11872
rect 20352 11756 20404 11762
rect 20352 11698 20404 11704
rect 20260 11144 20312 11150
rect 20260 11086 20312 11092
rect 20260 11008 20312 11014
rect 20260 10950 20312 10956
rect 20272 10130 20300 10950
rect 20260 10124 20312 10130
rect 20260 10066 20312 10072
rect 20260 9580 20312 9586
rect 20260 9522 20312 9528
rect 20272 8838 20300 9522
rect 20364 9217 20392 11698
rect 20456 11354 20484 13806
rect 20628 13728 20680 13734
rect 20628 13670 20680 13676
rect 20536 13184 20588 13190
rect 20536 13126 20588 13132
rect 20548 12782 20576 13126
rect 20536 12776 20588 12782
rect 20536 12718 20588 12724
rect 20640 12594 20668 13670
rect 20732 12889 20760 13874
rect 20718 12880 20774 12889
rect 20718 12815 20774 12824
rect 20548 12566 20668 12594
rect 20548 11558 20576 12566
rect 20626 12472 20682 12481
rect 20824 12442 20852 16050
rect 20904 15972 20956 15978
rect 20904 15914 20956 15920
rect 20916 14906 20944 15914
rect 20996 15904 21048 15910
rect 20996 15846 21048 15852
rect 21008 15706 21036 15846
rect 20996 15700 21048 15706
rect 20996 15642 21048 15648
rect 20916 14878 21036 14906
rect 20904 14816 20956 14822
rect 20904 14758 20956 14764
rect 20916 13841 20944 14758
rect 21008 14346 21036 14878
rect 20996 14340 21048 14346
rect 20996 14282 21048 14288
rect 20902 13832 20958 13841
rect 20902 13767 20958 13776
rect 20902 13424 20958 13433
rect 20902 13359 20904 13368
rect 20956 13359 20958 13368
rect 20904 13330 20956 13336
rect 20996 12980 21048 12986
rect 20996 12922 21048 12928
rect 20626 12407 20682 12416
rect 20812 12436 20864 12442
rect 20640 11898 20668 12407
rect 20812 12378 20864 12384
rect 20904 12436 20956 12442
rect 20904 12378 20956 12384
rect 20628 11892 20680 11898
rect 20628 11834 20680 11840
rect 20536 11552 20588 11558
rect 20812 11552 20864 11558
rect 20536 11494 20588 11500
rect 20640 11500 20812 11506
rect 20640 11494 20864 11500
rect 20444 11348 20496 11354
rect 20444 11290 20496 11296
rect 20456 11082 20484 11290
rect 20444 11076 20496 11082
rect 20444 11018 20496 11024
rect 20548 10962 20576 11494
rect 20640 11478 20852 11494
rect 20640 11354 20668 11478
rect 20628 11348 20680 11354
rect 20628 11290 20680 11296
rect 20916 11234 20944 12378
rect 21008 12306 21036 12922
rect 20996 12300 21048 12306
rect 20996 12242 21048 12248
rect 20996 12096 21048 12102
rect 20996 12038 21048 12044
rect 20824 11206 20944 11234
rect 21008 11218 21036 12038
rect 20996 11212 21048 11218
rect 20628 11144 20680 11150
rect 20628 11086 20680 11092
rect 20456 10934 20576 10962
rect 20456 10470 20484 10934
rect 20534 10840 20590 10849
rect 20534 10775 20590 10784
rect 20444 10464 20496 10470
rect 20444 10406 20496 10412
rect 20444 10192 20496 10198
rect 20444 10134 20496 10140
rect 20456 9518 20484 10134
rect 20444 9512 20496 9518
rect 20444 9454 20496 9460
rect 20350 9208 20406 9217
rect 20350 9143 20406 9152
rect 20352 9036 20404 9042
rect 20352 8978 20404 8984
rect 20260 8832 20312 8838
rect 20260 8774 20312 8780
rect 20258 8664 20314 8673
rect 20258 8599 20314 8608
rect 20076 7948 20128 7954
rect 20076 7890 20128 7896
rect 20074 7168 20130 7177
rect 20074 7103 20130 7112
rect 20088 3641 20116 7103
rect 20272 6934 20300 8599
rect 20364 8498 20392 8978
rect 20352 8492 20404 8498
rect 20352 8434 20404 8440
rect 20364 7342 20392 8434
rect 20548 8344 20576 10775
rect 20640 9058 20668 11086
rect 20640 9030 20760 9058
rect 20628 8968 20680 8974
rect 20628 8910 20680 8916
rect 20640 8498 20668 8910
rect 20628 8492 20680 8498
rect 20628 8434 20680 8440
rect 20456 8316 20576 8344
rect 20352 7336 20404 7342
rect 20352 7278 20404 7284
rect 20260 6928 20312 6934
rect 20260 6870 20312 6876
rect 20168 6860 20220 6866
rect 20168 6802 20220 6808
rect 20180 5574 20208 6802
rect 20260 6792 20312 6798
rect 20260 6734 20312 6740
rect 20350 6760 20406 6769
rect 20168 5568 20220 5574
rect 20168 5510 20220 5516
rect 20168 4616 20220 4622
rect 20168 4558 20220 4564
rect 20074 3632 20130 3641
rect 20074 3567 20130 3576
rect 20180 3194 20208 4558
rect 20272 3398 20300 6734
rect 20350 6695 20406 6704
rect 20364 5409 20392 6695
rect 20456 6610 20484 8316
rect 20534 8256 20590 8265
rect 20534 8191 20590 8200
rect 20548 7410 20576 8191
rect 20640 8090 20668 8434
rect 20628 8084 20680 8090
rect 20628 8026 20680 8032
rect 20732 7970 20760 9030
rect 20640 7942 20760 7970
rect 20536 7404 20588 7410
rect 20536 7346 20588 7352
rect 20456 6582 20576 6610
rect 20444 6452 20496 6458
rect 20444 6394 20496 6400
rect 20456 5846 20484 6394
rect 20444 5840 20496 5846
rect 20444 5782 20496 5788
rect 20444 5636 20496 5642
rect 20444 5578 20496 5584
rect 20350 5400 20406 5409
rect 20350 5335 20406 5344
rect 20456 5250 20484 5578
rect 20364 5222 20484 5250
rect 20364 4554 20392 5222
rect 20352 4548 20404 4554
rect 20352 4490 20404 4496
rect 20364 4214 20392 4490
rect 20352 4208 20404 4214
rect 20352 4150 20404 4156
rect 20548 4078 20576 6582
rect 20640 5166 20668 7942
rect 20720 7880 20772 7886
rect 20720 7822 20772 7828
rect 20732 6662 20760 7822
rect 20720 6656 20772 6662
rect 20720 6598 20772 6604
rect 20824 5658 20852 11206
rect 20996 11154 21048 11160
rect 20904 11144 20956 11150
rect 20904 11086 20956 11092
rect 20916 10062 20944 11086
rect 20904 10056 20956 10062
rect 20904 9998 20956 10004
rect 20916 9586 20944 9998
rect 20904 9580 20956 9586
rect 20904 9522 20956 9528
rect 20916 7954 20944 9522
rect 20904 7948 20956 7954
rect 20904 7890 20956 7896
rect 21008 7886 21036 11154
rect 20996 7880 21048 7886
rect 20996 7822 21048 7828
rect 20902 7576 20958 7585
rect 20902 7511 20958 7520
rect 20916 7478 20944 7511
rect 20904 7472 20956 7478
rect 20904 7414 20956 7420
rect 20904 7336 20956 7342
rect 20904 7278 20956 7284
rect 20916 6798 20944 7278
rect 20904 6792 20956 6798
rect 20904 6734 20956 6740
rect 20916 6254 20944 6734
rect 20904 6248 20956 6254
rect 20904 6190 20956 6196
rect 20996 6112 21048 6118
rect 20996 6054 21048 6060
rect 20904 5772 20956 5778
rect 20904 5714 20956 5720
rect 20732 5630 20852 5658
rect 20628 5160 20680 5166
rect 20628 5102 20680 5108
rect 20732 4842 20760 5630
rect 20812 5568 20864 5574
rect 20812 5510 20864 5516
rect 20824 5234 20852 5510
rect 20916 5370 20944 5714
rect 20904 5364 20956 5370
rect 20904 5306 20956 5312
rect 20902 5264 20958 5273
rect 20812 5228 20864 5234
rect 20902 5199 20904 5208
rect 20812 5170 20864 5176
rect 20956 5199 20958 5208
rect 20904 5170 20956 5176
rect 21008 5166 21036 6054
rect 20996 5160 21048 5166
rect 20996 5102 21048 5108
rect 20904 5092 20956 5098
rect 20904 5034 20956 5040
rect 20640 4814 20760 4842
rect 20640 4486 20668 4814
rect 20720 4752 20772 4758
rect 20718 4720 20720 4729
rect 20772 4720 20774 4729
rect 20718 4655 20774 4664
rect 20812 4684 20864 4690
rect 20812 4626 20864 4632
rect 20628 4480 20680 4486
rect 20628 4422 20680 4428
rect 20536 4072 20588 4078
rect 20536 4014 20588 4020
rect 20444 3936 20496 3942
rect 20444 3878 20496 3884
rect 20456 3398 20484 3878
rect 20260 3392 20312 3398
rect 20260 3334 20312 3340
rect 20444 3392 20496 3398
rect 20444 3334 20496 3340
rect 20168 3188 20220 3194
rect 20168 3130 20220 3136
rect 20180 2582 20208 3130
rect 20456 2990 20484 3334
rect 20824 2990 20852 4626
rect 20916 4078 20944 5034
rect 20996 4616 21048 4622
rect 20996 4558 21048 4564
rect 21008 4078 21036 4558
rect 20904 4072 20956 4078
rect 20904 4014 20956 4020
rect 20996 4072 21048 4078
rect 20996 4014 21048 4020
rect 21008 3890 21036 4014
rect 20916 3862 21036 3890
rect 20916 3534 20944 3862
rect 20904 3528 20956 3534
rect 20904 3470 20956 3476
rect 20444 2984 20496 2990
rect 20444 2926 20496 2932
rect 20812 2984 20864 2990
rect 20812 2926 20864 2932
rect 20824 2650 20852 2926
rect 20916 2922 20944 3470
rect 20904 2916 20956 2922
rect 20904 2858 20956 2864
rect 20812 2644 20864 2650
rect 20812 2586 20864 2592
rect 20168 2576 20220 2582
rect 20168 2518 20220 2524
rect 20916 2514 20944 2858
rect 21100 2582 21128 17750
rect 21192 17134 21220 18770
rect 21180 17128 21232 17134
rect 21180 17070 21232 17076
rect 21180 16992 21232 16998
rect 21180 16934 21232 16940
rect 21192 12442 21220 16934
rect 21284 14362 21312 21422
rect 21364 20936 21416 20942
rect 21364 20878 21416 20884
rect 21376 20602 21404 20878
rect 21364 20596 21416 20602
rect 21364 20538 21416 20544
rect 21468 20058 21496 23600
rect 21640 22092 21692 22098
rect 21640 22034 21692 22040
rect 21652 21622 21680 22034
rect 21640 21616 21692 21622
rect 21640 21558 21692 21564
rect 22008 21548 22060 21554
rect 22008 21490 22060 21496
rect 21732 21344 21784 21350
rect 21732 21286 21784 21292
rect 21548 20256 21600 20262
rect 21548 20198 21600 20204
rect 21456 20052 21508 20058
rect 21456 19994 21508 20000
rect 21456 19916 21508 19922
rect 21456 19858 21508 19864
rect 21364 18624 21416 18630
rect 21364 18566 21416 18572
rect 21376 18057 21404 18566
rect 21362 18048 21418 18057
rect 21362 17983 21418 17992
rect 21468 17882 21496 19858
rect 21560 19689 21588 20198
rect 21546 19680 21602 19689
rect 21546 19615 21602 19624
rect 21640 19508 21692 19514
rect 21640 19450 21692 19456
rect 21652 19417 21680 19450
rect 21638 19408 21694 19417
rect 21638 19343 21694 19352
rect 21640 19236 21692 19242
rect 21640 19178 21692 19184
rect 21652 18086 21680 19178
rect 21744 18970 21772 21286
rect 21916 20324 21968 20330
rect 21916 20266 21968 20272
rect 21824 19916 21876 19922
rect 21824 19858 21876 19864
rect 21732 18964 21784 18970
rect 21732 18906 21784 18912
rect 21640 18080 21692 18086
rect 21638 18048 21640 18057
rect 21692 18048 21694 18057
rect 21638 17983 21694 17992
rect 21456 17876 21508 17882
rect 21456 17818 21508 17824
rect 21468 16998 21496 17818
rect 21640 17060 21692 17066
rect 21640 17002 21692 17008
rect 21456 16992 21508 16998
rect 21652 16946 21680 17002
rect 21456 16934 21508 16940
rect 21560 16918 21680 16946
rect 21732 16992 21784 16998
rect 21732 16934 21784 16940
rect 21364 16652 21416 16658
rect 21364 16594 21416 16600
rect 21376 16182 21404 16594
rect 21456 16584 21508 16590
rect 21456 16526 21508 16532
rect 21364 16176 21416 16182
rect 21364 16118 21416 16124
rect 21364 16040 21416 16046
rect 21364 15982 21416 15988
rect 21376 15638 21404 15982
rect 21364 15632 21416 15638
rect 21468 15609 21496 16526
rect 21364 15574 21416 15580
rect 21454 15600 21510 15609
rect 21454 15535 21510 15544
rect 21364 14816 21416 14822
rect 21364 14758 21416 14764
rect 21376 14618 21404 14758
rect 21364 14612 21416 14618
rect 21364 14554 21416 14560
rect 21284 14334 21496 14362
rect 21364 14272 21416 14278
rect 21364 14214 21416 14220
rect 21270 13968 21326 13977
rect 21270 13903 21326 13912
rect 21284 13870 21312 13903
rect 21272 13864 21324 13870
rect 21272 13806 21324 13812
rect 21272 13728 21324 13734
rect 21272 13670 21324 13676
rect 21284 13569 21312 13670
rect 21270 13560 21326 13569
rect 21270 13495 21326 13504
rect 21376 13394 21404 14214
rect 21364 13388 21416 13394
rect 21364 13330 21416 13336
rect 21376 12986 21404 13330
rect 21364 12980 21416 12986
rect 21364 12922 21416 12928
rect 21272 12640 21324 12646
rect 21272 12582 21324 12588
rect 21180 12436 21232 12442
rect 21180 12378 21232 12384
rect 21284 12374 21312 12582
rect 21272 12368 21324 12374
rect 21192 12316 21272 12322
rect 21192 12310 21324 12316
rect 21192 12294 21312 12310
rect 21192 7818 21220 12294
rect 21284 12245 21312 12294
rect 21468 12152 21496 14334
rect 21284 12124 21496 12152
rect 21284 11694 21312 12124
rect 21362 12064 21418 12073
rect 21362 11999 21418 12008
rect 21272 11688 21324 11694
rect 21272 11630 21324 11636
rect 21284 10810 21312 11630
rect 21272 10804 21324 10810
rect 21272 10746 21324 10752
rect 21272 10464 21324 10470
rect 21272 10406 21324 10412
rect 21180 7812 21232 7818
rect 21180 7754 21232 7760
rect 21180 5160 21232 5166
rect 21180 5102 21232 5108
rect 21192 4622 21220 5102
rect 21180 4616 21232 4622
rect 21180 4558 21232 4564
rect 21088 2576 21140 2582
rect 21088 2518 21140 2524
rect 20904 2508 20956 2514
rect 20904 2450 20956 2456
rect 19984 2100 20036 2106
rect 19984 2042 20036 2048
rect 16856 1964 16908 1970
rect 16856 1906 16908 1912
rect 19892 1964 19944 1970
rect 19892 1906 19944 1912
rect 1674 0 1730 800
rect 5078 0 5134 800
rect 8574 0 8630 800
rect 12070 0 12126 800
rect 15566 0 15622 800
rect 19062 0 19118 800
rect 21284 377 21312 10406
rect 21376 1601 21404 11999
rect 21560 11608 21588 16918
rect 21744 15978 21772 16934
rect 21732 15972 21784 15978
rect 21732 15914 21784 15920
rect 21732 14884 21784 14890
rect 21732 14826 21784 14832
rect 21640 14612 21692 14618
rect 21640 14554 21692 14560
rect 21652 13394 21680 14554
rect 21640 13388 21692 13394
rect 21640 13330 21692 13336
rect 21468 11580 21588 11608
rect 21468 10266 21496 11580
rect 21548 10668 21600 10674
rect 21548 10610 21600 10616
rect 21456 10260 21508 10266
rect 21456 10202 21508 10208
rect 21560 9568 21588 10610
rect 21551 9540 21588 9568
rect 21551 9500 21579 9540
rect 21551 9472 21588 9500
rect 21456 8968 21508 8974
rect 21456 8910 21508 8916
rect 21468 6866 21496 8910
rect 21560 7274 21588 9472
rect 21548 7268 21600 7274
rect 21548 7210 21600 7216
rect 21456 6860 21508 6866
rect 21456 6802 21508 6808
rect 21468 6458 21496 6802
rect 21456 6452 21508 6458
rect 21456 6394 21508 6400
rect 21652 5896 21680 13330
rect 21744 12986 21772 14826
rect 21732 12980 21784 12986
rect 21732 12922 21784 12928
rect 21836 10470 21864 19858
rect 21928 19825 21956 20266
rect 21914 19816 21970 19825
rect 21914 19751 21970 19760
rect 22020 18766 22048 21490
rect 22112 19514 22140 23600
rect 22468 21004 22520 21010
rect 22468 20946 22520 20952
rect 22652 21004 22704 21010
rect 22652 20946 22704 20952
rect 22376 20256 22428 20262
rect 22376 20198 22428 20204
rect 22388 20097 22416 20198
rect 22374 20088 22430 20097
rect 22374 20023 22430 20032
rect 22100 19508 22152 19514
rect 22100 19450 22152 19456
rect 22192 19168 22244 19174
rect 22192 19110 22244 19116
rect 22008 18760 22060 18766
rect 22008 18702 22060 18708
rect 22100 18624 22152 18630
rect 22100 18566 22152 18572
rect 21916 18284 21968 18290
rect 21916 18226 21968 18232
rect 21928 11762 21956 18226
rect 22008 18080 22060 18086
rect 22008 18022 22060 18028
rect 21916 11756 21968 11762
rect 21916 11698 21968 11704
rect 22020 10577 22048 18022
rect 22112 17338 22140 18566
rect 22204 17814 22232 19110
rect 22284 18080 22336 18086
rect 22284 18022 22336 18028
rect 22376 18080 22428 18086
rect 22376 18022 22428 18028
rect 22192 17808 22244 17814
rect 22192 17750 22244 17756
rect 22100 17332 22152 17338
rect 22100 17274 22152 17280
rect 22192 17128 22244 17134
rect 22192 17070 22244 17076
rect 22100 16720 22152 16726
rect 22100 16662 22152 16668
rect 22112 14385 22140 16662
rect 22204 16046 22232 17070
rect 22192 16040 22244 16046
rect 22192 15982 22244 15988
rect 22296 15314 22324 18022
rect 22388 16250 22416 18022
rect 22376 16244 22428 16250
rect 22376 16186 22428 16192
rect 22204 15286 22324 15314
rect 22376 15360 22428 15366
rect 22376 15302 22428 15308
rect 22098 14376 22154 14385
rect 22098 14311 22154 14320
rect 22100 14272 22152 14278
rect 22100 14214 22152 14220
rect 22006 10568 22062 10577
rect 21916 10532 21968 10538
rect 22006 10503 22062 10512
rect 21916 10474 21968 10480
rect 21824 10464 21876 10470
rect 21824 10406 21876 10412
rect 21824 10260 21876 10266
rect 21824 10202 21876 10208
rect 21732 9104 21784 9110
rect 21732 9046 21784 9052
rect 21744 8294 21772 9046
rect 21732 8288 21784 8294
rect 21732 8230 21784 8236
rect 21744 7313 21772 8230
rect 21730 7304 21786 7313
rect 21730 7239 21786 7248
rect 21836 7206 21864 10202
rect 21928 9178 21956 10474
rect 22008 10464 22060 10470
rect 22008 10406 22060 10412
rect 21916 9172 21968 9178
rect 21916 9114 21968 9120
rect 21824 7200 21876 7206
rect 21824 7142 21876 7148
rect 21824 6316 21876 6322
rect 21824 6258 21876 6264
rect 21468 5868 21680 5896
rect 21468 2038 21496 5868
rect 21548 5772 21600 5778
rect 21548 5714 21600 5720
rect 21560 3738 21588 5714
rect 21836 5710 21864 6258
rect 22020 6254 22048 10406
rect 22008 6248 22060 6254
rect 22008 6190 22060 6196
rect 21916 6180 21968 6186
rect 21916 6122 21968 6128
rect 21732 5704 21784 5710
rect 21732 5646 21784 5652
rect 21824 5704 21876 5710
rect 21824 5646 21876 5652
rect 21640 5092 21692 5098
rect 21640 5034 21692 5040
rect 21652 4826 21680 5034
rect 21640 4820 21692 4826
rect 21640 4762 21692 4768
rect 21548 3732 21600 3738
rect 21548 3674 21600 3680
rect 21560 3618 21588 3674
rect 21744 3670 21772 5646
rect 21928 4690 21956 6122
rect 22008 6112 22060 6118
rect 22008 6054 22060 6060
rect 21916 4684 21968 4690
rect 21916 4626 21968 4632
rect 21824 4004 21876 4010
rect 21824 3946 21876 3952
rect 21732 3664 21784 3670
rect 21560 3590 21680 3618
rect 21732 3606 21784 3612
rect 21652 2582 21680 3590
rect 21744 3194 21772 3606
rect 21732 3188 21784 3194
rect 21732 3130 21784 3136
rect 21836 2650 21864 3946
rect 21928 3942 21956 4626
rect 22020 4078 22048 6054
rect 22112 5001 22140 14214
rect 22204 11354 22232 15286
rect 22284 14816 22336 14822
rect 22284 14758 22336 14764
rect 22296 14074 22324 14758
rect 22388 14550 22416 15302
rect 22376 14544 22428 14550
rect 22376 14486 22428 14492
rect 22480 14090 22508 20946
rect 22560 19712 22612 19718
rect 22560 19654 22612 19660
rect 22572 17066 22600 19654
rect 22560 17060 22612 17066
rect 22560 17002 22612 17008
rect 22284 14068 22336 14074
rect 22284 14010 22336 14016
rect 22388 14062 22508 14090
rect 22388 13818 22416 14062
rect 22468 13932 22520 13938
rect 22468 13874 22520 13880
rect 22296 13790 22416 13818
rect 22296 12730 22324 13790
rect 22376 13728 22428 13734
rect 22376 13670 22428 13676
rect 22388 13462 22416 13670
rect 22376 13456 22428 13462
rect 22376 13398 22428 13404
rect 22374 13152 22430 13161
rect 22480 13138 22508 13874
rect 22430 13110 22508 13138
rect 22374 13087 22430 13096
rect 22388 12850 22416 13087
rect 22376 12844 22428 12850
rect 22376 12786 22428 12792
rect 22296 12702 22508 12730
rect 22284 12640 22336 12646
rect 22284 12582 22336 12588
rect 22296 12345 22324 12582
rect 22282 12336 22338 12345
rect 22282 12271 22338 12280
rect 22282 11792 22338 11801
rect 22282 11727 22338 11736
rect 22296 11694 22324 11727
rect 22284 11688 22336 11694
rect 22284 11630 22336 11636
rect 22192 11348 22244 11354
rect 22192 11290 22244 11296
rect 22480 10266 22508 12702
rect 22468 10260 22520 10266
rect 22468 10202 22520 10208
rect 22192 9988 22244 9994
rect 22192 9930 22244 9936
rect 22204 9518 22232 9930
rect 22192 9512 22244 9518
rect 22192 9454 22244 9460
rect 22468 8968 22520 8974
rect 22468 8910 22520 8916
rect 22284 8832 22336 8838
rect 22284 8774 22336 8780
rect 22296 8498 22324 8774
rect 22284 8492 22336 8498
rect 22284 8434 22336 8440
rect 22480 8022 22508 8910
rect 22664 8634 22692 20946
rect 22756 17542 22784 23600
rect 22928 21548 22980 21554
rect 22928 21490 22980 21496
rect 22836 20800 22888 20806
rect 22836 20742 22888 20748
rect 22848 20097 22876 20742
rect 22834 20088 22890 20097
rect 22834 20023 22890 20032
rect 22836 19712 22888 19718
rect 22836 19654 22888 19660
rect 22848 19417 22876 19654
rect 22834 19408 22890 19417
rect 22834 19343 22890 19352
rect 22836 17672 22888 17678
rect 22836 17614 22888 17620
rect 22744 17536 22796 17542
rect 22744 17478 22796 17484
rect 22744 15904 22796 15910
rect 22744 15846 22796 15852
rect 22756 15570 22784 15846
rect 22744 15564 22796 15570
rect 22744 15506 22796 15512
rect 22848 11234 22876 17614
rect 22756 11206 22876 11234
rect 22652 8628 22704 8634
rect 22652 8570 22704 8576
rect 22652 8492 22704 8498
rect 22652 8434 22704 8440
rect 22560 8356 22612 8362
rect 22560 8298 22612 8304
rect 22468 8016 22520 8022
rect 22468 7958 22520 7964
rect 22376 7744 22428 7750
rect 22376 7686 22428 7692
rect 22190 7440 22246 7449
rect 22190 7375 22246 7384
rect 22098 4992 22154 5001
rect 22098 4927 22154 4936
rect 22204 4321 22232 7375
rect 22388 7274 22416 7686
rect 22480 7546 22508 7958
rect 22468 7540 22520 7546
rect 22468 7482 22520 7488
rect 22376 7268 22428 7274
rect 22376 7210 22428 7216
rect 22572 6866 22600 8298
rect 22664 7342 22692 8434
rect 22652 7336 22704 7342
rect 22652 7278 22704 7284
rect 22664 7002 22692 7278
rect 22652 6996 22704 7002
rect 22652 6938 22704 6944
rect 22560 6860 22612 6866
rect 22560 6802 22612 6808
rect 22558 6216 22614 6225
rect 22558 6151 22614 6160
rect 22572 5846 22600 6151
rect 22560 5840 22612 5846
rect 22560 5782 22612 5788
rect 22190 4312 22246 4321
rect 22190 4247 22246 4256
rect 22008 4072 22060 4078
rect 22008 4014 22060 4020
rect 21916 3936 21968 3942
rect 21916 3878 21968 3884
rect 22098 3496 22154 3505
rect 22098 3431 22154 3440
rect 22112 2990 22140 3431
rect 22100 2984 22152 2990
rect 22100 2926 22152 2932
rect 22560 2916 22612 2922
rect 22560 2858 22612 2864
rect 21824 2644 21876 2650
rect 21824 2586 21876 2592
rect 21640 2576 21692 2582
rect 21640 2518 21692 2524
rect 21456 2032 21508 2038
rect 21456 1974 21508 1980
rect 21362 1592 21418 1601
rect 21362 1527 21418 1536
rect 22572 800 22600 2858
rect 22756 2854 22784 11206
rect 22836 11076 22888 11082
rect 22836 11018 22888 11024
rect 22848 8945 22876 11018
rect 22940 9994 22968 21490
rect 23204 21344 23256 21350
rect 23204 21286 23256 21292
rect 23020 20936 23072 20942
rect 23020 20878 23072 20884
rect 23032 10198 23060 20878
rect 23112 16652 23164 16658
rect 23112 16594 23164 16600
rect 23020 10192 23072 10198
rect 23020 10134 23072 10140
rect 22928 9988 22980 9994
rect 22928 9930 22980 9936
rect 23124 9625 23152 16594
rect 23216 10810 23244 21286
rect 23400 20534 23428 23600
rect 24044 21690 24072 23600
rect 24032 21684 24084 21690
rect 24032 21626 24084 21632
rect 23388 20528 23440 20534
rect 23388 20470 23440 20476
rect 23204 10804 23256 10810
rect 23204 10746 23256 10752
rect 23110 9616 23166 9625
rect 23110 9551 23166 9560
rect 22834 8936 22890 8945
rect 22834 8871 22890 8880
rect 22848 5545 22876 8871
rect 22928 8628 22980 8634
rect 22928 8570 22980 8576
rect 22940 8294 22968 8570
rect 22928 8288 22980 8294
rect 22928 8230 22980 8236
rect 22834 5536 22890 5545
rect 22834 5471 22890 5480
rect 22744 2848 22796 2854
rect 22744 2790 22796 2796
rect 22940 921 22968 8230
rect 23386 6896 23442 6905
rect 23386 6831 23388 6840
rect 23440 6831 23442 6840
rect 23388 6802 23440 6808
rect 22926 912 22982 921
rect 22926 847 22982 856
rect 21270 368 21326 377
rect 21270 303 21326 312
rect 22558 0 22614 800
<< via2 >>
rect 19430 23976 19486 24032
rect 1858 19760 1914 19816
rect 2778 19760 2834 19816
rect 3238 20168 3294 20224
rect 1490 15408 1546 15464
rect 1858 15136 1914 15192
rect 1674 14320 1730 14376
rect 1582 12280 1638 12336
rect 1490 9016 1546 9072
rect 1950 3052 2006 3088
rect 1950 3032 1952 3052
rect 1952 3032 2004 3052
rect 2004 3032 2006 3052
rect 2870 13776 2926 13832
rect 3790 19896 3846 19952
rect 3330 16632 3386 16688
rect 4654 21786 4710 21788
rect 4734 21786 4790 21788
rect 4814 21786 4870 21788
rect 4894 21786 4950 21788
rect 4654 21734 4680 21786
rect 4680 21734 4710 21786
rect 4734 21734 4744 21786
rect 4744 21734 4790 21786
rect 4814 21734 4860 21786
rect 4860 21734 4870 21786
rect 4894 21734 4924 21786
rect 4924 21734 4950 21786
rect 4654 21732 4710 21734
rect 4734 21732 4790 21734
rect 4814 21732 4870 21734
rect 4894 21732 4950 21734
rect 4342 21392 4398 21448
rect 3790 15000 3846 15056
rect 4654 20698 4710 20700
rect 4734 20698 4790 20700
rect 4814 20698 4870 20700
rect 4894 20698 4950 20700
rect 4654 20646 4680 20698
rect 4680 20646 4710 20698
rect 4734 20646 4744 20698
rect 4744 20646 4790 20698
rect 4814 20646 4860 20698
rect 4860 20646 4870 20698
rect 4894 20646 4924 20698
rect 4924 20646 4950 20698
rect 4654 20644 4710 20646
rect 4734 20644 4790 20646
rect 4814 20644 4870 20646
rect 4894 20644 4950 20646
rect 4802 19760 4858 19816
rect 4654 19610 4710 19612
rect 4734 19610 4790 19612
rect 4814 19610 4870 19612
rect 4894 19610 4950 19612
rect 4654 19558 4680 19610
rect 4680 19558 4710 19610
rect 4734 19558 4744 19610
rect 4744 19558 4790 19610
rect 4814 19558 4860 19610
rect 4860 19558 4870 19610
rect 4894 19558 4924 19610
rect 4924 19558 4950 19610
rect 4654 19556 4710 19558
rect 4734 19556 4790 19558
rect 4814 19556 4870 19558
rect 4894 19556 4950 19558
rect 4654 18522 4710 18524
rect 4734 18522 4790 18524
rect 4814 18522 4870 18524
rect 4894 18522 4950 18524
rect 4654 18470 4680 18522
rect 4680 18470 4710 18522
rect 4734 18470 4744 18522
rect 4744 18470 4790 18522
rect 4814 18470 4860 18522
rect 4860 18470 4870 18522
rect 4894 18470 4924 18522
rect 4924 18470 4950 18522
rect 4654 18468 4710 18470
rect 4734 18468 4790 18470
rect 4814 18468 4870 18470
rect 4894 18468 4950 18470
rect 4894 17584 4950 17640
rect 4654 17434 4710 17436
rect 4734 17434 4790 17436
rect 4814 17434 4870 17436
rect 4894 17434 4950 17436
rect 4654 17382 4680 17434
rect 4680 17382 4710 17434
rect 4734 17382 4744 17434
rect 4744 17382 4790 17434
rect 4814 17382 4860 17434
rect 4860 17382 4870 17434
rect 4894 17382 4924 17434
rect 4924 17382 4950 17434
rect 4654 17380 4710 17382
rect 4734 17380 4790 17382
rect 4814 17380 4870 17382
rect 4894 17380 4950 17382
rect 4802 17176 4858 17232
rect 3974 13232 4030 13288
rect 3882 12416 3938 12472
rect 3606 10004 3608 10024
rect 3608 10004 3660 10024
rect 3660 10004 3662 10024
rect 3606 9968 3662 10004
rect 4654 16346 4710 16348
rect 4734 16346 4790 16348
rect 4814 16346 4870 16348
rect 4894 16346 4950 16348
rect 4654 16294 4680 16346
rect 4680 16294 4710 16346
rect 4734 16294 4744 16346
rect 4744 16294 4790 16346
rect 4814 16294 4860 16346
rect 4860 16294 4870 16346
rect 4894 16294 4924 16346
rect 4924 16294 4950 16346
rect 4654 16292 4710 16294
rect 4734 16292 4790 16294
rect 4814 16292 4870 16294
rect 4894 16292 4950 16294
rect 5262 16904 5318 16960
rect 4654 15258 4710 15260
rect 4734 15258 4790 15260
rect 4814 15258 4870 15260
rect 4894 15258 4950 15260
rect 4654 15206 4680 15258
rect 4680 15206 4710 15258
rect 4734 15206 4744 15258
rect 4744 15206 4790 15258
rect 4814 15206 4860 15258
rect 4860 15206 4870 15258
rect 4894 15206 4924 15258
rect 4924 15206 4950 15258
rect 4654 15204 4710 15206
rect 4734 15204 4790 15206
rect 4814 15204 4870 15206
rect 4894 15204 4950 15206
rect 4654 14170 4710 14172
rect 4734 14170 4790 14172
rect 4814 14170 4870 14172
rect 4894 14170 4950 14172
rect 4654 14118 4680 14170
rect 4680 14118 4710 14170
rect 4734 14118 4744 14170
rect 4744 14118 4790 14170
rect 4814 14118 4860 14170
rect 4860 14118 4870 14170
rect 4894 14118 4924 14170
rect 4924 14118 4950 14170
rect 4654 14116 4710 14118
rect 4734 14116 4790 14118
rect 4814 14116 4870 14118
rect 4894 14116 4950 14118
rect 4654 13082 4710 13084
rect 4734 13082 4790 13084
rect 4814 13082 4870 13084
rect 4894 13082 4950 13084
rect 4654 13030 4680 13082
rect 4680 13030 4710 13082
rect 4734 13030 4744 13082
rect 4744 13030 4790 13082
rect 4814 13030 4860 13082
rect 4860 13030 4870 13082
rect 4894 13030 4924 13082
rect 4924 13030 4950 13082
rect 4654 13028 4710 13030
rect 4734 13028 4790 13030
rect 4814 13028 4870 13030
rect 4894 13028 4950 13030
rect 4654 11994 4710 11996
rect 4734 11994 4790 11996
rect 4814 11994 4870 11996
rect 4894 11994 4950 11996
rect 4654 11942 4680 11994
rect 4680 11942 4710 11994
rect 4734 11942 4744 11994
rect 4744 11942 4790 11994
rect 4814 11942 4860 11994
rect 4860 11942 4870 11994
rect 4894 11942 4924 11994
rect 4924 11942 4950 11994
rect 4654 11940 4710 11942
rect 4734 11940 4790 11942
rect 4814 11940 4870 11942
rect 4894 11940 4950 11942
rect 4654 10906 4710 10908
rect 4734 10906 4790 10908
rect 4814 10906 4870 10908
rect 4894 10906 4950 10908
rect 4654 10854 4680 10906
rect 4680 10854 4710 10906
rect 4734 10854 4744 10906
rect 4744 10854 4790 10906
rect 4814 10854 4860 10906
rect 4860 10854 4870 10906
rect 4894 10854 4924 10906
rect 4924 10854 4950 10906
rect 4654 10852 4710 10854
rect 4734 10852 4790 10854
rect 4814 10852 4870 10854
rect 4894 10852 4950 10854
rect 4654 9818 4710 9820
rect 4734 9818 4790 9820
rect 4814 9818 4870 9820
rect 4894 9818 4950 9820
rect 4654 9766 4680 9818
rect 4680 9766 4710 9818
rect 4734 9766 4744 9818
rect 4744 9766 4790 9818
rect 4814 9766 4860 9818
rect 4860 9766 4870 9818
rect 4894 9766 4924 9818
rect 4924 9766 4950 9818
rect 4654 9764 4710 9766
rect 4734 9764 4790 9766
rect 4814 9764 4870 9766
rect 4894 9764 4950 9766
rect 4894 9560 4950 9616
rect 4654 8730 4710 8732
rect 4734 8730 4790 8732
rect 4814 8730 4870 8732
rect 4894 8730 4950 8732
rect 4654 8678 4680 8730
rect 4680 8678 4710 8730
rect 4734 8678 4744 8730
rect 4744 8678 4790 8730
rect 4814 8678 4860 8730
rect 4860 8678 4870 8730
rect 4894 8678 4924 8730
rect 4924 8678 4950 8730
rect 4654 8676 4710 8678
rect 4734 8676 4790 8678
rect 4814 8676 4870 8678
rect 4894 8676 4950 8678
rect 4710 8336 4766 8392
rect 5630 20204 5632 20224
rect 5632 20204 5684 20224
rect 5684 20204 5686 20224
rect 5630 20168 5686 20204
rect 6182 21936 6238 21992
rect 6090 21528 6146 21584
rect 5722 19760 5778 19816
rect 6642 19488 6698 19544
rect 6734 19216 6790 19272
rect 6550 18536 6606 18592
rect 6458 17720 6514 17776
rect 5170 9968 5226 10024
rect 4654 7642 4710 7644
rect 4734 7642 4790 7644
rect 4814 7642 4870 7644
rect 4894 7642 4950 7644
rect 4654 7590 4680 7642
rect 4680 7590 4710 7642
rect 4734 7590 4744 7642
rect 4744 7590 4790 7642
rect 4814 7590 4860 7642
rect 4860 7590 4870 7642
rect 4894 7590 4924 7642
rect 4924 7590 4950 7642
rect 4654 7588 4710 7590
rect 4734 7588 4790 7590
rect 4814 7588 4870 7590
rect 4894 7588 4950 7590
rect 4654 6554 4710 6556
rect 4734 6554 4790 6556
rect 4814 6554 4870 6556
rect 4894 6554 4950 6556
rect 4654 6502 4680 6554
rect 4680 6502 4710 6554
rect 4734 6502 4744 6554
rect 4744 6502 4790 6554
rect 4814 6502 4860 6554
rect 4860 6502 4870 6554
rect 4894 6502 4924 6554
rect 4924 6502 4950 6554
rect 4654 6500 4710 6502
rect 4734 6500 4790 6502
rect 4814 6500 4870 6502
rect 4894 6500 4950 6502
rect 4654 5466 4710 5468
rect 4734 5466 4790 5468
rect 4814 5466 4870 5468
rect 4894 5466 4950 5468
rect 4654 5414 4680 5466
rect 4680 5414 4710 5466
rect 4734 5414 4744 5466
rect 4744 5414 4790 5466
rect 4814 5414 4860 5466
rect 4860 5414 4870 5466
rect 4894 5414 4924 5466
rect 4924 5414 4950 5466
rect 4654 5412 4710 5414
rect 4734 5412 4790 5414
rect 4814 5412 4870 5414
rect 4894 5412 4950 5414
rect 4654 4378 4710 4380
rect 4734 4378 4790 4380
rect 4814 4378 4870 4380
rect 4894 4378 4950 4380
rect 4654 4326 4680 4378
rect 4680 4326 4710 4378
rect 4734 4326 4744 4378
rect 4744 4326 4790 4378
rect 4814 4326 4860 4378
rect 4860 4326 4870 4378
rect 4894 4326 4924 4378
rect 4924 4326 4950 4378
rect 4654 4324 4710 4326
rect 4734 4324 4790 4326
rect 4814 4324 4870 4326
rect 4894 4324 4950 4326
rect 5998 13368 6054 13424
rect 5446 8780 5448 8800
rect 5448 8780 5500 8800
rect 5500 8780 5502 8800
rect 5446 8744 5502 8780
rect 5354 8492 5410 8528
rect 5354 8472 5356 8492
rect 5356 8472 5408 8492
rect 5408 8472 5410 8492
rect 5722 9016 5778 9072
rect 6642 17176 6698 17232
rect 7010 20304 7066 20360
rect 7010 17176 7066 17232
rect 7194 17040 7250 17096
rect 6458 12824 6514 12880
rect 6366 12416 6422 12472
rect 6366 10512 6422 10568
rect 5630 7812 5686 7848
rect 5630 7792 5632 7812
rect 5632 7792 5684 7812
rect 5684 7792 5686 7812
rect 5262 4664 5318 4720
rect 4654 3290 4710 3292
rect 4734 3290 4790 3292
rect 4814 3290 4870 3292
rect 4894 3290 4950 3292
rect 4654 3238 4680 3290
rect 4680 3238 4710 3290
rect 4734 3238 4744 3290
rect 4744 3238 4790 3290
rect 4814 3238 4860 3290
rect 4860 3238 4870 3290
rect 4894 3238 4924 3290
rect 4924 3238 4950 3290
rect 4654 3236 4710 3238
rect 4734 3236 4790 3238
rect 4814 3236 4870 3238
rect 4894 3236 4950 3238
rect 4654 2202 4710 2204
rect 4734 2202 4790 2204
rect 4814 2202 4870 2204
rect 4894 2202 4950 2204
rect 4654 2150 4680 2202
rect 4680 2150 4710 2202
rect 4734 2150 4744 2202
rect 4744 2150 4790 2202
rect 4814 2150 4860 2202
rect 4860 2150 4870 2202
rect 4894 2150 4924 2202
rect 4924 2150 4950 2202
rect 4654 2148 4710 2150
rect 4734 2148 4790 2150
rect 4814 2148 4870 2150
rect 4894 2148 4950 2150
rect 6550 11464 6606 11520
rect 7102 15544 7158 15600
rect 6826 14184 6882 14240
rect 6826 12688 6882 12744
rect 6918 12164 6974 12200
rect 6918 12144 6920 12164
rect 6920 12144 6972 12164
rect 6972 12144 6974 12164
rect 7010 9988 7066 10024
rect 7010 9968 7012 9988
rect 7012 9968 7064 9988
rect 7064 9968 7066 9988
rect 6918 7384 6974 7440
rect 6826 6432 6882 6488
rect 8353 21242 8409 21244
rect 8433 21242 8489 21244
rect 8513 21242 8569 21244
rect 8593 21242 8649 21244
rect 8353 21190 8379 21242
rect 8379 21190 8409 21242
rect 8433 21190 8443 21242
rect 8443 21190 8489 21242
rect 8513 21190 8559 21242
rect 8559 21190 8569 21242
rect 8593 21190 8623 21242
rect 8623 21190 8649 21242
rect 8353 21188 8409 21190
rect 8433 21188 8489 21190
rect 8513 21188 8569 21190
rect 8593 21188 8649 21190
rect 8353 20154 8409 20156
rect 8433 20154 8489 20156
rect 8513 20154 8569 20156
rect 8593 20154 8649 20156
rect 8353 20102 8379 20154
rect 8379 20102 8409 20154
rect 8433 20102 8443 20154
rect 8443 20102 8489 20154
rect 8513 20102 8559 20154
rect 8559 20102 8569 20154
rect 8593 20102 8623 20154
rect 8623 20102 8649 20154
rect 8353 20100 8409 20102
rect 8433 20100 8489 20102
rect 8513 20100 8569 20102
rect 8593 20100 8649 20102
rect 7654 19352 7710 19408
rect 7378 18672 7434 18728
rect 7378 16496 7434 16552
rect 7286 13912 7342 13968
rect 7286 10104 7342 10160
rect 7194 8880 7250 8936
rect 7470 14456 7526 14512
rect 9034 21528 9090 21584
rect 8942 21428 8944 21448
rect 8944 21428 8996 21448
rect 8996 21428 8998 21448
rect 8942 21392 8998 21428
rect 8850 20340 8852 20360
rect 8852 20340 8904 20360
rect 8904 20340 8906 20360
rect 8850 20304 8906 20340
rect 8942 19760 8998 19816
rect 7930 19372 7986 19408
rect 7930 19352 7932 19372
rect 7932 19352 7984 19372
rect 7984 19352 7986 19372
rect 8353 19066 8409 19068
rect 8433 19066 8489 19068
rect 8513 19066 8569 19068
rect 8593 19066 8649 19068
rect 8353 19014 8379 19066
rect 8379 19014 8409 19066
rect 8433 19014 8443 19066
rect 8443 19014 8489 19066
rect 8513 19014 8559 19066
rect 8559 19014 8569 19066
rect 8593 19014 8623 19066
rect 8623 19014 8649 19066
rect 8353 19012 8409 19014
rect 8433 19012 8489 19014
rect 8513 19012 8569 19014
rect 8593 19012 8649 19014
rect 8482 18572 8484 18592
rect 8484 18572 8536 18592
rect 8536 18572 8538 18592
rect 8482 18536 8538 18572
rect 8353 17978 8409 17980
rect 8433 17978 8489 17980
rect 8513 17978 8569 17980
rect 8593 17978 8649 17980
rect 8353 17926 8379 17978
rect 8379 17926 8409 17978
rect 8433 17926 8443 17978
rect 8443 17926 8489 17978
rect 8513 17926 8559 17978
rect 8559 17926 8569 17978
rect 8593 17926 8623 17978
rect 8623 17926 8649 17978
rect 8353 17924 8409 17926
rect 8433 17924 8489 17926
rect 8513 17924 8569 17926
rect 8593 17924 8649 17926
rect 9126 20032 9182 20088
rect 9126 17584 9182 17640
rect 8353 16890 8409 16892
rect 8433 16890 8489 16892
rect 8513 16890 8569 16892
rect 8593 16890 8649 16892
rect 8353 16838 8379 16890
rect 8379 16838 8409 16890
rect 8433 16838 8443 16890
rect 8443 16838 8489 16890
rect 8513 16838 8559 16890
rect 8559 16838 8569 16890
rect 8593 16838 8623 16890
rect 8623 16838 8649 16890
rect 8353 16836 8409 16838
rect 8433 16836 8489 16838
rect 8513 16836 8569 16838
rect 8593 16836 8649 16838
rect 7470 9424 7526 9480
rect 7470 8608 7526 8664
rect 8353 15802 8409 15804
rect 8433 15802 8489 15804
rect 8513 15802 8569 15804
rect 8593 15802 8649 15804
rect 8353 15750 8379 15802
rect 8379 15750 8409 15802
rect 8433 15750 8443 15802
rect 8443 15750 8489 15802
rect 8513 15750 8559 15802
rect 8559 15750 8569 15802
rect 8593 15750 8623 15802
rect 8623 15750 8649 15802
rect 8353 15748 8409 15750
rect 8433 15748 8489 15750
rect 8513 15748 8569 15750
rect 8593 15748 8649 15750
rect 9678 21936 9734 21992
rect 9402 20168 9458 20224
rect 9586 20032 9642 20088
rect 9310 19760 9366 19816
rect 9402 19624 9458 19680
rect 9494 19488 9550 19544
rect 9310 17620 9312 17640
rect 9312 17620 9364 17640
rect 9364 17620 9366 17640
rect 9310 17584 9366 17620
rect 9586 19216 9642 19272
rect 9494 17992 9550 18048
rect 8942 16108 8998 16144
rect 8942 16088 8944 16108
rect 8944 16088 8996 16108
rect 8996 16088 8998 16108
rect 8353 14714 8409 14716
rect 8433 14714 8489 14716
rect 8513 14714 8569 14716
rect 8593 14714 8649 14716
rect 8353 14662 8379 14714
rect 8379 14662 8409 14714
rect 8433 14662 8443 14714
rect 8443 14662 8489 14714
rect 8513 14662 8559 14714
rect 8559 14662 8569 14714
rect 8593 14662 8623 14714
rect 8623 14662 8649 14714
rect 8353 14660 8409 14662
rect 8433 14660 8489 14662
rect 8513 14660 8569 14662
rect 8593 14660 8649 14662
rect 7930 9424 7986 9480
rect 7562 6724 7618 6760
rect 7562 6704 7564 6724
rect 7564 6704 7616 6724
rect 7616 6704 7618 6724
rect 8353 13626 8409 13628
rect 8433 13626 8489 13628
rect 8513 13626 8569 13628
rect 8593 13626 8649 13628
rect 8353 13574 8379 13626
rect 8379 13574 8409 13626
rect 8433 13574 8443 13626
rect 8443 13574 8489 13626
rect 8513 13574 8559 13626
rect 8559 13574 8569 13626
rect 8593 13574 8623 13626
rect 8623 13574 8649 13626
rect 8353 13572 8409 13574
rect 8433 13572 8489 13574
rect 8513 13572 8569 13574
rect 8593 13572 8649 13574
rect 8353 12538 8409 12540
rect 8433 12538 8489 12540
rect 8513 12538 8569 12540
rect 8593 12538 8649 12540
rect 8353 12486 8379 12538
rect 8379 12486 8409 12538
rect 8433 12486 8443 12538
rect 8443 12486 8489 12538
rect 8513 12486 8559 12538
rect 8559 12486 8569 12538
rect 8593 12486 8623 12538
rect 8623 12486 8649 12538
rect 8353 12484 8409 12486
rect 8433 12484 8489 12486
rect 8513 12484 8569 12486
rect 8593 12484 8649 12486
rect 8942 12280 8998 12336
rect 9402 15816 9458 15872
rect 9218 13132 9220 13152
rect 9220 13132 9272 13152
rect 9272 13132 9274 13152
rect 9218 13096 9274 13132
rect 8353 11450 8409 11452
rect 8433 11450 8489 11452
rect 8513 11450 8569 11452
rect 8593 11450 8649 11452
rect 8353 11398 8379 11450
rect 8379 11398 8409 11450
rect 8433 11398 8443 11450
rect 8443 11398 8489 11450
rect 8513 11398 8559 11450
rect 8559 11398 8569 11450
rect 8593 11398 8623 11450
rect 8623 11398 8649 11450
rect 8353 11396 8409 11398
rect 8433 11396 8489 11398
rect 8513 11396 8569 11398
rect 8593 11396 8649 11398
rect 8353 10362 8409 10364
rect 8433 10362 8489 10364
rect 8513 10362 8569 10364
rect 8593 10362 8649 10364
rect 8353 10310 8379 10362
rect 8379 10310 8409 10362
rect 8433 10310 8443 10362
rect 8443 10310 8489 10362
rect 8513 10310 8559 10362
rect 8559 10310 8569 10362
rect 8593 10310 8623 10362
rect 8623 10310 8649 10362
rect 8353 10308 8409 10310
rect 8433 10308 8489 10310
rect 8513 10308 8569 10310
rect 8593 10308 8649 10310
rect 8353 9274 8409 9276
rect 8433 9274 8489 9276
rect 8513 9274 8569 9276
rect 8593 9274 8649 9276
rect 8353 9222 8379 9274
rect 8379 9222 8409 9274
rect 8433 9222 8443 9274
rect 8443 9222 8489 9274
rect 8513 9222 8559 9274
rect 8559 9222 8569 9274
rect 8593 9222 8623 9274
rect 8623 9222 8649 9274
rect 8353 9220 8409 9222
rect 8433 9220 8489 9222
rect 8513 9220 8569 9222
rect 8593 9220 8649 9222
rect 10506 20848 10562 20904
rect 10414 20440 10470 20496
rect 9862 20052 9918 20088
rect 9862 20032 9864 20052
rect 9864 20032 9916 20052
rect 9916 20032 9918 20052
rect 10046 19352 10102 19408
rect 10046 19080 10102 19136
rect 9954 16224 10010 16280
rect 10598 19080 10654 19136
rect 11058 20168 11114 20224
rect 11150 19896 11206 19952
rect 11058 18264 11114 18320
rect 10598 17720 10654 17776
rect 9954 13776 10010 13832
rect 10322 16088 10378 16144
rect 9586 11600 9642 11656
rect 10598 14900 10600 14920
rect 10600 14900 10652 14920
rect 10652 14900 10654 14920
rect 10598 14864 10654 14900
rect 9862 10920 9918 10976
rect 9678 10648 9734 10704
rect 9862 10648 9918 10704
rect 9658 10260 9714 10296
rect 9658 10240 9680 10260
rect 9680 10240 9714 10260
rect 10046 10648 10102 10704
rect 10046 10376 10102 10432
rect 9218 9016 9274 9072
rect 9678 9696 9734 9752
rect 9862 9832 9918 9888
rect 9218 8744 9274 8800
rect 8353 8186 8409 8188
rect 8433 8186 8489 8188
rect 8513 8186 8569 8188
rect 8593 8186 8649 8188
rect 8353 8134 8379 8186
rect 8379 8134 8409 8186
rect 8433 8134 8443 8186
rect 8443 8134 8489 8186
rect 8513 8134 8559 8186
rect 8559 8134 8569 8186
rect 8593 8134 8623 8186
rect 8623 8134 8649 8186
rect 8353 8132 8409 8134
rect 8433 8132 8489 8134
rect 8513 8132 8569 8134
rect 8593 8132 8649 8134
rect 8353 7098 8409 7100
rect 8433 7098 8489 7100
rect 8513 7098 8569 7100
rect 8593 7098 8649 7100
rect 8353 7046 8379 7098
rect 8379 7046 8409 7098
rect 8433 7046 8443 7098
rect 8443 7046 8489 7098
rect 8513 7046 8559 7098
rect 8559 7046 8569 7098
rect 8593 7046 8623 7098
rect 8623 7046 8649 7098
rect 8353 7044 8409 7046
rect 8433 7044 8489 7046
rect 8513 7044 8569 7046
rect 8593 7044 8649 7046
rect 10782 16088 10838 16144
rect 10230 8064 10286 8120
rect 10690 8200 10746 8256
rect 8850 6976 8906 7032
rect 8482 6296 8538 6352
rect 8353 6010 8409 6012
rect 8433 6010 8489 6012
rect 8513 6010 8569 6012
rect 8593 6010 8649 6012
rect 8353 5958 8379 6010
rect 8379 5958 8409 6010
rect 8433 5958 8443 6010
rect 8443 5958 8489 6010
rect 8513 5958 8559 6010
rect 8559 5958 8569 6010
rect 8593 5958 8623 6010
rect 8623 5958 8649 6010
rect 8353 5956 8409 5958
rect 8433 5956 8489 5958
rect 8513 5956 8569 5958
rect 8593 5956 8649 5958
rect 9586 6996 9642 7032
rect 9586 6976 9588 6996
rect 9588 6976 9640 6996
rect 9640 6976 9642 6996
rect 9770 5772 9826 5808
rect 9770 5752 9772 5772
rect 9772 5752 9824 5772
rect 9824 5752 9826 5772
rect 8666 5208 8722 5264
rect 8353 4922 8409 4924
rect 8433 4922 8489 4924
rect 8513 4922 8569 4924
rect 8593 4922 8649 4924
rect 8353 4870 8379 4922
rect 8379 4870 8409 4922
rect 8433 4870 8443 4922
rect 8443 4870 8489 4922
rect 8513 4870 8559 4922
rect 8559 4870 8569 4922
rect 8593 4870 8623 4922
rect 8623 4870 8649 4922
rect 8353 4868 8409 4870
rect 8433 4868 8489 4870
rect 8513 4868 8569 4870
rect 8593 4868 8649 4870
rect 8353 3834 8409 3836
rect 8433 3834 8489 3836
rect 8513 3834 8569 3836
rect 8593 3834 8649 3836
rect 8353 3782 8379 3834
rect 8379 3782 8409 3834
rect 8433 3782 8443 3834
rect 8443 3782 8489 3834
rect 8513 3782 8559 3834
rect 8559 3782 8569 3834
rect 8593 3782 8623 3834
rect 8623 3782 8649 3834
rect 8353 3780 8409 3782
rect 8433 3780 8489 3782
rect 8513 3780 8569 3782
rect 8593 3780 8649 3782
rect 8353 2746 8409 2748
rect 8433 2746 8489 2748
rect 8513 2746 8569 2748
rect 8593 2746 8649 2748
rect 8353 2694 8379 2746
rect 8379 2694 8409 2746
rect 8433 2694 8443 2746
rect 8443 2694 8489 2746
rect 8513 2694 8559 2746
rect 8559 2694 8569 2746
rect 8593 2694 8623 2746
rect 8623 2694 8649 2746
rect 8353 2692 8409 2694
rect 8433 2692 8489 2694
rect 8513 2692 8569 2694
rect 8593 2692 8649 2694
rect 10414 6840 10470 6896
rect 10966 14864 11022 14920
rect 11058 14456 11114 14512
rect 11242 15952 11298 16008
rect 11150 14184 11206 14240
rect 11334 13504 11390 13560
rect 11058 12552 11114 12608
rect 10874 10648 10930 10704
rect 11518 12144 11574 12200
rect 12052 21786 12108 21788
rect 12132 21786 12188 21788
rect 12212 21786 12268 21788
rect 12292 21786 12348 21788
rect 12052 21734 12078 21786
rect 12078 21734 12108 21786
rect 12132 21734 12142 21786
rect 12142 21734 12188 21786
rect 12212 21734 12258 21786
rect 12258 21734 12268 21786
rect 12292 21734 12322 21786
rect 12322 21734 12348 21786
rect 12052 21732 12108 21734
rect 12132 21732 12188 21734
rect 12212 21732 12268 21734
rect 12292 21732 12348 21734
rect 11794 18672 11850 18728
rect 12052 20698 12108 20700
rect 12132 20698 12188 20700
rect 12212 20698 12268 20700
rect 12292 20698 12348 20700
rect 12052 20646 12078 20698
rect 12078 20646 12108 20698
rect 12132 20646 12142 20698
rect 12142 20646 12188 20698
rect 12212 20646 12258 20698
rect 12258 20646 12268 20698
rect 12292 20646 12322 20698
rect 12322 20646 12348 20698
rect 12052 20644 12108 20646
rect 12132 20644 12188 20646
rect 12212 20644 12268 20646
rect 12292 20644 12348 20646
rect 12052 19610 12108 19612
rect 12132 19610 12188 19612
rect 12212 19610 12268 19612
rect 12292 19610 12348 19612
rect 12052 19558 12078 19610
rect 12078 19558 12108 19610
rect 12132 19558 12142 19610
rect 12142 19558 12188 19610
rect 12212 19558 12258 19610
rect 12258 19558 12268 19610
rect 12292 19558 12322 19610
rect 12322 19558 12348 19610
rect 12052 19556 12108 19558
rect 12132 19556 12188 19558
rect 12212 19556 12268 19558
rect 12292 19556 12348 19558
rect 11794 17992 11850 18048
rect 11702 16224 11758 16280
rect 12070 18692 12126 18728
rect 12070 18672 12072 18692
rect 12072 18672 12124 18692
rect 12124 18672 12126 18692
rect 12052 18522 12108 18524
rect 12132 18522 12188 18524
rect 12212 18522 12268 18524
rect 12292 18522 12348 18524
rect 12052 18470 12078 18522
rect 12078 18470 12108 18522
rect 12132 18470 12142 18522
rect 12142 18470 12188 18522
rect 12212 18470 12258 18522
rect 12258 18470 12268 18522
rect 12292 18470 12322 18522
rect 12322 18470 12348 18522
rect 12052 18468 12108 18470
rect 12132 18468 12188 18470
rect 12212 18468 12268 18470
rect 12292 18468 12348 18470
rect 12530 17604 12586 17640
rect 12530 17584 12532 17604
rect 12532 17584 12584 17604
rect 12584 17584 12586 17604
rect 12052 17434 12108 17436
rect 12132 17434 12188 17436
rect 12212 17434 12268 17436
rect 12292 17434 12348 17436
rect 12052 17382 12078 17434
rect 12078 17382 12108 17434
rect 12132 17382 12142 17434
rect 12142 17382 12188 17434
rect 12212 17382 12258 17434
rect 12258 17382 12268 17434
rect 12292 17382 12322 17434
rect 12322 17382 12348 17434
rect 12052 17380 12108 17382
rect 12132 17380 12188 17382
rect 12212 17380 12268 17382
rect 12292 17380 12348 17382
rect 12438 17312 12494 17368
rect 11978 17076 11980 17096
rect 11980 17076 12032 17096
rect 12032 17076 12034 17096
rect 11978 17040 12034 17076
rect 12438 17076 12440 17096
rect 12440 17076 12492 17096
rect 12492 17076 12494 17096
rect 12438 17040 12494 17076
rect 12438 16360 12494 16416
rect 12052 16346 12108 16348
rect 12132 16346 12188 16348
rect 12212 16346 12268 16348
rect 12292 16346 12348 16348
rect 12052 16294 12078 16346
rect 12078 16294 12108 16346
rect 12132 16294 12142 16346
rect 12142 16294 12188 16346
rect 12212 16294 12258 16346
rect 12258 16294 12268 16346
rect 12292 16294 12322 16346
rect 12322 16294 12348 16346
rect 12052 16292 12108 16294
rect 12132 16292 12188 16294
rect 12212 16292 12268 16294
rect 12292 16292 12348 16294
rect 11794 15000 11850 15056
rect 11702 14864 11758 14920
rect 12052 15258 12108 15260
rect 12132 15258 12188 15260
rect 12212 15258 12268 15260
rect 12292 15258 12348 15260
rect 12052 15206 12078 15258
rect 12078 15206 12108 15258
rect 12132 15206 12142 15258
rect 12142 15206 12188 15258
rect 12212 15206 12258 15258
rect 12258 15206 12268 15258
rect 12292 15206 12322 15258
rect 12322 15206 12348 15258
rect 12052 15204 12108 15206
rect 12132 15204 12188 15206
rect 12212 15204 12268 15206
rect 12292 15204 12348 15206
rect 12346 15000 12402 15056
rect 11978 14728 12034 14784
rect 12052 14170 12108 14172
rect 12132 14170 12188 14172
rect 12212 14170 12268 14172
rect 12292 14170 12348 14172
rect 12052 14118 12078 14170
rect 12078 14118 12108 14170
rect 12132 14118 12142 14170
rect 12142 14118 12188 14170
rect 12212 14118 12258 14170
rect 12258 14118 12268 14170
rect 12292 14118 12322 14170
rect 12322 14118 12348 14170
rect 12052 14116 12108 14118
rect 12132 14116 12188 14118
rect 12212 14116 12268 14118
rect 12292 14116 12348 14118
rect 12070 13504 12126 13560
rect 12530 15136 12586 15192
rect 11886 13096 11942 13152
rect 12052 13082 12108 13084
rect 12132 13082 12188 13084
rect 12212 13082 12268 13084
rect 12292 13082 12348 13084
rect 12052 13030 12078 13082
rect 12078 13030 12108 13082
rect 12132 13030 12142 13082
rect 12142 13030 12188 13082
rect 12212 13030 12258 13082
rect 12258 13030 12268 13082
rect 12292 13030 12322 13082
rect 12322 13030 12348 13082
rect 12052 13028 12108 13030
rect 12132 13028 12188 13030
rect 12212 13028 12268 13030
rect 12292 13028 12348 13030
rect 12990 20032 13046 20088
rect 13082 19216 13138 19272
rect 12990 18672 13046 18728
rect 12714 16496 12770 16552
rect 12898 17176 12954 17232
rect 13174 17992 13230 18048
rect 12990 16244 13046 16280
rect 12990 16224 12992 16244
rect 12992 16224 13044 16244
rect 13044 16224 13046 16244
rect 12898 15952 12954 16008
rect 12806 15680 12862 15736
rect 12806 15272 12862 15328
rect 12806 14864 12862 14920
rect 12898 14184 12954 14240
rect 13358 17448 13414 17504
rect 13082 13504 13138 13560
rect 12052 11994 12108 11996
rect 12132 11994 12188 11996
rect 12212 11994 12268 11996
rect 12292 11994 12348 11996
rect 12052 11942 12078 11994
rect 12078 11942 12108 11994
rect 12132 11942 12142 11994
rect 12142 11942 12188 11994
rect 12212 11942 12258 11994
rect 12258 11942 12268 11994
rect 12292 11942 12322 11994
rect 12322 11942 12348 11994
rect 12052 11940 12108 11942
rect 12132 11940 12188 11942
rect 12212 11940 12268 11942
rect 12292 11940 12348 11942
rect 12052 10906 12108 10908
rect 12132 10906 12188 10908
rect 12212 10906 12268 10908
rect 12292 10906 12348 10908
rect 12052 10854 12078 10906
rect 12078 10854 12108 10906
rect 12132 10854 12142 10906
rect 12142 10854 12188 10906
rect 12212 10854 12258 10906
rect 12258 10854 12268 10906
rect 12292 10854 12322 10906
rect 12322 10854 12348 10906
rect 12052 10852 12108 10854
rect 12132 10852 12188 10854
rect 12212 10852 12268 10854
rect 12292 10852 12348 10854
rect 11518 10240 11574 10296
rect 12990 10784 13046 10840
rect 12052 9818 12108 9820
rect 12132 9818 12188 9820
rect 12212 9818 12268 9820
rect 12292 9818 12348 9820
rect 12052 9766 12078 9818
rect 12078 9766 12108 9818
rect 12132 9766 12142 9818
rect 12142 9766 12188 9818
rect 12212 9766 12258 9818
rect 12258 9766 12268 9818
rect 12292 9766 12322 9818
rect 12322 9766 12348 9818
rect 12052 9764 12108 9766
rect 12132 9764 12188 9766
rect 12212 9764 12268 9766
rect 12292 9764 12348 9766
rect 11886 9424 11942 9480
rect 10874 6976 10930 7032
rect 11058 7928 11114 7984
rect 10874 6452 10930 6488
rect 10874 6432 10876 6452
rect 10876 6432 10928 6452
rect 10928 6432 10930 6452
rect 11242 6160 11298 6216
rect 11610 8608 11666 8664
rect 12052 8730 12108 8732
rect 12132 8730 12188 8732
rect 12212 8730 12268 8732
rect 12292 8730 12348 8732
rect 12052 8678 12078 8730
rect 12078 8678 12108 8730
rect 12132 8678 12142 8730
rect 12142 8678 12188 8730
rect 12212 8678 12258 8730
rect 12258 8678 12268 8730
rect 12292 8678 12322 8730
rect 12322 8678 12348 8730
rect 12052 8676 12108 8678
rect 12132 8676 12188 8678
rect 12212 8676 12268 8678
rect 12292 8676 12348 8678
rect 13818 20576 13874 20632
rect 14002 20440 14058 20496
rect 14278 19624 14334 19680
rect 14278 19216 14334 19272
rect 14186 17720 14242 17776
rect 14554 19488 14610 19544
rect 14278 15272 14334 15328
rect 12990 7792 13046 7848
rect 12052 7642 12108 7644
rect 12132 7642 12188 7644
rect 12212 7642 12268 7644
rect 12292 7642 12348 7644
rect 12052 7590 12078 7642
rect 12078 7590 12108 7642
rect 12132 7590 12142 7642
rect 12142 7590 12188 7642
rect 12212 7590 12258 7642
rect 12258 7590 12268 7642
rect 12292 7590 12322 7642
rect 12322 7590 12348 7642
rect 12052 7588 12108 7590
rect 12132 7588 12188 7590
rect 12212 7588 12268 7590
rect 12292 7588 12348 7590
rect 12438 7520 12494 7576
rect 11518 6024 11574 6080
rect 11702 6296 11758 6352
rect 11610 4528 11666 4584
rect 12052 6554 12108 6556
rect 12132 6554 12188 6556
rect 12212 6554 12268 6556
rect 12292 6554 12348 6556
rect 12052 6502 12078 6554
rect 12078 6502 12108 6554
rect 12132 6502 12142 6554
rect 12142 6502 12188 6554
rect 12212 6502 12258 6554
rect 12258 6502 12268 6554
rect 12292 6502 12322 6554
rect 12322 6502 12348 6554
rect 12052 6500 12108 6502
rect 12132 6500 12188 6502
rect 12212 6500 12268 6502
rect 12292 6500 12348 6502
rect 12254 5616 12310 5672
rect 10322 3576 10378 3632
rect 12052 5466 12108 5468
rect 12132 5466 12188 5468
rect 12212 5466 12268 5468
rect 12292 5466 12348 5468
rect 12052 5414 12078 5466
rect 12078 5414 12108 5466
rect 12132 5414 12142 5466
rect 12142 5414 12188 5466
rect 12212 5414 12258 5466
rect 12258 5414 12268 5466
rect 12292 5414 12322 5466
rect 12322 5414 12348 5466
rect 12052 5412 12108 5414
rect 12132 5412 12188 5414
rect 12212 5412 12268 5414
rect 12292 5412 12348 5414
rect 12254 5108 12256 5128
rect 12256 5108 12308 5128
rect 12308 5108 12310 5128
rect 12254 5072 12310 5108
rect 12052 4378 12108 4380
rect 12132 4378 12188 4380
rect 12212 4378 12268 4380
rect 12292 4378 12348 4380
rect 12052 4326 12078 4378
rect 12078 4326 12108 4378
rect 12132 4326 12142 4378
rect 12142 4326 12188 4378
rect 12212 4326 12258 4378
rect 12258 4326 12268 4378
rect 12292 4326 12322 4378
rect 12322 4326 12348 4378
rect 12052 4324 12108 4326
rect 12132 4324 12188 4326
rect 12212 4324 12268 4326
rect 12292 4324 12348 4326
rect 12990 7384 13046 7440
rect 12052 3290 12108 3292
rect 12132 3290 12188 3292
rect 12212 3290 12268 3292
rect 12292 3290 12348 3292
rect 12052 3238 12078 3290
rect 12078 3238 12108 3290
rect 12132 3238 12142 3290
rect 12142 3238 12188 3290
rect 12212 3238 12258 3290
rect 12258 3238 12268 3290
rect 12292 3238 12322 3290
rect 12322 3238 12348 3290
rect 12052 3236 12108 3238
rect 12132 3236 12188 3238
rect 12212 3236 12268 3238
rect 12292 3236 12348 3238
rect 13450 8780 13452 8800
rect 13452 8780 13504 8800
rect 13504 8780 13506 8800
rect 13450 8744 13506 8780
rect 13358 8200 13414 8256
rect 14186 14456 14242 14512
rect 14186 13640 14242 13696
rect 13910 10956 13912 10976
rect 13912 10956 13964 10976
rect 13964 10956 13966 10976
rect 13910 10920 13966 10956
rect 14278 12280 14334 12336
rect 14370 11872 14426 11928
rect 13726 8200 13782 8256
rect 13358 7384 13414 7440
rect 13358 6976 13414 7032
rect 13634 6568 13690 6624
rect 14186 10376 14242 10432
rect 14186 9832 14242 9888
rect 13910 6704 13966 6760
rect 14370 9968 14426 10024
rect 15290 19352 15346 19408
rect 15106 18536 15162 18592
rect 14922 17176 14978 17232
rect 15750 21242 15806 21244
rect 15830 21242 15886 21244
rect 15910 21242 15966 21244
rect 15990 21242 16046 21244
rect 15750 21190 15776 21242
rect 15776 21190 15806 21242
rect 15830 21190 15840 21242
rect 15840 21190 15886 21242
rect 15910 21190 15956 21242
rect 15956 21190 15966 21242
rect 15990 21190 16020 21242
rect 16020 21190 16046 21242
rect 15750 21188 15806 21190
rect 15830 21188 15886 21190
rect 15910 21188 15966 21190
rect 15990 21188 16046 21190
rect 15750 20154 15806 20156
rect 15830 20154 15886 20156
rect 15910 20154 15966 20156
rect 15990 20154 16046 20156
rect 15750 20102 15776 20154
rect 15776 20102 15806 20154
rect 15830 20102 15840 20154
rect 15840 20102 15886 20154
rect 15910 20102 15956 20154
rect 15956 20102 15966 20154
rect 15990 20102 16020 20154
rect 16020 20102 16046 20154
rect 15750 20100 15806 20102
rect 15830 20100 15886 20102
rect 15910 20100 15966 20102
rect 15990 20100 16046 20102
rect 16026 19624 16082 19680
rect 16762 19488 16818 19544
rect 15750 19066 15806 19068
rect 15830 19066 15886 19068
rect 15910 19066 15966 19068
rect 15990 19066 16046 19068
rect 15750 19014 15776 19066
rect 15776 19014 15806 19066
rect 15830 19014 15840 19066
rect 15840 19014 15886 19066
rect 15910 19014 15956 19066
rect 15956 19014 15966 19066
rect 15990 19014 16020 19066
rect 16020 19014 16046 19066
rect 15750 19012 15806 19014
rect 15830 19012 15886 19014
rect 15910 19012 15966 19014
rect 15990 19012 16046 19014
rect 16026 18808 16082 18864
rect 15750 18708 15752 18728
rect 15752 18708 15804 18728
rect 15804 18708 15806 18728
rect 15750 18672 15806 18708
rect 14738 15816 14794 15872
rect 15106 15680 15162 15736
rect 14830 15136 14886 15192
rect 15198 15136 15254 15192
rect 14922 13096 14978 13152
rect 14830 12552 14886 12608
rect 14646 12044 14648 12064
rect 14648 12044 14700 12064
rect 14700 12044 14702 12064
rect 14646 12008 14702 12044
rect 14830 11056 14886 11112
rect 14646 10240 14702 10296
rect 14646 9152 14702 9208
rect 14370 6432 14426 6488
rect 14186 5752 14242 5808
rect 13818 5108 13820 5128
rect 13820 5108 13872 5128
rect 13872 5108 13874 5128
rect 13818 5072 13874 5108
rect 13174 4020 13176 4040
rect 13176 4020 13228 4040
rect 13228 4020 13230 4040
rect 13174 3984 13230 4020
rect 13174 3884 13176 3904
rect 13176 3884 13228 3904
rect 13228 3884 13230 3904
rect 13174 3848 13230 3884
rect 13542 3168 13598 3224
rect 14370 5244 14372 5264
rect 14372 5244 14424 5264
rect 14424 5244 14426 5264
rect 14370 5208 14426 5244
rect 14370 5072 14426 5128
rect 15290 14728 15346 14784
rect 15474 14728 15530 14784
rect 15750 17978 15806 17980
rect 15830 17978 15886 17980
rect 15910 17978 15966 17980
rect 15990 17978 16046 17980
rect 15750 17926 15776 17978
rect 15776 17926 15806 17978
rect 15830 17926 15840 17978
rect 15840 17926 15886 17978
rect 15910 17926 15956 17978
rect 15956 17926 15966 17978
rect 15990 17926 16020 17978
rect 16020 17926 16046 17978
rect 15750 17924 15806 17926
rect 15830 17924 15886 17926
rect 15910 17924 15966 17926
rect 15990 17924 16046 17926
rect 15750 16890 15806 16892
rect 15830 16890 15886 16892
rect 15910 16890 15966 16892
rect 15990 16890 16046 16892
rect 15750 16838 15776 16890
rect 15776 16838 15806 16890
rect 15830 16838 15840 16890
rect 15840 16838 15886 16890
rect 15910 16838 15956 16890
rect 15956 16838 15966 16890
rect 15990 16838 16020 16890
rect 16020 16838 16046 16890
rect 15750 16836 15806 16838
rect 15830 16836 15886 16838
rect 15910 16836 15966 16838
rect 15990 16836 16046 16838
rect 15842 16224 15898 16280
rect 16118 16496 16174 16552
rect 16026 15952 16082 16008
rect 15750 15802 15806 15804
rect 15830 15802 15886 15804
rect 15910 15802 15966 15804
rect 15990 15802 16046 15804
rect 15750 15750 15776 15802
rect 15776 15750 15806 15802
rect 15830 15750 15840 15802
rect 15840 15750 15886 15802
rect 15910 15750 15956 15802
rect 15956 15750 15966 15802
rect 15990 15750 16020 15802
rect 16020 15750 16046 15802
rect 15750 15748 15806 15750
rect 15830 15748 15886 15750
rect 15910 15748 15966 15750
rect 15990 15748 16046 15750
rect 15750 15408 15806 15464
rect 15750 15272 15806 15328
rect 15934 15136 15990 15192
rect 16026 14864 16082 14920
rect 16302 18672 16358 18728
rect 16486 18944 16542 19000
rect 16578 18400 16634 18456
rect 16302 16360 16358 16416
rect 15750 14714 15806 14716
rect 15830 14714 15886 14716
rect 15910 14714 15966 14716
rect 15990 14714 16046 14716
rect 15750 14662 15776 14714
rect 15776 14662 15806 14714
rect 15830 14662 15840 14714
rect 15840 14662 15886 14714
rect 15910 14662 15956 14714
rect 15956 14662 15966 14714
rect 15990 14662 16020 14714
rect 16020 14662 16046 14714
rect 15750 14660 15806 14662
rect 15830 14660 15886 14662
rect 15910 14660 15966 14662
rect 15990 14660 16046 14662
rect 16026 14184 16082 14240
rect 16026 14048 16082 14104
rect 16302 14048 16358 14104
rect 15750 13626 15806 13628
rect 15830 13626 15886 13628
rect 15910 13626 15966 13628
rect 15990 13626 16046 13628
rect 15750 13574 15776 13626
rect 15776 13574 15806 13626
rect 15830 13574 15840 13626
rect 15840 13574 15886 13626
rect 15910 13574 15956 13626
rect 15956 13574 15966 13626
rect 15990 13574 16020 13626
rect 16020 13574 16046 13626
rect 15750 13572 15806 13574
rect 15830 13572 15886 13574
rect 15910 13572 15966 13574
rect 15990 13572 16046 13574
rect 15658 12960 15714 13016
rect 15750 12538 15806 12540
rect 15830 12538 15886 12540
rect 15910 12538 15966 12540
rect 15990 12538 16046 12540
rect 15750 12486 15776 12538
rect 15776 12486 15806 12538
rect 15830 12486 15840 12538
rect 15840 12486 15886 12538
rect 15910 12486 15956 12538
rect 15956 12486 15966 12538
rect 15990 12486 16020 12538
rect 16020 12486 16046 12538
rect 15750 12484 15806 12486
rect 15830 12484 15886 12486
rect 15910 12484 15966 12486
rect 15990 12484 16046 12486
rect 15750 11450 15806 11452
rect 15830 11450 15886 11452
rect 15910 11450 15966 11452
rect 15990 11450 16046 11452
rect 15750 11398 15776 11450
rect 15776 11398 15806 11450
rect 15830 11398 15840 11450
rect 15840 11398 15886 11450
rect 15910 11398 15956 11450
rect 15956 11398 15966 11450
rect 15990 11398 16020 11450
rect 16020 11398 16046 11450
rect 15750 11396 15806 11398
rect 15830 11396 15886 11398
rect 15910 11396 15966 11398
rect 15990 11396 16046 11398
rect 15658 11212 15714 11248
rect 15658 11192 15660 11212
rect 15660 11192 15712 11212
rect 15712 11192 15714 11212
rect 15382 10240 15438 10296
rect 15750 10362 15806 10364
rect 15830 10362 15886 10364
rect 15910 10362 15966 10364
rect 15990 10362 16046 10364
rect 15750 10310 15776 10362
rect 15776 10310 15806 10362
rect 15830 10310 15840 10362
rect 15840 10310 15886 10362
rect 15910 10310 15956 10362
rect 15956 10310 15966 10362
rect 15990 10310 16020 10362
rect 16020 10310 16046 10362
rect 15750 10308 15806 10310
rect 15830 10308 15886 10310
rect 15910 10308 15966 10310
rect 15990 10308 16046 10310
rect 15198 9832 15254 9888
rect 14922 7248 14978 7304
rect 15014 6432 15070 6488
rect 14830 5208 14886 5264
rect 14922 4392 14978 4448
rect 16210 13504 16266 13560
rect 16486 17176 16542 17232
rect 16762 17756 16764 17776
rect 16764 17756 16816 17776
rect 16816 17756 16818 17776
rect 16762 17720 16818 17756
rect 17222 20440 17278 20496
rect 17130 18672 17186 18728
rect 17130 17176 17186 17232
rect 16762 16360 16818 16416
rect 16670 15952 16726 16008
rect 16578 15272 16634 15328
rect 16578 15136 16634 15192
rect 16762 13912 16818 13968
rect 16394 13640 16450 13696
rect 16210 12552 16266 12608
rect 16302 12008 16358 12064
rect 16302 11464 16358 11520
rect 15566 9696 15622 9752
rect 16118 9560 16174 9616
rect 15750 9274 15806 9276
rect 15830 9274 15886 9276
rect 15910 9274 15966 9276
rect 15990 9274 16046 9276
rect 15750 9222 15776 9274
rect 15776 9222 15806 9274
rect 15830 9222 15840 9274
rect 15840 9222 15886 9274
rect 15910 9222 15956 9274
rect 15956 9222 15966 9274
rect 15990 9222 16020 9274
rect 16020 9222 16046 9274
rect 15750 9220 15806 9222
rect 15830 9220 15886 9222
rect 15910 9220 15966 9222
rect 15990 9220 16046 9222
rect 15382 8200 15438 8256
rect 15382 8084 15438 8120
rect 15382 8064 15384 8084
rect 15384 8064 15436 8084
rect 15436 8064 15438 8084
rect 16118 9016 16174 9072
rect 15750 8608 15806 8664
rect 15750 8186 15806 8188
rect 15830 8186 15886 8188
rect 15910 8186 15966 8188
rect 15990 8186 16046 8188
rect 15750 8134 15776 8186
rect 15776 8134 15806 8186
rect 15830 8134 15840 8186
rect 15840 8134 15886 8186
rect 15910 8134 15956 8186
rect 15956 8134 15966 8186
rect 15990 8134 16020 8186
rect 16020 8134 16046 8186
rect 15750 8132 15806 8134
rect 15830 8132 15886 8134
rect 15910 8132 15966 8134
rect 15990 8132 16046 8134
rect 12052 2202 12108 2204
rect 12132 2202 12188 2204
rect 12212 2202 12268 2204
rect 12292 2202 12348 2204
rect 12052 2150 12078 2202
rect 12078 2150 12108 2202
rect 12132 2150 12142 2202
rect 12142 2150 12188 2202
rect 12212 2150 12258 2202
rect 12258 2150 12268 2202
rect 12292 2150 12322 2202
rect 12322 2150 12348 2202
rect 12052 2148 12108 2150
rect 12132 2148 12188 2150
rect 12212 2148 12268 2150
rect 12292 2148 12348 2150
rect 17038 16360 17094 16416
rect 16854 12416 16910 12472
rect 16670 12008 16726 12064
rect 16762 11212 16818 11248
rect 16762 11192 16764 11212
rect 16764 11192 16816 11212
rect 16816 11192 16818 11212
rect 16670 10648 16726 10704
rect 16854 10648 16910 10704
rect 16394 9016 16450 9072
rect 16486 8744 16542 8800
rect 16210 7384 16266 7440
rect 15750 7248 15806 7304
rect 15750 7098 15806 7100
rect 15830 7098 15886 7100
rect 15910 7098 15966 7100
rect 15990 7098 16046 7100
rect 15750 7046 15776 7098
rect 15776 7046 15806 7098
rect 15830 7046 15840 7098
rect 15840 7046 15886 7098
rect 15910 7046 15956 7098
rect 15956 7046 15966 7098
rect 15990 7046 16020 7098
rect 16020 7046 16046 7098
rect 15750 7044 15806 7046
rect 15830 7044 15886 7046
rect 15910 7044 15966 7046
rect 15990 7044 16046 7046
rect 16670 7520 16726 7576
rect 16118 6432 16174 6488
rect 15750 6010 15806 6012
rect 15830 6010 15886 6012
rect 15910 6010 15966 6012
rect 15990 6010 16046 6012
rect 15750 5958 15776 6010
rect 15776 5958 15806 6010
rect 15830 5958 15840 6010
rect 15840 5958 15886 6010
rect 15910 5958 15956 6010
rect 15956 5958 15966 6010
rect 15990 5958 16020 6010
rect 16020 5958 16046 6010
rect 15750 5956 15806 5958
rect 15830 5956 15886 5958
rect 15910 5956 15966 5958
rect 15990 5956 16046 5958
rect 16486 6840 16542 6896
rect 16302 5752 16358 5808
rect 15750 4922 15806 4924
rect 15830 4922 15886 4924
rect 15910 4922 15966 4924
rect 15990 4922 16046 4924
rect 15750 4870 15776 4922
rect 15776 4870 15806 4922
rect 15830 4870 15840 4922
rect 15840 4870 15886 4922
rect 15910 4870 15956 4922
rect 15956 4870 15966 4922
rect 15990 4870 16020 4922
rect 16020 4870 16046 4922
rect 15750 4868 15806 4870
rect 15830 4868 15886 4870
rect 15910 4868 15966 4870
rect 15990 4868 16046 4870
rect 16118 4120 16174 4176
rect 15750 3834 15806 3836
rect 15830 3834 15886 3836
rect 15910 3834 15966 3836
rect 15990 3834 16046 3836
rect 15750 3782 15776 3834
rect 15776 3782 15806 3834
rect 15830 3782 15840 3834
rect 15840 3782 15886 3834
rect 15910 3782 15956 3834
rect 15956 3782 15966 3834
rect 15990 3782 16020 3834
rect 16020 3782 16046 3834
rect 15750 3780 15806 3782
rect 15830 3780 15886 3782
rect 15910 3780 15966 3782
rect 15990 3780 16046 3782
rect 15750 2746 15806 2748
rect 15830 2746 15886 2748
rect 15910 2746 15966 2748
rect 15990 2746 16046 2748
rect 15750 2694 15776 2746
rect 15776 2694 15806 2746
rect 15830 2694 15840 2746
rect 15840 2694 15886 2746
rect 15910 2694 15956 2746
rect 15956 2694 15966 2746
rect 15990 2694 16020 2746
rect 16020 2694 16046 2746
rect 15750 2692 15806 2694
rect 15830 2692 15886 2694
rect 15910 2692 15966 2694
rect 15990 2692 16046 2694
rect 15934 2508 15990 2544
rect 15934 2488 15936 2508
rect 15936 2488 15988 2508
rect 15988 2488 15990 2508
rect 17314 14456 17370 14512
rect 17314 13640 17370 13696
rect 17130 13096 17186 13152
rect 17314 13232 17370 13288
rect 17222 12144 17278 12200
rect 17130 9968 17186 10024
rect 17038 8880 17094 8936
rect 17498 12844 17554 12880
rect 17498 12824 17500 12844
rect 17500 12824 17552 12844
rect 17552 12824 17554 12844
rect 17314 11736 17370 11792
rect 17314 11328 17370 11384
rect 17682 15272 17738 15328
rect 18234 20576 18290 20632
rect 18142 19760 18198 19816
rect 17958 17040 18014 17096
rect 18142 16904 18198 16960
rect 17866 15680 17922 15736
rect 18050 14048 18106 14104
rect 17958 13232 18014 13288
rect 17774 13096 17830 13152
rect 17590 12416 17646 12472
rect 17682 11328 17738 11384
rect 17406 9288 17462 9344
rect 17314 9152 17370 9208
rect 17038 8064 17094 8120
rect 16946 6296 17002 6352
rect 16946 4936 17002 4992
rect 17682 6024 17738 6080
rect 17958 12144 18014 12200
rect 17866 12008 17922 12064
rect 18510 20032 18566 20088
rect 18326 18944 18382 19000
rect 18234 13504 18290 13560
rect 18234 11600 18290 11656
rect 17958 11056 18014 11112
rect 17866 8608 17922 8664
rect 17866 8472 17922 8528
rect 17866 8236 17868 8256
rect 17868 8236 17920 8256
rect 17920 8236 17922 8256
rect 17866 8200 17922 8236
rect 18326 9968 18382 10024
rect 18326 9152 18382 9208
rect 17958 7248 18014 7304
rect 17958 6568 18014 6624
rect 19338 23296 19394 23352
rect 19798 22616 19854 22672
rect 18786 18944 18842 19000
rect 18510 16088 18566 16144
rect 18510 14456 18566 14512
rect 18510 12824 18566 12880
rect 18510 9424 18566 9480
rect 19449 21786 19505 21788
rect 19529 21786 19585 21788
rect 19609 21786 19665 21788
rect 19689 21786 19745 21788
rect 19449 21734 19475 21786
rect 19475 21734 19505 21786
rect 19529 21734 19539 21786
rect 19539 21734 19585 21786
rect 19609 21734 19655 21786
rect 19655 21734 19665 21786
rect 19689 21734 19719 21786
rect 19719 21734 19745 21786
rect 19449 21732 19505 21734
rect 19529 21732 19585 21734
rect 19609 21732 19665 21734
rect 19689 21732 19745 21734
rect 19338 21256 19394 21312
rect 19449 20698 19505 20700
rect 19529 20698 19585 20700
rect 19609 20698 19665 20700
rect 19689 20698 19745 20700
rect 19449 20646 19475 20698
rect 19475 20646 19505 20698
rect 19529 20646 19539 20698
rect 19539 20646 19585 20698
rect 19609 20646 19655 20698
rect 19655 20646 19665 20698
rect 19689 20646 19719 20698
rect 19719 20646 19745 20698
rect 19449 20644 19505 20646
rect 19529 20644 19585 20646
rect 19609 20644 19665 20646
rect 19689 20644 19745 20646
rect 20442 21936 20498 21992
rect 19890 20324 19946 20360
rect 19890 20304 19892 20324
rect 19892 20304 19944 20324
rect 19944 20304 19946 20324
rect 20166 20304 20222 20360
rect 19449 19610 19505 19612
rect 19529 19610 19585 19612
rect 19609 19610 19665 19612
rect 19689 19610 19745 19612
rect 19449 19558 19475 19610
rect 19475 19558 19505 19610
rect 19529 19558 19539 19610
rect 19539 19558 19585 19610
rect 19609 19558 19655 19610
rect 19655 19558 19665 19610
rect 19689 19558 19719 19610
rect 19719 19558 19745 19610
rect 19449 19556 19505 19558
rect 19529 19556 19585 19558
rect 19609 19556 19665 19558
rect 19689 19556 19745 19558
rect 20166 19760 20222 19816
rect 19154 18400 19210 18456
rect 19449 18522 19505 18524
rect 19529 18522 19585 18524
rect 19609 18522 19665 18524
rect 19689 18522 19745 18524
rect 19449 18470 19475 18522
rect 19475 18470 19505 18522
rect 19529 18470 19539 18522
rect 19539 18470 19585 18522
rect 19609 18470 19655 18522
rect 19655 18470 19665 18522
rect 19689 18470 19719 18522
rect 19719 18470 19745 18522
rect 19449 18468 19505 18470
rect 19529 18468 19585 18470
rect 19609 18468 19665 18470
rect 19689 18468 19745 18470
rect 18878 16496 18934 16552
rect 18786 15136 18842 15192
rect 18970 12960 19026 13016
rect 19062 12824 19118 12880
rect 18878 12008 18934 12064
rect 18878 11328 18934 11384
rect 18510 7656 18566 7712
rect 18694 7928 18750 7984
rect 18878 7948 18934 7984
rect 18878 7928 18880 7948
rect 18880 7928 18932 7948
rect 18932 7928 18934 7948
rect 18878 7792 18934 7848
rect 17866 5752 17922 5808
rect 18050 6024 18106 6080
rect 18142 5208 18198 5264
rect 17682 3168 17738 3224
rect 18694 5772 18750 5808
rect 18694 5752 18696 5772
rect 18696 5752 18748 5772
rect 18748 5752 18750 5772
rect 18694 5108 18696 5128
rect 18696 5108 18748 5128
rect 18748 5108 18750 5128
rect 18694 5072 18750 5108
rect 18694 4428 18696 4448
rect 18696 4428 18748 4448
rect 18748 4428 18750 4448
rect 18694 4392 18750 4428
rect 19522 17584 19578 17640
rect 19449 17434 19505 17436
rect 19529 17434 19585 17436
rect 19609 17434 19665 17436
rect 19689 17434 19745 17436
rect 19449 17382 19475 17434
rect 19475 17382 19505 17434
rect 19529 17382 19539 17434
rect 19539 17382 19585 17434
rect 19609 17382 19655 17434
rect 19655 17382 19665 17434
rect 19689 17382 19719 17434
rect 19719 17382 19745 17434
rect 19449 17380 19505 17382
rect 19529 17380 19585 17382
rect 19609 17380 19665 17382
rect 19689 17380 19745 17382
rect 19246 17040 19302 17096
rect 19449 16346 19505 16348
rect 19529 16346 19585 16348
rect 19609 16346 19665 16348
rect 19689 16346 19745 16348
rect 19449 16294 19475 16346
rect 19475 16294 19505 16346
rect 19529 16294 19539 16346
rect 19539 16294 19585 16346
rect 19609 16294 19655 16346
rect 19655 16294 19665 16346
rect 19689 16294 19719 16346
rect 19719 16294 19745 16346
rect 19449 16292 19505 16294
rect 19529 16292 19585 16294
rect 19609 16292 19665 16294
rect 19689 16292 19745 16294
rect 19246 16224 19302 16280
rect 19338 15408 19394 15464
rect 19449 15258 19505 15260
rect 19529 15258 19585 15260
rect 19609 15258 19665 15260
rect 19689 15258 19745 15260
rect 19449 15206 19475 15258
rect 19475 15206 19505 15258
rect 19529 15206 19539 15258
rect 19539 15206 19585 15258
rect 19609 15206 19655 15258
rect 19655 15206 19665 15258
rect 19689 15206 19719 15258
rect 19719 15206 19745 15258
rect 19449 15204 19505 15206
rect 19529 15204 19585 15206
rect 19609 15204 19665 15206
rect 19689 15204 19745 15206
rect 19338 14728 19394 14784
rect 19430 14476 19486 14512
rect 19430 14456 19432 14476
rect 19432 14456 19484 14476
rect 19484 14456 19486 14476
rect 19449 14170 19505 14172
rect 19529 14170 19585 14172
rect 19609 14170 19665 14172
rect 19689 14170 19745 14172
rect 19449 14118 19475 14170
rect 19475 14118 19505 14170
rect 19529 14118 19539 14170
rect 19539 14118 19585 14170
rect 19609 14118 19655 14170
rect 19655 14118 19665 14170
rect 19689 14118 19719 14170
rect 19719 14118 19745 14170
rect 19449 14116 19505 14118
rect 19529 14116 19585 14118
rect 19609 14116 19665 14118
rect 19689 14116 19745 14118
rect 19614 13504 19670 13560
rect 20166 18672 20222 18728
rect 20074 18400 20130 18456
rect 20166 18264 20222 18320
rect 19890 17720 19946 17776
rect 19890 17312 19946 17368
rect 19890 15680 19946 15736
rect 20258 17196 20314 17232
rect 20258 17176 20260 17196
rect 20260 17176 20312 17196
rect 20312 17176 20314 17196
rect 19449 13082 19505 13084
rect 19529 13082 19585 13084
rect 19609 13082 19665 13084
rect 19689 13082 19745 13084
rect 19449 13030 19475 13082
rect 19475 13030 19505 13082
rect 19529 13030 19539 13082
rect 19539 13030 19585 13082
rect 19609 13030 19655 13082
rect 19655 13030 19665 13082
rect 19689 13030 19719 13082
rect 19719 13030 19745 13082
rect 19449 13028 19505 13030
rect 19529 13028 19585 13030
rect 19609 13028 19665 13030
rect 19689 13028 19745 13030
rect 19890 13096 19946 13152
rect 20074 14864 20130 14920
rect 19338 12416 19394 12472
rect 19338 12280 19394 12336
rect 19246 11600 19302 11656
rect 19614 12144 19670 12200
rect 19449 11994 19505 11996
rect 19529 11994 19585 11996
rect 19609 11994 19665 11996
rect 19689 11994 19745 11996
rect 19449 11942 19475 11994
rect 19475 11942 19505 11994
rect 19529 11942 19539 11994
rect 19539 11942 19585 11994
rect 19609 11942 19655 11994
rect 19655 11942 19665 11994
rect 19689 11942 19719 11994
rect 19719 11942 19745 11994
rect 19449 11940 19505 11942
rect 19529 11940 19585 11942
rect 19609 11940 19665 11942
rect 19689 11940 19745 11942
rect 20074 12416 20130 12472
rect 19338 11464 19394 11520
rect 19449 10906 19505 10908
rect 19529 10906 19585 10908
rect 19609 10906 19665 10908
rect 19689 10906 19745 10908
rect 19449 10854 19475 10906
rect 19475 10854 19505 10906
rect 19529 10854 19539 10906
rect 19539 10854 19585 10906
rect 19609 10854 19655 10906
rect 19655 10854 19665 10906
rect 19689 10854 19719 10906
rect 19719 10854 19745 10906
rect 19449 10852 19505 10854
rect 19529 10852 19585 10854
rect 19609 10852 19665 10854
rect 19689 10852 19745 10854
rect 19246 10804 19302 10840
rect 19246 10784 19248 10804
rect 19248 10784 19300 10804
rect 19300 10784 19302 10804
rect 19614 10512 19670 10568
rect 19338 10104 19394 10160
rect 19449 9818 19505 9820
rect 19529 9818 19585 9820
rect 19609 9818 19665 9820
rect 19689 9818 19745 9820
rect 19449 9766 19475 9818
rect 19475 9766 19505 9818
rect 19529 9766 19539 9818
rect 19539 9766 19585 9818
rect 19609 9766 19655 9818
rect 19655 9766 19665 9818
rect 19689 9766 19719 9818
rect 19719 9766 19745 9818
rect 19449 9764 19505 9766
rect 19529 9764 19585 9766
rect 19609 9764 19665 9766
rect 19689 9764 19745 9766
rect 19449 8730 19505 8732
rect 19529 8730 19585 8732
rect 19609 8730 19665 8732
rect 19689 8730 19745 8732
rect 19449 8678 19475 8730
rect 19475 8678 19505 8730
rect 19529 8678 19539 8730
rect 19539 8678 19585 8730
rect 19609 8678 19655 8730
rect 19655 8678 19665 8730
rect 19689 8678 19719 8730
rect 19719 8678 19745 8730
rect 19449 8676 19505 8678
rect 19529 8676 19585 8678
rect 19609 8676 19665 8678
rect 19689 8676 19745 8678
rect 19062 8064 19118 8120
rect 19338 8336 19394 8392
rect 19338 8064 19394 8120
rect 19522 8336 19578 8392
rect 19706 7928 19762 7984
rect 19890 8200 19946 8256
rect 19798 7792 19854 7848
rect 19449 7642 19505 7644
rect 19529 7642 19585 7644
rect 19609 7642 19665 7644
rect 19689 7642 19745 7644
rect 19449 7590 19475 7642
rect 19475 7590 19505 7642
rect 19529 7590 19539 7642
rect 19539 7590 19585 7642
rect 19609 7590 19655 7642
rect 19655 7590 19665 7642
rect 19689 7590 19719 7642
rect 19719 7590 19745 7642
rect 19449 7588 19505 7590
rect 19529 7588 19585 7590
rect 19609 7588 19665 7590
rect 19689 7588 19745 7590
rect 19246 5616 19302 5672
rect 19449 6554 19505 6556
rect 19529 6554 19585 6556
rect 19609 6554 19665 6556
rect 19689 6554 19745 6556
rect 19449 6502 19475 6554
rect 19475 6502 19505 6554
rect 19529 6502 19539 6554
rect 19539 6502 19585 6554
rect 19609 6502 19655 6554
rect 19655 6502 19665 6554
rect 19689 6502 19719 6554
rect 19719 6502 19745 6554
rect 19449 6500 19505 6502
rect 19529 6500 19585 6502
rect 19609 6500 19665 6502
rect 19689 6500 19745 6502
rect 19449 5466 19505 5468
rect 19529 5466 19585 5468
rect 19609 5466 19665 5468
rect 19689 5466 19745 5468
rect 19449 5414 19475 5466
rect 19475 5414 19505 5466
rect 19529 5414 19539 5466
rect 19539 5414 19585 5466
rect 19609 5414 19655 5466
rect 19655 5414 19665 5466
rect 19689 5414 19719 5466
rect 19719 5414 19745 5466
rect 19449 5412 19505 5414
rect 19529 5412 19585 5414
rect 19609 5412 19665 5414
rect 19689 5412 19745 5414
rect 19890 6296 19946 6352
rect 19614 5228 19670 5264
rect 19614 5208 19616 5228
rect 19616 5208 19668 5228
rect 19668 5208 19670 5228
rect 19449 4378 19505 4380
rect 19529 4378 19585 4380
rect 19609 4378 19665 4380
rect 19689 4378 19745 4380
rect 19449 4326 19475 4378
rect 19475 4326 19505 4378
rect 19529 4326 19539 4378
rect 19539 4326 19585 4378
rect 19609 4326 19655 4378
rect 19655 4326 19665 4378
rect 19689 4326 19719 4378
rect 19719 4326 19745 4378
rect 19449 4324 19505 4326
rect 19529 4324 19585 4326
rect 19609 4324 19665 4326
rect 19689 4324 19745 4326
rect 19338 4120 19394 4176
rect 19449 3290 19505 3292
rect 19529 3290 19585 3292
rect 19609 3290 19665 3292
rect 19689 3290 19745 3292
rect 19449 3238 19475 3290
rect 19475 3238 19505 3290
rect 19529 3238 19539 3290
rect 19539 3238 19585 3290
rect 19609 3238 19655 3290
rect 19655 3238 19665 3290
rect 19689 3238 19719 3290
rect 19719 3238 19745 3290
rect 19449 3236 19505 3238
rect 19529 3236 19585 3238
rect 19609 3236 19665 3238
rect 19689 3236 19745 3238
rect 19890 2216 19946 2272
rect 19449 2202 19505 2204
rect 19529 2202 19585 2204
rect 19609 2202 19665 2204
rect 19689 2202 19745 2204
rect 19449 2150 19475 2202
rect 19475 2150 19505 2202
rect 19529 2150 19539 2202
rect 19539 2150 19585 2202
rect 19609 2150 19655 2202
rect 19655 2150 19665 2202
rect 19689 2150 19719 2202
rect 19719 2150 19745 2202
rect 19449 2148 19505 2150
rect 19529 2148 19585 2150
rect 19609 2148 19665 2150
rect 19689 2148 19745 2150
rect 20258 12552 20314 12608
rect 20166 12144 20222 12200
rect 20626 20576 20682 20632
rect 20534 19896 20590 19952
rect 21178 20848 21234 20904
rect 20902 19216 20958 19272
rect 20718 18672 20774 18728
rect 20994 17992 21050 18048
rect 20902 16632 20958 16688
rect 20626 15000 20682 15056
rect 20442 14592 20498 14648
rect 20626 14048 20682 14104
rect 20350 11872 20406 11928
rect 20718 12824 20774 12880
rect 20626 12416 20682 12472
rect 20902 13776 20958 13832
rect 20902 13388 20958 13424
rect 20902 13368 20904 13388
rect 20904 13368 20956 13388
rect 20956 13368 20958 13388
rect 20534 10784 20590 10840
rect 20350 9152 20406 9208
rect 20258 8608 20314 8664
rect 20074 7112 20130 7168
rect 20074 3576 20130 3632
rect 20350 6704 20406 6760
rect 20534 8200 20590 8256
rect 20350 5344 20406 5400
rect 20902 7520 20958 7576
rect 20902 5228 20958 5264
rect 20902 5208 20904 5228
rect 20904 5208 20956 5228
rect 20956 5208 20958 5228
rect 20718 4700 20720 4720
rect 20720 4700 20772 4720
rect 20772 4700 20774 4720
rect 20718 4664 20774 4700
rect 21362 17992 21418 18048
rect 21546 19624 21602 19680
rect 21638 19352 21694 19408
rect 21638 18028 21640 18048
rect 21640 18028 21692 18048
rect 21692 18028 21694 18048
rect 21638 17992 21694 18028
rect 21454 15544 21510 15600
rect 21270 13912 21326 13968
rect 21270 13504 21326 13560
rect 21362 12008 21418 12064
rect 21914 19760 21970 19816
rect 22374 20032 22430 20088
rect 22098 14320 22154 14376
rect 22006 10512 22062 10568
rect 21730 7248 21786 7304
rect 22374 13096 22430 13152
rect 22282 12280 22338 12336
rect 22282 11736 22338 11792
rect 22834 20032 22890 20088
rect 22834 19352 22890 19408
rect 22190 7384 22246 7440
rect 22098 4936 22154 4992
rect 22558 6160 22614 6216
rect 22190 4256 22246 4312
rect 22098 3440 22154 3496
rect 21362 1536 21418 1592
rect 23110 9560 23166 9616
rect 22834 8880 22890 8936
rect 22834 5480 22890 5536
rect 23386 6860 23442 6896
rect 23386 6840 23388 6860
rect 23388 6840 23440 6860
rect 23440 6840 23442 6860
rect 22926 856 22982 912
rect 21270 312 21326 368
<< metal3 >>
rect 19425 24034 19491 24037
rect 23600 24034 24400 24064
rect 19425 24032 24400 24034
rect 19425 23976 19430 24032
rect 19486 23976 24400 24032
rect 19425 23974 24400 23976
rect 19425 23971 19491 23974
rect 23600 23944 24400 23974
rect 19333 23354 19399 23357
rect 23600 23354 24400 23384
rect 19333 23352 24400 23354
rect 19333 23296 19338 23352
rect 19394 23296 24400 23352
rect 19333 23294 24400 23296
rect 19333 23291 19399 23294
rect 23600 23264 24400 23294
rect 19793 22674 19859 22677
rect 23600 22674 24400 22704
rect 19793 22672 24400 22674
rect 19793 22616 19798 22672
rect 19854 22616 24400 22672
rect 19793 22614 24400 22616
rect 19793 22611 19859 22614
rect 23600 22584 24400 22614
rect 6177 21994 6243 21997
rect 9673 21994 9739 21997
rect 6177 21992 9739 21994
rect 6177 21936 6182 21992
rect 6238 21936 9678 21992
rect 9734 21936 9739 21992
rect 6177 21934 9739 21936
rect 6177 21931 6243 21934
rect 9673 21931 9739 21934
rect 20437 21994 20503 21997
rect 23600 21994 24400 22024
rect 20437 21992 24400 21994
rect 20437 21936 20442 21992
rect 20498 21936 24400 21992
rect 20437 21934 24400 21936
rect 20437 21931 20503 21934
rect 23600 21904 24400 21934
rect 4642 21792 4962 21793
rect 4642 21728 4650 21792
rect 4714 21728 4730 21792
rect 4794 21728 4810 21792
rect 4874 21728 4890 21792
rect 4954 21728 4962 21792
rect 4642 21727 4962 21728
rect 12040 21792 12360 21793
rect 12040 21728 12048 21792
rect 12112 21728 12128 21792
rect 12192 21728 12208 21792
rect 12272 21728 12288 21792
rect 12352 21728 12360 21792
rect 12040 21727 12360 21728
rect 19437 21792 19757 21793
rect 19437 21728 19445 21792
rect 19509 21728 19525 21792
rect 19589 21728 19605 21792
rect 19669 21728 19685 21792
rect 19749 21728 19757 21792
rect 19437 21727 19757 21728
rect 6085 21586 6151 21589
rect 9029 21586 9095 21589
rect 6085 21584 9095 21586
rect 6085 21528 6090 21584
rect 6146 21528 9034 21584
rect 9090 21528 9095 21584
rect 6085 21526 9095 21528
rect 6085 21523 6151 21526
rect 9029 21523 9095 21526
rect 4337 21450 4403 21453
rect 8937 21450 9003 21453
rect 4337 21448 9003 21450
rect 4337 21392 4342 21448
rect 4398 21392 8942 21448
rect 8998 21392 9003 21448
rect 4337 21390 9003 21392
rect 4337 21387 4403 21390
rect 8937 21387 9003 21390
rect 0 21224 800 21344
rect 19333 21314 19399 21317
rect 23600 21314 24400 21344
rect 19333 21312 24400 21314
rect 19333 21256 19338 21312
rect 19394 21256 24400 21312
rect 19333 21254 24400 21256
rect 19333 21251 19399 21254
rect 8341 21248 8661 21249
rect 8341 21184 8349 21248
rect 8413 21184 8429 21248
rect 8493 21184 8509 21248
rect 8573 21184 8589 21248
rect 8653 21184 8661 21248
rect 8341 21183 8661 21184
rect 15738 21248 16058 21249
rect 15738 21184 15746 21248
rect 15810 21184 15826 21248
rect 15890 21184 15906 21248
rect 15970 21184 15986 21248
rect 16050 21184 16058 21248
rect 23600 21224 24400 21254
rect 15738 21183 16058 21184
rect 10501 20906 10567 20909
rect 13118 20906 13124 20908
rect 10501 20904 13124 20906
rect 10501 20848 10506 20904
rect 10562 20848 13124 20904
rect 10501 20846 13124 20848
rect 10501 20843 10567 20846
rect 13118 20844 13124 20846
rect 13188 20844 13194 20908
rect 13302 20844 13308 20908
rect 13372 20906 13378 20908
rect 21173 20906 21239 20909
rect 13372 20904 21239 20906
rect 13372 20848 21178 20904
rect 21234 20848 21239 20904
rect 13372 20846 21239 20848
rect 13372 20844 13378 20846
rect 21173 20843 21239 20846
rect 4642 20704 4962 20705
rect 4642 20640 4650 20704
rect 4714 20640 4730 20704
rect 4794 20640 4810 20704
rect 4874 20640 4890 20704
rect 4954 20640 4962 20704
rect 4642 20639 4962 20640
rect 12040 20704 12360 20705
rect 12040 20640 12048 20704
rect 12112 20640 12128 20704
rect 12192 20640 12208 20704
rect 12272 20640 12288 20704
rect 12352 20640 12360 20704
rect 12040 20639 12360 20640
rect 19437 20704 19757 20705
rect 19437 20640 19445 20704
rect 19509 20640 19525 20704
rect 19589 20640 19605 20704
rect 19669 20640 19685 20704
rect 19749 20640 19757 20704
rect 19437 20639 19757 20640
rect 13813 20634 13879 20637
rect 18229 20634 18295 20637
rect 12574 20632 18295 20634
rect 12574 20576 13818 20632
rect 13874 20576 18234 20632
rect 18290 20576 18295 20632
rect 12574 20574 18295 20576
rect 10409 20498 10475 20501
rect 12574 20498 12634 20574
rect 13813 20571 13879 20574
rect 18229 20571 18295 20574
rect 20621 20634 20687 20637
rect 23600 20634 24400 20664
rect 20621 20632 24400 20634
rect 20621 20576 20626 20632
rect 20682 20576 24400 20632
rect 20621 20574 24400 20576
rect 20621 20571 20687 20574
rect 23600 20544 24400 20574
rect 10409 20496 12634 20498
rect 10409 20440 10414 20496
rect 10470 20440 12634 20496
rect 10409 20438 12634 20440
rect 13997 20498 14063 20501
rect 17217 20498 17283 20501
rect 13997 20496 17283 20498
rect 13997 20440 14002 20496
rect 14058 20440 17222 20496
rect 17278 20440 17283 20496
rect 13997 20438 17283 20440
rect 10409 20435 10475 20438
rect 13997 20435 14063 20438
rect 17217 20435 17283 20438
rect 7005 20362 7071 20365
rect 8845 20362 8911 20365
rect 7005 20360 8911 20362
rect 7005 20304 7010 20360
rect 7066 20304 8850 20360
rect 8906 20304 8911 20360
rect 7005 20302 8911 20304
rect 7005 20299 7071 20302
rect 8845 20299 8911 20302
rect 19885 20362 19951 20365
rect 20161 20362 20227 20365
rect 19885 20360 20227 20362
rect 19885 20304 19890 20360
rect 19946 20304 20166 20360
rect 20222 20304 20227 20360
rect 19885 20302 20227 20304
rect 19885 20299 19951 20302
rect 20161 20299 20227 20302
rect 3233 20226 3299 20229
rect 5625 20226 5691 20229
rect 3233 20224 5691 20226
rect 3233 20168 3238 20224
rect 3294 20168 5630 20224
rect 5686 20168 5691 20224
rect 3233 20166 5691 20168
rect 3233 20163 3299 20166
rect 5625 20163 5691 20166
rect 9397 20226 9463 20229
rect 11053 20226 11119 20229
rect 9397 20224 11119 20226
rect 9397 20168 9402 20224
rect 9458 20168 11058 20224
rect 11114 20168 11119 20224
rect 9397 20166 11119 20168
rect 9397 20163 9463 20166
rect 11053 20163 11119 20166
rect 8341 20160 8661 20161
rect 8341 20096 8349 20160
rect 8413 20096 8429 20160
rect 8493 20096 8509 20160
rect 8573 20096 8589 20160
rect 8653 20096 8661 20160
rect 8341 20095 8661 20096
rect 15738 20160 16058 20161
rect 15738 20096 15746 20160
rect 15810 20096 15826 20160
rect 15890 20096 15906 20160
rect 15970 20096 15986 20160
rect 16050 20096 16058 20160
rect 15738 20095 16058 20096
rect 9121 20090 9187 20093
rect 9581 20090 9647 20093
rect 9121 20088 9647 20090
rect 9121 20032 9126 20088
rect 9182 20032 9586 20088
rect 9642 20032 9647 20088
rect 9121 20030 9647 20032
rect 9121 20027 9187 20030
rect 9581 20027 9647 20030
rect 9857 20090 9923 20093
rect 12985 20090 13051 20093
rect 9857 20088 13051 20090
rect 9857 20032 9862 20088
rect 9918 20032 12990 20088
rect 13046 20032 13051 20088
rect 9857 20030 13051 20032
rect 9857 20027 9923 20030
rect 12985 20027 13051 20030
rect 18505 20090 18571 20093
rect 22369 20090 22435 20093
rect 18505 20088 22435 20090
rect 18505 20032 18510 20088
rect 18566 20032 22374 20088
rect 22430 20032 22435 20088
rect 18505 20030 22435 20032
rect 18505 20027 18571 20030
rect 22369 20027 22435 20030
rect 22829 20090 22895 20093
rect 23600 20090 24400 20120
rect 22829 20088 24400 20090
rect 22829 20032 22834 20088
rect 22890 20032 24400 20088
rect 22829 20030 24400 20032
rect 22829 20027 22895 20030
rect 23600 20000 24400 20030
rect 3785 19954 3851 19957
rect 11145 19954 11211 19957
rect 3785 19952 11211 19954
rect 3785 19896 3790 19952
rect 3846 19896 11150 19952
rect 11206 19896 11211 19952
rect 3785 19894 11211 19896
rect 3785 19891 3851 19894
rect 11145 19891 11211 19894
rect 20529 19954 20595 19957
rect 20662 19954 20668 19956
rect 20529 19952 20668 19954
rect 20529 19896 20534 19952
rect 20590 19896 20668 19952
rect 20529 19894 20668 19896
rect 20529 19891 20595 19894
rect 20662 19892 20668 19894
rect 20732 19892 20738 19956
rect 1853 19818 1919 19821
rect 2773 19818 2839 19821
rect 4797 19818 4863 19821
rect 1853 19816 4863 19818
rect 1853 19760 1858 19816
rect 1914 19760 2778 19816
rect 2834 19760 4802 19816
rect 4858 19760 4863 19816
rect 1853 19758 4863 19760
rect 1853 19755 1919 19758
rect 2773 19755 2839 19758
rect 4797 19755 4863 19758
rect 5717 19818 5783 19821
rect 8937 19818 9003 19821
rect 9305 19818 9371 19821
rect 5717 19816 9003 19818
rect 5717 19760 5722 19816
rect 5778 19760 8942 19816
rect 8998 19760 9003 19816
rect 5717 19758 9003 19760
rect 5717 19755 5783 19758
rect 8937 19755 9003 19758
rect 9262 19816 9371 19818
rect 9262 19760 9310 19816
rect 9366 19760 9371 19816
rect 9262 19755 9371 19760
rect 18137 19818 18203 19821
rect 20161 19818 20227 19821
rect 21909 19818 21975 19821
rect 18137 19816 19948 19818
rect 18137 19760 18142 19816
rect 18198 19760 19948 19816
rect 18137 19758 19948 19760
rect 18137 19755 18203 19758
rect 9262 19682 9322 19755
rect 9397 19682 9463 19685
rect 9262 19680 9463 19682
rect 9262 19624 9402 19680
rect 9458 19624 9463 19680
rect 9262 19622 9463 19624
rect 9397 19619 9463 19622
rect 14273 19682 14339 19685
rect 16021 19682 16087 19685
rect 14273 19680 16087 19682
rect 14273 19624 14278 19680
rect 14334 19624 16026 19680
rect 16082 19624 16087 19680
rect 14273 19622 16087 19624
rect 19888 19682 19948 19758
rect 20161 19816 21975 19818
rect 20161 19760 20166 19816
rect 20222 19760 21914 19816
rect 21970 19760 21975 19816
rect 20161 19758 21975 19760
rect 20161 19755 20227 19758
rect 21909 19755 21975 19758
rect 21541 19682 21607 19685
rect 19888 19680 21607 19682
rect 19888 19624 21546 19680
rect 21602 19624 21607 19680
rect 19888 19622 21607 19624
rect 14273 19619 14339 19622
rect 16021 19619 16087 19622
rect 21541 19619 21607 19622
rect 4642 19616 4962 19617
rect 4642 19552 4650 19616
rect 4714 19552 4730 19616
rect 4794 19552 4810 19616
rect 4874 19552 4890 19616
rect 4954 19552 4962 19616
rect 4642 19551 4962 19552
rect 12040 19616 12360 19617
rect 12040 19552 12048 19616
rect 12112 19552 12128 19616
rect 12192 19552 12208 19616
rect 12272 19552 12288 19616
rect 12352 19552 12360 19616
rect 12040 19551 12360 19552
rect 19437 19616 19757 19617
rect 19437 19552 19445 19616
rect 19509 19552 19525 19616
rect 19589 19552 19605 19616
rect 19669 19552 19685 19616
rect 19749 19552 19757 19616
rect 19437 19551 19757 19552
rect 6637 19546 6703 19549
rect 9489 19546 9555 19549
rect 6637 19544 9555 19546
rect 6637 19488 6642 19544
rect 6698 19488 9494 19544
rect 9550 19488 9555 19544
rect 6637 19486 9555 19488
rect 6637 19483 6703 19486
rect 9489 19483 9555 19486
rect 14549 19546 14615 19549
rect 16757 19546 16823 19549
rect 14549 19544 16823 19546
rect 14549 19488 14554 19544
rect 14610 19488 16762 19544
rect 16818 19488 16823 19544
rect 14549 19486 16823 19488
rect 14549 19483 14615 19486
rect 16757 19483 16823 19486
rect 7649 19410 7715 19413
rect 6870 19408 7715 19410
rect 6870 19352 7654 19408
rect 7710 19352 7715 19408
rect 6870 19350 7715 19352
rect 6729 19274 6795 19277
rect 6870 19274 6930 19350
rect 7649 19347 7715 19350
rect 7925 19410 7991 19413
rect 10041 19410 10107 19413
rect 7925 19408 10107 19410
rect 7925 19352 7930 19408
rect 7986 19352 10046 19408
rect 10102 19352 10107 19408
rect 7925 19350 10107 19352
rect 7925 19347 7991 19350
rect 10041 19347 10107 19350
rect 15285 19410 15351 19413
rect 21633 19410 21699 19413
rect 15285 19408 21699 19410
rect 15285 19352 15290 19408
rect 15346 19352 21638 19408
rect 21694 19352 21699 19408
rect 15285 19350 21699 19352
rect 15285 19347 15351 19350
rect 21633 19347 21699 19350
rect 22829 19410 22895 19413
rect 23600 19410 24400 19440
rect 22829 19408 24400 19410
rect 22829 19352 22834 19408
rect 22890 19352 24400 19408
rect 22829 19350 24400 19352
rect 22829 19347 22895 19350
rect 23600 19320 24400 19350
rect 6729 19272 6930 19274
rect 6729 19216 6734 19272
rect 6790 19216 6930 19272
rect 6729 19214 6930 19216
rect 9581 19274 9647 19277
rect 13077 19274 13143 19277
rect 13486 19274 13492 19276
rect 9581 19272 13492 19274
rect 9581 19216 9586 19272
rect 9642 19216 13082 19272
rect 13138 19216 13492 19272
rect 9581 19214 13492 19216
rect 6729 19211 6795 19214
rect 9581 19211 9647 19214
rect 13077 19211 13143 19214
rect 13486 19212 13492 19214
rect 13556 19212 13562 19276
rect 14273 19274 14339 19277
rect 20897 19274 20963 19277
rect 14273 19272 20963 19274
rect 14273 19216 14278 19272
rect 14334 19216 20902 19272
rect 20958 19216 20963 19272
rect 14273 19214 20963 19216
rect 14273 19211 14339 19214
rect 20897 19211 20963 19214
rect 10041 19138 10107 19141
rect 10593 19138 10659 19141
rect 10041 19136 10659 19138
rect 10041 19080 10046 19136
rect 10102 19080 10598 19136
rect 10654 19080 10659 19136
rect 10041 19078 10659 19080
rect 10041 19075 10107 19078
rect 10593 19075 10659 19078
rect 8341 19072 8661 19073
rect 8341 19008 8349 19072
rect 8413 19008 8429 19072
rect 8493 19008 8509 19072
rect 8573 19008 8589 19072
rect 8653 19008 8661 19072
rect 8341 19007 8661 19008
rect 15738 19072 16058 19073
rect 15738 19008 15746 19072
rect 15810 19008 15826 19072
rect 15890 19008 15906 19072
rect 15970 19008 15986 19072
rect 16050 19008 16058 19072
rect 15738 19007 16058 19008
rect 16481 19002 16547 19005
rect 18321 19002 18387 19005
rect 18781 19002 18847 19005
rect 16481 19000 18387 19002
rect 16481 18944 16486 19000
rect 16542 18944 18326 19000
rect 18382 18944 18387 19000
rect 16481 18942 18387 18944
rect 16481 18939 16547 18942
rect 18321 18939 18387 18942
rect 18462 19000 18847 19002
rect 18462 18944 18786 19000
rect 18842 18944 18847 19000
rect 18462 18942 18847 18944
rect 16021 18866 16087 18869
rect 18462 18866 18522 18942
rect 18781 18939 18847 18942
rect 16021 18864 18522 18866
rect 16021 18808 16026 18864
rect 16082 18808 18522 18864
rect 16021 18806 18522 18808
rect 16021 18803 16087 18806
rect 7373 18730 7439 18733
rect 11789 18730 11855 18733
rect 7373 18728 11855 18730
rect 7373 18672 7378 18728
rect 7434 18672 11794 18728
rect 11850 18672 11855 18728
rect 7373 18670 11855 18672
rect 7373 18667 7439 18670
rect 11789 18667 11855 18670
rect 12065 18730 12131 18733
rect 12985 18730 13051 18733
rect 12065 18728 13051 18730
rect 12065 18672 12070 18728
rect 12126 18672 12990 18728
rect 13046 18672 13051 18728
rect 12065 18670 13051 18672
rect 12065 18667 12131 18670
rect 12985 18667 13051 18670
rect 15745 18730 15811 18733
rect 16297 18730 16363 18733
rect 15745 18728 16363 18730
rect 15745 18672 15750 18728
rect 15806 18672 16302 18728
rect 16358 18672 16363 18728
rect 15745 18670 16363 18672
rect 15745 18667 15811 18670
rect 16297 18667 16363 18670
rect 16982 18668 16988 18732
rect 17052 18730 17058 18732
rect 17125 18730 17191 18733
rect 19006 18730 19012 18732
rect 17052 18728 17191 18730
rect 17052 18672 17130 18728
rect 17186 18672 17191 18728
rect 17052 18670 17191 18672
rect 17052 18668 17058 18670
rect 17125 18667 17191 18670
rect 17312 18670 19012 18730
rect 6545 18594 6611 18597
rect 8477 18594 8543 18597
rect 6545 18592 8543 18594
rect 6545 18536 6550 18592
rect 6606 18536 8482 18592
rect 8538 18536 8543 18592
rect 6545 18534 8543 18536
rect 6545 18531 6611 18534
rect 8477 18531 8543 18534
rect 15101 18594 15167 18597
rect 17312 18594 17372 18670
rect 19006 18668 19012 18670
rect 19076 18730 19082 18732
rect 20161 18730 20227 18733
rect 19076 18728 20227 18730
rect 19076 18672 20166 18728
rect 20222 18672 20227 18728
rect 19076 18670 20227 18672
rect 19076 18668 19082 18670
rect 20161 18667 20227 18670
rect 20713 18730 20779 18733
rect 23600 18730 24400 18760
rect 20713 18728 24400 18730
rect 20713 18672 20718 18728
rect 20774 18672 24400 18728
rect 20713 18670 24400 18672
rect 20713 18667 20779 18670
rect 23600 18640 24400 18670
rect 15101 18592 17372 18594
rect 15101 18536 15106 18592
rect 15162 18536 17372 18592
rect 15101 18534 17372 18536
rect 15101 18531 15167 18534
rect 4642 18528 4962 18529
rect 4642 18464 4650 18528
rect 4714 18464 4730 18528
rect 4794 18464 4810 18528
rect 4874 18464 4890 18528
rect 4954 18464 4962 18528
rect 4642 18463 4962 18464
rect 12040 18528 12360 18529
rect 12040 18464 12048 18528
rect 12112 18464 12128 18528
rect 12192 18464 12208 18528
rect 12272 18464 12288 18528
rect 12352 18464 12360 18528
rect 12040 18463 12360 18464
rect 19437 18528 19757 18529
rect 19437 18464 19445 18528
rect 19509 18464 19525 18528
rect 19589 18464 19605 18528
rect 19669 18464 19685 18528
rect 19749 18464 19757 18528
rect 19437 18463 19757 18464
rect 16573 18458 16639 18461
rect 19149 18458 19215 18461
rect 20069 18460 20135 18461
rect 20069 18458 20116 18460
rect 16573 18456 19215 18458
rect 16573 18400 16578 18456
rect 16634 18400 19154 18456
rect 19210 18400 19215 18456
rect 16573 18398 19215 18400
rect 20024 18456 20116 18458
rect 20024 18400 20074 18456
rect 20024 18398 20116 18400
rect 16573 18395 16639 18398
rect 19149 18395 19215 18398
rect 20069 18396 20116 18398
rect 20180 18396 20186 18460
rect 20069 18395 20135 18396
rect 11053 18322 11119 18325
rect 20161 18322 20227 18325
rect 11053 18320 20227 18322
rect 11053 18264 11058 18320
rect 11114 18264 20166 18320
rect 20222 18264 20227 18320
rect 11053 18262 20227 18264
rect 11053 18259 11119 18262
rect 20161 18259 20227 18262
rect 14222 18124 14228 18188
rect 14292 18186 14298 18188
rect 14292 18126 19626 18186
rect 14292 18124 14298 18126
rect 9489 18050 9555 18053
rect 11789 18050 11855 18053
rect 13169 18052 13235 18053
rect 9489 18048 11855 18050
rect 9489 17992 9494 18048
rect 9550 17992 11794 18048
rect 11850 17992 11855 18048
rect 9489 17990 11855 17992
rect 9489 17987 9555 17990
rect 11789 17987 11855 17990
rect 13118 17988 13124 18052
rect 13188 18050 13235 18052
rect 19566 18050 19626 18126
rect 19926 18124 19932 18188
rect 19996 18186 20002 18188
rect 19996 18126 23490 18186
rect 19996 18124 20002 18126
rect 20989 18050 21055 18053
rect 13188 18048 13280 18050
rect 13230 17992 13280 18048
rect 13188 17990 13280 17992
rect 19566 18048 21055 18050
rect 19566 17992 20994 18048
rect 21050 17992 21055 18048
rect 19566 17990 21055 17992
rect 13188 17988 13235 17990
rect 13169 17987 13235 17988
rect 20989 17987 21055 17990
rect 21357 18052 21423 18053
rect 21633 18052 21699 18053
rect 21357 18048 21404 18052
rect 21468 18050 21474 18052
rect 21357 17992 21362 18048
rect 21357 17988 21404 17992
rect 21468 17990 21514 18050
rect 21468 17988 21474 17990
rect 21582 17988 21588 18052
rect 21652 18050 21699 18052
rect 23430 18050 23490 18126
rect 23600 18050 24400 18080
rect 21652 18048 21744 18050
rect 21694 17992 21744 18048
rect 21652 17990 21744 17992
rect 23430 17990 24400 18050
rect 21652 17988 21699 17990
rect 21357 17987 21423 17988
rect 21633 17987 21699 17988
rect 8341 17984 8661 17985
rect 8341 17920 8349 17984
rect 8413 17920 8429 17984
rect 8493 17920 8509 17984
rect 8573 17920 8589 17984
rect 8653 17920 8661 17984
rect 8341 17919 8661 17920
rect 15738 17984 16058 17985
rect 15738 17920 15746 17984
rect 15810 17920 15826 17984
rect 15890 17920 15906 17984
rect 15970 17920 15986 17984
rect 16050 17920 16058 17984
rect 23600 17960 24400 17990
rect 15738 17919 16058 17920
rect 6453 17778 6519 17781
rect 10593 17778 10659 17781
rect 6453 17776 10659 17778
rect 6453 17720 6458 17776
rect 6514 17720 10598 17776
rect 10654 17720 10659 17776
rect 6453 17718 10659 17720
rect 6453 17715 6519 17718
rect 10593 17715 10659 17718
rect 14181 17778 14247 17781
rect 16757 17778 16823 17781
rect 14181 17776 16823 17778
rect 14181 17720 14186 17776
rect 14242 17720 16762 17776
rect 16818 17720 16823 17776
rect 14181 17718 16823 17720
rect 14181 17715 14247 17718
rect 16757 17715 16823 17718
rect 19190 17716 19196 17780
rect 19260 17778 19266 17780
rect 19885 17778 19951 17781
rect 19260 17776 19951 17778
rect 19260 17720 19890 17776
rect 19946 17720 19951 17776
rect 19260 17718 19951 17720
rect 19260 17716 19266 17718
rect 19885 17715 19951 17718
rect 4889 17642 4955 17645
rect 9121 17642 9187 17645
rect 4889 17640 9187 17642
rect 4889 17584 4894 17640
rect 4950 17584 9126 17640
rect 9182 17584 9187 17640
rect 4889 17582 9187 17584
rect 4889 17579 4955 17582
rect 9121 17579 9187 17582
rect 9305 17642 9371 17645
rect 12525 17642 12591 17645
rect 9305 17640 12591 17642
rect 9305 17584 9310 17640
rect 9366 17584 12530 17640
rect 12586 17584 12591 17640
rect 9305 17582 12591 17584
rect 9305 17579 9371 17582
rect 12525 17579 12591 17582
rect 16430 17580 16436 17644
rect 16500 17642 16506 17644
rect 19517 17642 19583 17645
rect 16500 17640 19583 17642
rect 16500 17584 19522 17640
rect 19578 17584 19583 17640
rect 16500 17582 19583 17584
rect 16500 17580 16506 17582
rect 19517 17579 19583 17582
rect 13118 17444 13124 17508
rect 13188 17506 13194 17508
rect 13353 17506 13419 17509
rect 13188 17504 13419 17506
rect 13188 17448 13358 17504
rect 13414 17448 13419 17504
rect 13188 17446 13419 17448
rect 13188 17444 13194 17446
rect 13353 17443 13419 17446
rect 4642 17440 4962 17441
rect 4642 17376 4650 17440
rect 4714 17376 4730 17440
rect 4794 17376 4810 17440
rect 4874 17376 4890 17440
rect 4954 17376 4962 17440
rect 4642 17375 4962 17376
rect 12040 17440 12360 17441
rect 12040 17376 12048 17440
rect 12112 17376 12128 17440
rect 12192 17376 12208 17440
rect 12272 17376 12288 17440
rect 12352 17376 12360 17440
rect 12040 17375 12360 17376
rect 19437 17440 19757 17441
rect 19437 17376 19445 17440
rect 19509 17376 19525 17440
rect 19589 17376 19605 17440
rect 19669 17376 19685 17440
rect 19749 17376 19757 17440
rect 19437 17375 19757 17376
rect 12433 17370 12499 17373
rect 19885 17370 19951 17373
rect 23600 17370 24400 17400
rect 12433 17368 13186 17370
rect 12433 17312 12438 17368
rect 12494 17312 13186 17368
rect 12433 17310 13186 17312
rect 12433 17307 12499 17310
rect 4797 17234 4863 17237
rect 6637 17234 6703 17237
rect 7005 17234 7071 17237
rect 12893 17234 12959 17237
rect 4797 17232 7071 17234
rect 4797 17176 4802 17232
rect 4858 17176 6642 17232
rect 6698 17176 7010 17232
rect 7066 17176 7071 17232
rect 4797 17174 7071 17176
rect 4797 17171 4863 17174
rect 6637 17171 6703 17174
rect 7005 17171 7071 17174
rect 7238 17232 12959 17234
rect 7238 17176 12898 17232
rect 12954 17176 12959 17232
rect 7238 17174 12959 17176
rect 13126 17234 13186 17310
rect 19885 17368 24400 17370
rect 19885 17312 19890 17368
rect 19946 17312 24400 17368
rect 19885 17310 24400 17312
rect 19885 17307 19951 17310
rect 23600 17280 24400 17310
rect 14917 17234 14983 17237
rect 16481 17234 16547 17237
rect 13126 17232 16547 17234
rect 13126 17176 14922 17232
rect 14978 17176 16486 17232
rect 16542 17176 16547 17232
rect 13126 17174 16547 17176
rect 7238 17101 7298 17174
rect 12893 17171 12959 17174
rect 14917 17171 14983 17174
rect 16481 17171 16547 17174
rect 17125 17234 17191 17237
rect 17902 17234 17908 17236
rect 17125 17232 17908 17234
rect 17125 17176 17130 17232
rect 17186 17176 17908 17232
rect 17125 17174 17908 17176
rect 17125 17171 17191 17174
rect 17902 17172 17908 17174
rect 17972 17234 17978 17236
rect 20253 17234 20319 17237
rect 17972 17232 20319 17234
rect 17972 17176 20258 17232
rect 20314 17176 20319 17232
rect 17972 17174 20319 17176
rect 17972 17172 17978 17174
rect 20253 17171 20319 17174
rect 7189 17096 7298 17101
rect 11973 17098 12039 17101
rect 7189 17040 7194 17096
rect 7250 17040 7298 17096
rect 7189 17038 7298 17040
rect 7790 17096 12039 17098
rect 7790 17040 11978 17096
rect 12034 17040 12039 17096
rect 7790 17038 12039 17040
rect 7189 17035 7255 17038
rect 5257 16962 5323 16965
rect 7790 16962 7850 17038
rect 11973 17035 12039 17038
rect 12433 17098 12499 17101
rect 17953 17098 18019 17101
rect 19241 17098 19307 17101
rect 12433 17096 19307 17098
rect 12433 17040 12438 17096
rect 12494 17040 17958 17096
rect 18014 17040 19246 17096
rect 19302 17040 19307 17096
rect 12433 17038 19307 17040
rect 12433 17035 12499 17038
rect 17953 17035 18019 17038
rect 19241 17035 19307 17038
rect 18137 16964 18203 16965
rect 5257 16960 7850 16962
rect 5257 16904 5262 16960
rect 5318 16904 7850 16960
rect 5257 16902 7850 16904
rect 5257 16899 5323 16902
rect 18086 16900 18092 16964
rect 18156 16962 18203 16964
rect 18156 16960 18248 16962
rect 18198 16904 18248 16960
rect 18156 16902 18248 16904
rect 18156 16900 18203 16902
rect 18137 16899 18203 16900
rect 8341 16896 8661 16897
rect 8341 16832 8349 16896
rect 8413 16832 8429 16896
rect 8493 16832 8509 16896
rect 8573 16832 8589 16896
rect 8653 16832 8661 16896
rect 8341 16831 8661 16832
rect 15738 16896 16058 16897
rect 15738 16832 15746 16896
rect 15810 16832 15826 16896
rect 15890 16832 15906 16896
rect 15970 16832 15986 16896
rect 16050 16832 16058 16896
rect 15738 16831 16058 16832
rect 17166 16764 17172 16828
rect 17236 16826 17242 16828
rect 17236 16766 23490 16826
rect 17236 16764 17242 16766
rect 3325 16690 3391 16693
rect 20897 16690 20963 16693
rect 3325 16688 20963 16690
rect 3325 16632 3330 16688
rect 3386 16632 20902 16688
rect 20958 16632 20963 16688
rect 3325 16630 20963 16632
rect 23430 16690 23490 16766
rect 23600 16690 24400 16720
rect 23430 16630 24400 16690
rect 3325 16627 3391 16630
rect 20897 16627 20963 16630
rect 23600 16600 24400 16630
rect 7373 16554 7439 16557
rect 12709 16554 12775 16557
rect 7373 16552 12775 16554
rect 7373 16496 7378 16552
rect 7434 16496 12714 16552
rect 12770 16496 12775 16552
rect 7373 16494 12775 16496
rect 7373 16491 7439 16494
rect 12709 16491 12775 16494
rect 16113 16554 16179 16557
rect 18873 16554 18939 16557
rect 16113 16552 18939 16554
rect 16113 16496 16118 16552
rect 16174 16496 18878 16552
rect 18934 16496 18939 16552
rect 16113 16494 18939 16496
rect 16113 16491 16179 16494
rect 18873 16491 18939 16494
rect 12433 16418 12499 16421
rect 16297 16418 16363 16421
rect 12433 16416 16363 16418
rect 12433 16360 12438 16416
rect 12494 16360 16302 16416
rect 16358 16360 16363 16416
rect 12433 16358 16363 16360
rect 12433 16355 12499 16358
rect 16297 16355 16363 16358
rect 16757 16418 16823 16421
rect 17033 16418 17099 16421
rect 16757 16416 17099 16418
rect 16757 16360 16762 16416
rect 16818 16360 17038 16416
rect 17094 16360 17099 16416
rect 16757 16358 17099 16360
rect 16757 16355 16823 16358
rect 17033 16355 17099 16358
rect 4642 16352 4962 16353
rect 4642 16288 4650 16352
rect 4714 16288 4730 16352
rect 4794 16288 4810 16352
rect 4874 16288 4890 16352
rect 4954 16288 4962 16352
rect 4642 16287 4962 16288
rect 12040 16352 12360 16353
rect 12040 16288 12048 16352
rect 12112 16288 12128 16352
rect 12192 16288 12208 16352
rect 12272 16288 12288 16352
rect 12352 16288 12360 16352
rect 12040 16287 12360 16288
rect 19437 16352 19757 16353
rect 19437 16288 19445 16352
rect 19509 16288 19525 16352
rect 19589 16288 19605 16352
rect 19669 16288 19685 16352
rect 19749 16288 19757 16352
rect 19437 16287 19757 16288
rect 9949 16282 10015 16285
rect 11697 16282 11763 16285
rect 9949 16280 11763 16282
rect 9949 16224 9954 16280
rect 10010 16224 11702 16280
rect 11758 16224 11763 16280
rect 9949 16222 11763 16224
rect 9949 16219 10015 16222
rect 11697 16219 11763 16222
rect 12985 16282 13051 16285
rect 15837 16282 15903 16285
rect 19241 16284 19307 16285
rect 12985 16280 15903 16282
rect 12985 16224 12990 16280
rect 13046 16224 15842 16280
rect 15898 16224 15903 16280
rect 12985 16222 15903 16224
rect 12985 16219 13051 16222
rect 15837 16219 15903 16222
rect 19190 16220 19196 16284
rect 19260 16282 19307 16284
rect 19260 16280 19352 16282
rect 19302 16224 19352 16280
rect 19260 16222 19352 16224
rect 19260 16220 19307 16222
rect 19241 16219 19307 16220
rect 8937 16146 9003 16149
rect 10317 16146 10383 16149
rect 8937 16144 10383 16146
rect 8937 16088 8942 16144
rect 8998 16088 10322 16144
rect 10378 16088 10383 16144
rect 8937 16086 10383 16088
rect 8937 16083 9003 16086
rect 10317 16083 10383 16086
rect 10777 16146 10843 16149
rect 18505 16146 18571 16149
rect 10777 16144 18571 16146
rect 10777 16088 10782 16144
rect 10838 16088 18510 16144
rect 18566 16088 18571 16144
rect 10777 16086 18571 16088
rect 10777 16083 10843 16086
rect 18505 16083 18571 16086
rect 19190 16084 19196 16148
rect 19260 16146 19266 16148
rect 23600 16146 24400 16176
rect 19260 16086 24400 16146
rect 19260 16084 19266 16086
rect 23600 16056 24400 16086
rect 11237 16010 11303 16013
rect 12893 16010 12959 16013
rect 11237 16008 12959 16010
rect 11237 15952 11242 16008
rect 11298 15952 12898 16008
rect 12954 15952 12959 16008
rect 11237 15950 12959 15952
rect 11237 15947 11303 15950
rect 12893 15947 12959 15950
rect 16021 16010 16087 16013
rect 16665 16010 16731 16013
rect 16021 16008 16731 16010
rect 16021 15952 16026 16008
rect 16082 15952 16670 16008
rect 16726 15952 16731 16008
rect 16021 15950 16731 15952
rect 16021 15947 16087 15950
rect 16665 15947 16731 15950
rect 9397 15874 9463 15877
rect 14733 15874 14799 15877
rect 9397 15872 14799 15874
rect 9397 15816 9402 15872
rect 9458 15816 14738 15872
rect 14794 15816 14799 15872
rect 9397 15814 14799 15816
rect 9397 15811 9463 15814
rect 14733 15811 14799 15814
rect 8341 15808 8661 15809
rect 8341 15744 8349 15808
rect 8413 15744 8429 15808
rect 8493 15744 8509 15808
rect 8573 15744 8589 15808
rect 8653 15744 8661 15808
rect 8341 15743 8661 15744
rect 15738 15808 16058 15809
rect 15738 15744 15746 15808
rect 15810 15744 15826 15808
rect 15890 15744 15906 15808
rect 15970 15744 15986 15808
rect 16050 15744 16058 15808
rect 15738 15743 16058 15744
rect 12801 15738 12867 15741
rect 15101 15738 15167 15741
rect 12801 15736 15167 15738
rect 12801 15680 12806 15736
rect 12862 15680 15106 15736
rect 15162 15680 15167 15736
rect 12801 15678 15167 15680
rect 12801 15675 12867 15678
rect 15101 15675 15167 15678
rect 17861 15738 17927 15741
rect 19885 15738 19951 15741
rect 17861 15736 19951 15738
rect 17861 15680 17866 15736
rect 17922 15680 19890 15736
rect 19946 15680 19951 15736
rect 17861 15678 19951 15680
rect 17861 15675 17927 15678
rect 19885 15675 19951 15678
rect 7097 15602 7163 15605
rect 21449 15602 21515 15605
rect 7097 15600 21515 15602
rect 7097 15544 7102 15600
rect 7158 15544 21454 15600
rect 21510 15544 21515 15600
rect 7097 15542 21515 15544
rect 7097 15539 7163 15542
rect 21449 15539 21515 15542
rect 1485 15466 1551 15469
rect 15745 15466 15811 15469
rect 1485 15464 15811 15466
rect 1485 15408 1490 15464
rect 1546 15408 15750 15464
rect 15806 15408 15811 15464
rect 1485 15406 15811 15408
rect 1485 15403 1551 15406
rect 15745 15403 15811 15406
rect 19333 15466 19399 15469
rect 23600 15466 24400 15496
rect 19333 15464 24400 15466
rect 19333 15408 19338 15464
rect 19394 15408 24400 15464
rect 19333 15406 24400 15408
rect 19333 15403 19399 15406
rect 23600 15376 24400 15406
rect 12801 15330 12867 15333
rect 14273 15330 14339 15333
rect 12801 15328 14339 15330
rect 12801 15272 12806 15328
rect 12862 15272 14278 15328
rect 14334 15272 14339 15328
rect 12801 15270 14339 15272
rect 12801 15267 12867 15270
rect 14273 15267 14339 15270
rect 15745 15330 15811 15333
rect 16573 15330 16639 15333
rect 15745 15328 16639 15330
rect 15745 15272 15750 15328
rect 15806 15272 16578 15328
rect 16634 15272 16639 15328
rect 15745 15270 16639 15272
rect 15745 15267 15811 15270
rect 16573 15267 16639 15270
rect 16798 15268 16804 15332
rect 16868 15330 16874 15332
rect 17677 15330 17743 15333
rect 16868 15328 17743 15330
rect 16868 15272 17682 15328
rect 17738 15272 17743 15328
rect 16868 15270 17743 15272
rect 16868 15268 16874 15270
rect 17677 15267 17743 15270
rect 4642 15264 4962 15265
rect 0 15194 800 15224
rect 4642 15200 4650 15264
rect 4714 15200 4730 15264
rect 4794 15200 4810 15264
rect 4874 15200 4890 15264
rect 4954 15200 4962 15264
rect 4642 15199 4962 15200
rect 12040 15264 12360 15265
rect 12040 15200 12048 15264
rect 12112 15200 12128 15264
rect 12192 15200 12208 15264
rect 12272 15200 12288 15264
rect 12352 15200 12360 15264
rect 12040 15199 12360 15200
rect 19437 15264 19757 15265
rect 19437 15200 19445 15264
rect 19509 15200 19525 15264
rect 19589 15200 19605 15264
rect 19669 15200 19685 15264
rect 19749 15200 19757 15264
rect 19437 15199 19757 15200
rect 1853 15194 1919 15197
rect 0 15192 1919 15194
rect 0 15136 1858 15192
rect 1914 15136 1919 15192
rect 0 15134 1919 15136
rect 0 15104 800 15134
rect 1853 15131 1919 15134
rect 12525 15194 12591 15197
rect 14825 15194 14891 15197
rect 12525 15192 14891 15194
rect 12525 15136 12530 15192
rect 12586 15136 14830 15192
rect 14886 15136 14891 15192
rect 12525 15134 14891 15136
rect 12525 15131 12591 15134
rect 14825 15131 14891 15134
rect 15193 15194 15259 15197
rect 15929 15194 15995 15197
rect 15193 15192 15995 15194
rect 15193 15136 15198 15192
rect 15254 15136 15934 15192
rect 15990 15136 15995 15192
rect 15193 15134 15995 15136
rect 15193 15131 15259 15134
rect 15929 15131 15995 15134
rect 16573 15194 16639 15197
rect 18781 15194 18847 15197
rect 16573 15192 18847 15194
rect 16573 15136 16578 15192
rect 16634 15136 18786 15192
rect 18842 15136 18847 15192
rect 16573 15134 18847 15136
rect 16573 15131 16639 15134
rect 18781 15131 18847 15134
rect 3785 15058 3851 15061
rect 11789 15058 11855 15061
rect 3785 15056 11855 15058
rect 3785 15000 3790 15056
rect 3846 15000 11794 15056
rect 11850 15000 11855 15056
rect 3785 14998 11855 15000
rect 3785 14995 3851 14998
rect 11789 14995 11855 14998
rect 12341 15058 12407 15061
rect 20621 15058 20687 15061
rect 12341 15056 20687 15058
rect 12341 15000 12346 15056
rect 12402 15000 20626 15056
rect 20682 15000 20687 15056
rect 12341 14998 20687 15000
rect 12341 14995 12407 14998
rect 20621 14995 20687 14998
rect 10593 14922 10659 14925
rect 10961 14922 11027 14925
rect 10593 14920 11027 14922
rect 10593 14864 10598 14920
rect 10654 14864 10966 14920
rect 11022 14864 11027 14920
rect 10593 14862 11027 14864
rect 10593 14859 10659 14862
rect 10961 14859 11027 14862
rect 11697 14922 11763 14925
rect 12801 14922 12867 14925
rect 16021 14922 16087 14925
rect 11697 14920 12867 14922
rect 11697 14864 11702 14920
rect 11758 14864 12806 14920
rect 12862 14864 12867 14920
rect 11697 14862 12867 14864
rect 11697 14859 11763 14862
rect 12801 14859 12867 14862
rect 15518 14920 16087 14922
rect 15518 14864 16026 14920
rect 16082 14864 16087 14920
rect 15518 14862 16087 14864
rect 15518 14789 15578 14862
rect 16021 14859 16087 14862
rect 16614 14860 16620 14924
rect 16684 14922 16690 14924
rect 20069 14922 20135 14925
rect 16684 14920 20135 14922
rect 16684 14864 20074 14920
rect 20130 14864 20135 14920
rect 16684 14862 20135 14864
rect 16684 14860 16690 14862
rect 20069 14859 20135 14862
rect 11973 14786 12039 14789
rect 15285 14786 15351 14789
rect 11973 14784 15351 14786
rect 11973 14728 11978 14784
rect 12034 14728 15290 14784
rect 15346 14728 15351 14784
rect 11973 14726 15351 14728
rect 11973 14723 12039 14726
rect 15285 14723 15351 14726
rect 15469 14784 15578 14789
rect 15469 14728 15474 14784
rect 15530 14728 15578 14784
rect 15469 14726 15578 14728
rect 19333 14786 19399 14789
rect 23600 14786 24400 14816
rect 19333 14784 24400 14786
rect 19333 14728 19338 14784
rect 19394 14728 24400 14784
rect 19333 14726 24400 14728
rect 15469 14723 15535 14726
rect 19333 14723 19399 14726
rect 8341 14720 8661 14721
rect 8341 14656 8349 14720
rect 8413 14656 8429 14720
rect 8493 14656 8509 14720
rect 8573 14656 8589 14720
rect 8653 14656 8661 14720
rect 8341 14655 8661 14656
rect 15738 14720 16058 14721
rect 15738 14656 15746 14720
rect 15810 14656 15826 14720
rect 15890 14656 15906 14720
rect 15970 14656 15986 14720
rect 16050 14656 16058 14720
rect 23600 14696 24400 14726
rect 15738 14655 16058 14656
rect 9078 14590 14474 14650
rect 7465 14514 7531 14517
rect 9078 14514 9138 14590
rect 7465 14512 9138 14514
rect 7465 14456 7470 14512
rect 7526 14456 9138 14512
rect 7465 14454 9138 14456
rect 11053 14514 11119 14517
rect 14181 14514 14247 14517
rect 11053 14512 14247 14514
rect 11053 14456 11058 14512
rect 11114 14456 14186 14512
rect 14242 14456 14247 14512
rect 11053 14454 14247 14456
rect 14414 14514 14474 14590
rect 16246 14588 16252 14652
rect 16316 14650 16322 14652
rect 20437 14650 20503 14653
rect 16316 14648 20503 14650
rect 16316 14592 20442 14648
rect 20498 14592 20503 14648
rect 16316 14590 20503 14592
rect 16316 14588 16322 14590
rect 20437 14587 20503 14590
rect 17309 14514 17375 14517
rect 14414 14512 17375 14514
rect 14414 14456 17314 14512
rect 17370 14456 17375 14512
rect 14414 14454 17375 14456
rect 7465 14451 7531 14454
rect 11053 14451 11119 14454
rect 14181 14451 14247 14454
rect 17309 14451 17375 14454
rect 18505 14514 18571 14517
rect 19425 14514 19491 14517
rect 18505 14512 19491 14514
rect 18505 14456 18510 14512
rect 18566 14456 19430 14512
rect 19486 14456 19491 14512
rect 18505 14454 19491 14456
rect 18505 14451 18571 14454
rect 19425 14451 19491 14454
rect 1669 14378 1735 14381
rect 22093 14378 22159 14381
rect 1669 14376 22159 14378
rect 1669 14320 1674 14376
rect 1730 14320 22098 14376
rect 22154 14320 22159 14376
rect 1669 14318 22159 14320
rect 1669 14315 1735 14318
rect 22093 14315 22159 14318
rect 6821 14242 6887 14245
rect 11145 14242 11211 14245
rect 6821 14240 11211 14242
rect 6821 14184 6826 14240
rect 6882 14184 11150 14240
rect 11206 14184 11211 14240
rect 6821 14182 11211 14184
rect 6821 14179 6887 14182
rect 11145 14179 11211 14182
rect 12893 14242 12959 14245
rect 16021 14242 16087 14245
rect 12893 14240 16087 14242
rect 12893 14184 12898 14240
rect 12954 14184 16026 14240
rect 16082 14184 16087 14240
rect 12893 14182 16087 14184
rect 12893 14179 12959 14182
rect 16021 14179 16087 14182
rect 4642 14176 4962 14177
rect 4642 14112 4650 14176
rect 4714 14112 4730 14176
rect 4794 14112 4810 14176
rect 4874 14112 4890 14176
rect 4954 14112 4962 14176
rect 4642 14111 4962 14112
rect 12040 14176 12360 14177
rect 12040 14112 12048 14176
rect 12112 14112 12128 14176
rect 12192 14112 12208 14176
rect 12272 14112 12288 14176
rect 12352 14112 12360 14176
rect 12040 14111 12360 14112
rect 19437 14176 19757 14177
rect 19437 14112 19445 14176
rect 19509 14112 19525 14176
rect 19589 14112 19605 14176
rect 19669 14112 19685 14176
rect 19749 14112 19757 14176
rect 19437 14111 19757 14112
rect 13486 14044 13492 14108
rect 13556 14106 13562 14108
rect 16021 14106 16087 14109
rect 13556 14104 16087 14106
rect 13556 14048 16026 14104
rect 16082 14048 16087 14104
rect 13556 14046 16087 14048
rect 13556 14044 13562 14046
rect 16021 14043 16087 14046
rect 16297 14106 16363 14109
rect 18045 14106 18111 14109
rect 16297 14104 18111 14106
rect 16297 14048 16302 14104
rect 16358 14048 18050 14104
rect 18106 14048 18111 14104
rect 16297 14046 18111 14048
rect 16297 14043 16363 14046
rect 18045 14043 18111 14046
rect 20621 14106 20687 14109
rect 23600 14106 24400 14136
rect 20621 14104 24400 14106
rect 20621 14048 20626 14104
rect 20682 14048 24400 14104
rect 20621 14046 24400 14048
rect 20621 14043 20687 14046
rect 23600 14016 24400 14046
rect 7281 13970 7347 13973
rect 16757 13970 16823 13973
rect 7281 13968 16823 13970
rect 7281 13912 7286 13968
rect 7342 13912 16762 13968
rect 16818 13912 16823 13968
rect 7281 13910 16823 13912
rect 7281 13907 7347 13910
rect 16757 13907 16823 13910
rect 16982 13908 16988 13972
rect 17052 13970 17058 13972
rect 21265 13970 21331 13973
rect 17052 13968 21331 13970
rect 17052 13912 21270 13968
rect 21326 13912 21331 13968
rect 17052 13910 21331 13912
rect 17052 13908 17058 13910
rect 21265 13907 21331 13910
rect 2865 13834 2931 13837
rect 9949 13834 10015 13837
rect 20897 13834 20963 13837
rect 2865 13832 9322 13834
rect 2865 13776 2870 13832
rect 2926 13776 9322 13832
rect 2865 13774 9322 13776
rect 2865 13771 2931 13774
rect 9262 13698 9322 13774
rect 9949 13832 20963 13834
rect 9949 13776 9954 13832
rect 10010 13776 20902 13832
rect 20958 13776 20963 13832
rect 9949 13774 20963 13776
rect 9949 13771 10015 13774
rect 20897 13771 20963 13774
rect 14181 13698 14247 13701
rect 9262 13696 14247 13698
rect 9262 13640 14186 13696
rect 14242 13640 14247 13696
rect 9262 13638 14247 13640
rect 14181 13635 14247 13638
rect 16389 13698 16455 13701
rect 16798 13698 16804 13700
rect 16389 13696 16804 13698
rect 16389 13640 16394 13696
rect 16450 13640 16804 13696
rect 16389 13638 16804 13640
rect 16389 13635 16455 13638
rect 16798 13636 16804 13638
rect 16868 13636 16874 13700
rect 17309 13698 17375 13701
rect 19926 13698 19932 13700
rect 17309 13696 19932 13698
rect 17309 13640 17314 13696
rect 17370 13640 19932 13696
rect 17309 13638 19932 13640
rect 17309 13635 17375 13638
rect 19926 13636 19932 13638
rect 19996 13636 20002 13700
rect 8341 13632 8661 13633
rect 8341 13568 8349 13632
rect 8413 13568 8429 13632
rect 8493 13568 8509 13632
rect 8573 13568 8589 13632
rect 8653 13568 8661 13632
rect 8341 13567 8661 13568
rect 15738 13632 16058 13633
rect 15738 13568 15746 13632
rect 15810 13568 15826 13632
rect 15890 13568 15906 13632
rect 15970 13568 15986 13632
rect 16050 13568 16058 13632
rect 15738 13567 16058 13568
rect 11329 13562 11395 13565
rect 12065 13562 12131 13565
rect 13077 13564 13143 13565
rect 13077 13562 13124 13564
rect 11329 13560 12131 13562
rect 11329 13504 11334 13560
rect 11390 13504 12070 13560
rect 12126 13504 12131 13560
rect 11329 13502 12131 13504
rect 13032 13560 13124 13562
rect 13032 13504 13082 13560
rect 13032 13502 13124 13504
rect 11329 13499 11395 13502
rect 12065 13499 12131 13502
rect 13077 13500 13124 13502
rect 13188 13500 13194 13564
rect 16205 13562 16271 13565
rect 18229 13562 18295 13565
rect 16205 13560 18295 13562
rect 16205 13504 16210 13560
rect 16266 13504 18234 13560
rect 18290 13504 18295 13560
rect 16205 13502 18295 13504
rect 13077 13499 13143 13500
rect 16205 13499 16271 13502
rect 18229 13499 18295 13502
rect 19609 13562 19675 13565
rect 21265 13562 21331 13565
rect 19609 13560 21331 13562
rect 19609 13504 19614 13560
rect 19670 13504 21270 13560
rect 21326 13504 21331 13560
rect 19609 13502 21331 13504
rect 19609 13499 19675 13502
rect 21265 13499 21331 13502
rect 5993 13426 6059 13429
rect 20897 13426 20963 13429
rect 23600 13426 24400 13456
rect 5993 13424 20963 13426
rect 5993 13368 5998 13424
rect 6054 13368 20902 13424
rect 20958 13368 20963 13424
rect 5993 13366 20963 13368
rect 5993 13363 6059 13366
rect 20897 13363 20963 13366
rect 23430 13366 24400 13426
rect 3969 13290 4035 13293
rect 17309 13290 17375 13293
rect 3969 13288 17375 13290
rect 3969 13232 3974 13288
rect 4030 13232 17314 13288
rect 17370 13232 17375 13288
rect 3969 13230 17375 13232
rect 3969 13227 4035 13230
rect 17309 13227 17375 13230
rect 17953 13290 18019 13293
rect 23430 13290 23490 13366
rect 23600 13336 24400 13366
rect 17953 13288 23490 13290
rect 17953 13232 17958 13288
rect 18014 13232 23490 13288
rect 17953 13230 23490 13232
rect 17953 13227 18019 13230
rect 9213 13154 9279 13157
rect 11881 13154 11947 13157
rect 9213 13152 11947 13154
rect 9213 13096 9218 13152
rect 9274 13096 11886 13152
rect 11942 13096 11947 13152
rect 9213 13094 11947 13096
rect 9213 13091 9279 13094
rect 11881 13091 11947 13094
rect 14917 13154 14983 13157
rect 17125 13154 17191 13157
rect 14917 13152 17191 13154
rect 14917 13096 14922 13152
rect 14978 13096 17130 13152
rect 17186 13096 17191 13152
rect 14917 13094 17191 13096
rect 14917 13091 14983 13094
rect 17125 13091 17191 13094
rect 17769 13154 17835 13157
rect 17902 13154 17908 13156
rect 17769 13152 17908 13154
rect 17769 13096 17774 13152
rect 17830 13096 17908 13152
rect 17769 13094 17908 13096
rect 17769 13091 17835 13094
rect 17902 13092 17908 13094
rect 17972 13092 17978 13156
rect 19885 13154 19951 13157
rect 22369 13154 22435 13157
rect 19885 13152 22435 13154
rect 19885 13096 19890 13152
rect 19946 13096 22374 13152
rect 22430 13096 22435 13152
rect 19885 13094 22435 13096
rect 19885 13091 19951 13094
rect 22369 13091 22435 13094
rect 4642 13088 4962 13089
rect 4642 13024 4650 13088
rect 4714 13024 4730 13088
rect 4794 13024 4810 13088
rect 4874 13024 4890 13088
rect 4954 13024 4962 13088
rect 4642 13023 4962 13024
rect 12040 13088 12360 13089
rect 12040 13024 12048 13088
rect 12112 13024 12128 13088
rect 12192 13024 12208 13088
rect 12272 13024 12288 13088
rect 12352 13024 12360 13088
rect 12040 13023 12360 13024
rect 19437 13088 19757 13089
rect 19437 13024 19445 13088
rect 19509 13024 19525 13088
rect 19589 13024 19605 13088
rect 19669 13024 19685 13088
rect 19749 13024 19757 13088
rect 19437 13023 19757 13024
rect 15653 13018 15719 13021
rect 18965 13018 19031 13021
rect 15653 13016 19031 13018
rect 15653 12960 15658 13016
rect 15714 12960 18970 13016
rect 19026 12960 19031 13016
rect 15653 12958 19031 12960
rect 15653 12955 15719 12958
rect 18965 12955 19031 12958
rect 6453 12882 6519 12885
rect 17166 12882 17172 12884
rect 6453 12880 17172 12882
rect 6453 12824 6458 12880
rect 6514 12824 17172 12880
rect 6453 12822 17172 12824
rect 6453 12819 6519 12822
rect 17166 12820 17172 12822
rect 17236 12820 17242 12884
rect 17493 12882 17559 12885
rect 18505 12882 18571 12885
rect 17493 12880 18571 12882
rect 17493 12824 17498 12880
rect 17554 12824 18510 12880
rect 18566 12824 18571 12880
rect 17493 12822 18571 12824
rect 17493 12819 17559 12822
rect 18505 12819 18571 12822
rect 18638 12820 18644 12884
rect 18708 12882 18714 12884
rect 19057 12882 19123 12885
rect 18708 12880 19123 12882
rect 18708 12824 19062 12880
rect 19118 12824 19123 12880
rect 18708 12822 19123 12824
rect 18708 12820 18714 12822
rect 19057 12819 19123 12822
rect 19926 12820 19932 12884
rect 19996 12882 20002 12884
rect 20713 12882 20779 12885
rect 19996 12880 20779 12882
rect 19996 12824 20718 12880
rect 20774 12824 20779 12880
rect 19996 12822 20779 12824
rect 19996 12820 20002 12822
rect 20713 12819 20779 12822
rect 6821 12746 6887 12749
rect 23600 12746 24400 12776
rect 6821 12744 24400 12746
rect 6821 12688 6826 12744
rect 6882 12688 24400 12744
rect 6821 12686 24400 12688
rect 6821 12683 6887 12686
rect 23600 12656 24400 12686
rect 11053 12610 11119 12613
rect 14825 12610 14891 12613
rect 11053 12608 14891 12610
rect 11053 12552 11058 12608
rect 11114 12552 14830 12608
rect 14886 12552 14891 12608
rect 11053 12550 14891 12552
rect 11053 12547 11119 12550
rect 14825 12547 14891 12550
rect 16205 12610 16271 12613
rect 20253 12612 20319 12613
rect 16430 12610 16436 12612
rect 16205 12608 16436 12610
rect 16205 12552 16210 12608
rect 16266 12552 16436 12608
rect 16205 12550 16436 12552
rect 16205 12547 16271 12550
rect 16430 12548 16436 12550
rect 16500 12548 16506 12612
rect 20253 12608 20300 12612
rect 20364 12610 20370 12612
rect 20253 12552 20258 12608
rect 20253 12548 20300 12552
rect 20364 12550 20410 12610
rect 20364 12548 20370 12550
rect 20253 12547 20319 12548
rect 8341 12544 8661 12545
rect 8341 12480 8349 12544
rect 8413 12480 8429 12544
rect 8493 12480 8509 12544
rect 8573 12480 8589 12544
rect 8653 12480 8661 12544
rect 8341 12479 8661 12480
rect 15738 12544 16058 12545
rect 15738 12480 15746 12544
rect 15810 12480 15826 12544
rect 15890 12480 15906 12544
rect 15970 12480 15986 12544
rect 16050 12480 16058 12544
rect 15738 12479 16058 12480
rect 3877 12474 3943 12477
rect 6361 12474 6427 12477
rect 3877 12472 6427 12474
rect 3877 12416 3882 12472
rect 3938 12416 6366 12472
rect 6422 12416 6427 12472
rect 3877 12414 6427 12416
rect 3877 12411 3943 12414
rect 6361 12411 6427 12414
rect 16849 12474 16915 12477
rect 16982 12474 16988 12476
rect 16849 12472 16988 12474
rect 16849 12416 16854 12472
rect 16910 12416 16988 12472
rect 16849 12414 16988 12416
rect 16849 12411 16915 12414
rect 16982 12412 16988 12414
rect 17052 12412 17058 12476
rect 17585 12474 17651 12477
rect 17718 12474 17724 12476
rect 17585 12472 17724 12474
rect 17585 12416 17590 12472
rect 17646 12416 17724 12472
rect 17585 12414 17724 12416
rect 17585 12411 17651 12414
rect 17718 12412 17724 12414
rect 17788 12412 17794 12476
rect 19333 12474 19399 12477
rect 20069 12476 20135 12477
rect 20621 12476 20687 12477
rect 20069 12474 20116 12476
rect 19333 12472 19580 12474
rect 19333 12416 19338 12472
rect 19394 12416 19580 12472
rect 19333 12414 19580 12416
rect 20024 12472 20116 12474
rect 20024 12416 20074 12472
rect 20024 12414 20116 12416
rect 19333 12411 19399 12414
rect 1577 12338 1643 12341
rect 8937 12338 9003 12341
rect 1577 12336 9003 12338
rect 1577 12280 1582 12336
rect 1638 12280 8942 12336
rect 8998 12280 9003 12336
rect 1577 12278 9003 12280
rect 1577 12275 1643 12278
rect 8937 12275 9003 12278
rect 14273 12338 14339 12341
rect 18638 12338 18644 12340
rect 14273 12336 18644 12338
rect 14273 12280 14278 12336
rect 14334 12280 18644 12336
rect 14273 12278 18644 12280
rect 14273 12275 14339 12278
rect 18638 12276 18644 12278
rect 18708 12276 18714 12340
rect 19190 12276 19196 12340
rect 19260 12338 19266 12340
rect 19333 12338 19399 12341
rect 19260 12336 19399 12338
rect 19260 12280 19338 12336
rect 19394 12280 19399 12336
rect 19260 12278 19399 12280
rect 19520 12338 19580 12414
rect 20069 12412 20116 12414
rect 20180 12412 20186 12476
rect 20621 12474 20668 12476
rect 20576 12472 20668 12474
rect 20576 12416 20626 12472
rect 20576 12414 20668 12416
rect 20621 12412 20668 12414
rect 20732 12412 20738 12476
rect 20069 12411 20135 12412
rect 20621 12411 20687 12412
rect 22277 12338 22343 12341
rect 19520 12336 22343 12338
rect 19520 12280 22282 12336
rect 22338 12280 22343 12336
rect 19520 12278 22343 12280
rect 19260 12276 19266 12278
rect 19333 12275 19399 12278
rect 22277 12275 22343 12278
rect 6913 12202 6979 12205
rect 11513 12202 11579 12205
rect 6913 12200 11579 12202
rect 6913 12144 6918 12200
rect 6974 12144 11518 12200
rect 11574 12144 11579 12200
rect 6913 12142 11579 12144
rect 6913 12139 6979 12142
rect 11513 12139 11579 12142
rect 17217 12202 17283 12205
rect 17953 12202 18019 12205
rect 17217 12200 18019 12202
rect 17217 12144 17222 12200
rect 17278 12144 17958 12200
rect 18014 12144 18019 12200
rect 17217 12142 18019 12144
rect 17217 12139 17283 12142
rect 17953 12139 18019 12142
rect 19609 12202 19675 12205
rect 20161 12202 20227 12205
rect 23600 12202 24400 12232
rect 19609 12200 19948 12202
rect 19609 12144 19614 12200
rect 19670 12144 19948 12200
rect 19609 12142 19948 12144
rect 19609 12139 19675 12142
rect 14641 12066 14707 12069
rect 16297 12066 16363 12069
rect 14641 12064 16363 12066
rect 14641 12008 14646 12064
rect 14702 12008 16302 12064
rect 16358 12008 16363 12064
rect 14641 12006 16363 12008
rect 14641 12003 14707 12006
rect 16297 12003 16363 12006
rect 16665 12066 16731 12069
rect 17861 12066 17927 12069
rect 18873 12066 18939 12069
rect 16665 12064 18939 12066
rect 16665 12008 16670 12064
rect 16726 12008 17866 12064
rect 17922 12008 18878 12064
rect 18934 12008 18939 12064
rect 16665 12006 18939 12008
rect 19888 12066 19948 12142
rect 20161 12200 24400 12202
rect 20161 12144 20166 12200
rect 20222 12144 24400 12200
rect 20161 12142 24400 12144
rect 20161 12139 20227 12142
rect 23600 12112 24400 12142
rect 21357 12066 21423 12069
rect 19888 12064 21423 12066
rect 19888 12008 21362 12064
rect 21418 12008 21423 12064
rect 19888 12006 21423 12008
rect 16665 12003 16731 12006
rect 17861 12003 17927 12006
rect 18873 12003 18939 12006
rect 21357 12003 21423 12006
rect 4642 12000 4962 12001
rect 4642 11936 4650 12000
rect 4714 11936 4730 12000
rect 4794 11936 4810 12000
rect 4874 11936 4890 12000
rect 4954 11936 4962 12000
rect 4642 11935 4962 11936
rect 12040 12000 12360 12001
rect 12040 11936 12048 12000
rect 12112 11936 12128 12000
rect 12192 11936 12208 12000
rect 12272 11936 12288 12000
rect 12352 11936 12360 12000
rect 12040 11935 12360 11936
rect 19437 12000 19757 12001
rect 19437 11936 19445 12000
rect 19509 11936 19525 12000
rect 19589 11936 19605 12000
rect 19669 11936 19685 12000
rect 19749 11936 19757 12000
rect 19437 11935 19757 11936
rect 14365 11930 14431 11933
rect 14365 11928 17602 11930
rect 14365 11872 14370 11928
rect 14426 11872 17602 11928
rect 14365 11870 17602 11872
rect 14365 11867 14431 11870
rect 17309 11794 17375 11797
rect 6824 11792 17375 11794
rect 6824 11736 17314 11792
rect 17370 11736 17375 11792
rect 6824 11734 17375 11736
rect 17542 11794 17602 11870
rect 20110 11868 20116 11932
rect 20180 11930 20186 11932
rect 20345 11930 20411 11933
rect 20180 11928 20411 11930
rect 20180 11872 20350 11928
rect 20406 11872 20411 11928
rect 20180 11870 20411 11872
rect 20180 11868 20186 11870
rect 20345 11867 20411 11870
rect 22277 11794 22343 11797
rect 17542 11792 22343 11794
rect 17542 11736 22282 11792
rect 22338 11736 22343 11792
rect 17542 11734 22343 11736
rect 6545 11522 6611 11525
rect 6824 11522 6884 11734
rect 17309 11731 17375 11734
rect 22277 11731 22343 11734
rect 9581 11658 9647 11661
rect 18229 11658 18295 11661
rect 19241 11658 19307 11661
rect 9581 11656 18295 11658
rect 9581 11600 9586 11656
rect 9642 11600 18234 11656
rect 18290 11600 18295 11656
rect 9581 11598 18295 11600
rect 9581 11595 9647 11598
rect 18229 11595 18295 11598
rect 18462 11656 19307 11658
rect 18462 11600 19246 11656
rect 19302 11600 19307 11656
rect 18462 11598 19307 11600
rect 6545 11520 6884 11522
rect 6545 11464 6550 11520
rect 6606 11464 6884 11520
rect 6545 11462 6884 11464
rect 16297 11522 16363 11525
rect 18462 11522 18522 11598
rect 19241 11595 19307 11598
rect 16297 11520 18522 11522
rect 16297 11464 16302 11520
rect 16358 11464 18522 11520
rect 16297 11462 18522 11464
rect 19333 11522 19399 11525
rect 23600 11522 24400 11552
rect 19333 11520 24400 11522
rect 19333 11464 19338 11520
rect 19394 11464 24400 11520
rect 19333 11462 24400 11464
rect 6545 11459 6611 11462
rect 16297 11459 16363 11462
rect 19333 11459 19399 11462
rect 8341 11456 8661 11457
rect 8341 11392 8349 11456
rect 8413 11392 8429 11456
rect 8493 11392 8509 11456
rect 8573 11392 8589 11456
rect 8653 11392 8661 11456
rect 8341 11391 8661 11392
rect 15738 11456 16058 11457
rect 15738 11392 15746 11456
rect 15810 11392 15826 11456
rect 15890 11392 15906 11456
rect 15970 11392 15986 11456
rect 16050 11392 16058 11456
rect 23600 11432 24400 11462
rect 15738 11391 16058 11392
rect 17309 11386 17375 11389
rect 17677 11386 17743 11389
rect 17309 11384 17743 11386
rect 17309 11328 17314 11384
rect 17370 11328 17682 11384
rect 17738 11328 17743 11384
rect 17309 11326 17743 11328
rect 17309 11323 17375 11326
rect 17677 11323 17743 11326
rect 18873 11384 18939 11389
rect 18873 11328 18878 11384
rect 18934 11328 18939 11384
rect 18873 11323 18939 11328
rect 15653 11250 15719 11253
rect 16757 11250 16823 11253
rect 15653 11248 16823 11250
rect 15653 11192 15658 11248
rect 15714 11192 16762 11248
rect 16818 11192 16823 11248
rect 15653 11190 16823 11192
rect 15653 11187 15719 11190
rect 16757 11187 16823 11190
rect 14825 11114 14891 11117
rect 17953 11114 18019 11117
rect 14825 11112 18019 11114
rect 14825 11056 14830 11112
rect 14886 11056 17958 11112
rect 18014 11056 18019 11112
rect 14825 11054 18019 11056
rect 14825 11051 14891 11054
rect 17953 11051 18019 11054
rect 9857 10980 9923 10981
rect 9806 10916 9812 10980
rect 9876 10978 9923 10980
rect 13905 10978 13971 10981
rect 18876 10978 18936 11323
rect 9876 10976 9968 10978
rect 9918 10920 9968 10976
rect 9876 10918 9968 10920
rect 13905 10976 18936 10978
rect 13905 10920 13910 10976
rect 13966 10920 18936 10976
rect 13905 10918 18936 10920
rect 9876 10916 9923 10918
rect 9857 10915 9923 10916
rect 13905 10915 13971 10918
rect 4642 10912 4962 10913
rect 4642 10848 4650 10912
rect 4714 10848 4730 10912
rect 4794 10848 4810 10912
rect 4874 10848 4890 10912
rect 4954 10848 4962 10912
rect 4642 10847 4962 10848
rect 12040 10912 12360 10913
rect 12040 10848 12048 10912
rect 12112 10848 12128 10912
rect 12192 10848 12208 10912
rect 12272 10848 12288 10912
rect 12352 10848 12360 10912
rect 12040 10847 12360 10848
rect 19437 10912 19757 10913
rect 19437 10848 19445 10912
rect 19509 10848 19525 10912
rect 19589 10848 19605 10912
rect 19669 10848 19685 10912
rect 19749 10848 19757 10912
rect 19437 10847 19757 10848
rect 12985 10842 13051 10845
rect 19241 10842 19307 10845
rect 12985 10840 19307 10842
rect 12985 10784 12990 10840
rect 13046 10784 19246 10840
rect 19302 10784 19307 10840
rect 12985 10782 19307 10784
rect 12985 10779 13051 10782
rect 19241 10779 19307 10782
rect 20529 10842 20595 10845
rect 23600 10842 24400 10872
rect 20529 10840 24400 10842
rect 20529 10784 20534 10840
rect 20590 10784 24400 10840
rect 20529 10782 24400 10784
rect 20529 10779 20595 10782
rect 23600 10752 24400 10782
rect 9673 10708 9739 10709
rect 9622 10644 9628 10708
rect 9692 10706 9739 10708
rect 9857 10706 9923 10709
rect 10041 10706 10107 10709
rect 9692 10704 9784 10706
rect 9734 10648 9784 10704
rect 9692 10646 9784 10648
rect 9857 10704 10107 10706
rect 9857 10648 9862 10704
rect 9918 10648 10046 10704
rect 10102 10648 10107 10704
rect 9857 10646 10107 10648
rect 9692 10644 9739 10646
rect 9673 10643 9739 10644
rect 9857 10643 9923 10646
rect 10041 10643 10107 10646
rect 10869 10706 10935 10709
rect 16665 10706 16731 10709
rect 10869 10704 16731 10706
rect 10869 10648 10874 10704
rect 10930 10648 16670 10704
rect 16726 10648 16731 10704
rect 10869 10646 16731 10648
rect 10869 10643 10935 10646
rect 16665 10643 16731 10646
rect 16849 10706 16915 10709
rect 16982 10706 16988 10708
rect 16849 10704 16988 10706
rect 16849 10648 16854 10704
rect 16910 10648 16988 10704
rect 16849 10646 16988 10648
rect 16849 10643 16915 10646
rect 16982 10644 16988 10646
rect 17052 10644 17058 10708
rect 6361 10570 6427 10573
rect 19609 10570 19675 10573
rect 22001 10570 22067 10573
rect 6361 10568 19675 10570
rect 6361 10512 6366 10568
rect 6422 10512 19614 10568
rect 19670 10512 19675 10568
rect 6361 10510 19675 10512
rect 6361 10507 6427 10510
rect 19609 10507 19675 10510
rect 19934 10568 22067 10570
rect 19934 10512 22006 10568
rect 22062 10512 22067 10568
rect 19934 10510 22067 10512
rect 10041 10434 10107 10437
rect 14181 10434 14247 10437
rect 10041 10432 14247 10434
rect 10041 10376 10046 10432
rect 10102 10376 14186 10432
rect 14242 10376 14247 10432
rect 10041 10374 14247 10376
rect 10041 10371 10107 10374
rect 14181 10371 14247 10374
rect 8341 10368 8661 10369
rect 8341 10304 8349 10368
rect 8413 10304 8429 10368
rect 8493 10304 8509 10368
rect 8573 10304 8589 10368
rect 8653 10304 8661 10368
rect 8341 10303 8661 10304
rect 15738 10368 16058 10369
rect 15738 10304 15746 10368
rect 15810 10304 15826 10368
rect 15890 10304 15906 10368
rect 15970 10304 15986 10368
rect 16050 10304 16058 10368
rect 15738 10303 16058 10304
rect 9653 10298 9719 10301
rect 11513 10298 11579 10301
rect 9653 10296 11579 10298
rect 9653 10240 9658 10296
rect 9714 10240 11518 10296
rect 11574 10240 11579 10296
rect 9653 10238 11579 10240
rect 9653 10235 9719 10238
rect 11513 10235 11579 10238
rect 14641 10298 14707 10301
rect 15377 10298 15443 10301
rect 19934 10298 19994 10510
rect 22001 10507 22067 10510
rect 14641 10296 15443 10298
rect 14641 10240 14646 10296
rect 14702 10240 15382 10296
rect 15438 10240 15443 10296
rect 14641 10238 15443 10240
rect 14641 10235 14707 10238
rect 15377 10235 15443 10238
rect 17174 10238 19994 10298
rect 7281 10162 7347 10165
rect 17174 10162 17234 10238
rect 7281 10160 17234 10162
rect 7281 10104 7286 10160
rect 7342 10104 17234 10160
rect 7281 10102 17234 10104
rect 19333 10162 19399 10165
rect 23600 10162 24400 10192
rect 19333 10160 24400 10162
rect 19333 10104 19338 10160
rect 19394 10104 24400 10160
rect 19333 10102 24400 10104
rect 7281 10099 7347 10102
rect 19333 10099 19399 10102
rect 23600 10072 24400 10102
rect 3601 10026 3667 10029
rect 5165 10026 5231 10029
rect 3601 10024 5231 10026
rect 3601 9968 3606 10024
rect 3662 9968 5170 10024
rect 5226 9968 5231 10024
rect 3601 9966 5231 9968
rect 3601 9963 3667 9966
rect 5165 9963 5231 9966
rect 7005 10026 7071 10029
rect 14365 10026 14431 10029
rect 16246 10026 16252 10028
rect 7005 10024 16252 10026
rect 7005 9968 7010 10024
rect 7066 9968 14370 10024
rect 14426 9968 16252 10024
rect 7005 9966 16252 9968
rect 7005 9963 7071 9966
rect 14365 9963 14431 9966
rect 16246 9964 16252 9966
rect 16316 9964 16322 10028
rect 17125 10026 17191 10029
rect 18321 10026 18387 10029
rect 17125 10024 18387 10026
rect 17125 9968 17130 10024
rect 17186 9968 18326 10024
rect 18382 9968 18387 10024
rect 17125 9966 18387 9968
rect 17125 9963 17191 9966
rect 18321 9963 18387 9966
rect 9857 9892 9923 9893
rect 9806 9890 9812 9892
rect 9766 9830 9812 9890
rect 9876 9888 9923 9892
rect 14181 9892 14247 9893
rect 14181 9890 14228 9892
rect 9918 9832 9923 9888
rect 9806 9828 9812 9830
rect 9876 9828 9923 9832
rect 14136 9888 14228 9890
rect 14136 9832 14186 9888
rect 14136 9830 14228 9832
rect 9857 9827 9923 9828
rect 14181 9828 14228 9830
rect 14292 9828 14298 9892
rect 15193 9890 15259 9893
rect 18086 9890 18092 9892
rect 15193 9888 18092 9890
rect 15193 9832 15198 9888
rect 15254 9832 18092 9888
rect 15193 9830 18092 9832
rect 14181 9827 14247 9828
rect 15193 9827 15259 9830
rect 18086 9828 18092 9830
rect 18156 9828 18162 9892
rect 4642 9824 4962 9825
rect 4642 9760 4650 9824
rect 4714 9760 4730 9824
rect 4794 9760 4810 9824
rect 4874 9760 4890 9824
rect 4954 9760 4962 9824
rect 4642 9759 4962 9760
rect 12040 9824 12360 9825
rect 12040 9760 12048 9824
rect 12112 9760 12128 9824
rect 12192 9760 12208 9824
rect 12272 9760 12288 9824
rect 12352 9760 12360 9824
rect 12040 9759 12360 9760
rect 19437 9824 19757 9825
rect 19437 9760 19445 9824
rect 19509 9760 19525 9824
rect 19589 9760 19605 9824
rect 19669 9760 19685 9824
rect 19749 9760 19757 9824
rect 19437 9759 19757 9760
rect 9673 9756 9739 9757
rect 9622 9692 9628 9756
rect 9692 9754 9739 9756
rect 15561 9754 15627 9757
rect 16614 9754 16620 9756
rect 9692 9752 9784 9754
rect 9734 9696 9784 9752
rect 9692 9694 9784 9696
rect 15561 9752 16620 9754
rect 15561 9696 15566 9752
rect 15622 9696 16620 9752
rect 15561 9694 16620 9696
rect 9692 9692 9739 9694
rect 9673 9691 9739 9692
rect 15561 9691 15627 9694
rect 16614 9692 16620 9694
rect 16684 9692 16690 9756
rect 4889 9618 4955 9621
rect 16113 9618 16179 9621
rect 23105 9618 23171 9621
rect 4889 9616 15578 9618
rect 4889 9560 4894 9616
rect 4950 9560 15578 9616
rect 4889 9558 15578 9560
rect 4889 9555 4955 9558
rect 7465 9482 7531 9485
rect 7925 9482 7991 9485
rect 11881 9482 11947 9485
rect 7465 9480 11947 9482
rect 7465 9424 7470 9480
rect 7526 9424 7930 9480
rect 7986 9424 11886 9480
rect 11942 9424 11947 9480
rect 7465 9422 11947 9424
rect 15518 9482 15578 9558
rect 16113 9616 23171 9618
rect 16113 9560 16118 9616
rect 16174 9560 23110 9616
rect 23166 9560 23171 9616
rect 16113 9558 23171 9560
rect 16113 9555 16179 9558
rect 23105 9555 23171 9558
rect 18505 9482 18571 9485
rect 23600 9482 24400 9512
rect 15518 9480 18571 9482
rect 15518 9424 18510 9480
rect 18566 9424 18571 9480
rect 15518 9422 18571 9424
rect 7465 9419 7531 9422
rect 7925 9419 7991 9422
rect 11881 9419 11947 9422
rect 18505 9419 18571 9422
rect 22878 9422 24400 9482
rect 17401 9346 17467 9349
rect 22878 9346 22938 9422
rect 23600 9392 24400 9422
rect 17401 9344 22938 9346
rect 17401 9288 17406 9344
rect 17462 9288 22938 9344
rect 17401 9286 22938 9288
rect 17401 9283 17467 9286
rect 8341 9280 8661 9281
rect 8341 9216 8349 9280
rect 8413 9216 8429 9280
rect 8493 9216 8509 9280
rect 8573 9216 8589 9280
rect 8653 9216 8661 9280
rect 8341 9215 8661 9216
rect 15738 9280 16058 9281
rect 15738 9216 15746 9280
rect 15810 9216 15826 9280
rect 15890 9216 15906 9280
rect 15970 9216 15986 9280
rect 16050 9216 16058 9280
rect 15738 9215 16058 9216
rect 14641 9210 14707 9213
rect 9078 9208 14707 9210
rect 9078 9152 14646 9208
rect 14702 9152 14707 9208
rect 9078 9150 14707 9152
rect 0 9074 800 9104
rect 1485 9074 1551 9077
rect 0 9072 1551 9074
rect 0 9016 1490 9072
rect 1546 9016 1551 9072
rect 0 9014 1551 9016
rect 0 8984 800 9014
rect 1485 9011 1551 9014
rect 5717 9074 5783 9077
rect 9078 9074 9138 9150
rect 14641 9147 14707 9150
rect 17309 9210 17375 9213
rect 18321 9210 18387 9213
rect 17309 9208 18387 9210
rect 17309 9152 17314 9208
rect 17370 9152 18326 9208
rect 18382 9152 18387 9208
rect 17309 9150 18387 9152
rect 17309 9147 17375 9150
rect 18321 9147 18387 9150
rect 20345 9210 20411 9213
rect 20478 9210 20484 9212
rect 20345 9208 20484 9210
rect 20345 9152 20350 9208
rect 20406 9152 20484 9208
rect 20345 9150 20484 9152
rect 20345 9147 20411 9150
rect 20478 9148 20484 9150
rect 20548 9148 20554 9212
rect 5717 9072 9138 9074
rect 5717 9016 5722 9072
rect 5778 9016 9138 9072
rect 5717 9014 9138 9016
rect 9213 9074 9279 9077
rect 16113 9074 16179 9077
rect 9213 9072 16179 9074
rect 9213 9016 9218 9072
rect 9274 9016 16118 9072
rect 16174 9016 16179 9072
rect 9213 9014 16179 9016
rect 5717 9011 5783 9014
rect 9213 9011 9279 9014
rect 16113 9011 16179 9014
rect 16389 9074 16455 9077
rect 20294 9074 20300 9076
rect 16389 9072 20300 9074
rect 16389 9016 16394 9072
rect 16450 9016 20300 9072
rect 16389 9014 20300 9016
rect 16389 9011 16455 9014
rect 20294 9012 20300 9014
rect 20364 9012 20370 9076
rect 7189 8938 7255 8941
rect 17033 8938 17099 8941
rect 7189 8936 17099 8938
rect 7189 8880 7194 8936
rect 7250 8880 17038 8936
rect 17094 8880 17099 8936
rect 7189 8878 17099 8880
rect 7189 8875 7255 8878
rect 17033 8875 17099 8878
rect 17166 8876 17172 8940
rect 17236 8938 17242 8940
rect 22829 8938 22895 8941
rect 17236 8936 22895 8938
rect 17236 8880 22834 8936
rect 22890 8880 22895 8936
rect 17236 8878 22895 8880
rect 17236 8876 17242 8878
rect 22829 8875 22895 8878
rect 5441 8802 5507 8805
rect 9213 8802 9279 8805
rect 5441 8800 9279 8802
rect 5441 8744 5446 8800
rect 5502 8744 9218 8800
rect 9274 8744 9279 8800
rect 5441 8742 9279 8744
rect 5441 8739 5507 8742
rect 9213 8739 9279 8742
rect 13445 8802 13511 8805
rect 16481 8802 16547 8805
rect 23600 8802 24400 8832
rect 13445 8800 16547 8802
rect 13445 8744 13450 8800
rect 13506 8744 16486 8800
rect 16542 8744 16547 8800
rect 13445 8742 16547 8744
rect 13445 8739 13511 8742
rect 16481 8739 16547 8742
rect 22878 8742 24400 8802
rect 4642 8736 4962 8737
rect 4642 8672 4650 8736
rect 4714 8672 4730 8736
rect 4794 8672 4810 8736
rect 4874 8672 4890 8736
rect 4954 8672 4962 8736
rect 4642 8671 4962 8672
rect 12040 8736 12360 8737
rect 12040 8672 12048 8736
rect 12112 8672 12128 8736
rect 12192 8672 12208 8736
rect 12272 8672 12288 8736
rect 12352 8672 12360 8736
rect 12040 8671 12360 8672
rect 19437 8736 19757 8737
rect 19437 8672 19445 8736
rect 19509 8672 19525 8736
rect 19589 8672 19605 8736
rect 19669 8672 19685 8736
rect 19749 8672 19757 8736
rect 19437 8671 19757 8672
rect 7465 8666 7531 8669
rect 11605 8666 11671 8669
rect 7465 8664 11671 8666
rect 7465 8608 7470 8664
rect 7526 8608 11610 8664
rect 11666 8608 11671 8664
rect 7465 8606 11671 8608
rect 7465 8603 7531 8606
rect 11605 8603 11671 8606
rect 15745 8666 15811 8669
rect 17861 8666 17927 8669
rect 15745 8664 17927 8666
rect 15745 8608 15750 8664
rect 15806 8608 17866 8664
rect 17922 8608 17927 8664
rect 15745 8606 17927 8608
rect 15745 8603 15811 8606
rect 17861 8603 17927 8606
rect 19926 8604 19932 8668
rect 19996 8666 20002 8668
rect 20253 8666 20319 8669
rect 19996 8664 20319 8666
rect 19996 8608 20258 8664
rect 20314 8608 20319 8664
rect 19996 8606 20319 8608
rect 19996 8604 20002 8606
rect 20253 8603 20319 8606
rect 5349 8530 5415 8533
rect 17166 8530 17172 8532
rect 5349 8528 17172 8530
rect 5349 8472 5354 8528
rect 5410 8472 17172 8528
rect 5349 8470 17172 8472
rect 5349 8467 5415 8470
rect 17166 8468 17172 8470
rect 17236 8468 17242 8532
rect 17861 8530 17927 8533
rect 22878 8530 22938 8742
rect 23600 8712 24400 8742
rect 17861 8528 22938 8530
rect 17861 8472 17866 8528
rect 17922 8472 22938 8528
rect 17861 8470 22938 8472
rect 17861 8467 17927 8470
rect 4705 8394 4771 8397
rect 19333 8394 19399 8397
rect 4705 8392 19399 8394
rect 4705 8336 4710 8392
rect 4766 8336 19338 8392
rect 19394 8336 19399 8392
rect 4705 8334 19399 8336
rect 4705 8331 4771 8334
rect 19333 8331 19399 8334
rect 19517 8394 19583 8397
rect 20110 8394 20116 8396
rect 19517 8392 20116 8394
rect 19517 8336 19522 8392
rect 19578 8336 20116 8392
rect 19517 8334 20116 8336
rect 19517 8331 19583 8334
rect 20110 8332 20116 8334
rect 20180 8332 20186 8396
rect 10685 8258 10751 8261
rect 13353 8258 13419 8261
rect 10685 8256 13419 8258
rect 10685 8200 10690 8256
rect 10746 8200 13358 8256
rect 13414 8200 13419 8256
rect 10685 8198 13419 8200
rect 10685 8195 10751 8198
rect 13353 8195 13419 8198
rect 13721 8258 13787 8261
rect 15377 8258 15443 8261
rect 13721 8256 15443 8258
rect 13721 8200 13726 8256
rect 13782 8200 15382 8256
rect 15438 8200 15443 8256
rect 13721 8198 15443 8200
rect 13721 8195 13787 8198
rect 15377 8195 15443 8198
rect 17861 8258 17927 8261
rect 19885 8258 19951 8261
rect 17861 8256 19951 8258
rect 17861 8200 17866 8256
rect 17922 8200 19890 8256
rect 19946 8200 19951 8256
rect 17861 8198 19951 8200
rect 17861 8195 17927 8198
rect 19885 8195 19951 8198
rect 20529 8258 20595 8261
rect 23600 8258 24400 8288
rect 20529 8256 24400 8258
rect 20529 8200 20534 8256
rect 20590 8200 24400 8256
rect 20529 8198 24400 8200
rect 20529 8195 20595 8198
rect 8341 8192 8661 8193
rect 8341 8128 8349 8192
rect 8413 8128 8429 8192
rect 8493 8128 8509 8192
rect 8573 8128 8589 8192
rect 8653 8128 8661 8192
rect 8341 8127 8661 8128
rect 15738 8192 16058 8193
rect 15738 8128 15746 8192
rect 15810 8128 15826 8192
rect 15890 8128 15906 8192
rect 15970 8128 15986 8192
rect 16050 8128 16058 8192
rect 23600 8168 24400 8198
rect 15738 8127 16058 8128
rect 10225 8122 10291 8125
rect 15377 8122 15443 8125
rect 10225 8120 15443 8122
rect 10225 8064 10230 8120
rect 10286 8064 15382 8120
rect 15438 8064 15443 8120
rect 10225 8062 15443 8064
rect 10225 8059 10291 8062
rect 15377 8059 15443 8062
rect 17033 8122 17099 8125
rect 19057 8122 19123 8125
rect 17033 8120 19123 8122
rect 17033 8064 17038 8120
rect 17094 8064 19062 8120
rect 19118 8064 19123 8120
rect 17033 8062 19123 8064
rect 17033 8059 17099 8062
rect 19057 8059 19123 8062
rect 19333 8122 19399 8125
rect 20478 8122 20484 8124
rect 19333 8120 20484 8122
rect 19333 8064 19338 8120
rect 19394 8064 20484 8120
rect 19333 8062 20484 8064
rect 19333 8059 19399 8062
rect 20478 8060 20484 8062
rect 20548 8060 20554 8124
rect 11053 7986 11119 7989
rect 18689 7986 18755 7989
rect 11053 7984 18755 7986
rect 11053 7928 11058 7984
rect 11114 7928 18694 7984
rect 18750 7928 18755 7984
rect 11053 7926 18755 7928
rect 11053 7923 11119 7926
rect 18689 7923 18755 7926
rect 18873 7986 18939 7989
rect 19701 7986 19767 7989
rect 18873 7984 19767 7986
rect 18873 7928 18878 7984
rect 18934 7928 19706 7984
rect 19762 7928 19767 7984
rect 18873 7926 19767 7928
rect 18873 7923 18939 7926
rect 19701 7923 19767 7926
rect 5625 7850 5691 7853
rect 12985 7850 13051 7853
rect 18873 7850 18939 7853
rect 19793 7850 19859 7853
rect 5625 7848 12818 7850
rect 5625 7792 5630 7848
rect 5686 7792 12818 7848
rect 5625 7790 12818 7792
rect 5625 7787 5691 7790
rect 12758 7714 12818 7790
rect 12985 7848 18939 7850
rect 12985 7792 12990 7848
rect 13046 7792 18878 7848
rect 18934 7792 18939 7848
rect 12985 7790 18939 7792
rect 12985 7787 13051 7790
rect 18873 7787 18939 7790
rect 19014 7848 19859 7850
rect 19014 7792 19798 7848
rect 19854 7792 19859 7848
rect 19014 7790 19859 7792
rect 17718 7714 17724 7716
rect 12758 7654 17724 7714
rect 17718 7652 17724 7654
rect 17788 7652 17794 7716
rect 18505 7714 18571 7717
rect 19014 7714 19074 7790
rect 19793 7787 19859 7790
rect 18505 7712 19074 7714
rect 18505 7656 18510 7712
rect 18566 7656 19074 7712
rect 18505 7654 19074 7656
rect 18505 7651 18571 7654
rect 4642 7648 4962 7649
rect 4642 7584 4650 7648
rect 4714 7584 4730 7648
rect 4794 7584 4810 7648
rect 4874 7584 4890 7648
rect 4954 7584 4962 7648
rect 4642 7583 4962 7584
rect 12040 7648 12360 7649
rect 12040 7584 12048 7648
rect 12112 7584 12128 7648
rect 12192 7584 12208 7648
rect 12272 7584 12288 7648
rect 12352 7584 12360 7648
rect 12040 7583 12360 7584
rect 19437 7648 19757 7649
rect 19437 7584 19445 7648
rect 19509 7584 19525 7648
rect 19589 7584 19605 7648
rect 19669 7584 19685 7648
rect 19749 7584 19757 7648
rect 19437 7583 19757 7584
rect 12433 7578 12499 7581
rect 16665 7578 16731 7581
rect 12433 7576 16731 7578
rect 12433 7520 12438 7576
rect 12494 7520 16670 7576
rect 16726 7520 16731 7576
rect 12433 7518 16731 7520
rect 12433 7515 12499 7518
rect 16665 7515 16731 7518
rect 20897 7578 20963 7581
rect 23600 7578 24400 7608
rect 20897 7576 24400 7578
rect 20897 7520 20902 7576
rect 20958 7520 24400 7576
rect 20897 7518 24400 7520
rect 20897 7515 20963 7518
rect 23600 7488 24400 7518
rect 6913 7442 6979 7445
rect 12985 7442 13051 7445
rect 6913 7440 13051 7442
rect 6913 7384 6918 7440
rect 6974 7384 12990 7440
rect 13046 7384 13051 7440
rect 6913 7382 13051 7384
rect 6913 7379 6979 7382
rect 12985 7379 13051 7382
rect 13353 7442 13419 7445
rect 16205 7442 16271 7445
rect 13353 7440 16271 7442
rect 13353 7384 13358 7440
rect 13414 7384 16210 7440
rect 16266 7384 16271 7440
rect 13353 7382 16271 7384
rect 13353 7379 13419 7382
rect 16205 7379 16271 7382
rect 17718 7380 17724 7444
rect 17788 7442 17794 7444
rect 22185 7442 22251 7445
rect 17788 7440 22251 7442
rect 17788 7384 22190 7440
rect 22246 7384 22251 7440
rect 17788 7382 22251 7384
rect 17788 7380 17794 7382
rect 22185 7379 22251 7382
rect 14917 7306 14983 7309
rect 15745 7306 15811 7309
rect 14917 7304 15811 7306
rect 14917 7248 14922 7304
rect 14978 7248 15750 7304
rect 15806 7248 15811 7304
rect 14917 7246 15811 7248
rect 14917 7243 14983 7246
rect 15745 7243 15811 7246
rect 17953 7306 18019 7309
rect 21725 7306 21791 7309
rect 17953 7304 21791 7306
rect 17953 7248 17958 7304
rect 18014 7248 21730 7304
rect 21786 7248 21791 7304
rect 17953 7246 21791 7248
rect 17953 7243 18019 7246
rect 21725 7243 21791 7246
rect 19006 7108 19012 7172
rect 19076 7170 19082 7172
rect 20069 7170 20135 7173
rect 19076 7168 20135 7170
rect 19076 7112 20074 7168
rect 20130 7112 20135 7168
rect 19076 7110 20135 7112
rect 19076 7108 19082 7110
rect 20069 7107 20135 7110
rect 8341 7104 8661 7105
rect 8341 7040 8349 7104
rect 8413 7040 8429 7104
rect 8493 7040 8509 7104
rect 8573 7040 8589 7104
rect 8653 7040 8661 7104
rect 8341 7039 8661 7040
rect 15738 7104 16058 7105
rect 15738 7040 15746 7104
rect 15810 7040 15826 7104
rect 15890 7040 15906 7104
rect 15970 7040 15986 7104
rect 16050 7040 16058 7104
rect 15738 7039 16058 7040
rect 8845 7034 8911 7037
rect 9581 7034 9647 7037
rect 8845 7032 9647 7034
rect 8845 6976 8850 7032
rect 8906 6976 9586 7032
rect 9642 6976 9647 7032
rect 8845 6974 9647 6976
rect 8845 6971 8911 6974
rect 9581 6971 9647 6974
rect 10869 7034 10935 7037
rect 13353 7034 13419 7037
rect 10869 7032 13419 7034
rect 10869 6976 10874 7032
rect 10930 6976 13358 7032
rect 13414 6976 13419 7032
rect 10869 6974 13419 6976
rect 10869 6971 10935 6974
rect 13353 6971 13419 6974
rect 10409 6898 10475 6901
rect 16481 6898 16547 6901
rect 10409 6896 16547 6898
rect 10409 6840 10414 6896
rect 10470 6840 16486 6896
rect 16542 6840 16547 6896
rect 10409 6838 16547 6840
rect 10409 6835 10475 6838
rect 16481 6835 16547 6838
rect 23381 6898 23447 6901
rect 23600 6898 24400 6928
rect 23381 6896 24400 6898
rect 23381 6840 23386 6896
rect 23442 6840 24400 6896
rect 23381 6838 24400 6840
rect 23381 6835 23447 6838
rect 23600 6808 24400 6838
rect 7557 6762 7623 6765
rect 13905 6762 13971 6765
rect 20345 6762 20411 6765
rect 7557 6760 20411 6762
rect 7557 6704 7562 6760
rect 7618 6704 13910 6760
rect 13966 6704 20350 6760
rect 20406 6704 20411 6760
rect 7557 6702 20411 6704
rect 7557 6699 7623 6702
rect 13905 6699 13971 6702
rect 20345 6699 20411 6702
rect 13629 6626 13695 6629
rect 17953 6626 18019 6629
rect 13629 6624 18019 6626
rect 13629 6568 13634 6624
rect 13690 6568 17958 6624
rect 18014 6568 18019 6624
rect 13629 6566 18019 6568
rect 13629 6563 13695 6566
rect 17953 6563 18019 6566
rect 4642 6560 4962 6561
rect 4642 6496 4650 6560
rect 4714 6496 4730 6560
rect 4794 6496 4810 6560
rect 4874 6496 4890 6560
rect 4954 6496 4962 6560
rect 4642 6495 4962 6496
rect 12040 6560 12360 6561
rect 12040 6496 12048 6560
rect 12112 6496 12128 6560
rect 12192 6496 12208 6560
rect 12272 6496 12288 6560
rect 12352 6496 12360 6560
rect 12040 6495 12360 6496
rect 19437 6560 19757 6561
rect 19437 6496 19445 6560
rect 19509 6496 19525 6560
rect 19589 6496 19605 6560
rect 19669 6496 19685 6560
rect 19749 6496 19757 6560
rect 19437 6495 19757 6496
rect 6821 6490 6887 6493
rect 10869 6490 10935 6493
rect 6821 6488 10935 6490
rect 6821 6432 6826 6488
rect 6882 6432 10874 6488
rect 10930 6432 10935 6488
rect 6821 6430 10935 6432
rect 6821 6427 6887 6430
rect 10869 6427 10935 6430
rect 14365 6490 14431 6493
rect 15009 6490 15075 6493
rect 16113 6490 16179 6493
rect 14365 6488 16179 6490
rect 14365 6432 14370 6488
rect 14426 6432 15014 6488
rect 15070 6432 16118 6488
rect 16174 6432 16179 6488
rect 14365 6430 16179 6432
rect 14365 6427 14431 6430
rect 15009 6427 15075 6430
rect 16113 6427 16179 6430
rect 8477 6354 8543 6357
rect 11697 6354 11763 6357
rect 16941 6354 17007 6357
rect 8477 6352 17007 6354
rect 8477 6296 8482 6352
rect 8538 6296 11702 6352
rect 11758 6296 16946 6352
rect 17002 6296 17007 6352
rect 8477 6294 17007 6296
rect 8477 6291 8543 6294
rect 11697 6291 11763 6294
rect 16941 6291 17007 6294
rect 19885 6356 19951 6357
rect 19885 6352 19932 6356
rect 19996 6354 20002 6356
rect 19885 6296 19890 6352
rect 19885 6292 19932 6296
rect 19996 6294 20042 6354
rect 19996 6292 20002 6294
rect 19885 6291 19951 6292
rect 11237 6218 11303 6221
rect 22553 6218 22619 6221
rect 23600 6218 24400 6248
rect 11237 6216 11346 6218
rect 11237 6160 11242 6216
rect 11298 6160 11346 6216
rect 11237 6155 11346 6160
rect 22553 6216 24400 6218
rect 22553 6160 22558 6216
rect 22614 6160 24400 6216
rect 22553 6158 24400 6160
rect 22553 6155 22619 6158
rect 11286 6082 11346 6155
rect 23600 6128 24400 6158
rect 11513 6082 11579 6085
rect 11286 6080 11579 6082
rect 11286 6024 11518 6080
rect 11574 6024 11579 6080
rect 11286 6022 11579 6024
rect 11513 6019 11579 6022
rect 17677 6082 17743 6085
rect 18045 6082 18111 6085
rect 17677 6080 18111 6082
rect 17677 6024 17682 6080
rect 17738 6024 18050 6080
rect 18106 6024 18111 6080
rect 17677 6022 18111 6024
rect 17677 6019 17743 6022
rect 18045 6019 18111 6022
rect 8341 6016 8661 6017
rect 8341 5952 8349 6016
rect 8413 5952 8429 6016
rect 8493 5952 8509 6016
rect 8573 5952 8589 6016
rect 8653 5952 8661 6016
rect 8341 5951 8661 5952
rect 15738 6016 16058 6017
rect 15738 5952 15746 6016
rect 15810 5952 15826 6016
rect 15890 5952 15906 6016
rect 15970 5952 15986 6016
rect 16050 5952 16058 6016
rect 15738 5951 16058 5952
rect 9765 5810 9831 5813
rect 14181 5810 14247 5813
rect 9765 5808 14247 5810
rect 9765 5752 9770 5808
rect 9826 5752 14186 5808
rect 14242 5752 14247 5808
rect 9765 5750 14247 5752
rect 9765 5747 9831 5750
rect 14181 5747 14247 5750
rect 16297 5810 16363 5813
rect 17861 5810 17927 5813
rect 18689 5810 18755 5813
rect 16297 5808 18755 5810
rect 16297 5752 16302 5808
rect 16358 5752 17866 5808
rect 17922 5752 18694 5808
rect 18750 5752 18755 5808
rect 16297 5750 18755 5752
rect 16297 5747 16363 5750
rect 17861 5747 17927 5750
rect 18689 5747 18755 5750
rect 12249 5674 12315 5677
rect 19241 5674 19307 5677
rect 12249 5672 19307 5674
rect 12249 5616 12254 5672
rect 12310 5616 19246 5672
rect 19302 5616 19307 5672
rect 12249 5614 19307 5616
rect 12249 5611 12315 5614
rect 19241 5611 19307 5614
rect 22829 5538 22895 5541
rect 23600 5538 24400 5568
rect 22829 5536 24400 5538
rect 22829 5480 22834 5536
rect 22890 5480 24400 5536
rect 22829 5478 24400 5480
rect 22829 5475 22895 5478
rect 4642 5472 4962 5473
rect 4642 5408 4650 5472
rect 4714 5408 4730 5472
rect 4794 5408 4810 5472
rect 4874 5408 4890 5472
rect 4954 5408 4962 5472
rect 4642 5407 4962 5408
rect 12040 5472 12360 5473
rect 12040 5408 12048 5472
rect 12112 5408 12128 5472
rect 12192 5408 12208 5472
rect 12272 5408 12288 5472
rect 12352 5408 12360 5472
rect 12040 5407 12360 5408
rect 19437 5472 19757 5473
rect 19437 5408 19445 5472
rect 19509 5408 19525 5472
rect 19589 5408 19605 5472
rect 19669 5408 19685 5472
rect 19749 5408 19757 5472
rect 23600 5448 24400 5478
rect 19437 5407 19757 5408
rect 20345 5402 20411 5405
rect 20345 5400 22938 5402
rect 20345 5344 20350 5400
rect 20406 5344 22938 5400
rect 20345 5342 22938 5344
rect 20345 5339 20411 5342
rect 8661 5266 8727 5269
rect 14365 5266 14431 5269
rect 8661 5264 14431 5266
rect 8661 5208 8666 5264
rect 8722 5208 14370 5264
rect 14426 5208 14431 5264
rect 8661 5206 14431 5208
rect 8661 5203 8727 5206
rect 14365 5203 14431 5206
rect 14825 5266 14891 5269
rect 18137 5266 18203 5269
rect 14825 5264 18203 5266
rect 14825 5208 14830 5264
rect 14886 5208 18142 5264
rect 18198 5208 18203 5264
rect 14825 5206 18203 5208
rect 14825 5203 14891 5206
rect 18137 5203 18203 5206
rect 19609 5266 19675 5269
rect 20897 5266 20963 5269
rect 19609 5264 20963 5266
rect 19609 5208 19614 5264
rect 19670 5208 20902 5264
rect 20958 5208 20963 5264
rect 19609 5206 20963 5208
rect 19609 5203 19675 5206
rect 20897 5203 20963 5206
rect 12249 5130 12315 5133
rect 13813 5130 13879 5133
rect 12249 5128 13879 5130
rect 12249 5072 12254 5128
rect 12310 5072 13818 5128
rect 13874 5072 13879 5128
rect 12249 5070 13879 5072
rect 12249 5067 12315 5070
rect 13813 5067 13879 5070
rect 14365 5130 14431 5133
rect 18689 5130 18755 5133
rect 14365 5128 18755 5130
rect 14365 5072 14370 5128
rect 14426 5072 18694 5128
rect 18750 5072 18755 5128
rect 14365 5070 18755 5072
rect 14365 5067 14431 5070
rect 18689 5067 18755 5070
rect 16941 4994 17007 4997
rect 22093 4994 22159 4997
rect 16941 4992 22159 4994
rect 16941 4936 16946 4992
rect 17002 4936 22098 4992
rect 22154 4936 22159 4992
rect 16941 4934 22159 4936
rect 16941 4931 17007 4934
rect 22093 4931 22159 4934
rect 8341 4928 8661 4929
rect 8341 4864 8349 4928
rect 8413 4864 8429 4928
rect 8493 4864 8509 4928
rect 8573 4864 8589 4928
rect 8653 4864 8661 4928
rect 8341 4863 8661 4864
rect 15738 4928 16058 4929
rect 15738 4864 15746 4928
rect 15810 4864 15826 4928
rect 15890 4864 15906 4928
rect 15970 4864 15986 4928
rect 16050 4864 16058 4928
rect 15738 4863 16058 4864
rect 22878 4858 22938 5342
rect 23600 4858 24400 4888
rect 22878 4798 24400 4858
rect 23600 4768 24400 4798
rect 5257 4722 5323 4725
rect 20713 4722 20779 4725
rect 5257 4720 20779 4722
rect 5257 4664 5262 4720
rect 5318 4664 20718 4720
rect 20774 4664 20779 4720
rect 5257 4662 20779 4664
rect 5257 4659 5323 4662
rect 20713 4659 20779 4662
rect 11605 4586 11671 4589
rect 16982 4586 16988 4588
rect 11605 4584 16988 4586
rect 11605 4528 11610 4584
rect 11666 4528 16988 4584
rect 11605 4526 16988 4528
rect 11605 4523 11671 4526
rect 16982 4524 16988 4526
rect 17052 4524 17058 4588
rect 14917 4450 14983 4453
rect 18689 4450 18755 4453
rect 14917 4448 18755 4450
rect 14917 4392 14922 4448
rect 14978 4392 18694 4448
rect 18750 4392 18755 4448
rect 14917 4390 18755 4392
rect 14917 4387 14983 4390
rect 18689 4387 18755 4390
rect 4642 4384 4962 4385
rect 4642 4320 4650 4384
rect 4714 4320 4730 4384
rect 4794 4320 4810 4384
rect 4874 4320 4890 4384
rect 4954 4320 4962 4384
rect 4642 4319 4962 4320
rect 12040 4384 12360 4385
rect 12040 4320 12048 4384
rect 12112 4320 12128 4384
rect 12192 4320 12208 4384
rect 12272 4320 12288 4384
rect 12352 4320 12360 4384
rect 12040 4319 12360 4320
rect 19437 4384 19757 4385
rect 19437 4320 19445 4384
rect 19509 4320 19525 4384
rect 19589 4320 19605 4384
rect 19669 4320 19685 4384
rect 19749 4320 19757 4384
rect 19437 4319 19757 4320
rect 22185 4314 22251 4317
rect 23600 4314 24400 4344
rect 22185 4312 24400 4314
rect 22185 4256 22190 4312
rect 22246 4256 24400 4312
rect 22185 4254 24400 4256
rect 22185 4251 22251 4254
rect 23600 4224 24400 4254
rect 16113 4178 16179 4181
rect 19333 4178 19399 4181
rect 16113 4176 19399 4178
rect 16113 4120 16118 4176
rect 16174 4120 19338 4176
rect 19394 4120 19399 4176
rect 16113 4118 19399 4120
rect 16113 4115 16179 4118
rect 19333 4115 19399 4118
rect 13169 4042 13235 4045
rect 13302 4042 13308 4044
rect 13169 4040 13308 4042
rect 13169 3984 13174 4040
rect 13230 3984 13308 4040
rect 13169 3982 13308 3984
rect 13169 3979 13235 3982
rect 13302 3980 13308 3982
rect 13372 3980 13378 4044
rect 21398 4042 21404 4044
rect 13494 3982 21404 4042
rect 13169 3906 13235 3909
rect 13494 3906 13554 3982
rect 21398 3980 21404 3982
rect 21468 3980 21474 4044
rect 13169 3904 13554 3906
rect 13169 3848 13174 3904
rect 13230 3848 13554 3904
rect 13169 3846 13554 3848
rect 13169 3843 13235 3846
rect 8341 3840 8661 3841
rect 8341 3776 8349 3840
rect 8413 3776 8429 3840
rect 8493 3776 8509 3840
rect 8573 3776 8589 3840
rect 8653 3776 8661 3840
rect 8341 3775 8661 3776
rect 15738 3840 16058 3841
rect 15738 3776 15746 3840
rect 15810 3776 15826 3840
rect 15890 3776 15906 3840
rect 15970 3776 15986 3840
rect 16050 3776 16058 3840
rect 15738 3775 16058 3776
rect 10317 3634 10383 3637
rect 19926 3634 19932 3636
rect 10317 3632 19932 3634
rect 10317 3576 10322 3632
rect 10378 3576 19932 3632
rect 10317 3574 19932 3576
rect 10317 3571 10383 3574
rect 19926 3572 19932 3574
rect 19996 3572 20002 3636
rect 20069 3634 20135 3637
rect 23600 3634 24400 3664
rect 20069 3632 24400 3634
rect 20069 3576 20074 3632
rect 20130 3576 24400 3632
rect 20069 3574 24400 3576
rect 19934 3498 19994 3572
rect 20069 3571 20135 3574
rect 23600 3544 24400 3574
rect 22093 3498 22159 3501
rect 19934 3496 22159 3498
rect 19934 3440 22098 3496
rect 22154 3440 22159 3496
rect 19934 3438 22159 3440
rect 22093 3435 22159 3438
rect 4642 3296 4962 3297
rect 4642 3232 4650 3296
rect 4714 3232 4730 3296
rect 4794 3232 4810 3296
rect 4874 3232 4890 3296
rect 4954 3232 4962 3296
rect 4642 3231 4962 3232
rect 12040 3296 12360 3297
rect 12040 3232 12048 3296
rect 12112 3232 12128 3296
rect 12192 3232 12208 3296
rect 12272 3232 12288 3296
rect 12352 3232 12360 3296
rect 12040 3231 12360 3232
rect 19437 3296 19757 3297
rect 19437 3232 19445 3296
rect 19509 3232 19525 3296
rect 19589 3232 19605 3296
rect 19669 3232 19685 3296
rect 19749 3232 19757 3296
rect 19437 3231 19757 3232
rect 13537 3226 13603 3229
rect 17677 3226 17743 3229
rect 13537 3224 17743 3226
rect 13537 3168 13542 3224
rect 13598 3168 17682 3224
rect 17738 3168 17743 3224
rect 13537 3166 17743 3168
rect 13537 3163 13603 3166
rect 17677 3163 17743 3166
rect 0 3090 800 3120
rect 1945 3090 2011 3093
rect 0 3088 2011 3090
rect 0 3032 1950 3088
rect 2006 3032 2011 3088
rect 0 3030 2011 3032
rect 0 3000 800 3030
rect 1945 3027 2011 3030
rect 20294 2892 20300 2956
rect 20364 2954 20370 2956
rect 23600 2954 24400 2984
rect 20364 2894 24400 2954
rect 20364 2892 20370 2894
rect 23600 2864 24400 2894
rect 8341 2752 8661 2753
rect 8341 2688 8349 2752
rect 8413 2688 8429 2752
rect 8493 2688 8509 2752
rect 8573 2688 8589 2752
rect 8653 2688 8661 2752
rect 8341 2687 8661 2688
rect 15738 2752 16058 2753
rect 15738 2688 15746 2752
rect 15810 2688 15826 2752
rect 15890 2688 15906 2752
rect 15970 2688 15986 2752
rect 16050 2688 16058 2752
rect 15738 2687 16058 2688
rect 15929 2546 15995 2549
rect 21582 2546 21588 2548
rect 15929 2544 21588 2546
rect 15929 2488 15934 2544
rect 15990 2488 21588 2544
rect 15929 2486 21588 2488
rect 15929 2483 15995 2486
rect 21582 2484 21588 2486
rect 21652 2484 21658 2548
rect 19885 2274 19951 2277
rect 23600 2274 24400 2304
rect 19885 2272 24400 2274
rect 19885 2216 19890 2272
rect 19946 2216 24400 2272
rect 19885 2214 24400 2216
rect 19885 2211 19951 2214
rect 4642 2208 4962 2209
rect 4642 2144 4650 2208
rect 4714 2144 4730 2208
rect 4794 2144 4810 2208
rect 4874 2144 4890 2208
rect 4954 2144 4962 2208
rect 4642 2143 4962 2144
rect 12040 2208 12360 2209
rect 12040 2144 12048 2208
rect 12112 2144 12128 2208
rect 12192 2144 12208 2208
rect 12272 2144 12288 2208
rect 12352 2144 12360 2208
rect 12040 2143 12360 2144
rect 19437 2208 19757 2209
rect 19437 2144 19445 2208
rect 19509 2144 19525 2208
rect 19589 2144 19605 2208
rect 19669 2144 19685 2208
rect 19749 2144 19757 2208
rect 23600 2184 24400 2214
rect 19437 2143 19757 2144
rect 21357 1594 21423 1597
rect 23600 1594 24400 1624
rect 21357 1592 24400 1594
rect 21357 1536 21362 1592
rect 21418 1536 24400 1592
rect 21357 1534 24400 1536
rect 21357 1531 21423 1534
rect 23600 1504 24400 1534
rect 22921 914 22987 917
rect 23600 914 24400 944
rect 22921 912 24400 914
rect 22921 856 22926 912
rect 22982 856 24400 912
rect 22921 854 24400 856
rect 22921 851 22987 854
rect 23600 824 24400 854
rect 21265 370 21331 373
rect 23600 370 24400 400
rect 21265 368 24400 370
rect 21265 312 21270 368
rect 21326 312 24400 368
rect 21265 310 24400 312
rect 21265 307 21331 310
rect 23600 280 24400 310
<< via3 >>
rect 4650 21788 4714 21792
rect 4650 21732 4654 21788
rect 4654 21732 4710 21788
rect 4710 21732 4714 21788
rect 4650 21728 4714 21732
rect 4730 21788 4794 21792
rect 4730 21732 4734 21788
rect 4734 21732 4790 21788
rect 4790 21732 4794 21788
rect 4730 21728 4794 21732
rect 4810 21788 4874 21792
rect 4810 21732 4814 21788
rect 4814 21732 4870 21788
rect 4870 21732 4874 21788
rect 4810 21728 4874 21732
rect 4890 21788 4954 21792
rect 4890 21732 4894 21788
rect 4894 21732 4950 21788
rect 4950 21732 4954 21788
rect 4890 21728 4954 21732
rect 12048 21788 12112 21792
rect 12048 21732 12052 21788
rect 12052 21732 12108 21788
rect 12108 21732 12112 21788
rect 12048 21728 12112 21732
rect 12128 21788 12192 21792
rect 12128 21732 12132 21788
rect 12132 21732 12188 21788
rect 12188 21732 12192 21788
rect 12128 21728 12192 21732
rect 12208 21788 12272 21792
rect 12208 21732 12212 21788
rect 12212 21732 12268 21788
rect 12268 21732 12272 21788
rect 12208 21728 12272 21732
rect 12288 21788 12352 21792
rect 12288 21732 12292 21788
rect 12292 21732 12348 21788
rect 12348 21732 12352 21788
rect 12288 21728 12352 21732
rect 19445 21788 19509 21792
rect 19445 21732 19449 21788
rect 19449 21732 19505 21788
rect 19505 21732 19509 21788
rect 19445 21728 19509 21732
rect 19525 21788 19589 21792
rect 19525 21732 19529 21788
rect 19529 21732 19585 21788
rect 19585 21732 19589 21788
rect 19525 21728 19589 21732
rect 19605 21788 19669 21792
rect 19605 21732 19609 21788
rect 19609 21732 19665 21788
rect 19665 21732 19669 21788
rect 19605 21728 19669 21732
rect 19685 21788 19749 21792
rect 19685 21732 19689 21788
rect 19689 21732 19745 21788
rect 19745 21732 19749 21788
rect 19685 21728 19749 21732
rect 8349 21244 8413 21248
rect 8349 21188 8353 21244
rect 8353 21188 8409 21244
rect 8409 21188 8413 21244
rect 8349 21184 8413 21188
rect 8429 21244 8493 21248
rect 8429 21188 8433 21244
rect 8433 21188 8489 21244
rect 8489 21188 8493 21244
rect 8429 21184 8493 21188
rect 8509 21244 8573 21248
rect 8509 21188 8513 21244
rect 8513 21188 8569 21244
rect 8569 21188 8573 21244
rect 8509 21184 8573 21188
rect 8589 21244 8653 21248
rect 8589 21188 8593 21244
rect 8593 21188 8649 21244
rect 8649 21188 8653 21244
rect 8589 21184 8653 21188
rect 15746 21244 15810 21248
rect 15746 21188 15750 21244
rect 15750 21188 15806 21244
rect 15806 21188 15810 21244
rect 15746 21184 15810 21188
rect 15826 21244 15890 21248
rect 15826 21188 15830 21244
rect 15830 21188 15886 21244
rect 15886 21188 15890 21244
rect 15826 21184 15890 21188
rect 15906 21244 15970 21248
rect 15906 21188 15910 21244
rect 15910 21188 15966 21244
rect 15966 21188 15970 21244
rect 15906 21184 15970 21188
rect 15986 21244 16050 21248
rect 15986 21188 15990 21244
rect 15990 21188 16046 21244
rect 16046 21188 16050 21244
rect 15986 21184 16050 21188
rect 13124 20844 13188 20908
rect 13308 20844 13372 20908
rect 4650 20700 4714 20704
rect 4650 20644 4654 20700
rect 4654 20644 4710 20700
rect 4710 20644 4714 20700
rect 4650 20640 4714 20644
rect 4730 20700 4794 20704
rect 4730 20644 4734 20700
rect 4734 20644 4790 20700
rect 4790 20644 4794 20700
rect 4730 20640 4794 20644
rect 4810 20700 4874 20704
rect 4810 20644 4814 20700
rect 4814 20644 4870 20700
rect 4870 20644 4874 20700
rect 4810 20640 4874 20644
rect 4890 20700 4954 20704
rect 4890 20644 4894 20700
rect 4894 20644 4950 20700
rect 4950 20644 4954 20700
rect 4890 20640 4954 20644
rect 12048 20700 12112 20704
rect 12048 20644 12052 20700
rect 12052 20644 12108 20700
rect 12108 20644 12112 20700
rect 12048 20640 12112 20644
rect 12128 20700 12192 20704
rect 12128 20644 12132 20700
rect 12132 20644 12188 20700
rect 12188 20644 12192 20700
rect 12128 20640 12192 20644
rect 12208 20700 12272 20704
rect 12208 20644 12212 20700
rect 12212 20644 12268 20700
rect 12268 20644 12272 20700
rect 12208 20640 12272 20644
rect 12288 20700 12352 20704
rect 12288 20644 12292 20700
rect 12292 20644 12348 20700
rect 12348 20644 12352 20700
rect 12288 20640 12352 20644
rect 19445 20700 19509 20704
rect 19445 20644 19449 20700
rect 19449 20644 19505 20700
rect 19505 20644 19509 20700
rect 19445 20640 19509 20644
rect 19525 20700 19589 20704
rect 19525 20644 19529 20700
rect 19529 20644 19585 20700
rect 19585 20644 19589 20700
rect 19525 20640 19589 20644
rect 19605 20700 19669 20704
rect 19605 20644 19609 20700
rect 19609 20644 19665 20700
rect 19665 20644 19669 20700
rect 19605 20640 19669 20644
rect 19685 20700 19749 20704
rect 19685 20644 19689 20700
rect 19689 20644 19745 20700
rect 19745 20644 19749 20700
rect 19685 20640 19749 20644
rect 8349 20156 8413 20160
rect 8349 20100 8353 20156
rect 8353 20100 8409 20156
rect 8409 20100 8413 20156
rect 8349 20096 8413 20100
rect 8429 20156 8493 20160
rect 8429 20100 8433 20156
rect 8433 20100 8489 20156
rect 8489 20100 8493 20156
rect 8429 20096 8493 20100
rect 8509 20156 8573 20160
rect 8509 20100 8513 20156
rect 8513 20100 8569 20156
rect 8569 20100 8573 20156
rect 8509 20096 8573 20100
rect 8589 20156 8653 20160
rect 8589 20100 8593 20156
rect 8593 20100 8649 20156
rect 8649 20100 8653 20156
rect 8589 20096 8653 20100
rect 15746 20156 15810 20160
rect 15746 20100 15750 20156
rect 15750 20100 15806 20156
rect 15806 20100 15810 20156
rect 15746 20096 15810 20100
rect 15826 20156 15890 20160
rect 15826 20100 15830 20156
rect 15830 20100 15886 20156
rect 15886 20100 15890 20156
rect 15826 20096 15890 20100
rect 15906 20156 15970 20160
rect 15906 20100 15910 20156
rect 15910 20100 15966 20156
rect 15966 20100 15970 20156
rect 15906 20096 15970 20100
rect 15986 20156 16050 20160
rect 15986 20100 15990 20156
rect 15990 20100 16046 20156
rect 16046 20100 16050 20156
rect 15986 20096 16050 20100
rect 20668 19892 20732 19956
rect 4650 19612 4714 19616
rect 4650 19556 4654 19612
rect 4654 19556 4710 19612
rect 4710 19556 4714 19612
rect 4650 19552 4714 19556
rect 4730 19612 4794 19616
rect 4730 19556 4734 19612
rect 4734 19556 4790 19612
rect 4790 19556 4794 19612
rect 4730 19552 4794 19556
rect 4810 19612 4874 19616
rect 4810 19556 4814 19612
rect 4814 19556 4870 19612
rect 4870 19556 4874 19612
rect 4810 19552 4874 19556
rect 4890 19612 4954 19616
rect 4890 19556 4894 19612
rect 4894 19556 4950 19612
rect 4950 19556 4954 19612
rect 4890 19552 4954 19556
rect 12048 19612 12112 19616
rect 12048 19556 12052 19612
rect 12052 19556 12108 19612
rect 12108 19556 12112 19612
rect 12048 19552 12112 19556
rect 12128 19612 12192 19616
rect 12128 19556 12132 19612
rect 12132 19556 12188 19612
rect 12188 19556 12192 19612
rect 12128 19552 12192 19556
rect 12208 19612 12272 19616
rect 12208 19556 12212 19612
rect 12212 19556 12268 19612
rect 12268 19556 12272 19612
rect 12208 19552 12272 19556
rect 12288 19612 12352 19616
rect 12288 19556 12292 19612
rect 12292 19556 12348 19612
rect 12348 19556 12352 19612
rect 12288 19552 12352 19556
rect 19445 19612 19509 19616
rect 19445 19556 19449 19612
rect 19449 19556 19505 19612
rect 19505 19556 19509 19612
rect 19445 19552 19509 19556
rect 19525 19612 19589 19616
rect 19525 19556 19529 19612
rect 19529 19556 19585 19612
rect 19585 19556 19589 19612
rect 19525 19552 19589 19556
rect 19605 19612 19669 19616
rect 19605 19556 19609 19612
rect 19609 19556 19665 19612
rect 19665 19556 19669 19612
rect 19605 19552 19669 19556
rect 19685 19612 19749 19616
rect 19685 19556 19689 19612
rect 19689 19556 19745 19612
rect 19745 19556 19749 19612
rect 19685 19552 19749 19556
rect 13492 19212 13556 19276
rect 8349 19068 8413 19072
rect 8349 19012 8353 19068
rect 8353 19012 8409 19068
rect 8409 19012 8413 19068
rect 8349 19008 8413 19012
rect 8429 19068 8493 19072
rect 8429 19012 8433 19068
rect 8433 19012 8489 19068
rect 8489 19012 8493 19068
rect 8429 19008 8493 19012
rect 8509 19068 8573 19072
rect 8509 19012 8513 19068
rect 8513 19012 8569 19068
rect 8569 19012 8573 19068
rect 8509 19008 8573 19012
rect 8589 19068 8653 19072
rect 8589 19012 8593 19068
rect 8593 19012 8649 19068
rect 8649 19012 8653 19068
rect 8589 19008 8653 19012
rect 15746 19068 15810 19072
rect 15746 19012 15750 19068
rect 15750 19012 15806 19068
rect 15806 19012 15810 19068
rect 15746 19008 15810 19012
rect 15826 19068 15890 19072
rect 15826 19012 15830 19068
rect 15830 19012 15886 19068
rect 15886 19012 15890 19068
rect 15826 19008 15890 19012
rect 15906 19068 15970 19072
rect 15906 19012 15910 19068
rect 15910 19012 15966 19068
rect 15966 19012 15970 19068
rect 15906 19008 15970 19012
rect 15986 19068 16050 19072
rect 15986 19012 15990 19068
rect 15990 19012 16046 19068
rect 16046 19012 16050 19068
rect 15986 19008 16050 19012
rect 16988 18668 17052 18732
rect 19012 18668 19076 18732
rect 4650 18524 4714 18528
rect 4650 18468 4654 18524
rect 4654 18468 4710 18524
rect 4710 18468 4714 18524
rect 4650 18464 4714 18468
rect 4730 18524 4794 18528
rect 4730 18468 4734 18524
rect 4734 18468 4790 18524
rect 4790 18468 4794 18524
rect 4730 18464 4794 18468
rect 4810 18524 4874 18528
rect 4810 18468 4814 18524
rect 4814 18468 4870 18524
rect 4870 18468 4874 18524
rect 4810 18464 4874 18468
rect 4890 18524 4954 18528
rect 4890 18468 4894 18524
rect 4894 18468 4950 18524
rect 4950 18468 4954 18524
rect 4890 18464 4954 18468
rect 12048 18524 12112 18528
rect 12048 18468 12052 18524
rect 12052 18468 12108 18524
rect 12108 18468 12112 18524
rect 12048 18464 12112 18468
rect 12128 18524 12192 18528
rect 12128 18468 12132 18524
rect 12132 18468 12188 18524
rect 12188 18468 12192 18524
rect 12128 18464 12192 18468
rect 12208 18524 12272 18528
rect 12208 18468 12212 18524
rect 12212 18468 12268 18524
rect 12268 18468 12272 18524
rect 12208 18464 12272 18468
rect 12288 18524 12352 18528
rect 12288 18468 12292 18524
rect 12292 18468 12348 18524
rect 12348 18468 12352 18524
rect 12288 18464 12352 18468
rect 19445 18524 19509 18528
rect 19445 18468 19449 18524
rect 19449 18468 19505 18524
rect 19505 18468 19509 18524
rect 19445 18464 19509 18468
rect 19525 18524 19589 18528
rect 19525 18468 19529 18524
rect 19529 18468 19585 18524
rect 19585 18468 19589 18524
rect 19525 18464 19589 18468
rect 19605 18524 19669 18528
rect 19605 18468 19609 18524
rect 19609 18468 19665 18524
rect 19665 18468 19669 18524
rect 19605 18464 19669 18468
rect 19685 18524 19749 18528
rect 19685 18468 19689 18524
rect 19689 18468 19745 18524
rect 19745 18468 19749 18524
rect 19685 18464 19749 18468
rect 20116 18456 20180 18460
rect 20116 18400 20130 18456
rect 20130 18400 20180 18456
rect 20116 18396 20180 18400
rect 14228 18124 14292 18188
rect 13124 18048 13188 18052
rect 19932 18124 19996 18188
rect 13124 17992 13174 18048
rect 13174 17992 13188 18048
rect 13124 17988 13188 17992
rect 21404 18048 21468 18052
rect 21404 17992 21418 18048
rect 21418 17992 21468 18048
rect 21404 17988 21468 17992
rect 21588 18048 21652 18052
rect 21588 17992 21638 18048
rect 21638 17992 21652 18048
rect 21588 17988 21652 17992
rect 8349 17980 8413 17984
rect 8349 17924 8353 17980
rect 8353 17924 8409 17980
rect 8409 17924 8413 17980
rect 8349 17920 8413 17924
rect 8429 17980 8493 17984
rect 8429 17924 8433 17980
rect 8433 17924 8489 17980
rect 8489 17924 8493 17980
rect 8429 17920 8493 17924
rect 8509 17980 8573 17984
rect 8509 17924 8513 17980
rect 8513 17924 8569 17980
rect 8569 17924 8573 17980
rect 8509 17920 8573 17924
rect 8589 17980 8653 17984
rect 8589 17924 8593 17980
rect 8593 17924 8649 17980
rect 8649 17924 8653 17980
rect 8589 17920 8653 17924
rect 15746 17980 15810 17984
rect 15746 17924 15750 17980
rect 15750 17924 15806 17980
rect 15806 17924 15810 17980
rect 15746 17920 15810 17924
rect 15826 17980 15890 17984
rect 15826 17924 15830 17980
rect 15830 17924 15886 17980
rect 15886 17924 15890 17980
rect 15826 17920 15890 17924
rect 15906 17980 15970 17984
rect 15906 17924 15910 17980
rect 15910 17924 15966 17980
rect 15966 17924 15970 17980
rect 15906 17920 15970 17924
rect 15986 17980 16050 17984
rect 15986 17924 15990 17980
rect 15990 17924 16046 17980
rect 16046 17924 16050 17980
rect 15986 17920 16050 17924
rect 19196 17716 19260 17780
rect 16436 17580 16500 17644
rect 13124 17444 13188 17508
rect 4650 17436 4714 17440
rect 4650 17380 4654 17436
rect 4654 17380 4710 17436
rect 4710 17380 4714 17436
rect 4650 17376 4714 17380
rect 4730 17436 4794 17440
rect 4730 17380 4734 17436
rect 4734 17380 4790 17436
rect 4790 17380 4794 17436
rect 4730 17376 4794 17380
rect 4810 17436 4874 17440
rect 4810 17380 4814 17436
rect 4814 17380 4870 17436
rect 4870 17380 4874 17436
rect 4810 17376 4874 17380
rect 4890 17436 4954 17440
rect 4890 17380 4894 17436
rect 4894 17380 4950 17436
rect 4950 17380 4954 17436
rect 4890 17376 4954 17380
rect 12048 17436 12112 17440
rect 12048 17380 12052 17436
rect 12052 17380 12108 17436
rect 12108 17380 12112 17436
rect 12048 17376 12112 17380
rect 12128 17436 12192 17440
rect 12128 17380 12132 17436
rect 12132 17380 12188 17436
rect 12188 17380 12192 17436
rect 12128 17376 12192 17380
rect 12208 17436 12272 17440
rect 12208 17380 12212 17436
rect 12212 17380 12268 17436
rect 12268 17380 12272 17436
rect 12208 17376 12272 17380
rect 12288 17436 12352 17440
rect 12288 17380 12292 17436
rect 12292 17380 12348 17436
rect 12348 17380 12352 17436
rect 12288 17376 12352 17380
rect 19445 17436 19509 17440
rect 19445 17380 19449 17436
rect 19449 17380 19505 17436
rect 19505 17380 19509 17436
rect 19445 17376 19509 17380
rect 19525 17436 19589 17440
rect 19525 17380 19529 17436
rect 19529 17380 19585 17436
rect 19585 17380 19589 17436
rect 19525 17376 19589 17380
rect 19605 17436 19669 17440
rect 19605 17380 19609 17436
rect 19609 17380 19665 17436
rect 19665 17380 19669 17436
rect 19605 17376 19669 17380
rect 19685 17436 19749 17440
rect 19685 17380 19689 17436
rect 19689 17380 19745 17436
rect 19745 17380 19749 17436
rect 19685 17376 19749 17380
rect 17908 17172 17972 17236
rect 18092 16960 18156 16964
rect 18092 16904 18142 16960
rect 18142 16904 18156 16960
rect 18092 16900 18156 16904
rect 8349 16892 8413 16896
rect 8349 16836 8353 16892
rect 8353 16836 8409 16892
rect 8409 16836 8413 16892
rect 8349 16832 8413 16836
rect 8429 16892 8493 16896
rect 8429 16836 8433 16892
rect 8433 16836 8489 16892
rect 8489 16836 8493 16892
rect 8429 16832 8493 16836
rect 8509 16892 8573 16896
rect 8509 16836 8513 16892
rect 8513 16836 8569 16892
rect 8569 16836 8573 16892
rect 8509 16832 8573 16836
rect 8589 16892 8653 16896
rect 8589 16836 8593 16892
rect 8593 16836 8649 16892
rect 8649 16836 8653 16892
rect 8589 16832 8653 16836
rect 15746 16892 15810 16896
rect 15746 16836 15750 16892
rect 15750 16836 15806 16892
rect 15806 16836 15810 16892
rect 15746 16832 15810 16836
rect 15826 16892 15890 16896
rect 15826 16836 15830 16892
rect 15830 16836 15886 16892
rect 15886 16836 15890 16892
rect 15826 16832 15890 16836
rect 15906 16892 15970 16896
rect 15906 16836 15910 16892
rect 15910 16836 15966 16892
rect 15966 16836 15970 16892
rect 15906 16832 15970 16836
rect 15986 16892 16050 16896
rect 15986 16836 15990 16892
rect 15990 16836 16046 16892
rect 16046 16836 16050 16892
rect 15986 16832 16050 16836
rect 17172 16764 17236 16828
rect 4650 16348 4714 16352
rect 4650 16292 4654 16348
rect 4654 16292 4710 16348
rect 4710 16292 4714 16348
rect 4650 16288 4714 16292
rect 4730 16348 4794 16352
rect 4730 16292 4734 16348
rect 4734 16292 4790 16348
rect 4790 16292 4794 16348
rect 4730 16288 4794 16292
rect 4810 16348 4874 16352
rect 4810 16292 4814 16348
rect 4814 16292 4870 16348
rect 4870 16292 4874 16348
rect 4810 16288 4874 16292
rect 4890 16348 4954 16352
rect 4890 16292 4894 16348
rect 4894 16292 4950 16348
rect 4950 16292 4954 16348
rect 4890 16288 4954 16292
rect 12048 16348 12112 16352
rect 12048 16292 12052 16348
rect 12052 16292 12108 16348
rect 12108 16292 12112 16348
rect 12048 16288 12112 16292
rect 12128 16348 12192 16352
rect 12128 16292 12132 16348
rect 12132 16292 12188 16348
rect 12188 16292 12192 16348
rect 12128 16288 12192 16292
rect 12208 16348 12272 16352
rect 12208 16292 12212 16348
rect 12212 16292 12268 16348
rect 12268 16292 12272 16348
rect 12208 16288 12272 16292
rect 12288 16348 12352 16352
rect 12288 16292 12292 16348
rect 12292 16292 12348 16348
rect 12348 16292 12352 16348
rect 12288 16288 12352 16292
rect 19445 16348 19509 16352
rect 19445 16292 19449 16348
rect 19449 16292 19505 16348
rect 19505 16292 19509 16348
rect 19445 16288 19509 16292
rect 19525 16348 19589 16352
rect 19525 16292 19529 16348
rect 19529 16292 19585 16348
rect 19585 16292 19589 16348
rect 19525 16288 19589 16292
rect 19605 16348 19669 16352
rect 19605 16292 19609 16348
rect 19609 16292 19665 16348
rect 19665 16292 19669 16348
rect 19605 16288 19669 16292
rect 19685 16348 19749 16352
rect 19685 16292 19689 16348
rect 19689 16292 19745 16348
rect 19745 16292 19749 16348
rect 19685 16288 19749 16292
rect 19196 16280 19260 16284
rect 19196 16224 19246 16280
rect 19246 16224 19260 16280
rect 19196 16220 19260 16224
rect 19196 16084 19260 16148
rect 8349 15804 8413 15808
rect 8349 15748 8353 15804
rect 8353 15748 8409 15804
rect 8409 15748 8413 15804
rect 8349 15744 8413 15748
rect 8429 15804 8493 15808
rect 8429 15748 8433 15804
rect 8433 15748 8489 15804
rect 8489 15748 8493 15804
rect 8429 15744 8493 15748
rect 8509 15804 8573 15808
rect 8509 15748 8513 15804
rect 8513 15748 8569 15804
rect 8569 15748 8573 15804
rect 8509 15744 8573 15748
rect 8589 15804 8653 15808
rect 8589 15748 8593 15804
rect 8593 15748 8649 15804
rect 8649 15748 8653 15804
rect 8589 15744 8653 15748
rect 15746 15804 15810 15808
rect 15746 15748 15750 15804
rect 15750 15748 15806 15804
rect 15806 15748 15810 15804
rect 15746 15744 15810 15748
rect 15826 15804 15890 15808
rect 15826 15748 15830 15804
rect 15830 15748 15886 15804
rect 15886 15748 15890 15804
rect 15826 15744 15890 15748
rect 15906 15804 15970 15808
rect 15906 15748 15910 15804
rect 15910 15748 15966 15804
rect 15966 15748 15970 15804
rect 15906 15744 15970 15748
rect 15986 15804 16050 15808
rect 15986 15748 15990 15804
rect 15990 15748 16046 15804
rect 16046 15748 16050 15804
rect 15986 15744 16050 15748
rect 16804 15268 16868 15332
rect 4650 15260 4714 15264
rect 4650 15204 4654 15260
rect 4654 15204 4710 15260
rect 4710 15204 4714 15260
rect 4650 15200 4714 15204
rect 4730 15260 4794 15264
rect 4730 15204 4734 15260
rect 4734 15204 4790 15260
rect 4790 15204 4794 15260
rect 4730 15200 4794 15204
rect 4810 15260 4874 15264
rect 4810 15204 4814 15260
rect 4814 15204 4870 15260
rect 4870 15204 4874 15260
rect 4810 15200 4874 15204
rect 4890 15260 4954 15264
rect 4890 15204 4894 15260
rect 4894 15204 4950 15260
rect 4950 15204 4954 15260
rect 4890 15200 4954 15204
rect 12048 15260 12112 15264
rect 12048 15204 12052 15260
rect 12052 15204 12108 15260
rect 12108 15204 12112 15260
rect 12048 15200 12112 15204
rect 12128 15260 12192 15264
rect 12128 15204 12132 15260
rect 12132 15204 12188 15260
rect 12188 15204 12192 15260
rect 12128 15200 12192 15204
rect 12208 15260 12272 15264
rect 12208 15204 12212 15260
rect 12212 15204 12268 15260
rect 12268 15204 12272 15260
rect 12208 15200 12272 15204
rect 12288 15260 12352 15264
rect 12288 15204 12292 15260
rect 12292 15204 12348 15260
rect 12348 15204 12352 15260
rect 12288 15200 12352 15204
rect 19445 15260 19509 15264
rect 19445 15204 19449 15260
rect 19449 15204 19505 15260
rect 19505 15204 19509 15260
rect 19445 15200 19509 15204
rect 19525 15260 19589 15264
rect 19525 15204 19529 15260
rect 19529 15204 19585 15260
rect 19585 15204 19589 15260
rect 19525 15200 19589 15204
rect 19605 15260 19669 15264
rect 19605 15204 19609 15260
rect 19609 15204 19665 15260
rect 19665 15204 19669 15260
rect 19605 15200 19669 15204
rect 19685 15260 19749 15264
rect 19685 15204 19689 15260
rect 19689 15204 19745 15260
rect 19745 15204 19749 15260
rect 19685 15200 19749 15204
rect 16620 14860 16684 14924
rect 8349 14716 8413 14720
rect 8349 14660 8353 14716
rect 8353 14660 8409 14716
rect 8409 14660 8413 14716
rect 8349 14656 8413 14660
rect 8429 14716 8493 14720
rect 8429 14660 8433 14716
rect 8433 14660 8489 14716
rect 8489 14660 8493 14716
rect 8429 14656 8493 14660
rect 8509 14716 8573 14720
rect 8509 14660 8513 14716
rect 8513 14660 8569 14716
rect 8569 14660 8573 14716
rect 8509 14656 8573 14660
rect 8589 14716 8653 14720
rect 8589 14660 8593 14716
rect 8593 14660 8649 14716
rect 8649 14660 8653 14716
rect 8589 14656 8653 14660
rect 15746 14716 15810 14720
rect 15746 14660 15750 14716
rect 15750 14660 15806 14716
rect 15806 14660 15810 14716
rect 15746 14656 15810 14660
rect 15826 14716 15890 14720
rect 15826 14660 15830 14716
rect 15830 14660 15886 14716
rect 15886 14660 15890 14716
rect 15826 14656 15890 14660
rect 15906 14716 15970 14720
rect 15906 14660 15910 14716
rect 15910 14660 15966 14716
rect 15966 14660 15970 14716
rect 15906 14656 15970 14660
rect 15986 14716 16050 14720
rect 15986 14660 15990 14716
rect 15990 14660 16046 14716
rect 16046 14660 16050 14716
rect 15986 14656 16050 14660
rect 16252 14588 16316 14652
rect 4650 14172 4714 14176
rect 4650 14116 4654 14172
rect 4654 14116 4710 14172
rect 4710 14116 4714 14172
rect 4650 14112 4714 14116
rect 4730 14172 4794 14176
rect 4730 14116 4734 14172
rect 4734 14116 4790 14172
rect 4790 14116 4794 14172
rect 4730 14112 4794 14116
rect 4810 14172 4874 14176
rect 4810 14116 4814 14172
rect 4814 14116 4870 14172
rect 4870 14116 4874 14172
rect 4810 14112 4874 14116
rect 4890 14172 4954 14176
rect 4890 14116 4894 14172
rect 4894 14116 4950 14172
rect 4950 14116 4954 14172
rect 4890 14112 4954 14116
rect 12048 14172 12112 14176
rect 12048 14116 12052 14172
rect 12052 14116 12108 14172
rect 12108 14116 12112 14172
rect 12048 14112 12112 14116
rect 12128 14172 12192 14176
rect 12128 14116 12132 14172
rect 12132 14116 12188 14172
rect 12188 14116 12192 14172
rect 12128 14112 12192 14116
rect 12208 14172 12272 14176
rect 12208 14116 12212 14172
rect 12212 14116 12268 14172
rect 12268 14116 12272 14172
rect 12208 14112 12272 14116
rect 12288 14172 12352 14176
rect 12288 14116 12292 14172
rect 12292 14116 12348 14172
rect 12348 14116 12352 14172
rect 12288 14112 12352 14116
rect 19445 14172 19509 14176
rect 19445 14116 19449 14172
rect 19449 14116 19505 14172
rect 19505 14116 19509 14172
rect 19445 14112 19509 14116
rect 19525 14172 19589 14176
rect 19525 14116 19529 14172
rect 19529 14116 19585 14172
rect 19585 14116 19589 14172
rect 19525 14112 19589 14116
rect 19605 14172 19669 14176
rect 19605 14116 19609 14172
rect 19609 14116 19665 14172
rect 19665 14116 19669 14172
rect 19605 14112 19669 14116
rect 19685 14172 19749 14176
rect 19685 14116 19689 14172
rect 19689 14116 19745 14172
rect 19745 14116 19749 14172
rect 19685 14112 19749 14116
rect 13492 14044 13556 14108
rect 16988 13908 17052 13972
rect 16804 13636 16868 13700
rect 19932 13636 19996 13700
rect 8349 13628 8413 13632
rect 8349 13572 8353 13628
rect 8353 13572 8409 13628
rect 8409 13572 8413 13628
rect 8349 13568 8413 13572
rect 8429 13628 8493 13632
rect 8429 13572 8433 13628
rect 8433 13572 8489 13628
rect 8489 13572 8493 13628
rect 8429 13568 8493 13572
rect 8509 13628 8573 13632
rect 8509 13572 8513 13628
rect 8513 13572 8569 13628
rect 8569 13572 8573 13628
rect 8509 13568 8573 13572
rect 8589 13628 8653 13632
rect 8589 13572 8593 13628
rect 8593 13572 8649 13628
rect 8649 13572 8653 13628
rect 8589 13568 8653 13572
rect 15746 13628 15810 13632
rect 15746 13572 15750 13628
rect 15750 13572 15806 13628
rect 15806 13572 15810 13628
rect 15746 13568 15810 13572
rect 15826 13628 15890 13632
rect 15826 13572 15830 13628
rect 15830 13572 15886 13628
rect 15886 13572 15890 13628
rect 15826 13568 15890 13572
rect 15906 13628 15970 13632
rect 15906 13572 15910 13628
rect 15910 13572 15966 13628
rect 15966 13572 15970 13628
rect 15906 13568 15970 13572
rect 15986 13628 16050 13632
rect 15986 13572 15990 13628
rect 15990 13572 16046 13628
rect 16046 13572 16050 13628
rect 15986 13568 16050 13572
rect 13124 13560 13188 13564
rect 13124 13504 13138 13560
rect 13138 13504 13188 13560
rect 13124 13500 13188 13504
rect 17908 13092 17972 13156
rect 4650 13084 4714 13088
rect 4650 13028 4654 13084
rect 4654 13028 4710 13084
rect 4710 13028 4714 13084
rect 4650 13024 4714 13028
rect 4730 13084 4794 13088
rect 4730 13028 4734 13084
rect 4734 13028 4790 13084
rect 4790 13028 4794 13084
rect 4730 13024 4794 13028
rect 4810 13084 4874 13088
rect 4810 13028 4814 13084
rect 4814 13028 4870 13084
rect 4870 13028 4874 13084
rect 4810 13024 4874 13028
rect 4890 13084 4954 13088
rect 4890 13028 4894 13084
rect 4894 13028 4950 13084
rect 4950 13028 4954 13084
rect 4890 13024 4954 13028
rect 12048 13084 12112 13088
rect 12048 13028 12052 13084
rect 12052 13028 12108 13084
rect 12108 13028 12112 13084
rect 12048 13024 12112 13028
rect 12128 13084 12192 13088
rect 12128 13028 12132 13084
rect 12132 13028 12188 13084
rect 12188 13028 12192 13084
rect 12128 13024 12192 13028
rect 12208 13084 12272 13088
rect 12208 13028 12212 13084
rect 12212 13028 12268 13084
rect 12268 13028 12272 13084
rect 12208 13024 12272 13028
rect 12288 13084 12352 13088
rect 12288 13028 12292 13084
rect 12292 13028 12348 13084
rect 12348 13028 12352 13084
rect 12288 13024 12352 13028
rect 19445 13084 19509 13088
rect 19445 13028 19449 13084
rect 19449 13028 19505 13084
rect 19505 13028 19509 13084
rect 19445 13024 19509 13028
rect 19525 13084 19589 13088
rect 19525 13028 19529 13084
rect 19529 13028 19585 13084
rect 19585 13028 19589 13084
rect 19525 13024 19589 13028
rect 19605 13084 19669 13088
rect 19605 13028 19609 13084
rect 19609 13028 19665 13084
rect 19665 13028 19669 13084
rect 19605 13024 19669 13028
rect 19685 13084 19749 13088
rect 19685 13028 19689 13084
rect 19689 13028 19745 13084
rect 19745 13028 19749 13084
rect 19685 13024 19749 13028
rect 17172 12820 17236 12884
rect 18644 12820 18708 12884
rect 19932 12820 19996 12884
rect 16436 12548 16500 12612
rect 20300 12608 20364 12612
rect 20300 12552 20314 12608
rect 20314 12552 20364 12608
rect 20300 12548 20364 12552
rect 8349 12540 8413 12544
rect 8349 12484 8353 12540
rect 8353 12484 8409 12540
rect 8409 12484 8413 12540
rect 8349 12480 8413 12484
rect 8429 12540 8493 12544
rect 8429 12484 8433 12540
rect 8433 12484 8489 12540
rect 8489 12484 8493 12540
rect 8429 12480 8493 12484
rect 8509 12540 8573 12544
rect 8509 12484 8513 12540
rect 8513 12484 8569 12540
rect 8569 12484 8573 12540
rect 8509 12480 8573 12484
rect 8589 12540 8653 12544
rect 8589 12484 8593 12540
rect 8593 12484 8649 12540
rect 8649 12484 8653 12540
rect 8589 12480 8653 12484
rect 15746 12540 15810 12544
rect 15746 12484 15750 12540
rect 15750 12484 15806 12540
rect 15806 12484 15810 12540
rect 15746 12480 15810 12484
rect 15826 12540 15890 12544
rect 15826 12484 15830 12540
rect 15830 12484 15886 12540
rect 15886 12484 15890 12540
rect 15826 12480 15890 12484
rect 15906 12540 15970 12544
rect 15906 12484 15910 12540
rect 15910 12484 15966 12540
rect 15966 12484 15970 12540
rect 15906 12480 15970 12484
rect 15986 12540 16050 12544
rect 15986 12484 15990 12540
rect 15990 12484 16046 12540
rect 16046 12484 16050 12540
rect 15986 12480 16050 12484
rect 16988 12412 17052 12476
rect 17724 12412 17788 12476
rect 20116 12472 20180 12476
rect 20116 12416 20130 12472
rect 20130 12416 20180 12472
rect 18644 12276 18708 12340
rect 19196 12276 19260 12340
rect 20116 12412 20180 12416
rect 20668 12472 20732 12476
rect 20668 12416 20682 12472
rect 20682 12416 20732 12472
rect 20668 12412 20732 12416
rect 4650 11996 4714 12000
rect 4650 11940 4654 11996
rect 4654 11940 4710 11996
rect 4710 11940 4714 11996
rect 4650 11936 4714 11940
rect 4730 11996 4794 12000
rect 4730 11940 4734 11996
rect 4734 11940 4790 11996
rect 4790 11940 4794 11996
rect 4730 11936 4794 11940
rect 4810 11996 4874 12000
rect 4810 11940 4814 11996
rect 4814 11940 4870 11996
rect 4870 11940 4874 11996
rect 4810 11936 4874 11940
rect 4890 11996 4954 12000
rect 4890 11940 4894 11996
rect 4894 11940 4950 11996
rect 4950 11940 4954 11996
rect 4890 11936 4954 11940
rect 12048 11996 12112 12000
rect 12048 11940 12052 11996
rect 12052 11940 12108 11996
rect 12108 11940 12112 11996
rect 12048 11936 12112 11940
rect 12128 11996 12192 12000
rect 12128 11940 12132 11996
rect 12132 11940 12188 11996
rect 12188 11940 12192 11996
rect 12128 11936 12192 11940
rect 12208 11996 12272 12000
rect 12208 11940 12212 11996
rect 12212 11940 12268 11996
rect 12268 11940 12272 11996
rect 12208 11936 12272 11940
rect 12288 11996 12352 12000
rect 12288 11940 12292 11996
rect 12292 11940 12348 11996
rect 12348 11940 12352 11996
rect 12288 11936 12352 11940
rect 19445 11996 19509 12000
rect 19445 11940 19449 11996
rect 19449 11940 19505 11996
rect 19505 11940 19509 11996
rect 19445 11936 19509 11940
rect 19525 11996 19589 12000
rect 19525 11940 19529 11996
rect 19529 11940 19585 11996
rect 19585 11940 19589 11996
rect 19525 11936 19589 11940
rect 19605 11996 19669 12000
rect 19605 11940 19609 11996
rect 19609 11940 19665 11996
rect 19665 11940 19669 11996
rect 19605 11936 19669 11940
rect 19685 11996 19749 12000
rect 19685 11940 19689 11996
rect 19689 11940 19745 11996
rect 19745 11940 19749 11996
rect 19685 11936 19749 11940
rect 20116 11868 20180 11932
rect 8349 11452 8413 11456
rect 8349 11396 8353 11452
rect 8353 11396 8409 11452
rect 8409 11396 8413 11452
rect 8349 11392 8413 11396
rect 8429 11452 8493 11456
rect 8429 11396 8433 11452
rect 8433 11396 8489 11452
rect 8489 11396 8493 11452
rect 8429 11392 8493 11396
rect 8509 11452 8573 11456
rect 8509 11396 8513 11452
rect 8513 11396 8569 11452
rect 8569 11396 8573 11452
rect 8509 11392 8573 11396
rect 8589 11452 8653 11456
rect 8589 11396 8593 11452
rect 8593 11396 8649 11452
rect 8649 11396 8653 11452
rect 8589 11392 8653 11396
rect 15746 11452 15810 11456
rect 15746 11396 15750 11452
rect 15750 11396 15806 11452
rect 15806 11396 15810 11452
rect 15746 11392 15810 11396
rect 15826 11452 15890 11456
rect 15826 11396 15830 11452
rect 15830 11396 15886 11452
rect 15886 11396 15890 11452
rect 15826 11392 15890 11396
rect 15906 11452 15970 11456
rect 15906 11396 15910 11452
rect 15910 11396 15966 11452
rect 15966 11396 15970 11452
rect 15906 11392 15970 11396
rect 15986 11452 16050 11456
rect 15986 11396 15990 11452
rect 15990 11396 16046 11452
rect 16046 11396 16050 11452
rect 15986 11392 16050 11396
rect 9812 10976 9876 10980
rect 9812 10920 9862 10976
rect 9862 10920 9876 10976
rect 9812 10916 9876 10920
rect 4650 10908 4714 10912
rect 4650 10852 4654 10908
rect 4654 10852 4710 10908
rect 4710 10852 4714 10908
rect 4650 10848 4714 10852
rect 4730 10908 4794 10912
rect 4730 10852 4734 10908
rect 4734 10852 4790 10908
rect 4790 10852 4794 10908
rect 4730 10848 4794 10852
rect 4810 10908 4874 10912
rect 4810 10852 4814 10908
rect 4814 10852 4870 10908
rect 4870 10852 4874 10908
rect 4810 10848 4874 10852
rect 4890 10908 4954 10912
rect 4890 10852 4894 10908
rect 4894 10852 4950 10908
rect 4950 10852 4954 10908
rect 4890 10848 4954 10852
rect 12048 10908 12112 10912
rect 12048 10852 12052 10908
rect 12052 10852 12108 10908
rect 12108 10852 12112 10908
rect 12048 10848 12112 10852
rect 12128 10908 12192 10912
rect 12128 10852 12132 10908
rect 12132 10852 12188 10908
rect 12188 10852 12192 10908
rect 12128 10848 12192 10852
rect 12208 10908 12272 10912
rect 12208 10852 12212 10908
rect 12212 10852 12268 10908
rect 12268 10852 12272 10908
rect 12208 10848 12272 10852
rect 12288 10908 12352 10912
rect 12288 10852 12292 10908
rect 12292 10852 12348 10908
rect 12348 10852 12352 10908
rect 12288 10848 12352 10852
rect 19445 10908 19509 10912
rect 19445 10852 19449 10908
rect 19449 10852 19505 10908
rect 19505 10852 19509 10908
rect 19445 10848 19509 10852
rect 19525 10908 19589 10912
rect 19525 10852 19529 10908
rect 19529 10852 19585 10908
rect 19585 10852 19589 10908
rect 19525 10848 19589 10852
rect 19605 10908 19669 10912
rect 19605 10852 19609 10908
rect 19609 10852 19665 10908
rect 19665 10852 19669 10908
rect 19605 10848 19669 10852
rect 19685 10908 19749 10912
rect 19685 10852 19689 10908
rect 19689 10852 19745 10908
rect 19745 10852 19749 10908
rect 19685 10848 19749 10852
rect 9628 10704 9692 10708
rect 9628 10648 9678 10704
rect 9678 10648 9692 10704
rect 9628 10644 9692 10648
rect 16988 10644 17052 10708
rect 8349 10364 8413 10368
rect 8349 10308 8353 10364
rect 8353 10308 8409 10364
rect 8409 10308 8413 10364
rect 8349 10304 8413 10308
rect 8429 10364 8493 10368
rect 8429 10308 8433 10364
rect 8433 10308 8489 10364
rect 8489 10308 8493 10364
rect 8429 10304 8493 10308
rect 8509 10364 8573 10368
rect 8509 10308 8513 10364
rect 8513 10308 8569 10364
rect 8569 10308 8573 10364
rect 8509 10304 8573 10308
rect 8589 10364 8653 10368
rect 8589 10308 8593 10364
rect 8593 10308 8649 10364
rect 8649 10308 8653 10364
rect 8589 10304 8653 10308
rect 15746 10364 15810 10368
rect 15746 10308 15750 10364
rect 15750 10308 15806 10364
rect 15806 10308 15810 10364
rect 15746 10304 15810 10308
rect 15826 10364 15890 10368
rect 15826 10308 15830 10364
rect 15830 10308 15886 10364
rect 15886 10308 15890 10364
rect 15826 10304 15890 10308
rect 15906 10364 15970 10368
rect 15906 10308 15910 10364
rect 15910 10308 15966 10364
rect 15966 10308 15970 10364
rect 15906 10304 15970 10308
rect 15986 10364 16050 10368
rect 15986 10308 15990 10364
rect 15990 10308 16046 10364
rect 16046 10308 16050 10364
rect 15986 10304 16050 10308
rect 16252 9964 16316 10028
rect 9812 9888 9876 9892
rect 9812 9832 9862 9888
rect 9862 9832 9876 9888
rect 9812 9828 9876 9832
rect 14228 9888 14292 9892
rect 14228 9832 14242 9888
rect 14242 9832 14292 9888
rect 14228 9828 14292 9832
rect 18092 9828 18156 9892
rect 4650 9820 4714 9824
rect 4650 9764 4654 9820
rect 4654 9764 4710 9820
rect 4710 9764 4714 9820
rect 4650 9760 4714 9764
rect 4730 9820 4794 9824
rect 4730 9764 4734 9820
rect 4734 9764 4790 9820
rect 4790 9764 4794 9820
rect 4730 9760 4794 9764
rect 4810 9820 4874 9824
rect 4810 9764 4814 9820
rect 4814 9764 4870 9820
rect 4870 9764 4874 9820
rect 4810 9760 4874 9764
rect 4890 9820 4954 9824
rect 4890 9764 4894 9820
rect 4894 9764 4950 9820
rect 4950 9764 4954 9820
rect 4890 9760 4954 9764
rect 12048 9820 12112 9824
rect 12048 9764 12052 9820
rect 12052 9764 12108 9820
rect 12108 9764 12112 9820
rect 12048 9760 12112 9764
rect 12128 9820 12192 9824
rect 12128 9764 12132 9820
rect 12132 9764 12188 9820
rect 12188 9764 12192 9820
rect 12128 9760 12192 9764
rect 12208 9820 12272 9824
rect 12208 9764 12212 9820
rect 12212 9764 12268 9820
rect 12268 9764 12272 9820
rect 12208 9760 12272 9764
rect 12288 9820 12352 9824
rect 12288 9764 12292 9820
rect 12292 9764 12348 9820
rect 12348 9764 12352 9820
rect 12288 9760 12352 9764
rect 19445 9820 19509 9824
rect 19445 9764 19449 9820
rect 19449 9764 19505 9820
rect 19505 9764 19509 9820
rect 19445 9760 19509 9764
rect 19525 9820 19589 9824
rect 19525 9764 19529 9820
rect 19529 9764 19585 9820
rect 19585 9764 19589 9820
rect 19525 9760 19589 9764
rect 19605 9820 19669 9824
rect 19605 9764 19609 9820
rect 19609 9764 19665 9820
rect 19665 9764 19669 9820
rect 19605 9760 19669 9764
rect 19685 9820 19749 9824
rect 19685 9764 19689 9820
rect 19689 9764 19745 9820
rect 19745 9764 19749 9820
rect 19685 9760 19749 9764
rect 9628 9752 9692 9756
rect 9628 9696 9678 9752
rect 9678 9696 9692 9752
rect 9628 9692 9692 9696
rect 16620 9692 16684 9756
rect 8349 9276 8413 9280
rect 8349 9220 8353 9276
rect 8353 9220 8409 9276
rect 8409 9220 8413 9276
rect 8349 9216 8413 9220
rect 8429 9276 8493 9280
rect 8429 9220 8433 9276
rect 8433 9220 8489 9276
rect 8489 9220 8493 9276
rect 8429 9216 8493 9220
rect 8509 9276 8573 9280
rect 8509 9220 8513 9276
rect 8513 9220 8569 9276
rect 8569 9220 8573 9276
rect 8509 9216 8573 9220
rect 8589 9276 8653 9280
rect 8589 9220 8593 9276
rect 8593 9220 8649 9276
rect 8649 9220 8653 9276
rect 8589 9216 8653 9220
rect 15746 9276 15810 9280
rect 15746 9220 15750 9276
rect 15750 9220 15806 9276
rect 15806 9220 15810 9276
rect 15746 9216 15810 9220
rect 15826 9276 15890 9280
rect 15826 9220 15830 9276
rect 15830 9220 15886 9276
rect 15886 9220 15890 9276
rect 15826 9216 15890 9220
rect 15906 9276 15970 9280
rect 15906 9220 15910 9276
rect 15910 9220 15966 9276
rect 15966 9220 15970 9276
rect 15906 9216 15970 9220
rect 15986 9276 16050 9280
rect 15986 9220 15990 9276
rect 15990 9220 16046 9276
rect 16046 9220 16050 9276
rect 15986 9216 16050 9220
rect 20484 9148 20548 9212
rect 20300 9012 20364 9076
rect 17172 8876 17236 8940
rect 4650 8732 4714 8736
rect 4650 8676 4654 8732
rect 4654 8676 4710 8732
rect 4710 8676 4714 8732
rect 4650 8672 4714 8676
rect 4730 8732 4794 8736
rect 4730 8676 4734 8732
rect 4734 8676 4790 8732
rect 4790 8676 4794 8732
rect 4730 8672 4794 8676
rect 4810 8732 4874 8736
rect 4810 8676 4814 8732
rect 4814 8676 4870 8732
rect 4870 8676 4874 8732
rect 4810 8672 4874 8676
rect 4890 8732 4954 8736
rect 4890 8676 4894 8732
rect 4894 8676 4950 8732
rect 4950 8676 4954 8732
rect 4890 8672 4954 8676
rect 12048 8732 12112 8736
rect 12048 8676 12052 8732
rect 12052 8676 12108 8732
rect 12108 8676 12112 8732
rect 12048 8672 12112 8676
rect 12128 8732 12192 8736
rect 12128 8676 12132 8732
rect 12132 8676 12188 8732
rect 12188 8676 12192 8732
rect 12128 8672 12192 8676
rect 12208 8732 12272 8736
rect 12208 8676 12212 8732
rect 12212 8676 12268 8732
rect 12268 8676 12272 8732
rect 12208 8672 12272 8676
rect 12288 8732 12352 8736
rect 12288 8676 12292 8732
rect 12292 8676 12348 8732
rect 12348 8676 12352 8732
rect 12288 8672 12352 8676
rect 19445 8732 19509 8736
rect 19445 8676 19449 8732
rect 19449 8676 19505 8732
rect 19505 8676 19509 8732
rect 19445 8672 19509 8676
rect 19525 8732 19589 8736
rect 19525 8676 19529 8732
rect 19529 8676 19585 8732
rect 19585 8676 19589 8732
rect 19525 8672 19589 8676
rect 19605 8732 19669 8736
rect 19605 8676 19609 8732
rect 19609 8676 19665 8732
rect 19665 8676 19669 8732
rect 19605 8672 19669 8676
rect 19685 8732 19749 8736
rect 19685 8676 19689 8732
rect 19689 8676 19745 8732
rect 19745 8676 19749 8732
rect 19685 8672 19749 8676
rect 19932 8604 19996 8668
rect 17172 8468 17236 8532
rect 20116 8332 20180 8396
rect 8349 8188 8413 8192
rect 8349 8132 8353 8188
rect 8353 8132 8409 8188
rect 8409 8132 8413 8188
rect 8349 8128 8413 8132
rect 8429 8188 8493 8192
rect 8429 8132 8433 8188
rect 8433 8132 8489 8188
rect 8489 8132 8493 8188
rect 8429 8128 8493 8132
rect 8509 8188 8573 8192
rect 8509 8132 8513 8188
rect 8513 8132 8569 8188
rect 8569 8132 8573 8188
rect 8509 8128 8573 8132
rect 8589 8188 8653 8192
rect 8589 8132 8593 8188
rect 8593 8132 8649 8188
rect 8649 8132 8653 8188
rect 8589 8128 8653 8132
rect 15746 8188 15810 8192
rect 15746 8132 15750 8188
rect 15750 8132 15806 8188
rect 15806 8132 15810 8188
rect 15746 8128 15810 8132
rect 15826 8188 15890 8192
rect 15826 8132 15830 8188
rect 15830 8132 15886 8188
rect 15886 8132 15890 8188
rect 15826 8128 15890 8132
rect 15906 8188 15970 8192
rect 15906 8132 15910 8188
rect 15910 8132 15966 8188
rect 15966 8132 15970 8188
rect 15906 8128 15970 8132
rect 15986 8188 16050 8192
rect 15986 8132 15990 8188
rect 15990 8132 16046 8188
rect 16046 8132 16050 8188
rect 15986 8128 16050 8132
rect 20484 8060 20548 8124
rect 17724 7652 17788 7716
rect 4650 7644 4714 7648
rect 4650 7588 4654 7644
rect 4654 7588 4710 7644
rect 4710 7588 4714 7644
rect 4650 7584 4714 7588
rect 4730 7644 4794 7648
rect 4730 7588 4734 7644
rect 4734 7588 4790 7644
rect 4790 7588 4794 7644
rect 4730 7584 4794 7588
rect 4810 7644 4874 7648
rect 4810 7588 4814 7644
rect 4814 7588 4870 7644
rect 4870 7588 4874 7644
rect 4810 7584 4874 7588
rect 4890 7644 4954 7648
rect 4890 7588 4894 7644
rect 4894 7588 4950 7644
rect 4950 7588 4954 7644
rect 4890 7584 4954 7588
rect 12048 7644 12112 7648
rect 12048 7588 12052 7644
rect 12052 7588 12108 7644
rect 12108 7588 12112 7644
rect 12048 7584 12112 7588
rect 12128 7644 12192 7648
rect 12128 7588 12132 7644
rect 12132 7588 12188 7644
rect 12188 7588 12192 7644
rect 12128 7584 12192 7588
rect 12208 7644 12272 7648
rect 12208 7588 12212 7644
rect 12212 7588 12268 7644
rect 12268 7588 12272 7644
rect 12208 7584 12272 7588
rect 12288 7644 12352 7648
rect 12288 7588 12292 7644
rect 12292 7588 12348 7644
rect 12348 7588 12352 7644
rect 12288 7584 12352 7588
rect 19445 7644 19509 7648
rect 19445 7588 19449 7644
rect 19449 7588 19505 7644
rect 19505 7588 19509 7644
rect 19445 7584 19509 7588
rect 19525 7644 19589 7648
rect 19525 7588 19529 7644
rect 19529 7588 19585 7644
rect 19585 7588 19589 7644
rect 19525 7584 19589 7588
rect 19605 7644 19669 7648
rect 19605 7588 19609 7644
rect 19609 7588 19665 7644
rect 19665 7588 19669 7644
rect 19605 7584 19669 7588
rect 19685 7644 19749 7648
rect 19685 7588 19689 7644
rect 19689 7588 19745 7644
rect 19745 7588 19749 7644
rect 19685 7584 19749 7588
rect 17724 7380 17788 7444
rect 19012 7108 19076 7172
rect 8349 7100 8413 7104
rect 8349 7044 8353 7100
rect 8353 7044 8409 7100
rect 8409 7044 8413 7100
rect 8349 7040 8413 7044
rect 8429 7100 8493 7104
rect 8429 7044 8433 7100
rect 8433 7044 8489 7100
rect 8489 7044 8493 7100
rect 8429 7040 8493 7044
rect 8509 7100 8573 7104
rect 8509 7044 8513 7100
rect 8513 7044 8569 7100
rect 8569 7044 8573 7100
rect 8509 7040 8573 7044
rect 8589 7100 8653 7104
rect 8589 7044 8593 7100
rect 8593 7044 8649 7100
rect 8649 7044 8653 7100
rect 8589 7040 8653 7044
rect 15746 7100 15810 7104
rect 15746 7044 15750 7100
rect 15750 7044 15806 7100
rect 15806 7044 15810 7100
rect 15746 7040 15810 7044
rect 15826 7100 15890 7104
rect 15826 7044 15830 7100
rect 15830 7044 15886 7100
rect 15886 7044 15890 7100
rect 15826 7040 15890 7044
rect 15906 7100 15970 7104
rect 15906 7044 15910 7100
rect 15910 7044 15966 7100
rect 15966 7044 15970 7100
rect 15906 7040 15970 7044
rect 15986 7100 16050 7104
rect 15986 7044 15990 7100
rect 15990 7044 16046 7100
rect 16046 7044 16050 7100
rect 15986 7040 16050 7044
rect 4650 6556 4714 6560
rect 4650 6500 4654 6556
rect 4654 6500 4710 6556
rect 4710 6500 4714 6556
rect 4650 6496 4714 6500
rect 4730 6556 4794 6560
rect 4730 6500 4734 6556
rect 4734 6500 4790 6556
rect 4790 6500 4794 6556
rect 4730 6496 4794 6500
rect 4810 6556 4874 6560
rect 4810 6500 4814 6556
rect 4814 6500 4870 6556
rect 4870 6500 4874 6556
rect 4810 6496 4874 6500
rect 4890 6556 4954 6560
rect 4890 6500 4894 6556
rect 4894 6500 4950 6556
rect 4950 6500 4954 6556
rect 4890 6496 4954 6500
rect 12048 6556 12112 6560
rect 12048 6500 12052 6556
rect 12052 6500 12108 6556
rect 12108 6500 12112 6556
rect 12048 6496 12112 6500
rect 12128 6556 12192 6560
rect 12128 6500 12132 6556
rect 12132 6500 12188 6556
rect 12188 6500 12192 6556
rect 12128 6496 12192 6500
rect 12208 6556 12272 6560
rect 12208 6500 12212 6556
rect 12212 6500 12268 6556
rect 12268 6500 12272 6556
rect 12208 6496 12272 6500
rect 12288 6556 12352 6560
rect 12288 6500 12292 6556
rect 12292 6500 12348 6556
rect 12348 6500 12352 6556
rect 12288 6496 12352 6500
rect 19445 6556 19509 6560
rect 19445 6500 19449 6556
rect 19449 6500 19505 6556
rect 19505 6500 19509 6556
rect 19445 6496 19509 6500
rect 19525 6556 19589 6560
rect 19525 6500 19529 6556
rect 19529 6500 19585 6556
rect 19585 6500 19589 6556
rect 19525 6496 19589 6500
rect 19605 6556 19669 6560
rect 19605 6500 19609 6556
rect 19609 6500 19665 6556
rect 19665 6500 19669 6556
rect 19605 6496 19669 6500
rect 19685 6556 19749 6560
rect 19685 6500 19689 6556
rect 19689 6500 19745 6556
rect 19745 6500 19749 6556
rect 19685 6496 19749 6500
rect 19932 6352 19996 6356
rect 19932 6296 19946 6352
rect 19946 6296 19996 6352
rect 19932 6292 19996 6296
rect 8349 6012 8413 6016
rect 8349 5956 8353 6012
rect 8353 5956 8409 6012
rect 8409 5956 8413 6012
rect 8349 5952 8413 5956
rect 8429 6012 8493 6016
rect 8429 5956 8433 6012
rect 8433 5956 8489 6012
rect 8489 5956 8493 6012
rect 8429 5952 8493 5956
rect 8509 6012 8573 6016
rect 8509 5956 8513 6012
rect 8513 5956 8569 6012
rect 8569 5956 8573 6012
rect 8509 5952 8573 5956
rect 8589 6012 8653 6016
rect 8589 5956 8593 6012
rect 8593 5956 8649 6012
rect 8649 5956 8653 6012
rect 8589 5952 8653 5956
rect 15746 6012 15810 6016
rect 15746 5956 15750 6012
rect 15750 5956 15806 6012
rect 15806 5956 15810 6012
rect 15746 5952 15810 5956
rect 15826 6012 15890 6016
rect 15826 5956 15830 6012
rect 15830 5956 15886 6012
rect 15886 5956 15890 6012
rect 15826 5952 15890 5956
rect 15906 6012 15970 6016
rect 15906 5956 15910 6012
rect 15910 5956 15966 6012
rect 15966 5956 15970 6012
rect 15906 5952 15970 5956
rect 15986 6012 16050 6016
rect 15986 5956 15990 6012
rect 15990 5956 16046 6012
rect 16046 5956 16050 6012
rect 15986 5952 16050 5956
rect 4650 5468 4714 5472
rect 4650 5412 4654 5468
rect 4654 5412 4710 5468
rect 4710 5412 4714 5468
rect 4650 5408 4714 5412
rect 4730 5468 4794 5472
rect 4730 5412 4734 5468
rect 4734 5412 4790 5468
rect 4790 5412 4794 5468
rect 4730 5408 4794 5412
rect 4810 5468 4874 5472
rect 4810 5412 4814 5468
rect 4814 5412 4870 5468
rect 4870 5412 4874 5468
rect 4810 5408 4874 5412
rect 4890 5468 4954 5472
rect 4890 5412 4894 5468
rect 4894 5412 4950 5468
rect 4950 5412 4954 5468
rect 4890 5408 4954 5412
rect 12048 5468 12112 5472
rect 12048 5412 12052 5468
rect 12052 5412 12108 5468
rect 12108 5412 12112 5468
rect 12048 5408 12112 5412
rect 12128 5468 12192 5472
rect 12128 5412 12132 5468
rect 12132 5412 12188 5468
rect 12188 5412 12192 5468
rect 12128 5408 12192 5412
rect 12208 5468 12272 5472
rect 12208 5412 12212 5468
rect 12212 5412 12268 5468
rect 12268 5412 12272 5468
rect 12208 5408 12272 5412
rect 12288 5468 12352 5472
rect 12288 5412 12292 5468
rect 12292 5412 12348 5468
rect 12348 5412 12352 5468
rect 12288 5408 12352 5412
rect 19445 5468 19509 5472
rect 19445 5412 19449 5468
rect 19449 5412 19505 5468
rect 19505 5412 19509 5468
rect 19445 5408 19509 5412
rect 19525 5468 19589 5472
rect 19525 5412 19529 5468
rect 19529 5412 19585 5468
rect 19585 5412 19589 5468
rect 19525 5408 19589 5412
rect 19605 5468 19669 5472
rect 19605 5412 19609 5468
rect 19609 5412 19665 5468
rect 19665 5412 19669 5468
rect 19605 5408 19669 5412
rect 19685 5468 19749 5472
rect 19685 5412 19689 5468
rect 19689 5412 19745 5468
rect 19745 5412 19749 5468
rect 19685 5408 19749 5412
rect 8349 4924 8413 4928
rect 8349 4868 8353 4924
rect 8353 4868 8409 4924
rect 8409 4868 8413 4924
rect 8349 4864 8413 4868
rect 8429 4924 8493 4928
rect 8429 4868 8433 4924
rect 8433 4868 8489 4924
rect 8489 4868 8493 4924
rect 8429 4864 8493 4868
rect 8509 4924 8573 4928
rect 8509 4868 8513 4924
rect 8513 4868 8569 4924
rect 8569 4868 8573 4924
rect 8509 4864 8573 4868
rect 8589 4924 8653 4928
rect 8589 4868 8593 4924
rect 8593 4868 8649 4924
rect 8649 4868 8653 4924
rect 8589 4864 8653 4868
rect 15746 4924 15810 4928
rect 15746 4868 15750 4924
rect 15750 4868 15806 4924
rect 15806 4868 15810 4924
rect 15746 4864 15810 4868
rect 15826 4924 15890 4928
rect 15826 4868 15830 4924
rect 15830 4868 15886 4924
rect 15886 4868 15890 4924
rect 15826 4864 15890 4868
rect 15906 4924 15970 4928
rect 15906 4868 15910 4924
rect 15910 4868 15966 4924
rect 15966 4868 15970 4924
rect 15906 4864 15970 4868
rect 15986 4924 16050 4928
rect 15986 4868 15990 4924
rect 15990 4868 16046 4924
rect 16046 4868 16050 4924
rect 15986 4864 16050 4868
rect 16988 4524 17052 4588
rect 4650 4380 4714 4384
rect 4650 4324 4654 4380
rect 4654 4324 4710 4380
rect 4710 4324 4714 4380
rect 4650 4320 4714 4324
rect 4730 4380 4794 4384
rect 4730 4324 4734 4380
rect 4734 4324 4790 4380
rect 4790 4324 4794 4380
rect 4730 4320 4794 4324
rect 4810 4380 4874 4384
rect 4810 4324 4814 4380
rect 4814 4324 4870 4380
rect 4870 4324 4874 4380
rect 4810 4320 4874 4324
rect 4890 4380 4954 4384
rect 4890 4324 4894 4380
rect 4894 4324 4950 4380
rect 4950 4324 4954 4380
rect 4890 4320 4954 4324
rect 12048 4380 12112 4384
rect 12048 4324 12052 4380
rect 12052 4324 12108 4380
rect 12108 4324 12112 4380
rect 12048 4320 12112 4324
rect 12128 4380 12192 4384
rect 12128 4324 12132 4380
rect 12132 4324 12188 4380
rect 12188 4324 12192 4380
rect 12128 4320 12192 4324
rect 12208 4380 12272 4384
rect 12208 4324 12212 4380
rect 12212 4324 12268 4380
rect 12268 4324 12272 4380
rect 12208 4320 12272 4324
rect 12288 4380 12352 4384
rect 12288 4324 12292 4380
rect 12292 4324 12348 4380
rect 12348 4324 12352 4380
rect 12288 4320 12352 4324
rect 19445 4380 19509 4384
rect 19445 4324 19449 4380
rect 19449 4324 19505 4380
rect 19505 4324 19509 4380
rect 19445 4320 19509 4324
rect 19525 4380 19589 4384
rect 19525 4324 19529 4380
rect 19529 4324 19585 4380
rect 19585 4324 19589 4380
rect 19525 4320 19589 4324
rect 19605 4380 19669 4384
rect 19605 4324 19609 4380
rect 19609 4324 19665 4380
rect 19665 4324 19669 4380
rect 19605 4320 19669 4324
rect 19685 4380 19749 4384
rect 19685 4324 19689 4380
rect 19689 4324 19745 4380
rect 19745 4324 19749 4380
rect 19685 4320 19749 4324
rect 13308 3980 13372 4044
rect 21404 3980 21468 4044
rect 8349 3836 8413 3840
rect 8349 3780 8353 3836
rect 8353 3780 8409 3836
rect 8409 3780 8413 3836
rect 8349 3776 8413 3780
rect 8429 3836 8493 3840
rect 8429 3780 8433 3836
rect 8433 3780 8489 3836
rect 8489 3780 8493 3836
rect 8429 3776 8493 3780
rect 8509 3836 8573 3840
rect 8509 3780 8513 3836
rect 8513 3780 8569 3836
rect 8569 3780 8573 3836
rect 8509 3776 8573 3780
rect 8589 3836 8653 3840
rect 8589 3780 8593 3836
rect 8593 3780 8649 3836
rect 8649 3780 8653 3836
rect 8589 3776 8653 3780
rect 15746 3836 15810 3840
rect 15746 3780 15750 3836
rect 15750 3780 15806 3836
rect 15806 3780 15810 3836
rect 15746 3776 15810 3780
rect 15826 3836 15890 3840
rect 15826 3780 15830 3836
rect 15830 3780 15886 3836
rect 15886 3780 15890 3836
rect 15826 3776 15890 3780
rect 15906 3836 15970 3840
rect 15906 3780 15910 3836
rect 15910 3780 15966 3836
rect 15966 3780 15970 3836
rect 15906 3776 15970 3780
rect 15986 3836 16050 3840
rect 15986 3780 15990 3836
rect 15990 3780 16046 3836
rect 16046 3780 16050 3836
rect 15986 3776 16050 3780
rect 19932 3572 19996 3636
rect 4650 3292 4714 3296
rect 4650 3236 4654 3292
rect 4654 3236 4710 3292
rect 4710 3236 4714 3292
rect 4650 3232 4714 3236
rect 4730 3292 4794 3296
rect 4730 3236 4734 3292
rect 4734 3236 4790 3292
rect 4790 3236 4794 3292
rect 4730 3232 4794 3236
rect 4810 3292 4874 3296
rect 4810 3236 4814 3292
rect 4814 3236 4870 3292
rect 4870 3236 4874 3292
rect 4810 3232 4874 3236
rect 4890 3292 4954 3296
rect 4890 3236 4894 3292
rect 4894 3236 4950 3292
rect 4950 3236 4954 3292
rect 4890 3232 4954 3236
rect 12048 3292 12112 3296
rect 12048 3236 12052 3292
rect 12052 3236 12108 3292
rect 12108 3236 12112 3292
rect 12048 3232 12112 3236
rect 12128 3292 12192 3296
rect 12128 3236 12132 3292
rect 12132 3236 12188 3292
rect 12188 3236 12192 3292
rect 12128 3232 12192 3236
rect 12208 3292 12272 3296
rect 12208 3236 12212 3292
rect 12212 3236 12268 3292
rect 12268 3236 12272 3292
rect 12208 3232 12272 3236
rect 12288 3292 12352 3296
rect 12288 3236 12292 3292
rect 12292 3236 12348 3292
rect 12348 3236 12352 3292
rect 12288 3232 12352 3236
rect 19445 3292 19509 3296
rect 19445 3236 19449 3292
rect 19449 3236 19505 3292
rect 19505 3236 19509 3292
rect 19445 3232 19509 3236
rect 19525 3292 19589 3296
rect 19525 3236 19529 3292
rect 19529 3236 19585 3292
rect 19585 3236 19589 3292
rect 19525 3232 19589 3236
rect 19605 3292 19669 3296
rect 19605 3236 19609 3292
rect 19609 3236 19665 3292
rect 19665 3236 19669 3292
rect 19605 3232 19669 3236
rect 19685 3292 19749 3296
rect 19685 3236 19689 3292
rect 19689 3236 19745 3292
rect 19745 3236 19749 3292
rect 19685 3232 19749 3236
rect 20300 2892 20364 2956
rect 8349 2748 8413 2752
rect 8349 2692 8353 2748
rect 8353 2692 8409 2748
rect 8409 2692 8413 2748
rect 8349 2688 8413 2692
rect 8429 2748 8493 2752
rect 8429 2692 8433 2748
rect 8433 2692 8489 2748
rect 8489 2692 8493 2748
rect 8429 2688 8493 2692
rect 8509 2748 8573 2752
rect 8509 2692 8513 2748
rect 8513 2692 8569 2748
rect 8569 2692 8573 2748
rect 8509 2688 8573 2692
rect 8589 2748 8653 2752
rect 8589 2692 8593 2748
rect 8593 2692 8649 2748
rect 8649 2692 8653 2748
rect 8589 2688 8653 2692
rect 15746 2748 15810 2752
rect 15746 2692 15750 2748
rect 15750 2692 15806 2748
rect 15806 2692 15810 2748
rect 15746 2688 15810 2692
rect 15826 2748 15890 2752
rect 15826 2692 15830 2748
rect 15830 2692 15886 2748
rect 15886 2692 15890 2748
rect 15826 2688 15890 2692
rect 15906 2748 15970 2752
rect 15906 2692 15910 2748
rect 15910 2692 15966 2748
rect 15966 2692 15970 2748
rect 15906 2688 15970 2692
rect 15986 2748 16050 2752
rect 15986 2692 15990 2748
rect 15990 2692 16046 2748
rect 16046 2692 16050 2748
rect 15986 2688 16050 2692
rect 21588 2484 21652 2548
rect 4650 2204 4714 2208
rect 4650 2148 4654 2204
rect 4654 2148 4710 2204
rect 4710 2148 4714 2204
rect 4650 2144 4714 2148
rect 4730 2204 4794 2208
rect 4730 2148 4734 2204
rect 4734 2148 4790 2204
rect 4790 2148 4794 2204
rect 4730 2144 4794 2148
rect 4810 2204 4874 2208
rect 4810 2148 4814 2204
rect 4814 2148 4870 2204
rect 4870 2148 4874 2204
rect 4810 2144 4874 2148
rect 4890 2204 4954 2208
rect 4890 2148 4894 2204
rect 4894 2148 4950 2204
rect 4950 2148 4954 2204
rect 4890 2144 4954 2148
rect 12048 2204 12112 2208
rect 12048 2148 12052 2204
rect 12052 2148 12108 2204
rect 12108 2148 12112 2204
rect 12048 2144 12112 2148
rect 12128 2204 12192 2208
rect 12128 2148 12132 2204
rect 12132 2148 12188 2204
rect 12188 2148 12192 2204
rect 12128 2144 12192 2148
rect 12208 2204 12272 2208
rect 12208 2148 12212 2204
rect 12212 2148 12268 2204
rect 12268 2148 12272 2204
rect 12208 2144 12272 2148
rect 12288 2204 12352 2208
rect 12288 2148 12292 2204
rect 12292 2148 12348 2204
rect 12348 2148 12352 2204
rect 12288 2144 12352 2148
rect 19445 2204 19509 2208
rect 19445 2148 19449 2204
rect 19449 2148 19505 2204
rect 19505 2148 19509 2204
rect 19445 2144 19509 2148
rect 19525 2204 19589 2208
rect 19525 2148 19529 2204
rect 19529 2148 19585 2204
rect 19585 2148 19589 2204
rect 19525 2144 19589 2148
rect 19605 2204 19669 2208
rect 19605 2148 19609 2204
rect 19609 2148 19665 2204
rect 19665 2148 19669 2204
rect 19605 2144 19669 2148
rect 19685 2204 19749 2208
rect 19685 2148 19689 2204
rect 19689 2148 19745 2204
rect 19745 2148 19749 2204
rect 19685 2144 19749 2148
<< metal4 >>
rect 4642 21792 4963 21808
rect 4642 21728 4650 21792
rect 4714 21728 4730 21792
rect 4794 21728 4810 21792
rect 4874 21728 4890 21792
rect 4954 21728 4963 21792
rect 4642 20704 4963 21728
rect 4642 20640 4650 20704
rect 4714 20640 4730 20704
rect 4794 20640 4810 20704
rect 4874 20640 4890 20704
rect 4954 20640 4963 20704
rect 4642 19616 4963 20640
rect 4642 19552 4650 19616
rect 4714 19552 4730 19616
rect 4794 19552 4810 19616
rect 4874 19552 4890 19616
rect 4954 19552 4963 19616
rect 4642 18528 4963 19552
rect 4642 18464 4650 18528
rect 4714 18464 4730 18528
rect 4794 18464 4810 18528
rect 4874 18464 4890 18528
rect 4954 18464 4963 18528
rect 4642 17440 4963 18464
rect 4642 17376 4650 17440
rect 4714 17376 4730 17440
rect 4794 17376 4810 17440
rect 4874 17376 4890 17440
rect 4954 17376 4963 17440
rect 4642 16352 4963 17376
rect 4642 16288 4650 16352
rect 4714 16288 4730 16352
rect 4794 16288 4810 16352
rect 4874 16288 4890 16352
rect 4954 16288 4963 16352
rect 4642 15264 4963 16288
rect 4642 15200 4650 15264
rect 4714 15200 4730 15264
rect 4794 15200 4810 15264
rect 4874 15200 4890 15264
rect 4954 15200 4963 15264
rect 4642 14176 4963 15200
rect 4642 14112 4650 14176
rect 4714 14112 4730 14176
rect 4794 14112 4810 14176
rect 4874 14112 4890 14176
rect 4954 14112 4963 14176
rect 4642 13088 4963 14112
rect 4642 13024 4650 13088
rect 4714 13024 4730 13088
rect 4794 13024 4810 13088
rect 4874 13024 4890 13088
rect 4954 13024 4963 13088
rect 4642 12000 4963 13024
rect 4642 11936 4650 12000
rect 4714 11936 4730 12000
rect 4794 11936 4810 12000
rect 4874 11936 4890 12000
rect 4954 11936 4963 12000
rect 4642 10912 4963 11936
rect 4642 10848 4650 10912
rect 4714 10848 4730 10912
rect 4794 10848 4810 10912
rect 4874 10848 4890 10912
rect 4954 10848 4963 10912
rect 4642 9824 4963 10848
rect 4642 9760 4650 9824
rect 4714 9760 4730 9824
rect 4794 9760 4810 9824
rect 4874 9760 4890 9824
rect 4954 9760 4963 9824
rect 4642 8736 4963 9760
rect 4642 8672 4650 8736
rect 4714 8672 4730 8736
rect 4794 8672 4810 8736
rect 4874 8672 4890 8736
rect 4954 8672 4963 8736
rect 4642 7648 4963 8672
rect 4642 7584 4650 7648
rect 4714 7584 4730 7648
rect 4794 7584 4810 7648
rect 4874 7584 4890 7648
rect 4954 7584 4963 7648
rect 4642 6560 4963 7584
rect 4642 6496 4650 6560
rect 4714 6496 4730 6560
rect 4794 6496 4810 6560
rect 4874 6496 4890 6560
rect 4954 6496 4963 6560
rect 4642 5472 4963 6496
rect 4642 5408 4650 5472
rect 4714 5408 4730 5472
rect 4794 5408 4810 5472
rect 4874 5408 4890 5472
rect 4954 5408 4963 5472
rect 4642 4384 4963 5408
rect 4642 4320 4650 4384
rect 4714 4320 4730 4384
rect 4794 4320 4810 4384
rect 4874 4320 4890 4384
rect 4954 4320 4963 4384
rect 4642 3296 4963 4320
rect 4642 3232 4650 3296
rect 4714 3232 4730 3296
rect 4794 3232 4810 3296
rect 4874 3232 4890 3296
rect 4954 3232 4963 3296
rect 4642 2208 4963 3232
rect 4642 2144 4650 2208
rect 4714 2144 4730 2208
rect 4794 2144 4810 2208
rect 4874 2144 4890 2208
rect 4954 2144 4963 2208
rect 4642 2128 4963 2144
rect 8341 21248 8661 21808
rect 8341 21184 8349 21248
rect 8413 21184 8429 21248
rect 8493 21184 8509 21248
rect 8573 21184 8589 21248
rect 8653 21184 8661 21248
rect 8341 20160 8661 21184
rect 8341 20096 8349 20160
rect 8413 20096 8429 20160
rect 8493 20096 8509 20160
rect 8573 20096 8589 20160
rect 8653 20096 8661 20160
rect 8341 19072 8661 20096
rect 8341 19008 8349 19072
rect 8413 19008 8429 19072
rect 8493 19008 8509 19072
rect 8573 19008 8589 19072
rect 8653 19008 8661 19072
rect 8341 17984 8661 19008
rect 8341 17920 8349 17984
rect 8413 17920 8429 17984
rect 8493 17920 8509 17984
rect 8573 17920 8589 17984
rect 8653 17920 8661 17984
rect 8341 16896 8661 17920
rect 8341 16832 8349 16896
rect 8413 16832 8429 16896
rect 8493 16832 8509 16896
rect 8573 16832 8589 16896
rect 8653 16832 8661 16896
rect 8341 15808 8661 16832
rect 8341 15744 8349 15808
rect 8413 15744 8429 15808
rect 8493 15744 8509 15808
rect 8573 15744 8589 15808
rect 8653 15744 8661 15808
rect 8341 14720 8661 15744
rect 8341 14656 8349 14720
rect 8413 14656 8429 14720
rect 8493 14656 8509 14720
rect 8573 14656 8589 14720
rect 8653 14656 8661 14720
rect 8341 13632 8661 14656
rect 8341 13568 8349 13632
rect 8413 13568 8429 13632
rect 8493 13568 8509 13632
rect 8573 13568 8589 13632
rect 8653 13568 8661 13632
rect 8341 12544 8661 13568
rect 8341 12480 8349 12544
rect 8413 12480 8429 12544
rect 8493 12480 8509 12544
rect 8573 12480 8589 12544
rect 8653 12480 8661 12544
rect 8341 11456 8661 12480
rect 8341 11392 8349 11456
rect 8413 11392 8429 11456
rect 8493 11392 8509 11456
rect 8573 11392 8589 11456
rect 8653 11392 8661 11456
rect 8341 10368 8661 11392
rect 12040 21792 12360 21808
rect 12040 21728 12048 21792
rect 12112 21728 12128 21792
rect 12192 21728 12208 21792
rect 12272 21728 12288 21792
rect 12352 21728 12360 21792
rect 12040 20704 12360 21728
rect 15738 21248 16058 21808
rect 15738 21184 15746 21248
rect 15810 21184 15826 21248
rect 15890 21184 15906 21248
rect 15970 21184 15986 21248
rect 16050 21184 16058 21248
rect 13123 20908 13189 20909
rect 13123 20844 13124 20908
rect 13188 20844 13189 20908
rect 13123 20843 13189 20844
rect 13307 20908 13373 20909
rect 13307 20844 13308 20908
rect 13372 20844 13373 20908
rect 13307 20843 13373 20844
rect 12040 20640 12048 20704
rect 12112 20640 12128 20704
rect 12192 20640 12208 20704
rect 12272 20640 12288 20704
rect 12352 20640 12360 20704
rect 12040 19616 12360 20640
rect 12040 19552 12048 19616
rect 12112 19552 12128 19616
rect 12192 19552 12208 19616
rect 12272 19552 12288 19616
rect 12352 19552 12360 19616
rect 12040 18528 12360 19552
rect 12040 18464 12048 18528
rect 12112 18464 12128 18528
rect 12192 18464 12208 18528
rect 12272 18464 12288 18528
rect 12352 18464 12360 18528
rect 12040 17440 12360 18464
rect 13126 18053 13186 20843
rect 13123 18052 13189 18053
rect 13123 17988 13124 18052
rect 13188 17988 13189 18052
rect 13123 17987 13189 17988
rect 13123 17508 13189 17509
rect 13123 17444 13124 17508
rect 13188 17444 13189 17508
rect 13123 17443 13189 17444
rect 12040 17376 12048 17440
rect 12112 17376 12128 17440
rect 12192 17376 12208 17440
rect 12272 17376 12288 17440
rect 12352 17376 12360 17440
rect 12040 16352 12360 17376
rect 12040 16288 12048 16352
rect 12112 16288 12128 16352
rect 12192 16288 12208 16352
rect 12272 16288 12288 16352
rect 12352 16288 12360 16352
rect 12040 15264 12360 16288
rect 12040 15200 12048 15264
rect 12112 15200 12128 15264
rect 12192 15200 12208 15264
rect 12272 15200 12288 15264
rect 12352 15200 12360 15264
rect 12040 14176 12360 15200
rect 12040 14112 12048 14176
rect 12112 14112 12128 14176
rect 12192 14112 12208 14176
rect 12272 14112 12288 14176
rect 12352 14112 12360 14176
rect 12040 13088 12360 14112
rect 13126 13565 13186 17443
rect 13123 13564 13189 13565
rect 13123 13500 13124 13564
rect 13188 13500 13189 13564
rect 13123 13499 13189 13500
rect 12040 13024 12048 13088
rect 12112 13024 12128 13088
rect 12192 13024 12208 13088
rect 12272 13024 12288 13088
rect 12352 13024 12360 13088
rect 12040 12000 12360 13024
rect 12040 11936 12048 12000
rect 12112 11936 12128 12000
rect 12192 11936 12208 12000
rect 12272 11936 12288 12000
rect 12352 11936 12360 12000
rect 9811 10980 9877 10981
rect 9811 10916 9812 10980
rect 9876 10916 9877 10980
rect 9811 10915 9877 10916
rect 9627 10708 9693 10709
rect 9627 10644 9628 10708
rect 9692 10644 9693 10708
rect 9627 10643 9693 10644
rect 8341 10304 8349 10368
rect 8413 10304 8429 10368
rect 8493 10304 8509 10368
rect 8573 10304 8589 10368
rect 8653 10304 8661 10368
rect 8341 9280 8661 10304
rect 9630 9757 9690 10643
rect 9814 9893 9874 10915
rect 12040 10912 12360 11936
rect 12040 10848 12048 10912
rect 12112 10848 12128 10912
rect 12192 10848 12208 10912
rect 12272 10848 12288 10912
rect 12352 10848 12360 10912
rect 9811 9892 9877 9893
rect 9811 9828 9812 9892
rect 9876 9828 9877 9892
rect 9811 9827 9877 9828
rect 12040 9824 12360 10848
rect 12040 9760 12048 9824
rect 12112 9760 12128 9824
rect 12192 9760 12208 9824
rect 12272 9760 12288 9824
rect 12352 9760 12360 9824
rect 9627 9756 9693 9757
rect 9627 9692 9628 9756
rect 9692 9692 9693 9756
rect 9627 9691 9693 9692
rect 8341 9216 8349 9280
rect 8413 9216 8429 9280
rect 8493 9216 8509 9280
rect 8573 9216 8589 9280
rect 8653 9216 8661 9280
rect 8341 8192 8661 9216
rect 8341 8128 8349 8192
rect 8413 8128 8429 8192
rect 8493 8128 8509 8192
rect 8573 8128 8589 8192
rect 8653 8128 8661 8192
rect 8341 7104 8661 8128
rect 8341 7040 8349 7104
rect 8413 7040 8429 7104
rect 8493 7040 8509 7104
rect 8573 7040 8589 7104
rect 8653 7040 8661 7104
rect 8341 6016 8661 7040
rect 8341 5952 8349 6016
rect 8413 5952 8429 6016
rect 8493 5952 8509 6016
rect 8573 5952 8589 6016
rect 8653 5952 8661 6016
rect 8341 4928 8661 5952
rect 8341 4864 8349 4928
rect 8413 4864 8429 4928
rect 8493 4864 8509 4928
rect 8573 4864 8589 4928
rect 8653 4864 8661 4928
rect 8341 3840 8661 4864
rect 8341 3776 8349 3840
rect 8413 3776 8429 3840
rect 8493 3776 8509 3840
rect 8573 3776 8589 3840
rect 8653 3776 8661 3840
rect 8341 2752 8661 3776
rect 8341 2688 8349 2752
rect 8413 2688 8429 2752
rect 8493 2688 8509 2752
rect 8573 2688 8589 2752
rect 8653 2688 8661 2752
rect 8341 2128 8661 2688
rect 12040 8736 12360 9760
rect 12040 8672 12048 8736
rect 12112 8672 12128 8736
rect 12192 8672 12208 8736
rect 12272 8672 12288 8736
rect 12352 8672 12360 8736
rect 12040 7648 12360 8672
rect 12040 7584 12048 7648
rect 12112 7584 12128 7648
rect 12192 7584 12208 7648
rect 12272 7584 12288 7648
rect 12352 7584 12360 7648
rect 12040 6560 12360 7584
rect 12040 6496 12048 6560
rect 12112 6496 12128 6560
rect 12192 6496 12208 6560
rect 12272 6496 12288 6560
rect 12352 6496 12360 6560
rect 12040 5472 12360 6496
rect 12040 5408 12048 5472
rect 12112 5408 12128 5472
rect 12192 5408 12208 5472
rect 12272 5408 12288 5472
rect 12352 5408 12360 5472
rect 12040 4384 12360 5408
rect 12040 4320 12048 4384
rect 12112 4320 12128 4384
rect 12192 4320 12208 4384
rect 12272 4320 12288 4384
rect 12352 4320 12360 4384
rect 12040 3296 12360 4320
rect 13310 4045 13370 20843
rect 15738 20160 16058 21184
rect 15738 20096 15746 20160
rect 15810 20096 15826 20160
rect 15890 20096 15906 20160
rect 15970 20096 15986 20160
rect 16050 20096 16058 20160
rect 13491 19276 13557 19277
rect 13491 19212 13492 19276
rect 13556 19212 13557 19276
rect 13491 19211 13557 19212
rect 13494 14109 13554 19211
rect 15738 19072 16058 20096
rect 15738 19008 15746 19072
rect 15810 19008 15826 19072
rect 15890 19008 15906 19072
rect 15970 19008 15986 19072
rect 16050 19008 16058 19072
rect 14227 18188 14293 18189
rect 14227 18124 14228 18188
rect 14292 18124 14293 18188
rect 14227 18123 14293 18124
rect 13491 14108 13557 14109
rect 13491 14044 13492 14108
rect 13556 14044 13557 14108
rect 13491 14043 13557 14044
rect 14230 9893 14290 18123
rect 15738 17984 16058 19008
rect 19437 21792 19757 21808
rect 19437 21728 19445 21792
rect 19509 21728 19525 21792
rect 19589 21728 19605 21792
rect 19669 21728 19685 21792
rect 19749 21728 19757 21792
rect 19437 20704 19757 21728
rect 19437 20640 19445 20704
rect 19509 20640 19525 20704
rect 19589 20640 19605 20704
rect 19669 20640 19685 20704
rect 19749 20640 19757 20704
rect 19437 19616 19757 20640
rect 20667 19956 20733 19957
rect 20667 19892 20668 19956
rect 20732 19892 20733 19956
rect 20667 19891 20733 19892
rect 19437 19552 19445 19616
rect 19509 19552 19525 19616
rect 19589 19552 19605 19616
rect 19669 19552 19685 19616
rect 19749 19552 19757 19616
rect 16987 18732 17053 18733
rect 16987 18668 16988 18732
rect 17052 18668 17053 18732
rect 16987 18667 17053 18668
rect 19011 18732 19077 18733
rect 19011 18668 19012 18732
rect 19076 18668 19077 18732
rect 19011 18667 19077 18668
rect 15738 17920 15746 17984
rect 15810 17920 15826 17984
rect 15890 17920 15906 17984
rect 15970 17920 15986 17984
rect 16050 17920 16058 17984
rect 15738 16896 16058 17920
rect 16435 17644 16501 17645
rect 16435 17580 16436 17644
rect 16500 17580 16501 17644
rect 16435 17579 16501 17580
rect 15738 16832 15746 16896
rect 15810 16832 15826 16896
rect 15890 16832 15906 16896
rect 15970 16832 15986 16896
rect 16050 16832 16058 16896
rect 15738 15808 16058 16832
rect 15738 15744 15746 15808
rect 15810 15744 15826 15808
rect 15890 15744 15906 15808
rect 15970 15744 15986 15808
rect 16050 15744 16058 15808
rect 15738 14720 16058 15744
rect 15738 14656 15746 14720
rect 15810 14656 15826 14720
rect 15890 14656 15906 14720
rect 15970 14656 15986 14720
rect 16050 14656 16058 14720
rect 15738 13632 16058 14656
rect 16251 14652 16317 14653
rect 16251 14588 16252 14652
rect 16316 14588 16317 14652
rect 16251 14587 16317 14588
rect 15738 13568 15746 13632
rect 15810 13568 15826 13632
rect 15890 13568 15906 13632
rect 15970 13568 15986 13632
rect 16050 13568 16058 13632
rect 15738 12544 16058 13568
rect 15738 12480 15746 12544
rect 15810 12480 15826 12544
rect 15890 12480 15906 12544
rect 15970 12480 15986 12544
rect 16050 12480 16058 12544
rect 15738 11456 16058 12480
rect 15738 11392 15746 11456
rect 15810 11392 15826 11456
rect 15890 11392 15906 11456
rect 15970 11392 15986 11456
rect 16050 11392 16058 11456
rect 15738 10368 16058 11392
rect 15738 10304 15746 10368
rect 15810 10304 15826 10368
rect 15890 10304 15906 10368
rect 15970 10304 15986 10368
rect 16050 10304 16058 10368
rect 14227 9892 14293 9893
rect 14227 9828 14228 9892
rect 14292 9828 14293 9892
rect 14227 9827 14293 9828
rect 15738 9280 16058 10304
rect 16254 10029 16314 14587
rect 16438 12613 16498 17579
rect 16803 15332 16869 15333
rect 16803 15268 16804 15332
rect 16868 15268 16869 15332
rect 16803 15267 16869 15268
rect 16619 14924 16685 14925
rect 16619 14860 16620 14924
rect 16684 14860 16685 14924
rect 16619 14859 16685 14860
rect 16435 12612 16501 12613
rect 16435 12548 16436 12612
rect 16500 12548 16501 12612
rect 16435 12547 16501 12548
rect 16251 10028 16317 10029
rect 16251 9964 16252 10028
rect 16316 9964 16317 10028
rect 16251 9963 16317 9964
rect 16622 9757 16682 14859
rect 16806 13701 16866 15267
rect 16990 13973 17050 18667
rect 17907 17236 17973 17237
rect 17907 17172 17908 17236
rect 17972 17172 17973 17236
rect 17907 17171 17973 17172
rect 17171 16828 17237 16829
rect 17171 16764 17172 16828
rect 17236 16764 17237 16828
rect 17171 16763 17237 16764
rect 16987 13972 17053 13973
rect 16987 13908 16988 13972
rect 17052 13908 17053 13972
rect 16987 13907 17053 13908
rect 16803 13700 16869 13701
rect 16803 13636 16804 13700
rect 16868 13636 16869 13700
rect 16803 13635 16869 13636
rect 16990 12477 17050 13907
rect 17174 12885 17234 16763
rect 17910 13157 17970 17171
rect 18091 16964 18157 16965
rect 18091 16900 18092 16964
rect 18156 16900 18157 16964
rect 18091 16899 18157 16900
rect 17907 13156 17973 13157
rect 17907 13092 17908 13156
rect 17972 13092 17973 13156
rect 17907 13091 17973 13092
rect 17171 12884 17237 12885
rect 17171 12820 17172 12884
rect 17236 12820 17237 12884
rect 17171 12819 17237 12820
rect 16987 12476 17053 12477
rect 16987 12412 16988 12476
rect 17052 12412 17053 12476
rect 16987 12411 17053 12412
rect 17723 12476 17789 12477
rect 17723 12412 17724 12476
rect 17788 12412 17789 12476
rect 17723 12411 17789 12412
rect 16987 10708 17053 10709
rect 16987 10644 16988 10708
rect 17052 10644 17053 10708
rect 16987 10643 17053 10644
rect 16619 9756 16685 9757
rect 16619 9692 16620 9756
rect 16684 9692 16685 9756
rect 16619 9691 16685 9692
rect 15738 9216 15746 9280
rect 15810 9216 15826 9280
rect 15890 9216 15906 9280
rect 15970 9216 15986 9280
rect 16050 9216 16058 9280
rect 15738 8192 16058 9216
rect 15738 8128 15746 8192
rect 15810 8128 15826 8192
rect 15890 8128 15906 8192
rect 15970 8128 15986 8192
rect 16050 8128 16058 8192
rect 15738 7104 16058 8128
rect 15738 7040 15746 7104
rect 15810 7040 15826 7104
rect 15890 7040 15906 7104
rect 15970 7040 15986 7104
rect 16050 7040 16058 7104
rect 15738 6016 16058 7040
rect 15738 5952 15746 6016
rect 15810 5952 15826 6016
rect 15890 5952 15906 6016
rect 15970 5952 15986 6016
rect 16050 5952 16058 6016
rect 15738 4928 16058 5952
rect 15738 4864 15746 4928
rect 15810 4864 15826 4928
rect 15890 4864 15906 4928
rect 15970 4864 15986 4928
rect 16050 4864 16058 4928
rect 13307 4044 13373 4045
rect 13307 3980 13308 4044
rect 13372 3980 13373 4044
rect 13307 3979 13373 3980
rect 12040 3232 12048 3296
rect 12112 3232 12128 3296
rect 12192 3232 12208 3296
rect 12272 3232 12288 3296
rect 12352 3232 12360 3296
rect 12040 2208 12360 3232
rect 12040 2144 12048 2208
rect 12112 2144 12128 2208
rect 12192 2144 12208 2208
rect 12272 2144 12288 2208
rect 12352 2144 12360 2208
rect 12040 2128 12360 2144
rect 15738 3840 16058 4864
rect 16990 4589 17050 10643
rect 17171 8940 17237 8941
rect 17171 8876 17172 8940
rect 17236 8876 17237 8940
rect 17171 8875 17237 8876
rect 17174 8533 17234 8875
rect 17171 8532 17237 8533
rect 17171 8468 17172 8532
rect 17236 8468 17237 8532
rect 17171 8467 17237 8468
rect 17726 7717 17786 12411
rect 18094 9893 18154 16899
rect 18643 12884 18709 12885
rect 18643 12820 18644 12884
rect 18708 12820 18709 12884
rect 18643 12819 18709 12820
rect 18646 12341 18706 12819
rect 18643 12340 18709 12341
rect 18643 12276 18644 12340
rect 18708 12276 18709 12340
rect 18643 12275 18709 12276
rect 18091 9892 18157 9893
rect 18091 9828 18092 9892
rect 18156 9828 18157 9892
rect 18091 9827 18157 9828
rect 17723 7716 17789 7717
rect 17723 7652 17724 7716
rect 17788 7652 17789 7716
rect 17723 7651 17789 7652
rect 17726 7445 17786 7651
rect 17723 7444 17789 7445
rect 17723 7380 17724 7444
rect 17788 7380 17789 7444
rect 17723 7379 17789 7380
rect 19014 7173 19074 18667
rect 19437 18528 19757 19552
rect 19437 18464 19445 18528
rect 19509 18464 19525 18528
rect 19589 18464 19605 18528
rect 19669 18464 19685 18528
rect 19749 18464 19757 18528
rect 19195 17780 19261 17781
rect 19195 17716 19196 17780
rect 19260 17716 19261 17780
rect 19195 17715 19261 17716
rect 19198 16285 19258 17715
rect 19437 17440 19757 18464
rect 20115 18460 20181 18461
rect 20115 18396 20116 18460
rect 20180 18396 20181 18460
rect 20115 18395 20181 18396
rect 19931 18188 19997 18189
rect 19931 18124 19932 18188
rect 19996 18124 19997 18188
rect 19931 18123 19997 18124
rect 19437 17376 19445 17440
rect 19509 17376 19525 17440
rect 19589 17376 19605 17440
rect 19669 17376 19685 17440
rect 19749 17376 19757 17440
rect 19437 16352 19757 17376
rect 19437 16288 19445 16352
rect 19509 16288 19525 16352
rect 19589 16288 19605 16352
rect 19669 16288 19685 16352
rect 19749 16288 19757 16352
rect 19195 16284 19261 16285
rect 19195 16220 19196 16284
rect 19260 16220 19261 16284
rect 19195 16219 19261 16220
rect 19195 16148 19261 16149
rect 19195 16084 19196 16148
rect 19260 16084 19261 16148
rect 19195 16083 19261 16084
rect 19198 12341 19258 16083
rect 19437 15264 19757 16288
rect 19437 15200 19445 15264
rect 19509 15200 19525 15264
rect 19589 15200 19605 15264
rect 19669 15200 19685 15264
rect 19749 15200 19757 15264
rect 19437 14176 19757 15200
rect 19437 14112 19445 14176
rect 19509 14112 19525 14176
rect 19589 14112 19605 14176
rect 19669 14112 19685 14176
rect 19749 14112 19757 14176
rect 19437 13088 19757 14112
rect 19934 13701 19994 18123
rect 19931 13700 19997 13701
rect 19931 13636 19932 13700
rect 19996 13636 19997 13700
rect 19931 13635 19997 13636
rect 19437 13024 19445 13088
rect 19509 13024 19525 13088
rect 19589 13024 19605 13088
rect 19669 13024 19685 13088
rect 19749 13024 19757 13088
rect 19195 12340 19261 12341
rect 19195 12276 19196 12340
rect 19260 12276 19261 12340
rect 19195 12275 19261 12276
rect 19437 12000 19757 13024
rect 19931 12884 19997 12885
rect 19931 12820 19932 12884
rect 19996 12820 19997 12884
rect 19931 12819 19997 12820
rect 19437 11936 19445 12000
rect 19509 11936 19525 12000
rect 19589 11936 19605 12000
rect 19669 11936 19685 12000
rect 19749 11936 19757 12000
rect 19437 10912 19757 11936
rect 19437 10848 19445 10912
rect 19509 10848 19525 10912
rect 19589 10848 19605 10912
rect 19669 10848 19685 10912
rect 19749 10848 19757 10912
rect 19437 9824 19757 10848
rect 19437 9760 19445 9824
rect 19509 9760 19525 9824
rect 19589 9760 19605 9824
rect 19669 9760 19685 9824
rect 19749 9760 19757 9824
rect 19437 8736 19757 9760
rect 19437 8672 19445 8736
rect 19509 8672 19525 8736
rect 19589 8672 19605 8736
rect 19669 8672 19685 8736
rect 19749 8672 19757 8736
rect 19437 7648 19757 8672
rect 19934 8669 19994 12819
rect 20118 12477 20178 18395
rect 20299 12612 20365 12613
rect 20299 12548 20300 12612
rect 20364 12548 20365 12612
rect 20299 12547 20365 12548
rect 20115 12476 20181 12477
rect 20115 12412 20116 12476
rect 20180 12412 20181 12476
rect 20115 12411 20181 12412
rect 20115 11932 20181 11933
rect 20115 11868 20116 11932
rect 20180 11868 20181 11932
rect 20115 11867 20181 11868
rect 19931 8668 19997 8669
rect 19931 8604 19932 8668
rect 19996 8604 19997 8668
rect 19931 8603 19997 8604
rect 20118 8397 20178 11867
rect 20302 9077 20362 12547
rect 20670 12477 20730 19891
rect 21403 18052 21469 18053
rect 21403 17988 21404 18052
rect 21468 17988 21469 18052
rect 21403 17987 21469 17988
rect 21587 18052 21653 18053
rect 21587 17988 21588 18052
rect 21652 17988 21653 18052
rect 21587 17987 21653 17988
rect 20667 12476 20733 12477
rect 20667 12412 20668 12476
rect 20732 12412 20733 12476
rect 20667 12411 20733 12412
rect 20483 9212 20549 9213
rect 20483 9148 20484 9212
rect 20548 9148 20549 9212
rect 20483 9147 20549 9148
rect 20299 9076 20365 9077
rect 20299 9012 20300 9076
rect 20364 9012 20365 9076
rect 20299 9011 20365 9012
rect 20115 8396 20181 8397
rect 20115 8332 20116 8396
rect 20180 8332 20181 8396
rect 20115 8331 20181 8332
rect 19437 7584 19445 7648
rect 19509 7584 19525 7648
rect 19589 7584 19605 7648
rect 19669 7584 19685 7648
rect 19749 7584 19757 7648
rect 19011 7172 19077 7173
rect 19011 7108 19012 7172
rect 19076 7108 19077 7172
rect 19011 7107 19077 7108
rect 19437 6560 19757 7584
rect 19437 6496 19445 6560
rect 19509 6496 19525 6560
rect 19589 6496 19605 6560
rect 19669 6496 19685 6560
rect 19749 6496 19757 6560
rect 19437 5472 19757 6496
rect 19931 6356 19997 6357
rect 19931 6292 19932 6356
rect 19996 6292 19997 6356
rect 19931 6291 19997 6292
rect 19437 5408 19445 5472
rect 19509 5408 19525 5472
rect 19589 5408 19605 5472
rect 19669 5408 19685 5472
rect 19749 5408 19757 5472
rect 16987 4588 17053 4589
rect 16987 4524 16988 4588
rect 17052 4524 17053 4588
rect 16987 4523 17053 4524
rect 15738 3776 15746 3840
rect 15810 3776 15826 3840
rect 15890 3776 15906 3840
rect 15970 3776 15986 3840
rect 16050 3776 16058 3840
rect 15738 2752 16058 3776
rect 15738 2688 15746 2752
rect 15810 2688 15826 2752
rect 15890 2688 15906 2752
rect 15970 2688 15986 2752
rect 16050 2688 16058 2752
rect 15738 2128 16058 2688
rect 19437 4384 19757 5408
rect 19437 4320 19445 4384
rect 19509 4320 19525 4384
rect 19589 4320 19605 4384
rect 19669 4320 19685 4384
rect 19749 4320 19757 4384
rect 19437 3296 19757 4320
rect 19934 3637 19994 6291
rect 19931 3636 19997 3637
rect 19931 3572 19932 3636
rect 19996 3572 19997 3636
rect 19931 3571 19997 3572
rect 19437 3232 19445 3296
rect 19509 3232 19525 3296
rect 19589 3232 19605 3296
rect 19669 3232 19685 3296
rect 19749 3232 19757 3296
rect 19437 2208 19757 3232
rect 20302 2957 20362 9011
rect 20486 8125 20546 9147
rect 20483 8124 20549 8125
rect 20483 8060 20484 8124
rect 20548 8060 20549 8124
rect 20483 8059 20549 8060
rect 21406 4045 21466 17987
rect 21403 4044 21469 4045
rect 21403 3980 21404 4044
rect 21468 3980 21469 4044
rect 21403 3979 21469 3980
rect 20299 2956 20365 2957
rect 20299 2892 20300 2956
rect 20364 2892 20365 2956
rect 20299 2891 20365 2892
rect 21590 2549 21650 17987
rect 21587 2548 21653 2549
rect 21587 2484 21588 2548
rect 21652 2484 21653 2548
rect 21587 2483 21653 2484
rect 19437 2144 19445 2208
rect 19509 2144 19525 2208
rect 19589 2144 19605 2208
rect 19669 2144 19685 2208
rect 19749 2144 19757 2208
rect 19437 2128 19757 2144
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.mux_fabric_out_1.mux_l1_in_0_
timestamp 1608228718
transform 1 0 22172 0 1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1608228718
transform -1 0 23276 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_35_227
timestamp 1608228718
transform 1 0 21988 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _34_
timestamp 1608228718
transform 1 0 20608 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.mux_fabric_out_0.mux_l2_in_0_
timestamp 1608228718
transform 1 0 19596 0 1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_
timestamp 1608228718
transform 1 0 21160 0 1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_204
timestamp 1608228718
transform 1 0 21068 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_35_199
timestamp 1608228718
transform 1 0 19412 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_210
timestamp 1608228718
transform 1 0 20424 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_215
timestamp 1608228718
transform 1 0 20884 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _65_
timestamp 1608228718
transform 1 0 17480 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__buf_8  clk_0_FTB00
timestamp 1608228718
transform 1 0 18308 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_203
timestamp 1608228718
transform 1 0 18216 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_35_176
timestamp 1608228718
transform 1 0 17296 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_182
timestamp 1608228718
transform 1 0 17848 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_
timestamp 1608228718
transform 1 0 15456 0 1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0_
timestamp 1608228718
transform 1 0 16468 0 1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_202
timestamp 1608228718
transform 1 0 15364 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_35_153
timestamp 1608228718
transform 1 0 15180 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_165
timestamp 1608228718
transform 1 0 16284 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _70_
timestamp 1608228718
transform 1 0 14812 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.mux_fabric_out_1.mux_l2_in_0_
timestamp 1608228718
transform 1 0 13616 0 1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_35_134
timestamp 1608228718
transform 1 0 13432 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_145
timestamp 1608228718
transform 1 0 14444 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _53_
timestamp 1608228718
transform 1 0 12052 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.mux_fabric_out_1.mux_l1_in_0_
timestamp 1608228718
transform 1 0 12604 0 1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_201
timestamp 1608228718
transform 1 0 12512 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_35_117
timestamp 1608228718
transform 1 0 11868 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_122
timestamp 1608228718
transform 1 0 12328 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.mux_fabric_out_1.mux_l2_in_0_
timestamp 1608228718
transform 1 0 10028 0 1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.mux_fabric_out_0.mux_l2_in_0_
timestamp 1608228718
transform 1 0 11040 0 1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_200
timestamp 1608228718
transform 1 0 9660 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_89
timestamp 1608228718
transform 1 0 9292 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_35_94
timestamp 1608228718
transform 1 0 9752 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_35_106
timestamp 1608228718
transform 1 0 10856 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6_
timestamp 1608228718
transform 1 0 8924 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0_
timestamp 1608228718
transform 1 0 7912 0 1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_35_72
timestamp 1608228718
transform 1 0 7728 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_83
timestamp 1608228718
transform 1 0 8740 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _79_
timestamp 1608228718
transform 1 0 6072 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_
timestamp 1608228718
transform 1 0 6900 0 1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_199
timestamp 1608228718
transform 1 0 6808 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_35_52
timestamp 1608228718
transform 1 0 5888 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_58
timestamp 1608228718
transform 1 0 6440 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3_
timestamp 1608228718
transform 1 0 4048 0 1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_
timestamp 1608228718
transform 1 0 5060 0 1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_198
timestamp 1608228718
transform 1 0 3956 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_27
timestamp 1608228718
transform 1 0 3588 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_35_41
timestamp 1608228718
transform 1 0 4876 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_
timestamp 1608228718
transform 1 0 2760 0 1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2_
timestamp 1608228718
transform 1 0 1748 0 1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1608228718
transform 1 0 1104 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_35_3
timestamp 1608228718
transform 1 0 1380 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_35_16
timestamp 1608228718
transform 1 0 2576 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _68_
timestamp 1608228718
transform 1 0 22632 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.mux_fabric_out_1.mux_l1_in_0_
timestamp 1608228718
transform 1 0 21988 0 1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.mux_fabric_out_0.mux_l2_in_0_
timestamp 1608228718
transform 1 0 21804 0 -1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1608228718
transform -1 0 23276 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1608228718
transform -1 0 23276 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_33_236
timestamp 1608228718
transform 1 0 22816 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_34_224
timestamp 1608228718
transform 1 0 21712 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0_
timestamp 1608228718
transform 1 0 21160 0 1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608228718
transform 1 0 19688 0 1 20128
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.mux_fabric_out_0.mux_l1_in_0_
timestamp 1608228718
transform 1 0 19780 0 -1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.mux_fabric_out_1.mux_l2_in_0_
timestamp 1608228718
transform 1 0 20884 0 -1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_197
timestamp 1608228718
transform 1 0 20792 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_33_200
timestamp 1608228718
transform 1 0 19504 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_201
timestamp 1608228718
transform 1 0 19596 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_212
timestamp 1608228718
transform 1 0 20608 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608228718
transform 1 0 18032 0 1 20128
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608228718
transform 1 0 18124 0 -1 21216
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_193
timestamp 1608228718
transform 1 0 17940 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_178
timestamp 1608228718
transform 1 0 17480 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_182
timestamp 1608228718
transform 1 0 17848 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_181
timestamp 1608228718
transform 1 0 17756 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3_
timestamp 1608228718
transform 1 0 16928 0 -1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608228718
transform 1 0 15272 0 -1 21216
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608228718
transform 1 0 16008 0 1 20128
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_196
timestamp 1608228718
transform 1 0 15180 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_33_160
timestamp 1608228718
transform 1 0 15824 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_170
timestamp 1608228718
transform 1 0 16744 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _54_
timestamp 1608228718
transform 1 0 14720 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_16_
timestamp 1608228718
transform 1 0 14352 0 1 20128
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_33_142
timestamp 1608228718
transform 1 0 14168 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_146
timestamp 1608228718
transform 1 0 14536 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_151
timestamp 1608228718
transform 1 0 14996 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608228718
transform 1 0 11316 0 -1 21216
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_14_
timestamp 1608228718
transform 1 0 12696 0 1 20128
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_15_
timestamp 1608228718
transform 1 0 13064 0 -1 21216
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_192
timestamp 1608228718
transform 1 0 12328 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_118
timestamp 1608228718
transform 1 0 11960 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_33_123
timestamp 1608228718
transform 1 0 12420 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_34_127
timestamp 1608228718
transform 1 0 12788 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608228718
transform 1 0 9660 0 -1 21216
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608228718
transform 1 0 10488 0 1 20128
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_195
timestamp 1608228718
transform 1 0 9568 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_33_100
timestamp 1608228718
transform 1 0 10304 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_90
timestamp 1608228718
transform 1 0 9384 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_109
timestamp 1608228718
transform 1 0 11132 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608228718
transform 1 0 8832 0 1 20128
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.mux_fabric_out_0.mux_l2_in_0_
timestamp 1608228718
transform 1 0 8556 0 -1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_33_78
timestamp 1608228718
transform 1 0 8280 0 1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_34_77
timestamp 1608228718
transform 1 0 8188 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0_
timestamp 1608228718
transform 1 0 5704 0 -1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_
timestamp 1608228718
transform 1 0 6072 0 1 20128
box -38 -48 498 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608228718
transform 1 0 6808 0 1 20128
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608228718
transform 1 0 6716 0 -1 21216
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_191
timestamp 1608228718
transform 1 0 6716 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_33_52
timestamp 1608228718
transform 1 0 5888 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_59
timestamp 1608228718
transform 1 0 6532 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_48
timestamp 1608228718
transform 1 0 5520 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_59
timestamp 1608228718
transform 1 0 6532 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1_
timestamp 1608228718
transform 1 0 5060 0 1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_16_
timestamp 1608228718
transform 1 0 3404 0 1 20128
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608228718
transform 1 0 4048 0 -1 21216
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_194
timestamp 1608228718
transform 1 0 3956 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_33_23
timestamp 1608228718
transform 1 0 3220 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_41
timestamp 1608228718
transform 1 0 4876 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_27
timestamp 1608228718
transform 1 0 3588 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _75_
timestamp 1608228718
transform 1 0 1564 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_14_
timestamp 1608228718
transform 1 0 1748 0 1 20128
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_15_
timestamp 1608228718
transform 1 0 2116 0 -1 21216
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1608228718
transform 1 0 1104 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1608228718
transform 1 0 1104 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_33_3
timestamp 1608228718
transform 1 0 1380 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_34_3
timestamp 1608228718
transform 1 0 1380 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_9
timestamp 1608228718
transform 1 0 1932 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _67_
timestamp 1608228718
transform 1 0 22632 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1608228718
transform -1 0 23276 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_15_
timestamp 1608228718
transform 1 0 21160 0 -1 20128
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_190
timestamp 1608228718
transform 1 0 20792 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_212
timestamp 1608228718
transform 1 0 20608 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_32_215
timestamp 1608228718
transform 1 0 20884 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_
timestamp 1608228718
transform 1 0 18124 0 -1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608228718
transform 1 0 19136 0 -1 20128
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_32_183
timestamp 1608228718
transform 1 0 17940 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_194
timestamp 1608228718
transform 1 0 18952 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_
timestamp 1608228718
transform 1 0 15272 0 -1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608228718
transform 1 0 16468 0 -1 20128
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_189
timestamp 1608228718
transform 1 0 15180 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_163
timestamp 1608228718
transform 1 0 16100 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_
timestamp 1608228718
transform 1 0 14536 0 -1 20128
box -38 -48 498 592
use sky130_fd_sc_hd__decap_4  FILLER_32_142
timestamp 1608228718
transform 1 0 14168 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_32_151
timestamp 1608228718
transform 1 0 14996 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_13_
timestamp 1608228718
transform 1 0 12696 0 -1 20128
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_32_124
timestamp 1608228718
transform 1 0 12512 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__sdfxtp_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_clb_fle_ff_0.sky130_fd_sc_hd__sdfxtp_1_0_
timestamp 1608228718
transform 1 0 10580 0 -1 20128
box -38 -48 1970 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_1_
timestamp 1608228718
transform 1 0 9660 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_188
timestamp 1608228718
transform 1 0 9568 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_7_0_ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
timestamp 1608228718
transform 1 0 10212 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_32_88
timestamp 1608228718
transform 1 0 9200 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_32_97
timestamp 1608228718
transform 1 0 10028 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_32_102
timestamp 1608228718
transform 1 0 10488 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_
timestamp 1608228718
transform 1 0 8832 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608228718
transform 1 0 7176 0 -1 20128
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_32_82
timestamp 1608228718
transform 1 0 8648 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608228718
transform 1 0 5336 0 -1 20128
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_32_45
timestamp 1608228718
transform 1 0 5244 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_62
timestamp 1608228718
transform 1 0 6808 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _76_
timestamp 1608228718
transform 1 0 3220 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_
timestamp 1608228718
transform 1 0 4048 0 -1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_187
timestamp 1608228718
transform 1 0 3956 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_27
timestamp 1608228718
transform 1 0 3588 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_41
timestamp 1608228718
transform 1 0 4876 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_13_
timestamp 1608228718
transform 1 0 1564 0 -1 20128
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1608228718
transform 1 0 1104 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_32_3
timestamp 1608228718
transform 1 0 1380 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_21
timestamp 1608228718
transform 1 0 3036 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1608228718
transform -1 0 23276 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_31_231
timestamp 1608228718
transform 1 0 22356 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_237
timestamp 1608228718
transform 1 0 22908 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_
timestamp 1608228718
transform 1 0 20056 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_13_
timestamp 1608228718
transform 1 0 20884 0 1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_31_205
timestamp 1608228718
transform 1 0 19964 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _32_
timestamp 1608228718
transform 1 0 17480 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_clb_fle_ff_1.sky130_fd_sc_hd__sdfxtp_1_0_
timestamp 1608228718
transform 1 0 18032 0 1 19040
box -38 -48 1970 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_186
timestamp 1608228718
transform 1 0 17940 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_31_176
timestamp 1608228718
transform 1 0 17296 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_181
timestamp 1608228718
transform 1 0 17756 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_
timestamp 1608228718
transform 1 0 15456 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2_
timestamp 1608228718
transform 1 0 16468 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_31_154
timestamp 1608228718
transform 1 0 15272 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_165
timestamp 1608228718
transform 1 0 16284 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.mux_ff_0_D_0.mux_l1_in_0_
timestamp 1608228718
transform 1 0 13432 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_
timestamp 1608228718
transform 1 0 14444 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_31_132
timestamp 1608228718
transform 1 0 13248 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_143
timestamp 1608228718
transform 1 0 14260 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.mux_fabric_out_1.mux_l1_in_0_
timestamp 1608228718
transform 1 0 12420 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_185
timestamp 1608228718
transform 1 0 12328 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_31_120
timestamp 1608228718
transform 1 0 12144 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608228718
transform 1 0 10672 0 1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.mux_fabric_out_0.mux_l1_in_0_
timestamp 1608228718
transform 1 0 9660 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_31_91
timestamp 1608228718
transform 1 0 9476 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_102
timestamp 1608228718
transform 1 0 10488 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__sdfxtp_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_clb_fle_ff_1.sky130_fd_sc_hd__sdfxtp_1_0_
timestamp 1608228718
transform 1 0 7544 0 1 19040
box -38 -48 1970 592
use sky130_fd_sc_hd__decap_4  FILLER_31_66
timestamp 1608228718
transform 1 0 7176 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _56_
timestamp 1608228718
transform 1 0 6256 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _82_
timestamp 1608228718
transform 1 0 6808 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_184
timestamp 1608228718
transform 1 0 6716 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_31_54
timestamp 1608228718
transform 1 0 6072 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_59
timestamp 1608228718
transform 1 0 6532 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_
timestamp 1608228718
transform 1 0 3588 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608228718
transform 1 0 4600 0 1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_31_25
timestamp 1608228718
transform 1 0 3404 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_36
timestamp 1608228718
transform 1 0 4416 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_
timestamp 1608228718
transform 1 0 2576 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_
timestamp 1608228718
transform 1 0 1564 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1608228718
transform 1 0 1104 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_31_3
timestamp 1608228718
transform 1 0 1380 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_14
timestamp 1608228718
transform 1 0 2392 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _49_
timestamp 1608228718
transform 1 0 22540 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_
timestamp 1608228718
transform 1 0 21344 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1608228718
transform -1 0 23276 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_3
timestamp 1608228718
transform 1 0 22356 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_30_219
timestamp 1608228718
transform 1 0 21252 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_229
timestamp 1608228718
transform 1 0 22172 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_236
timestamp 1608228718
transform 1 0 22816 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _50_
timestamp 1608228718
transform 1 0 20332 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_183
timestamp 1608228718
transform 1 0 20792 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_5
timestamp 1608228718
transform 1 0 20148 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_205
timestamp 1608228718
transform 1 0 19964 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_212
timestamp 1608228718
transform 1 0 20608 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_215
timestamp 1608228718
transform 1 0 20884 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_
timestamp 1608228718
transform 1 0 19136 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_9_
timestamp 1608228718
transform 1 0 17664 0 -1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_15_0_ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
timestamp 1608228718
transform 1 0 17388 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_30_175
timestamp 1608228718
transform 1 0 17204 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _35_
timestamp 1608228718
transform 1 0 15272 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608228718
transform 1 0 15732 0 -1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_182
timestamp 1608228718
transform 1 0 15180 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_157
timestamp 1608228718
transform 1 0 15548 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _72_
timestamp 1608228718
transform 1 0 14628 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_30_141
timestamp 1608228718
transform 1 0 14076 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_30_151
timestamp 1608228718
transform 1 0 14996 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_
timestamp 1608228718
transform 1 0 11776 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_12_
timestamp 1608228718
transform 1 0 12604 0 -1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_30_114
timestamp 1608228718
transform 1 0 11592 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_120
timestamp 1608228718
transform 1 0 12144 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_124
timestamp 1608228718
transform 1 0 12512 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__sdfxtp_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_clb_fle_ff_1.sky130_fd_sc_hd__sdfxtp_1_0_
timestamp 1608228718
transform 1 0 9660 0 -1 19040
box -38 -48 1970 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_181
timestamp 1608228718
transform 1 0 9568 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_30_89
timestamp 1608228718
transform 1 0 9292 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_
timestamp 1608228718
transform 1 0 8464 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_30_78
timestamp 1608228718
transform 1 0 8280 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _81_
timestamp 1608228718
transform 1 0 6164 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_
timestamp 1608228718
transform 1 0 5152 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608228718
transform 1 0 6808 0 -1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_30_53
timestamp 1608228718
transform 1 0 5980 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_30_59
timestamp 1608228718
transform 1 0 6532 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _77_
timestamp 1608228718
transform 1 0 3220 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_
timestamp 1608228718
transform 1 0 4048 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_180
timestamp 1608228718
transform 1 0 3956 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_27
timestamp 1608228718
transform 1 0 3588 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_30_41
timestamp 1608228718
transform 1 0 4876 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_12_
timestamp 1608228718
transform 1 0 1564 0 -1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1608228718
transform 1 0 1104 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_30_3
timestamp 1608228718
transform 1 0 1380 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_21
timestamp 1608228718
transform 1 0 3036 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0_
timestamp 1608228718
transform 1 0 21896 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1608228718
transform -1 0 23276 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_29_223
timestamp 1608228718
transform 1 0 21620 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_29_235
timestamp 1608228718
transform 1 0 22724 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_12_
timestamp 1608228718
transform 1 0 20148 0 1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_29_205
timestamp 1608228718
transform 1 0 19964 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _33_
timestamp 1608228718
transform 1 0 18032 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_11_
timestamp 1608228718
transform 1 0 18492 0 1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_179
timestamp 1608228718
transform 1 0 17940 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_179
timestamp 1608228718
transform 1 0 17572 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_29_187
timestamp 1608228718
transform 1 0 18308 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__sdfxtp_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_clb_fle_ff_0.sky130_fd_sc_hd__sdfxtp_1_0_
timestamp 1608228718
transform 1 0 15640 0 1 17952
box -38 -48 1970 592
use sky130_fd_sc_hd__decap_3  FILLER_29_155
timestamp 1608228718
transform 1 0 15364 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_
timestamp 1608228718
transform 1 0 14536 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_29_144
timestamp 1608228718
transform 1 0 14352 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _55_
timestamp 1608228718
transform 1 0 12420 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_11_
timestamp 1608228718
transform 1 0 12880 0 1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_178
timestamp 1608228718
transform 1 0 12328 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_118
timestamp 1608228718
transform 1 0 11960 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_29_126
timestamp 1608228718
transform 1 0 12696 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.mux_fabric_out_0.mux_l1_in_0_
timestamp 1608228718
transform 1 0 9384 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608228718
transform 1 0 10488 0 1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_29_88
timestamp 1608228718
transform 1 0 9200 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_29_99
timestamp 1608228718
transform 1 0 10212 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_clb_fle_ff_0.sky130_fd_sc_hd__sdfxtp_1_0_
timestamp 1608228718
transform 1 0 7268 0 1 17952
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _52_
timestamp 1608228718
transform 1 0 6808 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _57_
timestamp 1608228718
transform 1 0 6256 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_
timestamp 1608228718
transform 1 0 5244 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_177
timestamp 1608228718
transform 1 0 6716 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_29_44
timestamp 1608228718
transform 1 0 5152 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_29_54
timestamp 1608228718
transform 1 0 6072 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_59
timestamp 1608228718
transform 1 0 6532 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_65
timestamp 1608228718
transform 1 0 7084 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_9_
timestamp 1608228718
transform 1 0 3312 0 1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_29_22
timestamp 1608228718
transform 1 0 3128 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_40
timestamp 1608228718
transform 1 0 4784 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_11_
timestamp 1608228718
transform 1 0 1656 0 1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1608228718
transform 1 0 1104 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_29_3
timestamp 1608228718
transform 1 0 1380 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _48_
timestamp 1608228718
transform 1 0 22540 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1608228718
transform -1 0 23276 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_28_231
timestamp 1608228718
transform 1 0 22356 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_236
timestamp 1608228718
transform 1 0 22816 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.mux_ff_0_D_0.mux_l1_in_0_
timestamp 1608228718
transform 1 0 19780 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_14_
timestamp 1608228718
transform 1 0 20884 0 -1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_176
timestamp 1608228718
transform 1 0 20792 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_28_201
timestamp 1608228718
transform 1 0 19596 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_212
timestamp 1608228718
transform 1 0 20608 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_10_
timestamp 1608228718
transform 1 0 18124 0 -1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_28_181
timestamp 1608228718
transform 1 0 17756 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0_
timestamp 1608228718
transform 1 0 16928 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_9_
timestamp 1608228718
transform 1 0 15272 0 -1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_175
timestamp 1608228718
transform 1 0 15180 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_28_170
timestamp 1608228718
transform 1 0 16744 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _74_
timestamp 1608228718
transform 1 0 14628 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_28_145
timestamp 1608228718
transform 1 0 14444 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_151
timestamp 1608228718
transform 1 0 14996 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.mux_ff_0_D_0.mux_l2_in_0_
timestamp 1608228718
transform 1 0 11408 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_
timestamp 1608228718
transform 1 0 12420 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_10_
timestamp 1608228718
transform 1 0 12972 0 -1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_28_110
timestamp 1608228718
transform 1 0 11224 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_121
timestamp 1608228718
transform 1 0 12236 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_127
timestamp 1608228718
transform 1 0 12788 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608228718
transform 1 0 9752 0 -1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_174
timestamp 1608228718
transform 1 0 9568 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_88
timestamp 1608228718
transform 1 0 9200 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_93
timestamp 1608228718
transform 1 0 9660 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0_
timestamp 1608228718
transform 1 0 8372 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_28_77
timestamp 1608228718
transform 1 0 8188 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608228718
transform 1 0 6716 0 -1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_28_58
timestamp 1608228718
transform 1 0 6440 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _78_
timestamp 1608228718
transform 1 0 3404 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _80_
timestamp 1608228718
transform 1 0 4048 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608228718
transform 1 0 4968 0 -1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_173
timestamp 1608228718
transform 1 0 3956 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_28_23
timestamp 1608228718
transform 1 0 3220 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_29
timestamp 1608228718
transform 1 0 3772 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_28_36
timestamp 1608228718
transform 1 0 4416 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_10_
timestamp 1608228718
transform 1 0 1748 0 -1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1608228718
transform 1 0 1104 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_28_3
timestamp 1608228718
transform 1 0 1380 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_
timestamp 1608228718
transform 1 0 21896 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_16_
timestamp 1608228718
transform 1 0 21344 0 1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1608228718
transform -1 0 23276 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1608228718
transform -1 0 23276 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_26_224
timestamp 1608228718
transform 1 0 21712 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_26_235
timestamp 1608228718
transform 1 0 22724 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_27_236
timestamp 1608228718
transform 1 0 22816 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1_
timestamp 1608228718
transform 1 0 19872 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.mux_ff_0_D_0.mux_l2_in_0_
timestamp 1608228718
transform 1 0 19688 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0_
timestamp 1608228718
transform 1 0 20884 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_
timestamp 1608228718
transform 1 0 20700 0 1 16864
box -38 -48 498 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_169
timestamp 1608228718
transform 1 0 20792 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_26_213
timestamp 1608228718
transform 1 0 20700 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_200
timestamp 1608228718
transform 1 0 19504 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_211
timestamp 1608228718
transform 1 0 20516 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_218
timestamp 1608228718
transform 1 0 21160 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _58_
timestamp 1608228718
transform 1 0 17480 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_7_
timestamp 1608228718
transform 1 0 18400 0 -1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_8_
timestamp 1608228718
transform 1 0 18032 0 1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_172
timestamp 1608228718
transform 1 0 17940 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_176
timestamp 1608228718
transform 1 0 17296 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_181
timestamp 1608228718
transform 1 0 17756 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.mux_fabric_out_1.mux_l2_in_0_
timestamp 1608228718
transform 1 0 15456 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_
timestamp 1608228718
transform 1 0 16468 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_7_
timestamp 1608228718
transform 1 0 15272 0 -1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_6_
timestamp 1608228718
transform 1 0 16928 0 -1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_168
timestamp 1608228718
transform 1 0 15180 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_170
timestamp 1608228718
transform 1 0 16744 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_154
timestamp 1608228718
transform 1 0 15272 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_165
timestamp 1608228718
transform 1 0 16284 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.mux_fabric_out_1.mux_l1_in_0_
timestamp 1608228718
transform 1 0 13984 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_8_
timestamp 1608228718
transform 1 0 13800 0 1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_13_0_ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
timestamp 1608228718
transform 1 0 13524 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_26_138
timestamp 1608228718
transform 1 0 13800 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_149
timestamp 1608228718
transform 1 0 14812 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_27_132
timestamp 1608228718
transform 1 0 13248 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.mux_ff_0_D_0.mux_l1_in_0_
timestamp 1608228718
transform 1 0 11316 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608228718
transform 1 0 12328 0 -1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.mux_fabric_out_0.mux_l2_in_0_
timestamp 1608228718
transform 1 0 12420 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_171
timestamp 1608228718
transform 1 0 12328 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_120
timestamp 1608228718
transform 1 0 12144 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_120
timestamp 1608228718
transform 1 0 12144 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_
timestamp 1608228718
transform 1 0 9660 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__sdfxtp_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_clb_fle_ff_1.sky130_fd_sc_hd__sdfxtp_1_0_
timestamp 1608228718
transform 1 0 10212 0 -1 16864
box -38 -48 1970 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608228718
transform 1 0 9660 0 1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_167
timestamp 1608228718
transform 1 0 9568 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_3_0_ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
timestamp 1608228718
transform 1 0 9292 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_26_97
timestamp 1608228718
transform 1 0 10028 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_91
timestamp 1608228718
transform 1 0 9476 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_109
timestamp 1608228718
transform 1 0 11132 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_1_
timestamp 1608228718
transform 1 0 8740 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608228718
transform 1 0 8004 0 1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_26_81
timestamp 1608228718
transform 1 0 8556 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_87
timestamp 1608228718
transform 1 0 9108 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_73
timestamp 1608228718
transform 1 0 7820 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__or2_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_
timestamp 1608228718
transform 1 0 6440 0 -1 16864
box -38 -48 498 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608228718
transform 1 0 7084 0 -1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0_
timestamp 1608228718
transform 1 0 6992 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_170
timestamp 1608228718
transform 1 0 6716 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_56
timestamp 1608228718
transform 1 0 6256 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_63
timestamp 1608228718
transform 1 0 6900 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_57
timestamp 1608228718
transform 1 0 6348 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_62
timestamp 1608228718
transform 1 0 6808 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608228718
transform 1 0 4876 0 1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608228718
transform 1 0 4784 0 -1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_0_
timestamp 1608228718
transform 1 0 4324 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_2_
timestamp 1608228718
transform 1 0 4232 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_38
timestamp 1608228718
transform 1 0 4600 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_39
timestamp 1608228718
transform 1 0 4692 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_166
timestamp 1608228718
transform 1 0 3956 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_5_0_ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
timestamp 1608228718
transform 1 0 4048 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_26_27
timestamp 1608228718
transform 1 0 3588 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_32
timestamp 1608228718
transform 1 0 4048 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_27_29
timestamp 1608228718
transform 1 0 3772 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_7_
timestamp 1608228718
transform 1 0 2116 0 -1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_8_
timestamp 1608228718
transform 1 0 2300 0 1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_27_11
timestamp 1608228718
transform 1 0 2116 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_3_
timestamp 1608228718
transform 1 0 1748 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_4_
timestamp 1608228718
transform 1 0 1564 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1608228718
transform 1 0 1104 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1608228718
transform 1 0 1104 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_26_3
timestamp 1608228718
transform 1 0 1380 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_9
timestamp 1608228718
transform 1 0 1932 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_3
timestamp 1608228718
transform 1 0 1380 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608228718
transform 1 0 21344 0 1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1608228718
transform -1 0 23276 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_25_236
timestamp 1608228718
transform 1 0 22816 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_
timestamp 1608228718
transform 1 0 19688 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_
timestamp 1608228718
transform 1 0 20516 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_7
timestamp 1608228718
transform 1 0 19504 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _73_
timestamp 1608228718
transform 1 0 17388 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_165
timestamp 1608228718
transform 1 0 17940 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_181
timestamp 1608228718
transform 1 0 17756 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_25_184
timestamp 1608228718
transform 1 0 18032 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_25_196
timestamp 1608228718
transform 1 0 19136 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_6_
timestamp 1608228718
transform 1 0 15456 0 1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_7_0_ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
timestamp 1608228718
transform 1 0 17112 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_25_154
timestamp 1608228718
transform 1 0 15272 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_172
timestamp 1608228718
transform 1 0 16928 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_4_
timestamp 1608228718
transform 1 0 13800 0 1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_6_0_ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
timestamp 1608228718
transform 1 0 13524 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_25_132
timestamp 1608228718
transform 1 0 13248 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_
timestamp 1608228718
transform 1 0 11776 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.mux_fabric_out_0.mux_l1_in_0_
timestamp 1608228718
transform 1 0 12420 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_164
timestamp 1608228718
transform 1 0 12328 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_114
timestamp 1608228718
transform 1 0 11592 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_120
timestamp 1608228718
transform 1 0 12144 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0_
timestamp 1608228718
transform 1 0 10764 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_25_103
timestamp 1608228718
transform 1 0 10580 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_
timestamp 1608228718
transform 1 0 7360 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__sdfxtp_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_clb_fle_ff_0.sky130_fd_sc_hd__sdfxtp_1_0_
timestamp 1608228718
transform 1 0 8648 0 1 15776
box -38 -48 1970 592
use sky130_fd_sc_hd__fill_2  FILLER_25_66
timestamp 1608228718
transform 1 0 7176 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_77
timestamp 1608228718
transform 1 0 8188 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_81
timestamp 1608228718
transform 1 0 8556 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_2_
timestamp 1608228718
transform 1 0 6808 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_163
timestamp 1608228718
transform 1 0 6716 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_2_0_ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
timestamp 1608228718
transform 1 0 6440 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_25_56
timestamp 1608228718
transform 1 0 6256 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2_
timestamp 1608228718
transform 1 0 3128 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_
timestamp 1608228718
transform 1 0 4232 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1608228718
transform 1 0 4784 0 1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_25_31
timestamp 1608228718
transform 1 0 3956 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_25_38
timestamp 1608228718
transform 1 0 4600 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_4_
timestamp 1608228718
transform 1 0 1472 0 1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1608228718
transform 1 0 1104 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_25_3
timestamp 1608228718
transform 1 0 1380 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_20
timestamp 1608228718
transform 1 0 2944 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1608228718
transform -1 0 23276 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_24_232
timestamp 1608228718
transform 1 0 22448 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _69_
timestamp 1608228718
transform 1 0 20424 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _71_
timestamp 1608228718
transform 1 0 20056 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608228718
transform 1 0 20976 0 -1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_162
timestamp 1608228718
transform 1 0 20792 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_24_215
timestamp 1608228718
transform 1 0 20884 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1608228718
transform 1 0 18584 0 -1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_24_188
timestamp 1608228718
transform 1 0 18400 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_5_
timestamp 1608228718
transform 1 0 15272 0 -1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_5_
timestamp 1608228718
transform 1 0 16928 0 -1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_161
timestamp 1608228718
transform 1 0 15180 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_170
timestamp 1608228718
transform 1 0 16744 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_
timestamp 1608228718
transform 1 0 14352 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_3_0_ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
timestamp 1608228718
transform 1 0 14904 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_24_142
timestamp 1608228718
transform 1 0 14168 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_148
timestamp 1608228718
transform 1 0 14720 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608228718
transform 1 0 12696 0 -1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_1_0_0_ltile_clb_mode__0.clb_clk
timestamp 1608228718
transform 1 0 12420 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_24_120
timestamp 1608228718
transform 1 0 12144 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.mux_ff_0_D_0.mux_l2_in_0_
timestamp 1608228718
transform 1 0 9660 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608228718
transform 1 0 10672 0 -1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_160
timestamp 1608228718
transform 1 0 9568 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_90
timestamp 1608228718
transform 1 0 9384 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_102
timestamp 1608228718
transform 1 0 10488 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_0_
timestamp 1608228718
transform 1 0 9016 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608228718
transform 1 0 7360 0 -1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_24_66
timestamp 1608228718
transform 1 0 7176 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_84
timestamp 1608228718
transform 1 0 8832 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_16_
timestamp 1608228718
transform 1 0 5704 0 -1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_24_47
timestamp 1608228718
transform 1 0 5428 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3_
timestamp 1608228718
transform 1 0 4600 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6_
timestamp 1608228718
transform 1 0 4048 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_
timestamp 1608228718
transform 1 0 3404 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_159
timestamp 1608228718
transform 1 0 3956 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_23
timestamp 1608228718
transform 1 0 3220 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_29
timestamp 1608228718
transform 1 0 3772 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_36
timestamp 1608228718
transform 1 0 4416 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_5_
timestamp 1608228718
transform 1 0 1748 0 -1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1608228718
transform 1 0 1104 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_24_3
timestamp 1608228718
transform 1 0 1380 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2_
timestamp 1608228718
transform 1 0 21896 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1608228718
transform -1 0 23276 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_23_224
timestamp 1608228718
transform 1 0 21712 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_23_235
timestamp 1608228718
transform 1 0 22724 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_
timestamp 1608228718
transform 1 0 19872 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3_
timestamp 1608228718
transform 1 0 20884 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_23_202
timestamp 1608228718
transform 1 0 19688 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_213
timestamp 1608228718
transform 1 0 20700 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608228718
transform 1 0 18216 0 1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_158
timestamp 1608228718
transform 1 0 17940 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_23_181
timestamp 1608228718
transform 1 0 17756 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_184
timestamp 1608228718
transform 1 0 18032 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_0_
timestamp 1608228718
transform 1 0 15732 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_4_
timestamp 1608228718
transform 1 0 16284 0 1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_23_157
timestamp 1608228718
transform 1 0 15548 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_163
timestamp 1608228718
transform 1 0 16100 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1608228718
transform 1 0 14076 0 1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_23_139
timestamp 1608228718
transform 1 0 13892 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608228718
transform 1 0 12420 0 1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_157
timestamp 1608228718
transform 1 0 12328 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_23_120
timestamp 1608228718
transform 1 0 12144 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608228718
transform 1 0 10672 0 1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_23_100
timestamp 1608228718
transform 1 0 10304 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0_
timestamp 1608228718
transform 1 0 7820 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608228718
transform 1 0 8832 0 1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_23_71
timestamp 1608228718
transform 1 0 7636 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_82
timestamp 1608228718
transform 1 0 8648 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_
timestamp 1608228718
transform 1 0 5612 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_
timestamp 1608228718
transform 1 0 6808 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_156
timestamp 1608228718
transform 1 0 6716 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_23_47
timestamp 1608228718
transform 1 0 5428 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_23_58
timestamp 1608228718
transform 1 0 6440 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_
timestamp 1608228718
transform 1 0 3588 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_
timestamp 1608228718
transform 1 0 4600 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_23_25
timestamp 1608228718
transform 1 0 3404 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_36
timestamp 1608228718
transform 1 0 4416 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5_
timestamp 1608228718
transform 1 0 1380 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_6_
timestamp 1608228718
transform 1 0 1932 0 1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1608228718
transform 1 0 1104 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_23_7
timestamp 1608228718
transform 1 0 1748 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1608228718
transform -1 0 23276 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_22_234
timestamp 1608228718
transform 1 0 22632 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_
timestamp 1608228718
transform 1 0 19504 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608228718
transform 1 0 21160 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_155
timestamp 1608228718
transform 1 0 20792 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_14_0_ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
timestamp 1608228718
transform 1 0 20516 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_22_198
timestamp 1608228718
transform 1 0 19320 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_209
timestamp 1608228718
transform 1 0 20332 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_22_215
timestamp 1608228718
transform 1 0 20884 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608228718
transform 1 0 17848 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_22_181
timestamp 1608228718
transform 1 0 17756 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0_
timestamp 1608228718
transform 1 0 15272 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.mux_ff_0_D_0.mux_l2_in_0_
timestamp 1608228718
transform 1 0 16100 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_
timestamp 1608228718
transform 1 0 16928 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_154
timestamp 1608228718
transform 1 0 15180 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_
timestamp 1608228718
transform 1 0 13432 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_
timestamp 1608228718
transform 1 0 14260 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_22_133
timestamp 1608228718
transform 1 0 13340 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_22_152
timestamp 1608228718
transform 1 0 15088 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_
timestamp 1608228718
transform 1 0 12972 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608228718
transform 1 0 11500 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608228718
transform 1 0 9660 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_153
timestamp 1608228718
transform 1 0 9568 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_88
timestamp 1608228718
transform 1 0 9200 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_109
timestamp 1608228718
transform 1 0 11132 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_
timestamp 1608228718
transform 1 0 7360 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0_
timestamp 1608228718
transform 1 0 8372 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_22_66
timestamp 1608228718
transform 1 0 7176 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_77
timestamp 1608228718
transform 1 0 8188 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_15_
timestamp 1608228718
transform 1 0 5704 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_22_48
timestamp 1608228718
transform 1 0 5520 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5_
timestamp 1608228718
transform 1 0 3404 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_13_
timestamp 1608228718
transform 1 0 4048 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_152
timestamp 1608228718
transform 1 0 3956 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_4_0_ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
timestamp 1608228718
transform 1 0 3128 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_22_29
timestamp 1608228718
transform 1 0 3772 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_9_
timestamp 1608228718
transform 1 0 1472 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1608228718
transform 1 0 1104 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_22_3
timestamp 1608228718
transform 1 0 1380 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_20
timestamp 1608228718
transform 1 0 2944 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_
timestamp 1608228718
transform 1 0 21896 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1608228718
transform -1 0 23276 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_21_224
timestamp 1608228718
transform 1 0 21712 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_21_235
timestamp 1608228718
transform 1 0 22724 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_clb_fle_ff_1.sky130_fd_sc_hd__sdfxtp_1_0_
timestamp 1608228718
transform 1 0 19780 0 1 13600
box -38 -48 1970 592
use sky130_fd_sc_hd__decap_3  FILLER_21_200
timestamp 1608228718
transform 1 0 19504 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _47_
timestamp 1608228718
transform 1 0 17664 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_1_
timestamp 1608228718
transform 1 0 17296 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608228718
transform 1 0 18032 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_151
timestamp 1608228718
transform 1 0 17940 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_21_175
timestamp 1608228718
transform 1 0 17204 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.mux_ff_0_D_0.mux_l1_in_0_
timestamp 1608228718
transform 1 0 15548 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_
timestamp 1608228718
transform 1 0 16376 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_ltile_clb_mode__0.clb_clk
timestamp 1608228718
transform 1 0 13708 0 1 13600
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_4  FILLER_21_132
timestamp 1608228718
transform 1 0 13248 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_136
timestamp 1608228718
transform 1 0 13616 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_
timestamp 1608228718
transform 1 0 12420 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_0_
timestamp 1608228718
transform 1 0 11776 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_150
timestamp 1608228718
transform 1 0 12328 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_114
timestamp 1608228718
transform 1 0 11592 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_120
timestamp 1608228718
transform 1 0 12144 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_
timestamp 1608228718
transform 1 0 10764 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3_
timestamp 1608228718
transform 1 0 9752 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_21_91
timestamp 1608228718
transform 1 0 9476 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_21_103
timestamp 1608228718
transform 1 0 10580 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_
timestamp 1608228718
transform 1 0 8648 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_21_80
timestamp 1608228718
transform 1 0 8464 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_
timestamp 1608228718
transform 1 0 5336 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608228718
transform 1 0 6992 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_149
timestamp 1608228718
transform 1 0 6716 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_44
timestamp 1608228718
transform 1 0 5152 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_21_55
timestamp 1608228718
transform 1 0 6164 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_21_62
timestamp 1608228718
transform 1 0 6808 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_12_
timestamp 1608228718
transform 1 0 3680 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_21_26
timestamp 1608228718
transform 1 0 3496 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_11_
timestamp 1608228718
transform 1 0 2024 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5_
timestamp 1608228718
transform 1 0 1472 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1608228718
transform 1 0 1104 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_21_3
timestamp 1608228718
transform 1 0 1380 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_8
timestamp 1608228718
transform 1 0 1840 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_
timestamp 1608228718
transform 1 0 21712 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608228718
transform 1 0 21344 0 -1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1608228718
transform -1 0 23276 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1608228718
transform -1 0 23276 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_19_233
timestamp 1608228718
transform 1 0 22540 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_237
timestamp 1608228718
transform 1 0 22908 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_236
timestamp 1608228718
transform 1 0 22816 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _46_
timestamp 1608228718
transform 1 0 20884 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608228718
transform 1 0 20240 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_148
timestamp 1608228718
transform 1 0 20792 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_1_1_0_ltile_clb_mode__0.clb_clk
timestamp 1608228718
transform 1 0 19872 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1
timestamp 1608228718
transform 1 0 21160 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_202
timestamp 1608228718
transform 1 0 19688 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_19_207
timestamp 1608228718
transform 1 0 20148 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_212
timestamp 1608228718
transform 1 0 20608 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_4_
timestamp 1608228718
transform 1 0 18584 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_
timestamp 1608228718
transform 1 0 18032 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_
timestamp 1608228718
transform 1 0 18860 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608228718
transform 1 0 19136 0 -1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_144
timestamp 1608228718
transform 1 0 17940 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_181
timestamp 1608228718
transform 1 0 17756 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_188
timestamp 1608228718
transform 1 0 18400 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_194
timestamp 1608228718
transform 1 0 18952 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_13_
timestamp 1608228718
transform 1 0 15272 0 -1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_14_
timestamp 1608228718
transform 1 0 16284 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_16_
timestamp 1608228718
transform 1 0 16928 0 -1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_147
timestamp 1608228718
transform 1 0 15180 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_163
timestamp 1608228718
transform 1 0 16100 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_170
timestamp 1608228718
transform 1 0 16744 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_11_
timestamp 1608228718
transform 1 0 13524 0 -1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_12_
timestamp 1608228718
transform 1 0 14628 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_19_145
timestamp 1608228718
transform 1 0 14444 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_151
timestamp 1608228718
transform 1 0 14996 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6_
timestamp 1608228718
transform 1 0 11960 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_
timestamp 1608228718
transform 1 0 12420 0 1 12512
box -38 -48 498 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_16_
timestamp 1608228718
transform 1 0 12052 0 -1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_10_
timestamp 1608228718
transform 1 0 12972 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_143
timestamp 1608228718
transform 1 0 12328 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_116
timestamp 1608228718
transform 1 0 11776 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_19_128
timestamp 1608228718
transform 1 0 12880 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_
timestamp 1608228718
transform 1 0 9752 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_1_
timestamp 1608228718
transform 1 0 9936 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_14_
timestamp 1608228718
transform 1 0 10304 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_15_
timestamp 1608228718
transform 1 0 10580 0 -1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_146
timestamp 1608228718
transform 1 0 9568 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_1_0_0_ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
timestamp 1608228718
transform 1 0 9660 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_19_91
timestamp 1608228718
transform 1 0 9476 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_90
timestamp 1608228718
transform 1 0 9384 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_20_93
timestamp 1608228718
transform 1 0 9660 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_
timestamp 1608228718
transform 1 0 8648 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_2_
timestamp 1608228718
transform 1 0 9016 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_1_0_ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
timestamp 1608228718
transform 1 0 8740 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_19_80
timestamp 1608228718
transform 1 0 8464 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_81
timestamp 1608228718
transform 1 0 8556 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_4_
timestamp 1608228718
transform 1 0 6164 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608228718
transform 1 0 7084 0 -1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608228718
transform 1 0 6992 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_142
timestamp 1608228718
transform 1 0 6716 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_1_0_ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
timestamp 1608228718
transform 1 0 6440 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_19_55
timestamp 1608228718
transform 1 0 6164 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_19_62
timestamp 1608228718
transform 1 0 6808 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_53
timestamp 1608228718
transform 1 0 5980 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_20_59
timestamp 1608228718
transform 1 0 6532 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_14_
timestamp 1608228718
transform 1 0 4508 0 -1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_7_
timestamp 1608228718
transform 1 0 4692 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_19_36
timestamp 1608228718
transform 1 0 4416 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_20_35
timestamp 1608228718
transform 1 0 4324 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _59_
timestamp 1608228718
transform 1 0 4048 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_
timestamp 1608228718
transform 1 0 3588 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_3_
timestamp 1608228718
transform 1 0 3404 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_145
timestamp 1608228718
transform 1 0 3956 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_25
timestamp 1608228718
transform 1 0 3404 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_20_22
timestamp 1608228718
transform 1 0 3128 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_20_29
timestamp 1608228718
transform 1 0 3772 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_10_
timestamp 1608228718
transform 1 0 1656 0 -1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_8_
timestamp 1608228718
transform 1 0 1380 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_2_
timestamp 1608228718
transform 1 0 3036 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1608228718
transform 1 0 1104 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1608228718
transform 1 0 1104 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_19_19
timestamp 1608228718
transform 1 0 2852 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_20_3
timestamp 1608228718
transform 1 0 1380 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1608228718
transform -1 0 23276 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_18_232
timestamp 1608228718
transform 1 0 22448 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_
timestamp 1608228718
transform 1 0 19412 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608228718
transform 1 0 20976 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_141
timestamp 1608228718
transform 1 0 20792 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_197
timestamp 1608228718
transform 1 0 19228 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_18_208
timestamp 1608228718
transform 1 0 20240 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_215
timestamp 1608228718
transform 1 0 20884 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608228718
transform 1 0 17756 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_18_178
timestamp 1608228718
transform 1 0 17480 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_2_
timestamp 1608228718
transform 1 0 15456 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_15_
timestamp 1608228718
transform 1 0 16008 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_140
timestamp 1608228718
transform 1 0 15180 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_154
timestamp 1608228718
transform 1 0 15272 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_160
timestamp 1608228718
transform 1 0 15824 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_3_
timestamp 1608228718
transform 1 0 14720 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_8_
timestamp 1608228718
transform 1 0 13248 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_18_152
timestamp 1608228718
transform 1 0 15088 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
timestamp 1608228718
transform 1 0 11408 0 -1 12512
box -38 -48 1878 592
use sky130_fd_sc_hd__fill_2  FILLER_18_110
timestamp 1608228718
transform 1 0 11224 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_4_
timestamp 1608228718
transform 1 0 9660 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_139
timestamp 1608228718
transform 1 0 9568 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_3_0_ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
timestamp 1608228718
transform 1 0 10212 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_6_0_ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
timestamp 1608228718
transform 1 0 9200 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_12_0_ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
timestamp 1608228718
transform 1 0 10948 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_18_91
timestamp 1608228718
transform 1 0 9476 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_97
timestamp 1608228718
transform 1 0 10028 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_102
timestamp 1608228718
transform 1 0 10488 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_106
timestamp 1608228718
transform 1 0 10856 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_3_
timestamp 1608228718
transform 1 0 8648 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_80
timestamp 1608228718
transform 1 0 8464 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_86
timestamp 1608228718
transform 1 0 9016 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1608228718
transform 1 0 6992 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_
timestamp 1608228718
transform 1 0 6440 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_54
timestamp 1608228718
transform 1 0 6072 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_62
timestamp 1608228718
transform 1 0 6808 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_6_
timestamp 1608228718
transform 1 0 4600 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_
timestamp 1608228718
transform 1 0 4048 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_138
timestamp 1608228718
transform 1 0 3956 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_26
timestamp 1608228718
transform 1 0 3496 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_30
timestamp 1608228718
transform 1 0 3864 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_36
timestamp 1608228718
transform 1 0 4416 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_
timestamp 1608228718
transform 1 0 2668 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_
timestamp 1608228718
transform 1 0 1656 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1608228718
transform 1 0 1104 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_18_3
timestamp 1608228718
transform 1 0 1380 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_18_15
timestamp 1608228718
transform 1 0 2484 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_
timestamp 1608228718
transform 1 0 22264 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1608228718
transform -1 0 23276 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_17_228
timestamp 1608228718
transform 1 0 22080 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_234
timestamp 1608228718
transform 1 0 22632 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__sdfxtp_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_clb_fle_ff_0.sky130_fd_sc_hd__sdfxtp_1_0_
timestamp 1608228718
transform 1 0 20148 0 1 11424
box -38 -48 1970 592
use sky130_fd_sc_hd__decap_4  FILLER_17_202
timestamp 1608228718
transform 1 0 19688 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_206
timestamp 1608228718
transform 1 0 20056 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608228718
transform 1 0 18216 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_137
timestamp 1608228718
transform 1 0 17940 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_181
timestamp 1608228718
transform 1 0 17756 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_184
timestamp 1608228718
transform 1 0 18032 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.mux_fabric_out_1.mux_l2_in_0_
timestamp 1608228718
transform 1 0 16928 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_
timestamp 1608228718
transform 1 0 16284 0 1 11424
box -38 -48 498 592
use sky130_fd_sc_hd__decap_4  FILLER_17_161
timestamp 1608228718
transform 1 0 15916 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_170
timestamp 1608228718
transform 1 0 16744 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_9_
timestamp 1608228718
transform 1 0 14444 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_17_143
timestamp 1608228718
transform 1 0 14260 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _43_
timestamp 1608228718
transform 1 0 11868 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_7_
timestamp 1608228718
transform 1 0 12788 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_136
timestamp 1608228718
transform 1 0 12328 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_115
timestamp 1608228718
transform 1 0 11684 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_120
timestamp 1608228718
transform 1 0 12144 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_123
timestamp 1608228718
transform 1 0 12420 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5_
timestamp 1608228718
transform 1 0 9660 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_13_
timestamp 1608228718
transform 1 0 10212 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_17_89
timestamp 1608228718
transform 1 0 9292 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_97
timestamp 1608228718
transform 1 0 10028 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_
timestamp 1608228718
transform 1 0 8464 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_17_78
timestamp 1608228718
transform 1 0 8280 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_4_
timestamp 1608228718
transform 1 0 6808 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_0_
timestamp 1608228718
transform 1 0 6164 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_135
timestamp 1608228718
transform 1 0 6716 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_17_52
timestamp 1608228718
transform 1 0 5888 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_17_59
timestamp 1608228718
transform 1 0 6532 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_5_
timestamp 1608228718
transform 1 0 4416 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_0_0_ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
timestamp 1608228718
transform 1 0 4140 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_17_31
timestamp 1608228718
transform 1 0 3956 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0_
timestamp 1608228718
transform 1 0 1472 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608228718
transform 1 0 2484 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1608228718
transform 1 0 1104 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_17_3
timestamp 1608228718
transform 1 0 1380 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_13
timestamp 1608228718
transform 1 0 2300 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608228718
transform 1 0 21344 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1608228718
transform -1 0 23276 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_16_236
timestamp 1608228718
transform 1 0 22816 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _44_
timestamp 1608228718
transform 1 0 20884 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_134
timestamp 1608228718
transform 1 0 20792 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_209
timestamp 1608228718
transform 1 0 20332 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_213
timestamp 1608228718
transform 1 0 20700 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_218
timestamp 1608228718
transform 1 0 21160 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608228718
transform 1 0 18860 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608228718
transform 1 0 17204 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_16_191
timestamp 1608228718
transform 1 0 18676 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1608228718
transform 1 0 15548 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_133
timestamp 1608228718
transform 1 0 15180 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_16_154
timestamp 1608228718
transform 1 0 15272 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_16_173
timestamp 1608228718
transform 1 0 17020 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_
timestamp 1608228718
transform 1 0 14168 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_16_140
timestamp 1608228718
transform 1 0 13984 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_151
timestamp 1608228718
transform 1 0 14996 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_
timestamp 1608228718
transform 1 0 11592 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_5_
timestamp 1608228718
transform 1 0 12512 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_1_1_0_ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
timestamp 1608228718
transform 1 0 12236 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_16_112
timestamp 1608228718
transform 1 0 11408 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_16_118
timestamp 1608228718
transform 1 0 11960 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_12_
timestamp 1608228718
transform 1 0 9936 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_132
timestamp 1608228718
transform 1 0 9568 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_90
timestamp 1608228718
transform 1 0 9384 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_16_93
timestamp 1608228718
transform 1 0 9660 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_
timestamp 1608228718
transform 1 0 8556 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_16_79
timestamp 1608228718
transform 1 0 8372 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_
timestamp 1608228718
transform 1 0 5704 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_6_
timestamp 1608228718
transform 1 0 6900 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_16_48
timestamp 1608228718
transform 1 0 5520 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_59
timestamp 1608228718
transform 1 0 6532 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_4_
timestamp 1608228718
transform 1 0 4048 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_131
timestamp 1608228718
transform 1 0 3956 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_16_25
timestamp 1608228718
transform 1 0 3404 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608228718
transform 1 0 1932 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_3_
timestamp 1608228718
transform 1 0 1380 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1608228718
transform 1 0 1104 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_16_7
timestamp 1608228718
transform 1 0 1748 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.mux_fabric_out_1.mux_l2_in_0_
timestamp 1608228718
transform 1 0 21620 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1608228718
transform -1 0 23276 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_15_219
timestamp 1608228718
transform 1 0 21252 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_15_232
timestamp 1608228718
transform 1 0 22448 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__sdfxtp_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_clb_fle_ff_1.sky130_fd_sc_hd__sdfxtp_1_0_
timestamp 1608228718
transform 1 0 19320 0 1 10336
box -38 -48 1970 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.mux_fabric_out_1.mux_l1_in_0_
timestamp 1608228718
transform 1 0 18032 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_130
timestamp 1608228718
transform 1 0 17940 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_11_0_ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
timestamp 1608228718
transform 1 0 19044 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_15_181
timestamp 1608228718
transform 1 0 17756 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_193
timestamp 1608228718
transform 1 0 18860 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.mux_fabric_out_0.mux_l2_in_0_
timestamp 1608228718
transform 1 0 16928 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608228718
transform 1 0 15180 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_15_169
timestamp 1608228718
transform 1 0 16652 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.mux_ff_0_D_0.mux_l2_in_0_
timestamp 1608228718
transform 1 0 14168 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_15_139
timestamp 1608228718
transform 1 0 13892 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_15_151
timestamp 1608228718
transform 1 0 14996 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_
timestamp 1608228718
transform 1 0 11408 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_4_
timestamp 1608228718
transform 1 0 12420 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_129
timestamp 1608228718
transform 1 0 12328 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_110
timestamp 1608228718
transform 1 0 11224 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_15_116
timestamp 1608228718
transform 1 0 11776 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_11_
timestamp 1608228718
transform 1 0 9752 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_0_0_ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
timestamp 1608228718
transform 1 0 9476 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_15_89
timestamp 1608228718
transform 1 0 9292 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_
timestamp 1608228718
transform 1 0 8464 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_15_78
timestamp 1608228718
transform 1 0 8280 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_5_
timestamp 1608228718
transform 1 0 6808 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_1_
timestamp 1608228718
transform 1 0 6164 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_128
timestamp 1608228718
transform 1 0 6716 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_0_0_ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
timestamp 1608228718
transform 1 0 5888 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_15_49
timestamp 1608228718
transform 1 0 5612 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_15_59
timestamp 1608228718
transform 1 0 6532 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1_
timestamp 1608228718
transform 1 0 4784 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1608228718
transform 1 0 3128 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_15_38
timestamp 1608228718
transform 1 0 4600 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_
timestamp 1608228718
transform 1 0 1564 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2_
timestamp 1608228718
transform 1 0 2116 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1608228718
transform 1 0 1104 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_0
timestamp 1608228718
transform 1 0 1380 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_9
timestamp 1608228718
transform 1 0 1932 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_20
timestamp 1608228718
transform 1 0 2944 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _45_
timestamp 1608228718
transform 1 0 22540 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608228718
transform 1 0 21344 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1608228718
transform -1 0 23276 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1608228718
transform -1 0 23276 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_13_236
timestamp 1608228718
transform 1 0 22816 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_231
timestamp 1608228718
transform 1 0 22356 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_236
timestamp 1608228718
transform 1 0 22816 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.mux_ff_0_D_0.mux_l2_in_0_
timestamp 1608228718
transform 1 0 20148 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608228718
transform 1 0 20884 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_127
timestamp 1608228718
transform 1 0 20792 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_205
timestamp 1608228718
transform 1 0 19964 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_216
timestamp 1608228718
transform 1 0 20976 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_212
timestamp 1608228718
transform 1 0 20608 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _39_
timestamp 1608228718
transform 1 0 18676 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_clb_fle_ff_0.sky130_fd_sc_hd__sdfxtp_1_0_
timestamp 1608228718
transform 1 0 18032 0 1 9248
box -38 -48 1970 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608228718
transform 1 0 19136 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_123
timestamp 1608228718
transform 1 0 17940 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_5_0_ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
timestamp 1608228718
transform 1 0 17664 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_13_178
timestamp 1608228718
transform 1 0 17480 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_189
timestamp 1608228718
transform 1 0 18492 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_194
timestamp 1608228718
transform 1 0 18952 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_
timestamp 1608228718
transform 1 0 17112 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.mux_fabric_out_0.mux_l1_in_0_
timestamp 1608228718
transform 1 0 16100 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608228718
transform 1 0 15272 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608228718
transform 1 0 17020 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_126
timestamp 1608228718
transform 1 0 15180 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_161
timestamp 1608228718
transform 1 0 15916 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_172
timestamp 1608228718
transform 1 0 16928 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_14_170
timestamp 1608228718
transform 1 0 16744 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5_
timestamp 1608228718
transform 1 0 14352 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.mux_ff_0_D_0.mux_l1_in_0_
timestamp 1608228718
transform 1 0 13432 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608228718
transform 1 0 14444 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_2_0_ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
timestamp 1608228718
transform 1 0 14904 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_13_132
timestamp 1608228718
transform 1 0 13248 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_143
timestamp 1608228718
transform 1 0 14260 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_142
timestamp 1608228718
transform 1 0 14168 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_148
timestamp 1608228718
transform 1 0 14720 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_
timestamp 1608228718
transform 1 0 11316 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_
timestamp 1608228718
transform 1 0 12420 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0_
timestamp 1608228718
transform 1 0 11316 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_6_
timestamp 1608228718
transform 1 0 12696 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_122
timestamp 1608228718
transform 1 0 12328 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_9_0_ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
timestamp 1608228718
transform 1 0 12420 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_13_110
timestamp 1608228718
transform 1 0 11224 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_120
timestamp 1608228718
transform 1 0 12144 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_14_120
timestamp 1608228718
transform 1 0 12144 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_10_
timestamp 1608228718
transform 1 0 9660 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_9_
timestamp 1608228718
transform 1 0 9384 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_125
timestamp 1608228718
transform 1 0 9568 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_88
timestamp 1608228718
transform 1 0 9200 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_106
timestamp 1608228718
transform 1 0 10856 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_90
timestamp 1608228718
transform 1 0 9384 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_109
timestamp 1608228718
transform 1 0 11132 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_8_
timestamp 1608228718
transform 1 0 7728 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_
timestamp 1608228718
transform 1 0 9016 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_
timestamp 1608228718
transform 1 0 7176 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_70
timestamp 1608228718
transform 1 0 7544 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_81
timestamp 1608228718
transform 1 0 8556 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_85
timestamp 1608228718
transform 1 0 8924 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_7_
timestamp 1608228718
transform 1 0 7084 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_121
timestamp 1608228718
transform 1 0 6716 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_59
timestamp 1608228718
transform 1 0 6532 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_62
timestamp 1608228718
transform 1 0 6808 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_63
timestamp 1608228718
transform 1 0 6900 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0_
timestamp 1608228718
transform 1 0 6072 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.mux_fabric_out_1.mux_l2_in_0_
timestamp 1608228718
transform 1 0 5704 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_2
timestamp 1608228718
transform 1 0 5520 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_46
timestamp 1608228718
transform 1 0 5336 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_52
timestamp 1608228718
transform 1 0 5888 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_
timestamp 1608228718
transform 1 0 3128 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.mux_ff_0_D_0.mux_l1_in_0_
timestamp 1608228718
transform 1 0 5060 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_
timestamp 1608228718
transform 1 0 4048 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_
timestamp 1608228718
transform 1 0 4508 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_
timestamp 1608228718
transform 1 0 3680 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_124
timestamp 1608228718
transform 1 0 3956 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_26
timestamp 1608228718
transform 1 0 3496 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_29
timestamp 1608228718
transform 1 0 3772 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_41
timestamp 1608228718
transform 1 0 4876 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608228718
transform 1 0 1380 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_
timestamp 1608228718
transform 1 0 2392 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0_
timestamp 1608228718
transform 1 0 2944 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_13_19
timestamp 1608228718
transform 1 0 2852 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_14_12
timestamp 1608228718
transform 1 0 2208 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_18
timestamp 1608228718
transform 1 0 2760 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_0_
timestamp 1608228718
transform 1 0 1840 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1608228718
transform 1 0 1104 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1608228718
transform 1 0 1104 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_14_3
timestamp 1608228718
transform 1 0 1380 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_7
timestamp 1608228718
transform 1 0 1748 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.mux_fabric_out_1.mux_l1_in_0_
timestamp 1608228718
transform 1 0 21896 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1608228718
transform -1 0 23276 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_12_224
timestamp 1608228718
transform 1 0 21712 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_12_235
timestamp 1608228718
transform 1 0 22724 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.mux_fabric_out_0.mux_l1_in_0_
timestamp 1608228718
transform 1 0 20884 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_120
timestamp 1608228718
transform 1 0 20792 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_12_208
timestamp 1608228718
transform 1 0 20240 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608228718
transform 1 0 18768 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_12_188
timestamp 1608228718
transform 1 0 18400 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_
timestamp 1608228718
transform 1 0 16284 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0_
timestamp 1608228718
transform 1 0 15272 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608228718
transform 1 0 16928 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_119
timestamp 1608228718
transform 1 0 15180 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_163
timestamp 1608228718
transform 1 0 16100 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_12_169
timestamp 1608228718
transform 1 0 16652 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608228718
transform 1 0 13524 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_12_133
timestamp 1608228718
transform 1 0 13340 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_151
timestamp 1608228718
transform 1 0 14996 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6_
timestamp 1608228718
transform 1 0 12972 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608228718
transform 1 0 11224 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_12_126
timestamp 1608228718
transform 1 0 12696 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2_
timestamp 1608228718
transform 1 0 9660 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_1_
timestamp 1608228718
transform 1 0 10672 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_118
timestamp 1608228718
transform 1 0 9568 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_90
timestamp 1608228718
transform 1 0 9384 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_102
timestamp 1608228718
transform 1 0 10488 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_108
timestamp 1608228718
transform 1 0 11040 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1_
timestamp 1608228718
transform 1 0 7728 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_4_
timestamp 1608228718
transform 1 0 9016 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_1_0_ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
timestamp 1608228718
transform 1 0 8740 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_12_70
timestamp 1608228718
transform 1 0 7544 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_81
timestamp 1608228718
transform 1 0 8556 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.mux_fabric_out_0.mux_l1_in_0_
timestamp 1608228718
transform 1 0 6716 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.mux_ff_0_D_0.mux_l2_in_0_
timestamp 1608228718
transform 1 0 5704 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_12_48
timestamp 1608228718
transform 1 0 5520 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_59
timestamp 1608228718
transform 1 0 6532 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6_
timestamp 1608228718
transform 1 0 4140 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_
timestamp 1608228718
transform 1 0 4692 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_
timestamp 1608228718
transform 1 0 3404 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_117
timestamp 1608228718
transform 1 0 3956 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_23
timestamp 1608228718
transform 1 0 3220 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_29
timestamp 1608228718
transform 1 0 3772 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_12_32
timestamp 1608228718
transform 1 0 4048 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_37
timestamp 1608228718
transform 1 0 4508 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _62_
timestamp 1608228718
transform 1 0 2944 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1608228718
transform 1 0 1104 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_12_3
timestamp 1608228718
transform 1 0 1380 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_12_15
timestamp 1608228718
transform 1 0 2484 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_19
timestamp 1608228718
transform 1 0 2852 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.mux_fabric_out_0.mux_l2_in_0_
timestamp 1608228718
transform 1 0 21988 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1608228718
transform -1 0 23276 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_11_225
timestamp 1608228718
transform 1 0 21804 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_236
timestamp 1608228718
transform 1 0 22816 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__sdfxtp_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_clb_fle_ff_1.sky130_fd_sc_hd__sdfxtp_1_0_
timestamp 1608228718
transform 1 0 19872 0 1 8160
box -38 -48 1970 592
use sky130_fd_sc_hd__fill_2  FILLER_11_202
timestamp 1608228718
transform 1 0 19688 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0_
timestamp 1608228718
transform 1 0 18860 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  prog_clk_0_N_FTB01
timestamp 1608228718
transform 1 0 18124 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_116
timestamp 1608228718
transform 1 0 17940 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_181
timestamp 1608228718
transform 1 0 17756 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_11_184
timestamp 1608228718
transform 1 0 18032 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_191
timestamp 1608228718
transform 1 0 18676 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__sdfxtp_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_clb_fle_ff_1.sky130_fd_sc_hd__sdfxtp_1_0_
timestamp 1608228718
transform 1 0 15824 0 1 8160
box -38 -48 1970 592
use sky130_fd_sc_hd__decap_3  FILLER_11_157
timestamp 1608228718
transform 1 0 15548 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608228718
transform 1 0 14076 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_11_139
timestamp 1608228718
transform 1 0 13892 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1608228718
transform 1 0 12420 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_115
timestamp 1608228718
transform 1 0 12328 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_120
timestamp 1608228718
transform 1 0 12144 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_3_
timestamp 1608228718
transform 1 0 10120 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608228718
transform 1 0 10672 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_11_95
timestamp 1608228718
transform 1 0 9844 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_11_102
timestamp 1608228718
transform 1 0 10488 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1_
timestamp 1608228718
transform 1 0 7360 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_4_
timestamp 1608228718
transform 1 0 8372 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_11_66
timestamp 1608228718
transform 1 0 7176 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_77
timestamp 1608228718
transform 1 0 8188 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_
timestamp 1608228718
transform 1 0 6808 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3_
timestamp 1608228718
transform 1 0 5704 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_114
timestamp 1608228718
transform 1 0 6716 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_48
timestamp 1608228718
transform 1 0 5520 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_59
timestamp 1608228718
transform 1 0 6532 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6_
timestamp 1608228718
transform 1 0 4140 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.mux_ff_0_D_0.mux_l2_in_0_
timestamp 1608228718
transform 1 0 4692 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_11_25
timestamp 1608228718
transform 1 0 3404 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_11_37
timestamp 1608228718
transform 1 0 4508 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  Test_en_W_FTB01
timestamp 1608228718
transform 1 0 1748 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1608228718
transform 1 0 1104 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_11_3
timestamp 1608228718
transform 1 0 1380 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_11_13
timestamp 1608228718
transform 1 0 2300 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608228718
transform 1 0 21252 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1608228718
transform -1 0 23276 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_235
timestamp 1608228718
transform 1 0 22724 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_113
timestamp 1608228718
transform 1 0 20792 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_10_211
timestamp 1608228718
transform 1 0 20516 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_10_215
timestamp 1608228718
transform 1 0 20884 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__sdfxtp_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_clb_fle_ff_0.sky130_fd_sc_hd__sdfxtp_1_0_
timestamp 1608228718
transform 1 0 18584 0 -1 8160
box -38 -48 1970 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.mux_ff_0_D_0.mux_l1_in_0_
timestamp 1608228718
transform 1 0 17572 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_10_175
timestamp 1608228718
transform 1 0 17204 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_10_188
timestamp 1608228718
transform 1 0 18400 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__sdfxtp_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_clb_fle_ff_0.sky130_fd_sc_hd__sdfxtp_1_0_
timestamp 1608228718
transform 1 0 15272 0 -1 8160
box -38 -48 1970 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_112
timestamp 1608228718
transform 1 0 15180 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_
timestamp 1608228718
transform 1 0 13800 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_4_0_ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
timestamp 1608228718
transform 1 0 14812 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_10_136
timestamp 1608228718
transform 1 0 13616 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_147
timestamp 1608228718
transform 1 0 14628 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_10_152
timestamp 1608228718
transform 1 0 15088 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_
timestamp 1608228718
transform 1 0 12788 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_10_125
timestamp 1608228718
transform 1 0 12604 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _42_
timestamp 1608228718
transform 1 0 10672 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_
timestamp 1608228718
transform 1 0 9660 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608228718
transform 1 0 11132 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_111
timestamp 1608228718
transform 1 0 9568 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_90
timestamp 1608228718
transform 1 0 9384 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_102
timestamp 1608228718
transform 1 0 10488 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_107
timestamp 1608228718
transform 1 0 10948 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_6_
timestamp 1608228718
transform 1 0 7912 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_10_72
timestamp 1608228718
transform 1 0 7728 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__buf_8  Test_en_FTB00
timestamp 1608228718
transform 1 0 6624 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.mux_fabric_out_1.mux_l2_in_0_
timestamp 1608228718
transform 1 0 5612 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_6
timestamp 1608228718
transform 1 0 5428 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_45
timestamp 1608228718
transform 1 0 5244 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_58
timestamp 1608228718
transform 1 0 6440 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _60_
timestamp 1608228718
transform 1 0 4600 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5_
timestamp 1608228718
transform 1 0 4876 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_110
timestamp 1608228718
transform 1 0 3956 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_27
timestamp 1608228718
transform 1 0 3588 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_10_32
timestamp 1608228718
transform 1 0 4048 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1608228718
transform 1 0 1104 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_10_3
timestamp 1608228718
transform 1 0 1380 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_15
timestamp 1608228718
transform 1 0 2484 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1608228718
transform -1 0 23276 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_9_234
timestamp 1608228718
transform 1 0 22632 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608228718
transform 1 0 21160 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_4  prog_clk_0_E_FTB01
timestamp 1608228718
transform 1 0 20424 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_9_208
timestamp 1608228718
transform 1 0 20240 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_216
timestamp 1608228718
transform 1 0 20976 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_1_
timestamp 1608228718
transform 1 0 18216 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608228718
transform 1 0 18768 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_109
timestamp 1608228718
transform 1 0 17940 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_181
timestamp 1608228718
transform 1 0 17756 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_184
timestamp 1608228718
transform 1 0 18032 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_190
timestamp 1608228718
transform 1 0 18584 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608228718
transform 1 0 16284 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_8_0_ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
timestamp 1608228718
transform 1 0 15916 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_9_159
timestamp 1608228718
transform 1 0 15732 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_9_164
timestamp 1608228718
transform 1 0 16192 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_
timestamp 1608228718
transform 1 0 13708 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608228718
transform 1 0 14260 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_10_0_ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
timestamp 1608228718
transform 1 0 13432 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_9_132
timestamp 1608228718
transform 1 0 13248 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_141
timestamp 1608228718
transform 1 0 14076 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _41_
timestamp 1608228718
transform 1 0 11868 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3_
timestamp 1608228718
transform 1 0 12420 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_108
timestamp 1608228718
transform 1 0 12328 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_115
timestamp 1608228718
transform 1 0 11684 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_120
timestamp 1608228718
transform 1 0 12144 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_7_
timestamp 1608228718
transform 1 0 10212 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_9_97
timestamp 1608228718
transform 1 0 10028 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_5_
timestamp 1608228718
transform 1 0 8556 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1_
timestamp 1608228718
transform 1 0 7544 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_9_68
timestamp 1608228718
transform 1 0 7360 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_79
timestamp 1608228718
transform 1 0 8372 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_4_
timestamp 1608228718
transform 1 0 6992 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_3_
timestamp 1608228718
transform 1 0 6164 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_
timestamp 1608228718
transform 1 0 5612 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_107
timestamp 1608228718
transform 1 0 6716 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_47
timestamp 1608228718
transform 1 0 5428 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_53
timestamp 1608228718
transform 1 0 5980 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_59
timestamp 1608228718
transform 1 0 6532 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_62
timestamp 1608228718
transform 1 0 6808 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_9_27
timestamp 1608228718
transform 1 0 3588 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_39
timestamp 1608228718
transform 1 0 4692 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1608228718
transform 1 0 1104 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_9_3
timestamp 1608228718
transform 1 0 1380 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_15
timestamp 1608228718
transform 1 0 2484 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _37_
timestamp 1608228718
transform 1 0 22540 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1608228718
transform -1 0 23276 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_8_231
timestamp 1608228718
transform 1 0 22356 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_236
timestamp 1608228718
transform 1 0 22816 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_
timestamp 1608228718
transform 1 0 19780 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608228718
transform 1 0 20884 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_106
timestamp 1608228718
transform 1 0 20792 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_201
timestamp 1608228718
transform 1 0 19596 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_212
timestamp 1608228718
transform 1 0 20608 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0_
timestamp 1608228718
transform 1 0 18768 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_8_188
timestamp 1608228718
transform 1 0 18400 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608228718
transform 1 0 15272 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608228718
transform 1 0 16928 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_105
timestamp 1608228718
transform 1 0 15180 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_170
timestamp 1608228718
transform 1 0 16744 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_
timestamp 1608228718
transform 1 0 13340 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_
timestamp 1608228718
transform 1 0 14352 0 -1 7072
box -38 -48 498 592
use sky130_fd_sc_hd__fill_2  FILLER_8_142
timestamp 1608228718
transform 1 0 14168 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_149
timestamp 1608228718
transform 1 0 14812 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_
timestamp 1608228718
transform 1 0 11316 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_
timestamp 1608228718
transform 1 0 12328 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_8_120
timestamp 1608228718
transform 1 0 12144 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_131
timestamp 1608228718
transform 1 0 13156 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_9_
timestamp 1608228718
transform 1 0 9660 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_104
timestamp 1608228718
transform 1 0 9568 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_90
timestamp 1608228718
transform 1 0 9384 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_109
timestamp 1608228718
transform 1 0 11132 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_
timestamp 1608228718
transform 1 0 8556 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.mux_fabric_out_0.mux_l2_in_0_
timestamp 1608228718
transform 1 0 7544 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_4
timestamp 1608228718
transform 1 0 7360 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_66
timestamp 1608228718
transform 1 0 7176 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_79
timestamp 1608228718
transform 1 0 8372 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_1_
timestamp 1608228718
transform 1 0 6808 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_
timestamp 1608228718
transform 1 0 6440 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_8_44
timestamp 1608228718
transform 1 0 5152 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_8_56
timestamp 1608228718
transform 1 0 6256 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_103
timestamp 1608228718
transform 1 0 3956 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_27
timestamp 1608228718
transform 1 0 3588 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_8_32
timestamp 1608228718
transform 1 0 4048 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1608228718
transform 1 0 1104 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_8_3
timestamp 1608228718
transform 1 0 1380 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_15
timestamp 1608228718
transform 1 0 2484 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_4  Test_en_E_FTB01
timestamp 1608228718
transform 1 0 22264 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__conb_1  _38_
timestamp 1608228718
transform 1 0 22540 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1608228718
transform -1 0 23276 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1608228718
transform -1 0 23276 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_6_236
timestamp 1608228718
transform 1 0 22816 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_231
timestamp 1608228718
transform 1 0 22356 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_236
timestamp 1608228718
transform 1 0 22816 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_
timestamp 1608228718
transform 1 0 21252 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_
timestamp 1608228718
transform 1 0 21528 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_6_228
timestamp 1608228718
transform 1 0 22080 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608228718
transform 1 0 19504 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_99
timestamp 1608228718
transform 1 0 20792 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_6_208
timestamp 1608228718
transform 1 0 20240 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_6_215
timestamp 1608228718
transform 1 0 20884 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_198
timestamp 1608228718
transform 1 0 19320 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_7_216
timestamp 1608228718
transform 1 0 20976 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__conb_1  _36_
timestamp 1608228718
transform 1 0 18032 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_
timestamp 1608228718
transform 1 0 17756 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_
timestamp 1608228718
transform 1 0 18492 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608228718
transform 1 0 18768 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_102
timestamp 1608228718
transform 1 0 17940 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_179
timestamp 1608228718
transform 1 0 17572 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_190
timestamp 1608228718
transform 1 0 18584 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_181
timestamp 1608228718
transform 1 0 17756 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_187
timestamp 1608228718
transform 1 0 18308 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_3_
timestamp 1608228718
transform 1 0 16376 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6_
timestamp 1608228718
transform 1 0 15548 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608228718
transform 1 0 16100 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_
timestamp 1608228718
transform 1 0 16928 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_98
timestamp 1608228718
transform 1 0 15180 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_6_154
timestamp 1608228718
transform 1 0 15272 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_6_161
timestamp 1608228718
transform 1 0 15916 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_162
timestamp 1608228718
transform 1 0 16008 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_170
timestamp 1608228718
transform 1 0 16744 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_
timestamp 1608228718
transform 1 0 14628 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608228718
transform 1 0 14536 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_6_145
timestamp 1608228718
transform 1 0 14444 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_151
timestamp 1608228718
transform 1 0 14996 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_144
timestamp 1608228718
transform 1 0 14352 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_12_
timestamp 1608228718
transform 1 0 11316 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_15_
timestamp 1608228718
transform 1 0 12972 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_16_
timestamp 1608228718
transform 1 0 12880 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _40_
timestamp 1608228718
transform 1 0 12420 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_101
timestamp 1608228718
transform 1 0 12328 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_127
timestamp 1608228718
transform 1 0 12788 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_126
timestamp 1608228718
transform 1 0 12696 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_
timestamp 1608228718
transform 1 0 11776 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_2_0_ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
timestamp 1608228718
transform 1 0 11408 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_7_110
timestamp 1608228718
transform 1 0 11224 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_7_115
timestamp 1608228718
transform 1 0 11684 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_120
timestamp 1608228718
transform 1 0 12144 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_
timestamp 1608228718
transform 1 0 10396 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_10_
timestamp 1608228718
transform 1 0 9660 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_97
timestamp 1608228718
transform 1 0 9568 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_90
timestamp 1608228718
transform 1 0 9384 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_109
timestamp 1608228718
transform 1 0 11132 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_99
timestamp 1608228718
transform 1 0 10212 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_8_
timestamp 1608228718
transform 1 0 8740 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_
timestamp 1608228718
transform 1 0 8188 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.mux_ff_0_D_0.mux_l1_in_0_
timestamp 1608228718
transform 1 0 8556 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_6_79
timestamp 1608228718
transform 1 0 8372 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_81
timestamp 1608228718
transform 1 0 8556 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _63_
timestamp 1608228718
transform 1 0 8096 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_
timestamp 1608228718
transform 1 0 7636 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_6_68
timestamp 1608228718
transform 1 0 7360 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_7_70
timestamp 1608228718
transform 1 0 7544 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_75
timestamp 1608228718
transform 1 0 8004 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_100
timestamp 1608228718
transform 1 0 6716 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_44
timestamp 1608228718
transform 1 0 5152 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_56
timestamp 1608228718
transform 1 0 6256 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_51
timestamp 1608228718
transform 1 0 5796 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_7_59
timestamp 1608228718
transform 1 0 6532 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_7_62
timestamp 1608228718
transform 1 0 6808 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_96
timestamp 1608228718
transform 1 0 3956 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_27
timestamp 1608228718
transform 1 0 3588 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_6_32
timestamp 1608228718
transform 1 0 4048 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_27
timestamp 1608228718
transform 1 0 3588 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_39
timestamp 1608228718
transform 1 0 4692 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1608228718
transform 1 0 1104 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1608228718
transform 1 0 1104 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_6_3
timestamp 1608228718
transform 1 0 1380 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_15
timestamp 1608228718
transform 1 0 2484 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_3
timestamp 1608228718
transform 1 0 1380 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_15
timestamp 1608228718
transform 1 0 2484 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608228718
transform 1 0 21344 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1608228718
transform -1 0 23276 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_5_236
timestamp 1608228718
transform 1 0 22816 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2_
timestamp 1608228718
transform 1 0 19228 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3_
timestamp 1608228718
transform 1 0 20332 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_5_206
timestamp 1608228718
transform 1 0 20056 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_5_218
timestamp 1608228718
transform 1 0 21160 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0_
timestamp 1608228718
transform 1 0 18032 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_95
timestamp 1608228718
transform 1 0 17940 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_181
timestamp 1608228718
transform 1 0 17756 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_193
timestamp 1608228718
transform 1 0 18860 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608228718
transform 1 0 16284 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_5_161
timestamp 1608228718
transform 1 0 15916 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0_
timestamp 1608228718
transform 1 0 14076 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_
timestamp 1608228718
transform 1 0 15088 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_5_139
timestamp 1608228718
transform 1 0 13892 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_150
timestamp 1608228718
transform 1 0 14904 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_
timestamp 1608228718
transform 1 0 11776 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_14_
timestamp 1608228718
transform 1 0 12420 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_94
timestamp 1608228718
transform 1 0 12328 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_112
timestamp 1608228718
transform 1 0 11408 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_5_120
timestamp 1608228718
transform 1 0 12144 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5_
timestamp 1608228718
transform 1 0 9384 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_11_
timestamp 1608228718
transform 1 0 9936 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_5_88
timestamp 1608228718
transform 1 0 9200 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_94
timestamp 1608228718
transform 1 0 9752 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _61_
timestamp 1608228718
transform 1 0 8924 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_5_74
timestamp 1608228718
transform 1 0 7912 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_5_82
timestamp 1608228718
transform 1 0 8648 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_93
timestamp 1608228718
transform 1 0 6716 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_5_51
timestamp 1608228718
transform 1 0 5796 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_5_59
timestamp 1608228718
transform 1 0 6532 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_5_62
timestamp 1608228718
transform 1 0 6808 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_27
timestamp 1608228718
transform 1 0 3588 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_39
timestamp 1608228718
transform 1 0 4692 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1608228718
transform 1 0 1104 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_5_3
timestamp 1608228718
transform 1 0 1380 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_15
timestamp 1608228718
transform 1 0 2484 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_16_
timestamp 1608228718
transform 1 0 21344 0 -1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1608228718
transform -1 0 23276 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_4_236
timestamp 1608228718
transform 1 0 22816 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _51_
timestamp 1608228718
transform 1 0 20884 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_
timestamp 1608228718
transform 1 0 19688 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_92
timestamp 1608228718
transform 1 0 20792 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_198
timestamp 1608228718
transform 1 0 19320 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_4_211
timestamp 1608228718
transform 1 0 20516 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_4_218
timestamp 1608228718
transform 1 0 21160 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_
timestamp 1608228718
transform 1 0 17480 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_
timestamp 1608228718
transform 1 0 18492 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_4_176
timestamp 1608228718
transform 1 0 17296 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_187
timestamp 1608228718
transform 1 0 18308 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_4_
timestamp 1608228718
transform 1 0 15272 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608228718
transform 1 0 15824 0 -1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_91
timestamp 1608228718
transform 1 0 15180 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_158
timestamp 1608228718
transform 1 0 15640 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1_
timestamp 1608228718
transform 1 0 13984 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_4_138
timestamp 1608228718
transform 1 0 13800 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_149
timestamp 1608228718
transform 1 0 14812 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_
timestamp 1608228718
transform 1 0 12972 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_13_
timestamp 1608228718
transform 1 0 11316 0 -1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_4_127
timestamp 1608228718
transform 1 0 12788 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2_
timestamp 1608228718
transform 1 0 10120 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_90
timestamp 1608228718
transform 1 0 9568 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_93
timestamp 1608228718
transform 1 0 9660 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_97
timestamp 1608228718
transform 1 0 10028 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_107
timestamp 1608228718
transform 1 0 10948 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_4_68
timestamp 1608228718
transform 1 0 7360 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_80
timestamp 1608228718
transform 1 0 8464 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_44
timestamp 1608228718
transform 1 0 5152 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_56
timestamp 1608228718
transform 1 0 6256 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_89
timestamp 1608228718
transform 1 0 3956 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_27
timestamp 1608228718
transform 1 0 3588 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_4_32
timestamp 1608228718
transform 1 0 4048 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1608228718
transform 1 0 1104 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_4_3
timestamp 1608228718
transform 1 0 1380 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_15
timestamp 1608228718
transform 1 0 2484 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_15_
timestamp 1608228718
transform 1 0 21344 0 1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1608228718
transform -1 0 23276 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_3_236
timestamp 1608228718
transform 1 0 22816 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_
timestamp 1608228718
transform 1 0 19688 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_
timestamp 1608228718
transform 1 0 20700 0 1 3808
box -38 -48 498 592
use sky130_fd_sc_hd__fill_2  FILLER_3_200
timestamp 1608228718
transform 1 0 19504 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_211
timestamp 1608228718
transform 1 0 20516 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_218
timestamp 1608228718
transform 1 0 21160 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_0_
timestamp 1608228718
transform 1 0 17388 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_8_
timestamp 1608228718
transform 1 0 18032 0 1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_88
timestamp 1608228718
transform 1 0 17940 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_175
timestamp 1608228718
transform 1 0 17204 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_181
timestamp 1608228718
transform 1 0 17756 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1608228718
transform 1 0 15732 0 1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_3_157
timestamp 1608228718
transform 1 0 15548 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1_
timestamp 1608228718
transform 1 0 14720 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_
timestamp 1608228718
transform 1 0 13708 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_3_135
timestamp 1608228718
transform 1 0 13524 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_146
timestamp 1608228718
transform 1 0 14536 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0_
timestamp 1608228718
transform 1 0 12696 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.mux_fabric_out_1.mux_l1_in_0_
timestamp 1608228718
transform 1 0 11316 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_87
timestamp 1608228718
transform 1 0 12328 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_120
timestamp 1608228718
transform 1 0 12144 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_3_123
timestamp 1608228718
transform 1 0 12420 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_
timestamp 1608228718
transform 1 0 10764 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_3_98
timestamp 1608228718
transform 1 0 10120 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_104
timestamp 1608228718
transform 1 0 10672 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_109
timestamp 1608228718
transform 1 0 11132 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_3_74
timestamp 1608228718
transform 1 0 7912 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_86
timestamp 1608228718
transform 1 0 9016 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_86
timestamp 1608228718
transform 1 0 6716 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_3_51
timestamp 1608228718
transform 1 0 5796 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_3_59
timestamp 1608228718
transform 1 0 6532 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_3_62
timestamp 1608228718
transform 1 0 6808 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_27
timestamp 1608228718
transform 1 0 3588 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_39
timestamp 1608228718
transform 1 0 4692 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1608228718
transform 1 0 1104 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_3_3
timestamp 1608228718
transform 1 0 1380 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_15
timestamp 1608228718
transform 1 0 2484 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1608228718
transform -1 0 23276 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_2_231
timestamp 1608228718
transform 1 0 22356 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_237
timestamp 1608228718
transform 1 0 22908 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_13_
timestamp 1608228718
transform 1 0 20884 0 -1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_85
timestamp 1608228718
transform 1 0 20792 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_212
timestamp 1608228718
transform 1 0 20608 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_7_
timestamp 1608228718
transform 1 0 17480 0 -1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_9_
timestamp 1608228718
transform 1 0 19136 0 -1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_2_176
timestamp 1608228718
transform 1 0 17296 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_194
timestamp 1608228718
transform 1 0 18952 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5_
timestamp 1608228718
transform 1 0 15272 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_4_
timestamp 1608228718
transform 1 0 15824 0 -1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_84
timestamp 1608228718
transform 1 0 15180 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_158
timestamp 1608228718
transform 1 0 15640 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_
timestamp 1608228718
transform 1 0 14168 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_2_140
timestamp 1608228718
transform 1 0 13984 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_151
timestamp 1608228718
transform 1 0 14996 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_2_
timestamp 1608228718
transform 1 0 12604 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6_
timestamp 1608228718
transform 1 0 11960 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0_
timestamp 1608228718
transform 1 0 13156 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_2_117
timestamp 1608228718
transform 1 0 11868 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_2_122
timestamp 1608228718
transform 1 0 12328 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_2_129
timestamp 1608228718
transform 1 0 12972 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_83
timestamp 1608228718
transform 1 0 9568 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_93
timestamp 1608228718
transform 1 0 9660 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_105
timestamp 1608228718
transform 1 0 10764 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_68
timestamp 1608228718
transform 1 0 7360 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_80
timestamp 1608228718
transform 1 0 8464 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_44
timestamp 1608228718
transform 1 0 5152 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_56
timestamp 1608228718
transform 1 0 6256 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_82
timestamp 1608228718
transform 1 0 3956 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_26
timestamp 1608228718
transform 1 0 3496 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_30
timestamp 1608228718
transform 1 0 3864 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_32
timestamp 1608228718
transform 1 0 4048 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  prog_clk_0_FTB00
timestamp 1608228718
transform 1 0 2392 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1608228718
transform 1 0 1104 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_2_3
timestamp 1608228718
transform 1 0 1380 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_2_11
timestamp 1608228718
transform 1 0 2116 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  prog_clk_0_S_FTB01
timestamp 1608228718
transform 1 0 22172 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1608228718
transform -1 0 23276 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1608228718
transform -1 0 23276 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_234
timestamp 1608228718
transform 1 0 22632 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_227
timestamp 1608228718
transform 1 0 21988 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_1_235
timestamp 1608228718
transform 1 0 22724 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_11_
timestamp 1608228718
transform 1 0 19320 0 -1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_12_
timestamp 1608228718
transform 1 0 20516 0 1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_14_
timestamp 1608228718
transform 1 0 21160 0 -1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_78
timestamp 1608228718
transform 1 0 21068 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_214
timestamp 1608228718
transform 1 0 20792 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_1_209
timestamp 1608228718
transform 1 0 20332 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_10_
timestamp 1608228718
transform 1 0 18860 0 1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_
timestamp 1608228718
transform 1 0 18308 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_2_
timestamp 1608228718
transform 1 0 18308 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_77
timestamp 1608228718
transform 1 0 18216 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_196
timestamp 1608228718
transform 1 0 19136 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_191
timestamp 1608228718
transform 1 0 18676 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_81
timestamp 1608228718
transform 1 0 17940 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_183
timestamp 1608228718
transform 1 0 17940 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_1_178
timestamp 1608228718
transform 1 0 17480 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_182
timestamp 1608228718
transform 1 0 17848 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_1_184
timestamp 1608228718
transform 1 0 18032 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_5_
timestamp 1608228718
transform 1 0 16008 0 1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_6_
timestamp 1608228718
transform 1 0 16468 0 -1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_
timestamp 1608228718
transform 1 0 15456 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_76
timestamp 1608228718
transform 1 0 15364 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_153
timestamp 1608228718
transform 1 0 15180 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_165
timestamp 1608228718
transform 1 0 16284 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_160
timestamp 1608228718
transform 1 0 15824 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_
timestamp 1608228718
transform 1 0 14996 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.mux_fabric_out_0.mux_l1_in_0_
timestamp 1608228718
transform 1 0 14352 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_0_142
timestamp 1608228718
transform 1 0 14168 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_149
timestamp 1608228718
transform 1 0 14812 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_0_
timestamp 1608228718
transform 1 0 13432 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_2_
timestamp 1608228718
transform 1 0 13800 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_
timestamp 1608228718
transform 1 0 13984 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_0_137
timestamp 1608228718
transform 1 0 13708 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_132
timestamp 1608228718
transform 1 0 13248 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_138
timestamp 1608228718
transform 1 0 13800 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_4_
timestamp 1608228718
transform 1 0 12880 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_75
timestamp 1608228718
transform 1 0 12512 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_80
timestamp 1608228718
transform 1 0 12328 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_118
timestamp 1608228718
transform 1 0 11960 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_0_125
timestamp 1608228718
transform 1 0 12604 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_110
timestamp 1608228718
transform 1 0 11224 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_123
timestamp 1608228718
transform 1 0 12420 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_127
timestamp 1608228718
transform 1 0 12788 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_74
timestamp 1608228718
transform 1 0 9660 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_0_94
timestamp 1608228718
transform 1 0 9752 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_106
timestamp 1608228718
transform 1 0 10856 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_98
timestamp 1608228718
transform 1 0 10120 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_75
timestamp 1608228718
transform 1 0 8004 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_87
timestamp 1608228718
transform 1 0 9108 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_1_74
timestamp 1608228718
transform 1 0 7912 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_86
timestamp 1608228718
transform 1 0 9016 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_73
timestamp 1608228718
transform 1 0 6808 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_79
timestamp 1608228718
transform 1 0 6716 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_0_44
timestamp 1608228718
transform 1 0 5152 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_56
timestamp 1608228718
transform 1 0 6256 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_0_63
timestamp 1608228718
transform 1 0 6900 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_44
timestamp 1608228718
transform 1 0 5152 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_56
timestamp 1608228718
transform 1 0 6256 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_60
timestamp 1608228718
transform 1 0 6624 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_62
timestamp 1608228718
transform 1 0 6808 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _64_
timestamp 1608228718
transform 1 0 4876 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_72
timestamp 1608228718
transform 1 0 3956 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27
timestamp 1608228718
transform 1 0 3588 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_0_32
timestamp 1608228718
transform 1 0 4048 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_31
timestamp 1608228718
transform 1 0 3956 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_39
timestamp 1608228718
transform 1 0 4692 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _66_
timestamp 1608228718
transform 1 0 2484 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  prog_clk_0_W_FTB01
timestamp 1608228718
transform 1 0 1748 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1608228718
transform 1 0 1104 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1608228718
transform 1 0 1104 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_0_3
timestamp 1608228718
transform 1 0 1380 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_15
timestamp 1608228718
transform 1 0 2484 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_3
timestamp 1608228718
transform 1 0 1380 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_13
timestamp 1608228718
transform 1 0 2300 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_1_19
timestamp 1608228718
transform 1 0 2852 0 1 2720
box -38 -48 1142 592
<< labels >>
rlabel metal2 s 8574 0 8630 800 4 SC_IN_BOT
port 1 nsew
rlabel metal2 s 16946 23600 17002 24400 4 SC_IN_TOP
port 2 nsew
rlabel metal2 s 12070 0 12126 800 4 SC_OUT_BOT
port 3 nsew
rlabel metal2 s 17590 23600 17646 24400 4 SC_OUT_TOP
port 4 nsew
rlabel metal3 s 23600 6808 24400 6928 4 Test_en_E_in
port 5 nsew
rlabel metal3 s 23600 6128 24400 6248 4 Test_en_E_out
port 6 nsew
rlabel metal3 s 0 21224 800 21344 4 Test_en_W_in
port 7 nsew
rlabel metal3 s 0 15104 800 15224 4 Test_en_W_out
port 8 nsew
rlabel metal2 s 1674 0 1730 800 4 bottom_width_0_height_0__pin_50_
port 9 nsew
rlabel metal2 s 5078 0 5134 800 4 bottom_width_0_height_0__pin_51_
port 10 nsew
rlabel metal3 s 0 8984 800 9104 4 ccff_head
port 11 nsew
rlabel metal3 s 23600 5448 24400 5568 4 ccff_tail
port 12 nsew
rlabel metal2 s 18234 23600 18290 24400 4 clk_0_N_in
port 13 nsew
rlabel metal2 s 15566 0 15622 800 4 clk_0_S_in
port 14 nsew
rlabel metal3 s 23600 8168 24400 8288 4 prog_clk_0_E_out
port 15 nsew
rlabel metal3 s 23600 7488 24400 7608 4 prog_clk_0_N_in
port 16 nsew
rlabel metal2 s 18878 23600 18934 24400 4 prog_clk_0_N_out
port 17 nsew
rlabel metal2 s 19062 0 19118 800 4 prog_clk_0_S_in
port 18 nsew
rlabel metal2 s 22558 0 22614 800 4 prog_clk_0_S_out
port 19 nsew
rlabel metal3 s 0 3000 800 3120 4 prog_clk_0_W_out
port 20 nsew
rlabel metal3 s 23600 8712 24400 8832 4 right_width_0_height_0__pin_16_
port 21 nsew
rlabel metal3 s 23600 9392 24400 9512 4 right_width_0_height_0__pin_17_
port 22 nsew
rlabel metal3 s 23600 10072 24400 10192 4 right_width_0_height_0__pin_18_
port 23 nsew
rlabel metal3 s 23600 10752 24400 10872 4 right_width_0_height_0__pin_19_
port 24 nsew
rlabel metal3 s 23600 11432 24400 11552 4 right_width_0_height_0__pin_20_
port 25 nsew
rlabel metal3 s 23600 12112 24400 12232 4 right_width_0_height_0__pin_21_
port 26 nsew
rlabel metal3 s 23600 12656 24400 12776 4 right_width_0_height_0__pin_22_
port 27 nsew
rlabel metal3 s 23600 13336 24400 13456 4 right_width_0_height_0__pin_23_
port 28 nsew
rlabel metal3 s 23600 14016 24400 14136 4 right_width_0_height_0__pin_24_
port 29 nsew
rlabel metal3 s 23600 14696 24400 14816 4 right_width_0_height_0__pin_25_
port 30 nsew
rlabel metal3 s 23600 15376 24400 15496 4 right_width_0_height_0__pin_26_
port 31 nsew
rlabel metal3 s 23600 16056 24400 16176 4 right_width_0_height_0__pin_27_
port 32 nsew
rlabel metal3 s 23600 16600 24400 16720 4 right_width_0_height_0__pin_28_
port 33 nsew
rlabel metal3 s 23600 17280 24400 17400 4 right_width_0_height_0__pin_29_
port 34 nsew
rlabel metal3 s 23600 17960 24400 18080 4 right_width_0_height_0__pin_30_
port 35 nsew
rlabel metal3 s 23600 18640 24400 18760 4 right_width_0_height_0__pin_31_
port 36 nsew
rlabel metal3 s 23600 280 24400 400 4 right_width_0_height_0__pin_42_lower
port 37 nsew
rlabel metal3 s 23600 19320 24400 19440 4 right_width_0_height_0__pin_42_upper
port 38 nsew
rlabel metal3 s 23600 824 24400 944 4 right_width_0_height_0__pin_43_lower
port 39 nsew
rlabel metal3 s 23600 20000 24400 20120 4 right_width_0_height_0__pin_43_upper
port 40 nsew
rlabel metal3 s 23600 1504 24400 1624 4 right_width_0_height_0__pin_44_lower
port 41 nsew
rlabel metal3 s 23600 20544 24400 20664 4 right_width_0_height_0__pin_44_upper
port 42 nsew
rlabel metal3 s 23600 2184 24400 2304 4 right_width_0_height_0__pin_45_lower
port 43 nsew
rlabel metal3 s 23600 21224 24400 21344 4 right_width_0_height_0__pin_45_upper
port 44 nsew
rlabel metal3 s 23600 2864 24400 2984 4 right_width_0_height_0__pin_46_lower
port 45 nsew
rlabel metal3 s 23600 21904 24400 22024 4 right_width_0_height_0__pin_46_upper
port 46 nsew
rlabel metal3 s 23600 3544 24400 3664 4 right_width_0_height_0__pin_47_lower
port 47 nsew
rlabel metal3 s 23600 22584 24400 22704 4 right_width_0_height_0__pin_47_upper
port 48 nsew
rlabel metal3 s 23600 4224 24400 4344 4 right_width_0_height_0__pin_48_lower
port 49 nsew
rlabel metal3 s 23600 23264 24400 23384 4 right_width_0_height_0__pin_48_upper
port 50 nsew
rlabel metal3 s 23600 4768 24400 4888 4 right_width_0_height_0__pin_49_lower
port 51 nsew
rlabel metal3 s 23600 23944 24400 24064 4 right_width_0_height_0__pin_49_upper
port 52 nsew
rlabel metal2 s 5354 23600 5410 24400 4 top_width_0_height_0__pin_0_
port 53 nsew
rlabel metal2 s 11794 23600 11850 24400 4 top_width_0_height_0__pin_10_
port 54 nsew
rlabel metal2 s 12438 23600 12494 24400 4 top_width_0_height_0__pin_11_
port 55 nsew
rlabel metal2 s 13082 23600 13138 24400 4 top_width_0_height_0__pin_12_
port 56 nsew
rlabel metal2 s 13726 23600 13782 24400 4 top_width_0_height_0__pin_13_
port 57 nsew
rlabel metal2 s 14370 23600 14426 24400 4 top_width_0_height_0__pin_14_
port 58 nsew
rlabel metal2 s 15014 23600 15070 24400 4 top_width_0_height_0__pin_15_
port 59 nsew
rlabel metal2 s 5998 23600 6054 24400 4 top_width_0_height_0__pin_1_
port 60 nsew
rlabel metal2 s 6642 23600 6698 24400 4 top_width_0_height_0__pin_2_
port 61 nsew
rlabel metal2 s 15658 23600 15714 24400 4 top_width_0_height_0__pin_32_
port 62 nsew
rlabel metal2 s 16302 23600 16358 24400 4 top_width_0_height_0__pin_33_
port 63 nsew
rlabel metal2 s 19522 23600 19578 24400 4 top_width_0_height_0__pin_34_lower
port 64 nsew
rlabel metal2 s 294 23600 350 24400 4 top_width_0_height_0__pin_34_upper
port 65 nsew
rlabel metal2 s 20166 23600 20222 24400 4 top_width_0_height_0__pin_35_lower
port 66 nsew
rlabel metal2 s 846 23600 902 24400 4 top_width_0_height_0__pin_35_upper
port 67 nsew
rlabel metal2 s 20810 23600 20866 24400 4 top_width_0_height_0__pin_36_lower
port 68 nsew
rlabel metal2 s 1490 23600 1546 24400 4 top_width_0_height_0__pin_36_upper
port 69 nsew
rlabel metal2 s 21454 23600 21510 24400 4 top_width_0_height_0__pin_37_lower
port 70 nsew
rlabel metal2 s 2134 23600 2190 24400 4 top_width_0_height_0__pin_37_upper
port 71 nsew
rlabel metal2 s 22098 23600 22154 24400 4 top_width_0_height_0__pin_38_lower
port 72 nsew
rlabel metal2 s 2778 23600 2834 24400 4 top_width_0_height_0__pin_38_upper
port 73 nsew
rlabel metal2 s 22742 23600 22798 24400 4 top_width_0_height_0__pin_39_lower
port 74 nsew
rlabel metal2 s 3422 23600 3478 24400 4 top_width_0_height_0__pin_39_upper
port 75 nsew
rlabel metal2 s 7286 23600 7342 24400 4 top_width_0_height_0__pin_3_
port 76 nsew
rlabel metal2 s 23386 23600 23442 24400 4 top_width_0_height_0__pin_40_lower
port 77 nsew
rlabel metal2 s 4066 23600 4122 24400 4 top_width_0_height_0__pin_40_upper
port 78 nsew
rlabel metal2 s 24030 23600 24086 24400 4 top_width_0_height_0__pin_41_lower
port 79 nsew
rlabel metal2 s 4710 23600 4766 24400 4 top_width_0_height_0__pin_41_upper
port 80 nsew
rlabel metal2 s 7930 23600 7986 24400 4 top_width_0_height_0__pin_4_
port 81 nsew
rlabel metal2 s 8574 23600 8630 24400 4 top_width_0_height_0__pin_5_
port 82 nsew
rlabel metal2 s 9218 23600 9274 24400 4 top_width_0_height_0__pin_6_
port 83 nsew
rlabel metal2 s 9862 23600 9918 24400 4 top_width_0_height_0__pin_7_
port 84 nsew
rlabel metal2 s 10506 23600 10562 24400 4 top_width_0_height_0__pin_8_
port 85 nsew
rlabel metal2 s 11150 23600 11206 24400 4 top_width_0_height_0__pin_9_
port 86 nsew
rlabel metal4 s 4643 2128 4963 21808 4 VPWR
port 87 nsew
rlabel metal4 s 8341 2128 8661 21808 4 VGND
port 88 nsew
<< properties >>
string FIXED_BBOX 0 0 24400 24400
string GDS_FILE /ef/openfpga/openlane/runs/grid_clb/results/magic/grid_clb.gds
string GDS_END 1854502
string GDS_START 101400
<< end >>
