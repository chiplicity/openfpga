* NGSPICE file created from sb_0__2_.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_12 abstract view
.subckt sky130_fd_sc_hd__decap_12 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_1 abstract view
.subckt sky130_fd_sc_hd__dfxtp_1 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
.subckt sky130_fd_sc_hd__conb_1 VGND VNB VPB VPWR HI LO
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_8 abstract view
.subckt sky130_fd_sc_hd__buf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

.subckt sb_0__2_ SC_IN_TOP SC_OUT_BOT bottom_left_grid_pin_1_ ccff_head ccff_tail
+ chanx_right_in[0] chanx_right_in[10] chanx_right_in[11] chanx_right_in[12] chanx_right_in[13]
+ chanx_right_in[14] chanx_right_in[15] chanx_right_in[16] chanx_right_in[17] chanx_right_in[18]
+ chanx_right_in[19] chanx_right_in[1] chanx_right_in[2] chanx_right_in[3] chanx_right_in[4]
+ chanx_right_in[5] chanx_right_in[6] chanx_right_in[7] chanx_right_in[8] chanx_right_in[9]
+ chanx_right_out[0] chanx_right_out[10] chanx_right_out[11] chanx_right_out[12] chanx_right_out[13]
+ chanx_right_out[14] chanx_right_out[15] chanx_right_out[16] chanx_right_out[17]
+ chanx_right_out[18] chanx_right_out[19] chanx_right_out[1] chanx_right_out[2] chanx_right_out[3]
+ chanx_right_out[4] chanx_right_out[5] chanx_right_out[6] chanx_right_out[7] chanx_right_out[8]
+ chanx_right_out[9] chany_bottom_in[0] chany_bottom_in[10] chany_bottom_in[11] chany_bottom_in[12]
+ chany_bottom_in[13] chany_bottom_in[14] chany_bottom_in[15] chany_bottom_in[16]
+ chany_bottom_in[17] chany_bottom_in[18] chany_bottom_in[19] chany_bottom_in[1] chany_bottom_in[2]
+ chany_bottom_in[3] chany_bottom_in[4] chany_bottom_in[5] chany_bottom_in[6] chany_bottom_in[7]
+ chany_bottom_in[8] chany_bottom_in[9] chany_bottom_out[0] chany_bottom_out[10] chany_bottom_out[11]
+ chany_bottom_out[12] chany_bottom_out[13] chany_bottom_out[14] chany_bottom_out[15]
+ chany_bottom_out[16] chany_bottom_out[17] chany_bottom_out[18] chany_bottom_out[19]
+ chany_bottom_out[1] chany_bottom_out[2] chany_bottom_out[3] chany_bottom_out[4]
+ chany_bottom_out[5] chany_bottom_out[6] chany_bottom_out[7] chany_bottom_out[8]
+ chany_bottom_out[9] prog_clk_0_E_in right_bottom_grid_pin_34_ right_bottom_grid_pin_35_
+ right_bottom_grid_pin_36_ right_bottom_grid_pin_37_ right_bottom_grid_pin_38_ right_bottom_grid_pin_39_
+ right_bottom_grid_pin_40_ right_bottom_grid_pin_41_ right_top_grid_pin_1_ VPWR VGND
XFILLER_22_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmem_right_track_20.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_2_3_0_mem_bottom_track_1.prog_clk/X
+ mux_right_track_20.mux_l1_in_0_/S VGND VGND VPWR VPWR mux_right_track_20.mux_l2_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
Xmem_right_track_2.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_2_2_0_mem_bottom_track_1.prog_clk/X
+ mux_right_track_0.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_right_track_2.mux_l1_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_13_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_83_ chanx_right_in[4] VGND VGND VPWR VPWR chany_bottom_out[14] sky130_fd_sc_hd__buf_2
XFILLER_8_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_66_ _66_/A VGND VGND VPWR VPWR chanx_right_out[17] sky130_fd_sc_hd__buf_2
XFILLER_5_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_right_track_36.sky130_fd_sc_hd__buf_4_0_ mux_right_track_36.mux_l2_in_0_/X VGND
+ VGND VPWR VPWR _67_/A sky130_fd_sc_hd__buf_4
XFILLER_23_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_right_track_4.mux_l1_in_0__A1 right_top_grid_pin_1_ VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
Xmem_right_track_8.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_2_0_0_mem_bottom_track_1.prog_clk/X
+ mux_right_track_8.mux_l1_in_0_/S VGND VGND VPWR VPWR mux_right_track_8.mux_l2_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_2_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_49_ _49_/A VGND VGND VPWR VPWR chanx_right_out[0] sky130_fd_sc_hd__buf_2
XFILLER_29_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_track_2.mux_l2_in_1__A1 chany_bottom_in[17] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XPHY_192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_right_track_38.mux_l1_in_0_ chany_bottom_in[19] right_bottom_grid_pin_40_ mux_right_track_38.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_right_track_38.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_22_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmem_right_track_20.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_2_3_0_mem_bottom_track_1.prog_clk/X
+ mux_right_track_18.mux_l2_in_0_/S VGND VGND VPWR VPWR mux_right_track_20.mux_l1_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_13_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_82_ chanx_right_in[5] VGND VGND VPWR VPWR chany_bottom_out[13] sky130_fd_sc_hd__buf_2
Xclkbuf_1_0_0_mem_bottom_track_1.prog_clk clkbuf_0_mem_bottom_track_1.prog_clk/X VGND
+ VGND VPWR VPWR clkbuf_2_1_0_mem_bottom_track_1.prog_clk/A sky130_fd_sc_hd__clkbuf_1
XFILLER_33_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_65_ _65_/A VGND VGND VPWR VPWR chanx_right_out[16] sky130_fd_sc_hd__buf_2
XFILLER_15_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmem_right_track_8.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_2_0_0_mem_bottom_track_1.prog_clk/X
+ mux_right_track_6.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_right_track_8.mux_l1_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
Xmem_right_track_26.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_2_0_0_mem_bottom_track_1.prog_clk/X
+ mux_right_track_26.mux_l1_in_0_/S VGND VGND VPWR VPWR mux_right_track_26.mux_l2_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
X_48_ SC_IN_TOP VGND VGND VPWR VPWR SC_OUT_BOT sky130_fd_sc_hd__buf_2
XFILLER_18_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_bottom_track_25.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_2_3_0_mem_bottom_track_1.prog_clk/X
+ mux_bottom_track_25.mux_l1_in_0_/S VGND VGND VPWR VPWR ccff_tail sky130_fd_sc_hd__dfxtp_1
XFILLER_29_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_right_track_6.mux_l1_in_1__A0 right_bottom_grid_pin_40_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_81_ _81_/A VGND VGND VPWR VPWR chany_bottom_out[12] sky130_fd_sc_hd__buf_2
XFILLER_12_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_64_ _64_/A VGND VGND VPWR VPWR chanx_right_out[15] sky130_fd_sc_hd__buf_2
XFILLER_5_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmem_right_track_26.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_2_0_0_mem_bottom_track_1.prog_clk/X
+ mux_right_track_24.mux_l2_in_0_/S VGND VGND VPWR VPWR mux_right_track_26.mux_l1_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
X_47_ VGND VGND VPWR VPWR _47_/HI _47_/LO sky130_fd_sc_hd__conb_1
XFILLER_18_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmem_bottom_track_25.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_2_3_0_mem_bottom_track_1.prog_clk/X
+ mux_bottom_track_9.mux_l2_in_0_/S VGND VGND VPWR VPWR mux_bottom_track_25.mux_l1_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_29_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mux_right_track_6.mux_l1_in_1__A1 right_bottom_grid_pin_38_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
X_80_ chanx_right_in[7] VGND VGND VPWR VPWR chany_bottom_out[11] sky130_fd_sc_hd__buf_2
XFILLER_3_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_63_ _63_/A VGND VGND VPWR VPWR chanx_right_out[14] sky130_fd_sc_hd__buf_2
Xprog_clk_0_FTB00 prog_clk_0_E_in VGND VGND VPWR VPWR prog_clk_0_FTB00/X sky130_fd_sc_hd__buf_8
XFILLER_0_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mux_right_track_14.mux_l1_in_0__A0 chany_bottom_in[11] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_29_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_46_ VGND VGND VPWR VPWR _46_/HI _46_/LO sky130_fd_sc_hd__conb_1
XFILLER_20_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_right_track_10.mux_l2_in_0_ _41_/HI mux_right_track_10.mux_l1_in_0_/X mux_right_track_10.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR mux_right_track_10.mux_l2_in_0_/X sky130_fd_sc_hd__mux2_1
X_29_ VGND VGND VPWR VPWR _29_/HI _29_/LO sky130_fd_sc_hd__conb_1
XFILLER_4_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_track_22.mux_l1_in_0__A0 chany_bottom_in[7] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
X_62_ _62_/A VGND VGND VPWR VPWR chanx_right_out[13] sky130_fd_sc_hd__buf_2
Xmem_bottom_track_9.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_2_3_0_mem_bottom_track_1.prog_clk/X
+ mux_bottom_track_9.mux_l1_in_0_/S VGND VGND VPWR VPWR mux_bottom_track_9.mux_l2_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA_mux_right_track_14.mux_l1_in_0__A1 right_bottom_grid_pin_36_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_45_ VGND VGND VPWR VPWR _45_/HI _45_/LO sky130_fd_sc_hd__conb_1
X_28_ VGND VGND VPWR VPWR _28_/HI _28_/LO sky130_fd_sc_hd__conb_1
XFILLER_28_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmem_right_track_12.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_2_0_0_mem_bottom_track_1.prog_clk/X
+ mux_right_track_12.mux_l1_in_0_/S VGND VGND VPWR VPWR mux_right_track_12.mux_l2_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XPHY_185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmux_right_track_10.mux_l1_in_0_ chany_bottom_in[13] right_bottom_grid_pin_34_ mux_right_track_10.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_right_track_10.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
Xmux_right_track_8.mux_l2_in_0_ mux_right_track_8.mux_l1_in_1_/X mux_right_track_8.mux_l1_in_0_/X
+ mux_right_track_8.mux_l2_in_0_/S VGND VGND VPWR VPWR mux_right_track_8.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
Xmux_right_track_22.mux_l2_in_0_ _24_/HI mux_right_track_22.mux_l1_in_0_/X mux_right_track_22.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR mux_right_track_22.mux_l2_in_0_/X sky130_fd_sc_hd__mux2_1
XANTENNA_mux_right_track_30.mux_l1_in_0__A0 chany_bottom_in[3] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_26_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mux_right_track_22.mux_l1_in_0__A1 right_bottom_grid_pin_40_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_right_track_8.mux_l1_in_1_ _35_/HI chany_bottom_in[14] mux_right_track_8.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_right_track_8.mux_l1_in_1_/X sky130_fd_sc_hd__mux2_1
X_61_ _61_/A VGND VGND VPWR VPWR chanx_right_out[12] sky130_fd_sc_hd__buf_2
XFILLER_5_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmem_bottom_track_9.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_2_3_0_mem_bottom_track_1.prog_clk/X
+ mux_bottom_track_5.mux_l2_in_0_/S VGND VGND VPWR VPWR mux_bottom_track_9.mux_l1_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_9_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_44_ VGND VGND VPWR VPWR _44_/HI _44_/LO sky130_fd_sc_hd__conb_1
XFILLER_1_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_right_track_10.sky130_fd_sc_hd__buf_4_0_ mux_right_track_10.mux_l2_in_0_/X VGND
+ VGND VPWR VPWR _54_/A sky130_fd_sc_hd__buf_4
XFILLER_1_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27_ VGND VGND VPWR VPWR _27_/HI _27_/LO sky130_fd_sc_hd__conb_1
XFILLER_28_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmem_right_track_12.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_2_0_0_mem_bottom_track_1.prog_clk/X
+ mux_right_track_10.mux_l2_in_0_/S VGND VGND VPWR VPWR mux_right_track_12.mux_l1_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XPHY_186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_0 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mux_right_track_30.mux_l1_in_0__A1 right_bottom_grid_pin_36_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_bottom_track_25.mux_l1_in_0__A0 bottom_left_grid_pin_1_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_right_track_8.mux_l1_in_0_ right_bottom_grid_pin_41_ right_top_grid_pin_1_ mux_right_track_8.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_right_track_8.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_32_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_60_ _60_/A VGND VGND VPWR VPWR chanx_right_out[11] sky130_fd_sc_hd__buf_2
Xmem_right_track_18.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_2_3_0_mem_bottom_track_1.prog_clk/X
+ mux_right_track_18.mux_l1_in_0_/S VGND VGND VPWR VPWR mux_right_track_18.mux_l2_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
Xmux_right_track_22.mux_l1_in_0_ chany_bottom_in[7] right_bottom_grid_pin_40_ mux_right_track_22.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_right_track_22.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_5_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_right_track_34.mux_l2_in_0_ _30_/HI mux_right_track_34.mux_l1_in_0_/X mux_right_track_34.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR mux_right_track_34.mux_l2_in_0_/X sky130_fd_sc_hd__mux2_1
Xmux_right_track_8.sky130_fd_sc_hd__buf_4_0_ mux_right_track_8.mux_l2_in_0_/X VGND
+ VGND VPWR VPWR _53_/A sky130_fd_sc_hd__buf_4
XFILLER_14_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_43_ VGND VGND VPWR VPWR _43_/HI _43_/LO sky130_fd_sc_hd__conb_1
XFILLER_1_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26_ VGND VGND VPWR VPWR _26_/HI _26_/LO sky130_fd_sc_hd__conb_1
XFILLER_28_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_right_track_32.sky130_fd_sc_hd__buf_4_0_ mux_right_track_32.mux_l2_in_0_/X VGND
+ VGND VPWR VPWR _65_/A sky130_fd_sc_hd__buf_4
XFILLER_25_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_bottom_track_25.mux_l1_in_0__A1 chanx_right_in[6] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_32_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_right_track_26.sky130_fd_sc_hd__buf_4_0_ mux_right_track_26.mux_l2_in_0_/X VGND
+ VGND VPWR VPWR _62_/A sky130_fd_sc_hd__buf_4
XFILLER_12_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmem_right_track_18.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_2_1_0_mem_bottom_track_1.prog_clk/X
+ mux_right_track_16.mux_l2_in_0_/S VGND VGND VPWR VPWR mux_right_track_18.mux_l1_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_32_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_bottom_track_25.mux_l2_in_0_ _37_/HI mux_bottom_track_25.mux_l1_in_0_/X ccff_tail
+ VGND VGND VPWR VPWR mux_bottom_track_25.mux_l2_in_0_/X sky130_fd_sc_hd__mux2_1
X_42_ VGND VGND VPWR VPWR _42_/HI _42_/LO sky130_fd_sc_hd__conb_1
XFILLER_18_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmem_right_track_30.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_2_1_0_mem_bottom_track_1.prog_clk/X
+ mux_right_track_30.mux_l1_in_0_/S VGND VGND VPWR VPWR mux_right_track_30.mux_l2_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__48__A SC_IN_TOP VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_right_track_34.mux_l1_in_0_ chany_bottom_in[1] right_bottom_grid_pin_38_ mux_right_track_34.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_right_track_34.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_29_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25_ VGND VGND VPWR VPWR _25_/HI _25_/LO sky130_fd_sc_hd__conb_1
XFILLER_29_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_bottom_track_9.mux_l2_in_0_ _39_/HI mux_bottom_track_9.mux_l1_in_0_/X mux_bottom_track_9.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR mux_bottom_track_9.mux_l2_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_19_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_right_track_24.mux_l1_in_1__A1 chany_bottom_in[6] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_31_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mux_right_track_0.mux_l1_in_0__A0 right_bottom_grid_pin_35_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_41_ VGND VGND VPWR VPWR _41_/HI _41_/LO sky130_fd_sc_hd__conb_1
XFILLER_20_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmem_right_track_30.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_2_0_0_mem_bottom_track_1.prog_clk/X
+ mux_right_track_28.mux_l2_in_0_/S VGND VGND VPWR VPWR mux_right_track_30.mux_l1_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
X_24_ VGND VGND VPWR VPWR _24_/HI _24_/LO sky130_fd_sc_hd__conb_1
XFILLER_29_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_bottom_track_25.mux_l1_in_0_ bottom_left_grid_pin_1_ chanx_right_in[6] mux_bottom_track_25.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_bottom_track_25.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_32_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmem_right_track_36.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_2_3_0_mem_bottom_track_1.prog_clk/X
+ mux_right_track_36.mux_l1_in_0_/S VGND VGND VPWR VPWR mux_right_track_36.mux_l2_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_16_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_mux_right_track_0.mux_l1_in_0__A1 right_top_grid_pin_1_ VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XPHY_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_bottom_track_9.mux_l1_in_0_ bottom_left_grid_pin_1_ chanx_right_in[14] mux_bottom_track_9.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_bottom_track_9.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XANTENNA__72__A chanx_right_in[15] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_bottom_track_9.sky130_fd_sc_hd__buf_4_0_ mux_bottom_track_9.mux_l2_in_0_/X VGND
+ VGND VPWR VPWR _73_/A sky130_fd_sc_hd__buf_4
XFILLER_5_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_right_track_28.mux_l1_in_0__A0 chany_bottom_in[4] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_4_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_40_ VGND VGND VPWR VPWR _40_/HI _40_/LO sky130_fd_sc_hd__conb_1
XANTENNA__80__A chanx_right_in[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__75__A chanx_right_in[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_bottom_track_25.mux_l2_in_0__S ccff_tail VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmem_right_track_36.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_2_3_0_mem_bottom_track_1.prog_clk/X
+ mux_right_track_34.mux_l2_in_0_/S VGND VGND VPWR VPWR mux_right_track_36.mux_l1_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XPHY_124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_right_track_36.mux_l1_in_0__A0 chany_bottom_in[0] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_17_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__83__A chanx_right_in[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_28.mux_l1_in_0__A1 right_bottom_grid_pin_35_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xmux_right_track_4.mux_l3_in_0_ mux_right_track_4.mux_l2_in_1_/X mux_right_track_4.mux_l2_in_0_/X
+ mux_right_track_4.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_right_track_4.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_4_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__78__A chanx_right_in[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_right_track_4.sky130_fd_sc_hd__dfxtp_1_2_ clkbuf_2_2_0_mem_bottom_track_1.prog_clk/X
+ mux_right_track_4.mux_l2_in_0_/S VGND VGND VPWR VPWR mux_right_track_4.mux_l3_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_6_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_right_track_4.mux_l2_in_1_ _33_/HI mux_right_track_4.mux_l1_in_2_/X mux_right_track_4.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR mux_right_track_4.mux_l2_in_1_/X sky130_fd_sc_hd__mux2_1
XANTENNA_mux_right_track_2.mux_l1_in_1__A0 right_bottom_grid_pin_40_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmux_right_track_4.mux_l1_in_2_ chany_bottom_in[16] right_bottom_grid_pin_41_ mux_right_track_4.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_right_track_4.mux_l1_in_2_/X sky130_fd_sc_hd__mux2_1
XFILLER_30_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__86__A chanx_right_in[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_right_track_36.mux_l1_in_0__A1 right_bottom_grid_pin_39_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmem_right_track_4.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_2_2_0_mem_bottom_track_1.prog_clk/X
+ mux_right_track_4.mux_l1_in_0_/S VGND VGND VPWR VPWR mux_right_track_4.mux_l2_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
Xmux_right_track_16.mux_l2_in_0_ _44_/HI mux_right_track_16.mux_l1_in_0_/X mux_right_track_16.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR mux_right_track_16.mux_l2_in_0_/X sky130_fd_sc_hd__mux2_1
XANTENNA_mux_right_track_2.mux_l1_in_1__A1 right_bottom_grid_pin_38_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xmux_right_track_4.mux_l2_in_0_ mux_right_track_4.mux_l1_in_1_/X mux_right_track_4.mux_l1_in_0_/X
+ mux_right_track_4.mux_l2_in_0_/S VGND VGND VPWR VPWR mux_right_track_4.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_28_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmux_right_track_4.mux_l1_in_1_ right_bottom_grid_pin_39_ right_bottom_grid_pin_37_
+ mux_right_track_4.mux_l1_in_0_/S VGND VGND VPWR VPWR mux_right_track_4.mux_l1_in_1_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_30_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_right_track_10.mux_l1_in_0__A0 chany_bottom_in[13] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XPHY_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmem_right_track_22.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_2_2_0_mem_bottom_track_1.prog_clk/X
+ mux_right_track_22.mux_l1_in_0_/S VGND VGND VPWR VPWR mux_right_track_22.mux_l2_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_9_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmem_right_track_4.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_2_2_0_mem_bottom_track_1.prog_clk/X
+ mux_right_track_2.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_right_track_4.mux_l1_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_10_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmux_right_track_16.mux_l1_in_0_ chany_bottom_in[10] right_bottom_grid_pin_37_ mux_right_track_16.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_right_track_16.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XPHY_105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_right_track_4.mux_l1_in_0_ right_bottom_grid_pin_35_ right_top_grid_pin_1_ mux_right_track_4.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_right_track_4.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_24_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmux_right_track_4.sky130_fd_sc_hd__buf_4_0_ mux_right_track_4.mux_l3_in_0_/X VGND
+ VGND VPWR VPWR _51_/A sky130_fd_sc_hd__buf_4
XPHY_138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_right_track_28.mux_l2_in_0_ _27_/HI mux_right_track_28.mux_l1_in_0_/X mux_right_track_28.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR mux_right_track_28.mux_l2_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_23_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_right_track_30.mux_l2_in_0_ _28_/HI mux_right_track_30.mux_l1_in_0_/X mux_right_track_30.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR mux_right_track_30.mux_l2_in_0_/X sky130_fd_sc_hd__mux2_1
XANTENNA_mux_right_track_10.mux_l1_in_0__A1 right_bottom_grid_pin_34_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_6.mux_l1_in_0__A0 right_bottom_grid_pin_36_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mux_right_track_4.mux_l1_in_2__A0 chany_bottom_in[16] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_32_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmem_right_track_22.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_2_2_0_mem_bottom_track_1.prog_clk/X
+ mux_right_track_20.mux_l2_in_0_/S VGND VGND VPWR VPWR mux_right_track_22.mux_l1_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_1_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_right_track_22.sky130_fd_sc_hd__buf_4_0_ mux_right_track_22.mux_l2_in_0_/X VGND
+ VGND VPWR VPWR _60_/A sky130_fd_sc_hd__buf_4
XFILLER_10_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_79_ chanx_right_in[8] VGND VGND VPWR VPWR chany_bottom_out[10] sky130_fd_sc_hd__buf_2
XFILLER_19_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmem_right_track_28.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_2_0_0_mem_bottom_track_1.prog_clk/X
+ mux_right_track_28.mux_l1_in_0_/S VGND VGND VPWR VPWR mux_right_track_28.mux_l2_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_24_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_right_track_16.sky130_fd_sc_hd__buf_4_0_ mux_right_track_16.mux_l2_in_0_/X VGND
+ VGND VPWR VPWR _57_/A sky130_fd_sc_hd__buf_4
XPHY_139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_right_track_6.mux_l1_in_0__A1 right_bottom_grid_pin_34_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_right_track_28.mux_l1_in_0_ chany_bottom_in[4] right_bottom_grid_pin_35_ mux_right_track_28.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_right_track_28.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_27_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_right_track_4.mux_l1_in_2__A1 right_bottom_grid_pin_41_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_right_track_30.mux_l1_in_0_ chany_bottom_in[3] right_bottom_grid_pin_36_ mux_right_track_30.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_right_track_30.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
Xmux_bottom_track_5.mux_l2_in_0_ _38_/HI mux_bottom_track_5.mux_l1_in_0_/X mux_bottom_track_5.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR mux_bottom_track_5.mux_l2_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_24_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_78_ chanx_right_in[9] VGND VGND VPWR VPWR chany_bottom_out[9] sky130_fd_sc_hd__buf_2
XFILLER_10_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmem_right_track_28.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_2_0_0_mem_bottom_track_1.prog_clk/X
+ mux_right_track_26.mux_l2_in_0_/S VGND VGND VPWR VPWR mux_right_track_28.mux_l1_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_24_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_2_3_0_mem_bottom_track_1.prog_clk clkbuf_2_3_0_mem_bottom_track_1.prog_clk/A
+ VGND VGND VPWR VPWR clkbuf_2_3_0_mem_bottom_track_1.prog_clk/X sky130_fd_sc_hd__clkbuf_1
XPHY_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_prog_clk_0_FTB00_A prog_clk_0_E_in VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_right_track_38.sky130_fd_sc_hd__buf_4_0_ mux_right_track_38.mux_l2_in_0_/X VGND
+ VGND VPWR VPWR _68_/A sky130_fd_sc_hd__buf_4
XFILLER_16_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_2_3_0_mem_bottom_track_1.prog_clk/X
+ mux_bottom_track_5.mux_l1_in_0_/S VGND VGND VPWR VPWR mux_bottom_track_5.mux_l2_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_24_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_bottom_track_5.sky130_fd_sc_hd__buf_4_0_ mux_bottom_track_5.mux_l2_in_0_/X VGND
+ VGND VPWR VPWR _71_/A sky130_fd_sc_hd__buf_4
X_77_ chanx_right_in[10] VGND VGND VPWR VPWR chany_bottom_out[8] sky130_fd_sc_hd__buf_2
Xmux_bottom_track_5.mux_l1_in_0_ bottom_left_grid_pin_1_ chanx_right_in[16] mux_bottom_track_5.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_bottom_track_5.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_33_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_2_3_0_mem_bottom_track_1.prog_clk/X
+ mux_bottom_track_1.mux_l2_in_0_/S VGND VGND VPWR VPWR mux_bottom_track_5.mux_l1_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_1_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_76_ chanx_right_in[11] VGND VGND VPWR VPWR chany_bottom_out[7] sky130_fd_sc_hd__buf_2
XFILLER_1_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_right_track_8.mux_l1_in_1__A1 chany_bottom_in[14] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_10_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_59_ _59_/A VGND VGND VPWR VPWR chanx_right_out[10] sky130_fd_sc_hd__buf_2
XPHY_109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_right_track_0.mux_l3_in_0_ mux_right_track_0.mux_l2_in_1_/X mux_right_track_0.mux_l2_in_0_/X
+ mux_right_track_0.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_right_track_0.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_32_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_bottom_track_9.mux_l1_in_0__A0 bottom_left_grid_pin_1_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_16.mux_l1_in_0__A0 chany_bottom_in[10] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_14_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_right_track_0.mux_l2_in_1_ _40_/HI mux_right_track_0.mux_l1_in_2_/X mux_right_track_0.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR mux_right_track_0.mux_l2_in_1_/X sky130_fd_sc_hd__mux2_1
XFILLER_31_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmem_right_track_14.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_2_1_0_mem_bottom_track_1.prog_clk/X
+ mux_right_track_14.mux_l1_in_0_/S VGND VGND VPWR VPWR mux_right_track_14.mux_l2_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_13_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_right_track_0.mux_l1_in_2_ chany_bottom_in[18] right_bottom_grid_pin_41_ mux_right_track_0.mux_l1_in_1_/S
+ VGND VGND VPWR VPWR mux_right_track_0.mux_l1_in_2_/X sky130_fd_sc_hd__mux2_1
XFILLER_14_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_75_ chanx_right_in[12] VGND VGND VPWR VPWR chany_bottom_out[6] sky130_fd_sc_hd__buf_2
XFILLER_27_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_58_ _58_/A VGND VGND VPWR VPWR chanx_right_out[9] sky130_fd_sc_hd__buf_2
XANTENNA_mux_right_track_24.mux_l1_in_0__A0 right_bottom_grid_pin_41_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XPHY_90 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_bottom_track_9.mux_l1_in_0__A1 chanx_right_in[14] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_16.mux_l1_in_0__A1 right_bottom_grid_pin_37_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_right_track_12.mux_l2_in_0_ _42_/HI mux_right_track_12.mux_l1_in_0_/X mux_right_track_12.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR mux_right_track_12.mux_l2_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_4_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_right_track_0.mux_l2_in_0_ mux_right_track_0.mux_l1_in_1_/X mux_right_track_0.mux_l1_in_0_/X
+ mux_right_track_0.mux_l2_in_0_/S VGND VGND VPWR VPWR mux_right_track_0.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
Xmem_right_track_14.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_2_0_0_mem_bottom_track_1.prog_clk/X
+ mux_right_track_12.mux_l2_in_0_/S VGND VGND VPWR VPWR mux_right_track_14.mux_l1_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_22_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_right_track_0.mux_l1_in_1_ right_bottom_grid_pin_39_ right_bottom_grid_pin_37_
+ mux_right_track_0.mux_l1_in_1_/S VGND VGND VPWR VPWR mux_right_track_0.mux_l1_in_1_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_5_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_74_ chanx_right_in[13] VGND VGND VPWR VPWR chany_bottom_out[5] sky130_fd_sc_hd__buf_2
XANTENNA_mux_right_track_32.mux_l1_in_0__A0 chany_bottom_in[2] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_27_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_mux_right_track_24.mux_l1_in_0__A1 right_top_grid_pin_1_ VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XPHY_80 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_91 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_57_ _57_/A VGND VGND VPWR VPWR chanx_right_out[8] sky130_fd_sc_hd__buf_2
XFILLER_24_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_right_track_0.sky130_fd_sc_hd__buf_4_0_ mux_right_track_0.mux_l3_in_0_/X VGND
+ VGND VPWR VPWR _49_/A sky130_fd_sc_hd__buf_4
XFILLER_13_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_right_track_12.mux_l1_in_0_ chany_bottom_in[12] right_bottom_grid_pin_35_ mux_right_track_12.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_right_track_12.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_5_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_right_track_0.mux_l1_in_0_ right_bottom_grid_pin_35_ right_top_grid_pin_1_ mux_right_track_0.mux_l1_in_1_/S
+ VGND VGND VPWR VPWR mux_right_track_0.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_10_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_right_track_24.mux_l2_in_0_ mux_right_track_24.mux_l1_in_1_/X mux_right_track_24.mux_l1_in_0_/X
+ mux_right_track_24.mux_l2_in_0_/S VGND VGND VPWR VPWR mux_right_track_24.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
Xclkbuf_2_2_0_mem_bottom_track_1.prog_clk clkbuf_2_3_0_mem_bottom_track_1.prog_clk/A
+ VGND VGND VPWR VPWR clkbuf_2_2_0_mem_bottom_track_1.prog_clk/X sky130_fd_sc_hd__clkbuf_1
XFILLER_14_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_right_track_32.mux_l1_in_0__A1 right_bottom_grid_pin_37_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
X_73_ _73_/A VGND VGND VPWR VPWR chany_bottom_out[4] sky130_fd_sc_hd__buf_2
XFILLER_27_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_70 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_81 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_92 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_56_ _56_/A VGND VGND VPWR VPWR chanx_right_out[7] sky130_fd_sc_hd__buf_2
XFILLER_24_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_right_track_24.mux_l1_in_1_ _25_/HI chany_bottom_in[6] mux_right_track_24.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_right_track_24.mux_l1_in_1_/X sky130_fd_sc_hd__mux2_1
X_39_ VGND VGND VPWR VPWR _39_/HI _39_/LO sky130_fd_sc_hd__conb_1
Xmem_right_track_32.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_2_1_0_mem_bottom_track_1.prog_clk/X
+ mux_right_track_32.mux_l1_in_0_/S VGND VGND VPWR VPWR mux_right_track_32.mux_l2_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_32_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_right_track_12.sky130_fd_sc_hd__buf_4_0_ mux_right_track_12.mux_l2_in_0_/X VGND
+ VGND VPWR VPWR _55_/A sky130_fd_sc_hd__buf_4
XFILLER_12_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__70__A chanx_right_in[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_72_ chanx_right_in[15] VGND VGND VPWR VPWR chany_bottom_out[3] sky130_fd_sc_hd__buf_2
XFILLER_27_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_71 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_82 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_93 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_55_ _55_/A VGND VGND VPWR VPWR chanx_right_out[6] sky130_fd_sc_hd__buf_2
XFILLER_24_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_right_track_24.mux_l1_in_0_ right_bottom_grid_pin_41_ right_top_grid_pin_1_ mux_right_track_24.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_right_track_24.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_23_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_right_track_36.mux_l2_in_0_ _31_/HI mux_right_track_36.mux_l1_in_0_/X mux_right_track_36.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR mux_right_track_36.mux_l2_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_11_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_right_track_32.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_2_1_0_mem_bottom_track_1.prog_clk/X
+ mux_right_track_30.mux_l2_in_0_/S VGND VGND VPWR VPWR mux_right_track_32.mux_l1_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_20_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_38_ VGND VGND VPWR VPWR _38_/HI _38_/LO sky130_fd_sc_hd__conb_1
XFILLER_19_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_bottom_track_1.mux_l2_in_0_ _36_/HI mux_bottom_track_1.mux_l1_in_0_/X mux_bottom_track_1.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR mux_bottom_track_1.mux_l2_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_11_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmem_right_track_38.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_2_3_0_mem_bottom_track_1.prog_clk/X
+ mux_right_track_38.mux_l1_in_0_/S VGND VGND VPWR VPWR mux_right_track_38.mux_l2_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_3_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_right_track_34.sky130_fd_sc_hd__buf_4_0_ mux_right_track_34.mux_l2_in_0_/X VGND
+ VGND VPWR VPWR _66_/A sky130_fd_sc_hd__buf_4
Xmem_right_track_0.sky130_fd_sc_hd__dfxtp_1_2_ clkbuf_2_2_0_mem_bottom_track_1.prog_clk/X
+ mux_right_track_0.mux_l2_in_0_/S VGND VGND VPWR VPWR mux_right_track_0.mux_l3_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA_mux_right_track_2.mux_l1_in_0__A0 right_bottom_grid_pin_36_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
X_71_ _71_/A VGND VGND VPWR VPWR chany_bottom_out[2] sky130_fd_sc_hd__buf_2
XFILLER_27_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_72 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_83 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_94 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_right_track_28.sky130_fd_sc_hd__buf_4_0_ mux_right_track_28.mux_l2_in_0_/X VGND
+ VGND VPWR VPWR _63_/A sky130_fd_sc_hd__buf_4
X_54_ _54_/A VGND VGND VPWR VPWR chanx_right_out[5] sky130_fd_sc_hd__buf_2
XFILLER_2_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mux_right_track_0.mux_l1_in_2__A0 chany_bottom_in[18] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_23_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__76__A chanx_right_in[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_37_ VGND VGND VPWR VPWR _37_/HI _37_/LO sky130_fd_sc_hd__conb_1
Xmux_bottom_track_1.sky130_fd_sc_hd__buf_4_0_ mux_bottom_track_1.mux_l2_in_0_/X VGND
+ VGND VPWR VPWR _69_/A sky130_fd_sc_hd__buf_4
XFILLER_11_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_right_track_36.mux_l1_in_0_ chany_bottom_in[0] right_bottom_grid_pin_39_ mux_right_track_36.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_right_track_36.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_31_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmem_right_track_38.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_2_3_0_mem_bottom_track_1.prog_clk/X
+ mux_right_track_36.mux_l2_in_0_/S VGND VGND VPWR VPWR mux_right_track_38.mux_l1_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
Xmux_bottom_track_1.mux_l1_in_0_ bottom_left_grid_pin_1_ chanx_right_in[18] mux_bottom_track_1.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_bottom_track_1.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__84__A chanx_right_in[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_right_track_0.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_2_2_0_mem_bottom_track_1.prog_clk/X
+ mux_right_track_0.mux_l1_in_1_/S VGND VGND VPWR VPWR mux_right_track_0.mux_l2_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__79__A chanx_right_in[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_2.mux_l1_in_0__A1 right_bottom_grid_pin_34_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_70_ chanx_right_in[17] VGND VGND VPWR VPWR chany_bottom_out[1] sky130_fd_sc_hd__buf_2
XFILLER_18_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_53_ _53_/A VGND VGND VPWR VPWR chanx_right_out[4] sky130_fd_sc_hd__buf_2
XPHY_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_track_0.mux_l1_in_2__A1 right_bottom_grid_pin_41_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XPHY_95 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_73 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_84 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_0_mem_bottom_track_1.prog_clk prog_clk_0_FTB00/X VGND VGND VPWR VPWR clkbuf_0_mem_bottom_track_1.prog_clk/X
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_14_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_right_track_6.sky130_fd_sc_hd__dfxtp_1_2_ clkbuf_2_0_0_mem_bottom_track_1.prog_clk/X
+ mux_right_track_6.mux_l2_in_1_/S VGND VGND VPWR VPWR mux_right_track_6.mux_l3_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_28_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_36_ VGND VGND VPWR VPWR _36_/HI _36_/LO sky130_fd_sc_hd__conb_1
XFILLER_11_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__87__A chanx_right_in[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_right_track_0.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_2_3_0_mem_bottom_track_1.prog_clk/X
+ ccff_head VGND VGND VPWR VPWR mux_right_track_0.mux_l1_in_1_/S sky130_fd_sc_hd__dfxtp_1
XFILLER_10_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_track_38.mux_l1_in_0__A0 chany_bottom_in[19] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XPHY_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_52_ _52_/A VGND VGND VPWR VPWR chanx_right_out[3] sky130_fd_sc_hd__buf_2
XFILLER_18_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_74 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_85 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_96 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_right_track_6.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_2_2_0_mem_bottom_track_1.prog_clk/X
+ mux_right_track_6.mux_l1_in_0_/S VGND VGND VPWR VPWR mux_right_track_6.mux_l2_in_1_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_14_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_35_ VGND VGND VPWR VPWR _35_/HI _35_/LO sky130_fd_sc_hd__conb_1
XFILLER_28_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_2_1_0_mem_bottom_track_1.prog_clk clkbuf_2_1_0_mem_bottom_track_1.prog_clk/A
+ VGND VGND VPWR VPWR clkbuf_2_1_0_mem_bottom_track_1.prog_clk/X sky130_fd_sc_hd__clkbuf_1
XANTENNA_mux_right_track_4.mux_l1_in_1__A0 right_bottom_grid_pin_39_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_right_track_38.mux_l1_in_0__A1 right_bottom_grid_pin_40_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XPHY_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_75 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_86 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_97 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_51_ _51_/A VGND VGND VPWR VPWR chanx_right_out[2] sky130_fd_sc_hd__buf_2
XFILLER_2_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmem_right_track_24.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_2_0_0_mem_bottom_track_1.prog_clk/X
+ mux_right_track_24.mux_l1_in_0_/S VGND VGND VPWR VPWR mux_right_track_24.mux_l2_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
Xmux_right_track_6.mux_l3_in_0_ mux_right_track_6.mux_l2_in_1_/X mux_right_track_6.mux_l2_in_0_/X
+ mux_right_track_6.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_right_track_6.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
Xmem_right_track_6.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_2_2_0_mem_bottom_track_1.prog_clk/X
+ mux_right_track_4.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_right_track_6.mux_l1_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
X_34_ VGND VGND VPWR VPWR _34_/HI _34_/LO sky130_fd_sc_hd__conb_1
XFILLER_9_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_right_track_6.mux_l2_in_1_ _34_/HI chany_bottom_in[15] mux_right_track_6.mux_l2_in_1_/S
+ VGND VGND VPWR VPWR mux_right_track_6.mux_l2_in_1_/X sky130_fd_sc_hd__mux2_1
XFILLER_6_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_track_4.mux_l1_in_1__A1 right_bottom_grid_pin_37_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_bottom_track_5.mux_l1_in_0__A0 bottom_left_grid_pin_1_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_12.mux_l1_in_0__A0 chany_bottom_in[12] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XPHY_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_76 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_87 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_98 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_50_ _50_/A VGND VGND VPWR VPWR chanx_right_out[1] sky130_fd_sc_hd__buf_2
Xmem_right_track_24.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_2_1_0_mem_bottom_track_1.prog_clk/X
+ mux_right_track_22.mux_l2_in_0_/S VGND VGND VPWR VPWR mux_right_track_24.mux_l1_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_23_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_33_ VGND VGND VPWR VPWR _33_/HI _33_/LO sky130_fd_sc_hd__conb_1
XFILLER_22_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_right_track_18.mux_l2_in_0_ _45_/HI mux_right_track_18.mux_l1_in_0_/X mux_right_track_18.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR mux_right_track_18.mux_l2_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_8_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmux_right_track_6.mux_l2_in_0_ mux_right_track_6.mux_l1_in_1_/X mux_right_track_6.mux_l1_in_0_/X
+ mux_right_track_6.mux_l2_in_1_/S VGND VGND VPWR VPWR mux_right_track_6.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_6_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_right_track_20.mux_l2_in_0_ _47_/HI mux_right_track_20.mux_l1_in_0_/X mux_right_track_20.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR mux_right_track_20.mux_l2_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_30_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_2_3_0_mem_bottom_track_1.prog_clk/X
+ mux_bottom_track_1.mux_l1_in_0_/S VGND VGND VPWR VPWR mux_bottom_track_1.mux_l2_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_12_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mux_right_track_20.mux_l1_in_0__A0 chany_bottom_in[8] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
Xmux_right_track_6.mux_l1_in_1_ right_bottom_grid_pin_40_ right_bottom_grid_pin_38_
+ mux_right_track_6.mux_l1_in_0_/S VGND VGND VPWR VPWR mux_right_track_6.mux_l1_in_1_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_30_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_bottom_track_5.mux_l1_in_0__A1 chanx_right_in[16] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_12.mux_l1_in_0__A1 right_bottom_grid_pin_35_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_8.mux_l1_in_0__A0 right_bottom_grid_pin_41_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XPHY_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_99 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_77 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_88 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_32_ VGND VGND VPWR VPWR _32_/HI _32_/LO sky130_fd_sc_hd__conb_1
XFILLER_20_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_right_track_20.mux_l1_in_0__A1 right_bottom_grid_pin_39_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xmux_right_track_18.mux_l1_in_0_ chany_bottom_in[9] right_bottom_grid_pin_38_ mux_right_track_18.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_right_track_18.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_5_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_2_3_0_mem_bottom_track_1.prog_clk/X
+ mux_right_track_38.mux_l2_in_0_/S VGND VGND VPWR VPWR mux_bottom_track_1.mux_l1_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
Xmux_right_track_20.mux_l1_in_0_ chany_bottom_in[8] right_bottom_grid_pin_39_ mux_right_track_20.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_right_track_20.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
Xmux_bottom_track_25.sky130_fd_sc_hd__buf_4_0_ mux_bottom_track_25.mux_l2_in_0_/X
+ VGND VGND VPWR VPWR _81_/A sky130_fd_sc_hd__buf_4
Xmux_right_track_6.mux_l1_in_0_ right_bottom_grid_pin_36_ right_bottom_grid_pin_34_
+ mux_right_track_6.mux_l1_in_0_/S VGND VGND VPWR VPWR mux_right_track_6.mux_l1_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_5_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_right_track_6.sky130_fd_sc_hd__buf_4_0_ mux_right_track_6.mux_l3_in_0_/X VGND
+ VGND VPWR VPWR _52_/A sky130_fd_sc_hd__buf_4
XFILLER_14_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_right_track_32.mux_l2_in_0_ _29_/HI mux_right_track_32.mux_l1_in_0_/X mux_right_track_32.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR mux_right_track_32.mux_l2_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_29_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_right_track_8.mux_l1_in_0__A1 right_top_grid_pin_1_ VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XPHY_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_78 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_89 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_31_ VGND VGND VPWR VPWR _31_/HI _31_/LO sky130_fd_sc_hd__conb_1
Xmux_right_track_30.sky130_fd_sc_hd__buf_4_0_ mux_right_track_30.mux_l2_in_0_/X VGND
+ VGND VPWR VPWR _64_/A sky130_fd_sc_hd__buf_4
XFILLER_22_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_right_track_6.mux_l2_in_1__A1 chany_bottom_in[15] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_33_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_right_track_24.sky130_fd_sc_hd__buf_4_0_ mux_right_track_24.mux_l2_in_0_/X VGND
+ VGND VPWR VPWR _61_/A sky130_fd_sc_hd__buf_4
Xmem_right_track_10.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_2_0_0_mem_bottom_track_1.prog_clk/X
+ mux_right_track_10.mux_l1_in_0_/S VGND VGND VPWR VPWR mux_right_track_10.mux_l2_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_28_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_right_track_18.sky130_fd_sc_hd__buf_4_0_ mux_right_track_18.mux_l2_in_0_/X VGND
+ VGND VPWR VPWR _58_/A sky130_fd_sc_hd__buf_4
XFILLER_29_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_68 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_79 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_right_track_32.mux_l1_in_0_ chany_bottom_in[2] right_bottom_grid_pin_37_ mux_right_track_32.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_right_track_32.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
Xclkbuf_2_0_0_mem_bottom_track_1.prog_clk clkbuf_2_1_0_mem_bottom_track_1.prog_clk/A
+ VGND VGND VPWR VPWR clkbuf_2_0_0_mem_bottom_track_1.prog_clk/X sky130_fd_sc_hd__clkbuf_1
XFILLER_20_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_30_ VGND VGND VPWR VPWR _30_/HI _30_/LO sky130_fd_sc_hd__conb_1
XFILLER_13_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmem_right_track_10.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_2_0_0_mem_bottom_track_1.prog_clk/X
+ mux_right_track_8.mux_l2_in_0_/S VGND VGND VPWR VPWR mux_right_track_10.mux_l1_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_28_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmem_right_track_16.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_2_1_0_mem_bottom_track_1.prog_clk/X
+ mux_right_track_16.mux_l1_in_0_/S VGND VGND VPWR VPWR mux_right_track_16.mux_l2_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_1_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_69 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_right_track_0.sky130_fd_sc_hd__dfxtp_1_0__D ccff_head VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mux_right_track_18.mux_l1_in_0__A0 chany_bottom_in[9] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
Xmem_right_track_16.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_2_1_0_mem_bottom_track_1.prog_clk/X
+ mux_right_track_14.mux_l2_in_0_/S VGND VGND VPWR VPWR mux_right_track_16.mux_l1_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XPHY_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_88_ chanx_right_in[19] VGND VGND VPWR VPWR chany_bottom_out[19] sky130_fd_sc_hd__buf_2
XFILLER_13_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_track_26.mux_l1_in_0__A0 chany_bottom_in[5] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_30_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_right_track_2.mux_l3_in_0_ mux_right_track_2.mux_l2_in_1_/X mux_right_track_2.mux_l2_in_0_/X
+ mux_right_track_2.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_right_track_2.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_20_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mux_right_track_18.mux_l1_in_0__A1 right_bottom_grid_pin_38_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XPHY_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_right_track_2.mux_l2_in_1_ _46_/HI chany_bottom_in[17] mux_right_track_2.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR mux_right_track_2.mux_l2_in_1_/X sky130_fd_sc_hd__mux2_1
XFILLER_14_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_87_ chanx_right_in[0] VGND VGND VPWR VPWR chany_bottom_out[18] sky130_fd_sc_hd__buf_2
XFILLER_6_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mux_right_track_34.mux_l1_in_0__A0 chany_bottom_in[1] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_9_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmem_right_track_34.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_2_1_0_mem_bottom_track_1.prog_clk/X
+ mux_right_track_34.mux_l1_in_0_/S VGND VGND VPWR VPWR mux_right_track_34.mux_l2_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
Xclkbuf_1_1_0_mem_bottom_track_1.prog_clk clkbuf_0_mem_bottom_track_1.prog_clk/X VGND
+ VGND VPWR VPWR clkbuf_2_3_0_mem_bottom_track_1.prog_clk/A sky130_fd_sc_hd__clkbuf_1
XFILLER_18_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_right_track_26.mux_l1_in_0__A1 right_bottom_grid_pin_34_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_right_track_14.mux_l2_in_0_ _43_/HI mux_right_track_14.mux_l1_in_0_/X mux_right_track_14.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR mux_right_track_14.mux_l2_in_0_/X sky130_fd_sc_hd__mux2_1
XANTENNA_mux_right_track_0.mux_l1_in_1__A0 right_bottom_grid_pin_39_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmux_right_track_2.mux_l2_in_0_ mux_right_track_2.mux_l1_in_1_/X mux_right_track_2.mux_l1_in_0_/X
+ mux_right_track_2.mux_l2_in_0_/S VGND VGND VPWR VPWR mux_right_track_2.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_26_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_86_ chanx_right_in[1] VGND VGND VPWR VPWR chany_bottom_out[17] sky130_fd_sc_hd__buf_2
XFILLER_27_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_right_track_2.mux_l1_in_1_ right_bottom_grid_pin_40_ right_bottom_grid_pin_38_
+ mux_right_track_2.mux_l1_in_0_/S VGND VGND VPWR VPWR mux_right_track_2.mux_l1_in_1_/X
+ sky130_fd_sc_hd__mux2_1
X_69_ _69_/A VGND VGND VPWR VPWR chany_bottom_out[0] sky130_fd_sc_hd__buf_2
XANTENNA_mux_right_track_34.mux_l1_in_0__A1 right_bottom_grid_pin_38_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_right_track_34.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_2_1_0_mem_bottom_track_1.prog_clk/X
+ mux_right_track_32.mux_l2_in_0_/S VGND VGND VPWR VPWR mux_right_track_34.mux_l1_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_9_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__74__A chanx_right_in[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_mux_right_track_0.mux_l1_in_1__A1 right_bottom_grid_pin_37_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmem_right_track_2.sky130_fd_sc_hd__dfxtp_1_2_ clkbuf_2_2_0_mem_bottom_track_1.prog_clk/X
+ mux_right_track_2.mux_l2_in_0_/S VGND VGND VPWR VPWR mux_right_track_2.mux_l3_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__82__A chanx_right_in[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_85_ chanx_right_in[2] VGND VGND VPWR VPWR chany_bottom_out[16] sky130_fd_sc_hd__buf_2
Xmux_right_track_2.sky130_fd_sc_hd__buf_4_0_ mux_right_track_2.mux_l3_in_0_/X VGND
+ VGND VPWR VPWR _50_/A sky130_fd_sc_hd__buf_4
XFILLER_12_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_right_track_14.mux_l1_in_0_ chany_bottom_in[11] right_bottom_grid_pin_36_ mux_right_track_14.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_right_track_14.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_6_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_bottom_track_1.mux_l1_in_0__A0 bottom_left_grid_pin_1_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA__77__A chanx_right_in[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_right_track_26.mux_l2_in_0_ _26_/HI mux_right_track_26.mux_l1_in_0_/X mux_right_track_26.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR mux_right_track_26.mux_l2_in_0_/X sky130_fd_sc_hd__mux2_1
Xmux_right_track_2.mux_l1_in_0_ right_bottom_grid_pin_36_ right_bottom_grid_pin_34_
+ mux_right_track_2.mux_l1_in_0_/S VGND VGND VPWR VPWR mux_right_track_2.mux_l1_in_0_/X
+ sky130_fd_sc_hd__mux2_1
X_68_ _68_/A VGND VGND VPWR VPWR chanx_right_out[19] sky130_fd_sc_hd__buf_2
XFILLER_23_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__85__A chanx_right_in[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmux_right_track_20.sky130_fd_sc_hd__buf_4_0_ mux_right_track_20.mux_l2_in_0_/X VGND
+ VGND VPWR VPWR _59_/A sky130_fd_sc_hd__buf_4
XFILLER_25_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmem_right_track_2.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_2_2_0_mem_bottom_track_1.prog_clk/X
+ mux_right_track_2.mux_l1_in_0_/S VGND VGND VPWR VPWR mux_right_track_2.mux_l2_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_13_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_84_ chanx_right_in[3] VGND VGND VPWR VPWR chany_bottom_out[15] sky130_fd_sc_hd__buf_2
XFILLER_27_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_right_track_14.sky130_fd_sc_hd__buf_4_0_ mux_right_track_14.mux_l2_in_0_/X VGND
+ VGND VPWR VPWR _56_/A sky130_fd_sc_hd__buf_4
XANTENNA_mux_bottom_track_1.mux_l1_in_0__A1 chanx_right_in[18] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_5_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_67_ _67_/A VGND VGND VPWR VPWR chanx_right_out[18] sky130_fd_sc_hd__buf_2
XFILLER_30_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__88__A chanx_right_in[19] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_track_4.mux_l1_in_0__A0 right_bottom_grid_pin_35_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmux_right_track_26.mux_l1_in_0_ chany_bottom_in[5] right_bottom_grid_pin_34_ mux_right_track_26.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_right_track_26.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
Xmux_right_track_38.mux_l2_in_0_ _32_/HI mux_right_track_38.mux_l1_in_0_/X mux_right_track_38.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR mux_right_track_38.mux_l2_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_29_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
.ends

