VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sb_3__3_
  CLASS BLOCK ;
  FOREIGN sb_3__3_ ;
  ORIGIN 0.000 0.000 ;
  SIZE 140.000 BY 140.000 ;
  PIN address[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 4.690 137.600 4.970 140.000 ;
    END
  END address[0]
  PIN address[1]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 4.800 140.000 5.400 ;
    END
  END address[1]
  PIN address[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 24.470 0.000 24.750 2.400 ;
    END
  END address[2]
  PIN address[3]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 15.000 140.000 15.600 ;
    END
  END address[3]
  PIN address[4]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 2.760 2.400 3.360 ;
    END
  END address[4]
  PIN address[5]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 25.880 140.000 26.480 ;
    END
  END address[5]
  PIN bottom_left_grid_pin_13_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 34.590 0.000 34.870 2.400 ;
    END
  END bottom_left_grid_pin_13_
  PIN bottom_right_grid_pin_11_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 54.370 0.000 54.650 2.400 ;
    END
  END bottom_right_grid_pin_11_
  PIN bottom_right_grid_pin_13_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 22.480 2.400 23.080 ;
    END
  END bottom_right_grid_pin_13_
  PIN bottom_right_grid_pin_15_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 47.640 140.000 48.240 ;
    END
  END bottom_right_grid_pin_15_
  PIN bottom_right_grid_pin_1_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 8.880 2.400 9.480 ;
    END
  END bottom_right_grid_pin_1_
  PIN bottom_right_grid_pin_3_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 36.760 140.000 37.360 ;
    END
  END bottom_right_grid_pin_3_
  PIN bottom_right_grid_pin_5_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 44.250 0.000 44.530 2.400 ;
    END
  END bottom_right_grid_pin_5_
  PIN bottom_right_grid_pin_7_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 14.350 137.600 14.630 140.000 ;
    END
  END bottom_right_grid_pin_7_
  PIN bottom_right_grid_pin_9_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 15.680 2.400 16.280 ;
    END
  END bottom_right_grid_pin_9_
  PIN chanx_left_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 24.470 137.600 24.750 140.000 ;
    END
  END chanx_left_in[0]
  PIN chanx_left_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 29.280 2.400 29.880 ;
    END
  END chanx_left_in[1]
  PIN chanx_left_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 36.080 2.400 36.680 ;
    END
  END chanx_left_in[2]
  PIN chanx_left_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 64.490 0.000 64.770 2.400 ;
    END
  END chanx_left_in[3]
  PIN chanx_left_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 58.520 140.000 59.120 ;
    END
  END chanx_left_in[4]
  PIN chanx_left_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 34.590 137.600 34.870 140.000 ;
    END
  END chanx_left_in[5]
  PIN chanx_left_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 69.400 140.000 70.000 ;
    END
  END chanx_left_in[6]
  PIN chanx_left_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 42.200 2.400 42.800 ;
    END
  END chanx_left_in[7]
  PIN chanx_left_in[8]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 49.000 2.400 49.600 ;
    END
  END chanx_left_in[8]
  PIN chanx_left_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 44.250 137.600 44.530 140.000 ;
    END
  END chanx_left_out[0]
  PIN chanx_left_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 54.370 137.600 54.650 140.000 ;
    END
  END chanx_left_out[1]
  PIN chanx_left_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 55.800 2.400 56.400 ;
    END
  END chanx_left_out[2]
  PIN chanx_left_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 137.600 79.600 140.000 80.200 ;
    END
  END chanx_left_out[3]
  PIN chanx_left_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 74.610 0.000 74.890 2.400 ;
    END
  END chanx_left_out[4]
  PIN chanx_left_out[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 62.600 2.400 63.200 ;
    END
  END chanx_left_out[5]
  PIN chanx_left_out[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 84.270 0.000 84.550 2.400 ;
    END
  END chanx_left_out[6]
  PIN chanx_left_out[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 64.490 137.600 64.770 140.000 ;
    END
  END chanx_left_out[7]
  PIN chanx_left_out[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 69.400 2.400 70.000 ;
    END
  END chanx_left_out[8]
  PIN chany_bottom_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 74.610 137.600 74.890 140.000 ;
    END
  END chany_bottom_in[0]
  PIN chany_bottom_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 94.390 0.000 94.670 2.400 ;
    END
  END chany_bottom_in[1]
  PIN chany_bottom_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 75.520 2.400 76.120 ;
    END
  END chany_bottom_in[2]
  PIN chany_bottom_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 82.320 2.400 82.920 ;
    END
  END chany_bottom_in[3]
  PIN chany_bottom_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 89.120 2.400 89.720 ;
    END
  END chany_bottom_in[4]
  PIN chany_bottom_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 84.270 137.600 84.550 140.000 ;
    END
  END chany_bottom_in[5]
  PIN chany_bottom_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 104.510 0.000 104.790 2.400 ;
    END
  END chany_bottom_in[6]
  PIN chany_bottom_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 94.390 137.600 94.670 140.000 ;
    END
  END chany_bottom_in[7]
  PIN chany_bottom_in[8]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 90.480 140.000 91.080 ;
    END
  END chany_bottom_in[8]
  PIN chany_bottom_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 95.920 2.400 96.520 ;
    END
  END chany_bottom_out[0]
  PIN chany_bottom_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 104.510 137.600 104.790 140.000 ;
    END
  END chany_bottom_out[1]
  PIN chany_bottom_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 114.170 137.600 114.450 140.000 ;
    END
  END chany_bottom_out[2]
  PIN chany_bottom_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 137.600 101.360 140.000 101.960 ;
    END
  END chany_bottom_out[3]
  PIN chany_bottom_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 137.600 112.240 140.000 112.840 ;
    END
  END chany_bottom_out[4]
  PIN chany_bottom_out[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 102.720 2.400 103.320 ;
    END
  END chany_bottom_out[5]
  PIN chany_bottom_out[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 108.840 2.400 109.440 ;
    END
  END chany_bottom_out[6]
  PIN chany_bottom_out[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 114.170 0.000 114.450 2.400 ;
    END
  END chany_bottom_out[7]
  PIN chany_bottom_out[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 124.290 137.600 124.570 140.000 ;
    END
  END chany_bottom_out[8]
  PIN data_in
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 14.350 0.000 14.630 2.400 ;
    END
  END data_in
  PIN enable
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 4.690 0.000 4.970 2.400 ;
    END
  END enable
  PIN left_bottom_grid_pin_12_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 115.640 2.400 116.240 ;
    END
  END left_bottom_grid_pin_12_
  PIN left_top_grid_pin_11_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 124.290 0.000 124.570 2.400 ;
    END
  END left_top_grid_pin_11_
  PIN left_top_grid_pin_13_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 134.410 0.000 134.690 2.400 ;
    END
  END left_top_grid_pin_13_
  PIN left_top_grid_pin_15_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 136.040 2.400 136.640 ;
    END
  END left_top_grid_pin_15_
  PIN left_top_grid_pin_1_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 134.410 137.600 134.690 140.000 ;
    END
  END left_top_grid_pin_1_
  PIN left_top_grid_pin_3_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 123.120 140.000 123.720 ;
    END
  END left_top_grid_pin_3_
  PIN left_top_grid_pin_5_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 122.440 2.400 123.040 ;
    END
  END left_top_grid_pin_5_
  PIN left_top_grid_pin_7_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 129.240 2.400 129.840 ;
    END
  END left_top_grid_pin_7_
  PIN left_top_grid_pin_9_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 134.000 140.000 134.600 ;
    END
  END left_top_grid_pin_9_
  PIN vpwr
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT 28.055 10.640 29.655 128.080 ;
    END
  END vpwr
  PIN vgnd
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT 51.385 10.640 52.985 128.080 ;
    END
  END vgnd
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 134.320 127.925 ;
      LAYER met1 ;
        RECT 0.530 0.380 138.390 128.080 ;
      LAYER met2 ;
        RECT 0.550 137.320 4.410 137.770 ;
        RECT 5.250 137.320 14.070 137.770 ;
        RECT 14.910 137.320 24.190 137.770 ;
        RECT 25.030 137.320 34.310 137.770 ;
        RECT 35.150 137.320 43.970 137.770 ;
        RECT 44.810 137.320 54.090 137.770 ;
        RECT 54.930 137.320 64.210 137.770 ;
        RECT 65.050 137.320 74.330 137.770 ;
        RECT 75.170 137.320 83.990 137.770 ;
        RECT 84.830 137.320 94.110 137.770 ;
        RECT 94.950 137.320 104.230 137.770 ;
        RECT 105.070 137.320 113.890 137.770 ;
        RECT 114.730 137.320 124.010 137.770 ;
        RECT 124.850 137.320 134.130 137.770 ;
        RECT 134.970 137.320 138.370 137.770 ;
        RECT 0.550 2.680 138.370 137.320 ;
        RECT 0.550 0.155 4.410 2.680 ;
        RECT 5.250 0.155 14.070 2.680 ;
        RECT 14.910 0.155 24.190 2.680 ;
        RECT 25.030 0.155 34.310 2.680 ;
        RECT 35.150 0.155 43.970 2.680 ;
        RECT 44.810 0.155 54.090 2.680 ;
        RECT 54.930 0.155 64.210 2.680 ;
        RECT 65.050 0.155 74.330 2.680 ;
        RECT 75.170 0.155 83.990 2.680 ;
        RECT 84.830 0.155 94.110 2.680 ;
        RECT 94.950 0.155 104.230 2.680 ;
        RECT 105.070 0.155 113.890 2.680 ;
        RECT 114.730 0.155 124.010 2.680 ;
        RECT 124.850 0.155 134.130 2.680 ;
        RECT 134.970 0.155 138.370 2.680 ;
      LAYER met3 ;
        RECT 2.800 135.640 138.610 136.040 ;
        RECT 0.270 135.000 138.610 135.640 ;
        RECT 0.270 133.600 137.200 135.000 ;
        RECT 0.270 130.240 138.610 133.600 ;
        RECT 2.800 128.840 138.610 130.240 ;
        RECT 0.270 124.120 138.610 128.840 ;
        RECT 0.270 123.440 137.200 124.120 ;
        RECT 2.800 122.720 137.200 123.440 ;
        RECT 2.800 122.040 138.610 122.720 ;
        RECT 0.270 116.640 138.610 122.040 ;
        RECT 2.800 115.240 138.610 116.640 ;
        RECT 0.270 113.240 138.610 115.240 ;
        RECT 0.270 111.840 137.200 113.240 ;
        RECT 0.270 109.840 138.610 111.840 ;
        RECT 2.800 108.440 138.610 109.840 ;
        RECT 0.270 103.720 138.610 108.440 ;
        RECT 2.800 102.360 138.610 103.720 ;
        RECT 2.800 102.320 137.200 102.360 ;
        RECT 0.270 100.960 137.200 102.320 ;
        RECT 0.270 96.920 138.610 100.960 ;
        RECT 2.800 95.520 138.610 96.920 ;
        RECT 0.270 91.480 138.610 95.520 ;
        RECT 0.270 90.120 137.200 91.480 ;
        RECT 2.800 90.080 137.200 90.120 ;
        RECT 2.800 88.720 138.610 90.080 ;
        RECT 0.270 83.320 138.610 88.720 ;
        RECT 2.800 81.920 138.610 83.320 ;
        RECT 0.270 80.600 138.610 81.920 ;
        RECT 0.270 79.200 137.200 80.600 ;
        RECT 0.270 76.520 138.610 79.200 ;
        RECT 2.800 75.120 138.610 76.520 ;
        RECT 0.270 70.400 138.610 75.120 ;
        RECT 2.800 69.000 137.200 70.400 ;
        RECT 0.270 63.600 138.610 69.000 ;
        RECT 2.800 62.200 138.610 63.600 ;
        RECT 0.270 59.520 138.610 62.200 ;
        RECT 0.270 58.120 137.200 59.520 ;
        RECT 0.270 56.800 138.610 58.120 ;
        RECT 2.800 55.400 138.610 56.800 ;
        RECT 0.270 50.000 138.610 55.400 ;
        RECT 2.800 48.640 138.610 50.000 ;
        RECT 2.800 48.600 137.200 48.640 ;
        RECT 0.270 47.240 137.200 48.600 ;
        RECT 0.270 43.200 138.610 47.240 ;
        RECT 2.800 41.800 138.610 43.200 ;
        RECT 0.270 37.760 138.610 41.800 ;
        RECT 0.270 37.080 137.200 37.760 ;
        RECT 2.800 36.360 137.200 37.080 ;
        RECT 2.800 35.680 138.610 36.360 ;
        RECT 0.270 30.280 138.610 35.680 ;
        RECT 2.800 28.880 138.610 30.280 ;
        RECT 0.270 26.880 138.610 28.880 ;
        RECT 0.270 25.480 137.200 26.880 ;
        RECT 0.270 23.480 138.610 25.480 ;
        RECT 2.800 22.080 138.610 23.480 ;
        RECT 0.270 16.680 138.610 22.080 ;
        RECT 2.800 16.000 138.610 16.680 ;
        RECT 2.800 15.280 137.200 16.000 ;
        RECT 0.270 14.600 137.200 15.280 ;
        RECT 0.270 9.880 138.610 14.600 ;
        RECT 2.800 8.480 138.610 9.880 ;
        RECT 0.270 5.800 138.610 8.480 ;
        RECT 0.270 4.400 137.200 5.800 ;
        RECT 0.270 3.760 138.610 4.400 ;
        RECT 2.800 2.360 138.610 3.760 ;
        RECT 0.270 0.175 138.610 2.360 ;
      LAYER met4 ;
        RECT 0.295 10.640 27.655 128.080 ;
        RECT 30.055 10.640 50.985 128.080 ;
        RECT 53.385 10.640 122.985 128.080 ;
  END
END sb_3__3_
END LIBRARY

