magic
tech EFS8A
magscale 1 2
timestamp 1604337736
<< locali >>
rect 31493 12631 31527 12733
rect 34069 12087 34103 12325
rect 4353 11611 4387 11781
rect 12541 7259 12575 7361
rect 25053 6715 25087 6953
rect 16129 4675 16163 4777
<< viali >>
rect 5365 13481 5399 13515
rect 7113 13481 7147 13515
rect 34437 13481 34471 13515
rect 2973 13413 3007 13447
rect 1409 13345 1443 13379
rect 2697 13345 2731 13379
rect 3433 13345 3467 13379
rect 4077 13345 4111 13379
rect 5181 13345 5215 13379
rect 6929 13345 6963 13379
rect 24041 13345 24075 13379
rect 24317 13345 24351 13379
rect 33149 13345 33183 13379
rect 33701 13345 33735 13379
rect 34253 13345 34287 13379
rect 35449 13345 35483 13379
rect 36559 13345 36593 13379
rect 33333 13209 33367 13243
rect 1593 13141 1627 13175
rect 4261 13141 4295 13175
rect 24869 13141 24903 13175
rect 34069 13141 34103 13175
rect 34897 13141 34931 13175
rect 35633 13141 35667 13175
rect 36737 13141 36771 13175
rect 1593 12937 1627 12971
rect 8309 12937 8343 12971
rect 36369 12937 36403 12971
rect 37105 12937 37139 12971
rect 4261 12869 4295 12903
rect 24593 12869 24627 12903
rect 32321 12869 32355 12903
rect 33333 12869 33367 12903
rect 2145 12801 2179 12835
rect 7113 12801 7147 12835
rect 13277 12801 13311 12835
rect 16497 12801 16531 12835
rect 19073 12801 19107 12835
rect 22109 12801 22143 12835
rect 25145 12801 25179 12835
rect 27629 12801 27663 12835
rect 31125 12801 31159 12835
rect 33793 12801 33827 12835
rect 34621 12801 34655 12835
rect 35173 12801 35207 12835
rect 1869 12733 1903 12767
rect 2605 12733 2639 12767
rect 3709 12733 3743 12767
rect 6653 12733 6687 12767
rect 6837 12733 6871 12767
rect 8125 12733 8159 12767
rect 8677 12733 8711 12767
rect 10333 12733 10367 12767
rect 13001 12733 13035 12767
rect 13737 12733 13771 12767
rect 16221 12733 16255 12767
rect 16957 12733 16991 12767
rect 18797 12733 18831 12767
rect 19533 12733 19567 12767
rect 21833 12733 21867 12767
rect 22661 12733 22695 12767
rect 27353 12733 27387 12767
rect 30849 12733 30883 12767
rect 31493 12733 31527 12767
rect 31585 12733 31619 12767
rect 32137 12733 32171 12767
rect 32689 12733 32723 12767
rect 34897 12733 34931 12767
rect 36185 12733 36219 12767
rect 36737 12733 36771 12767
rect 37289 12733 37323 12767
rect 37841 12733 37875 12767
rect 3341 12665 3375 12699
rect 4537 12665 4571 12699
rect 4813 12665 4847 12699
rect 5273 12665 5307 12699
rect 10609 12665 10643 12699
rect 11161 12665 11195 12699
rect 24041 12665 24075 12699
rect 24869 12665 24903 12699
rect 28181 12665 28215 12699
rect 33885 12665 33919 12699
rect 3985 12597 4019 12631
rect 4721 12597 4755 12631
rect 5549 12597 5583 12631
rect 5733 12597 5767 12631
rect 7573 12597 7607 12631
rect 23489 12597 23523 12631
rect 24409 12597 24443 12631
rect 25053 12597 25087 12631
rect 31493 12597 31527 12631
rect 33149 12597 33183 12631
rect 33793 12597 33827 12631
rect 34345 12597 34379 12631
rect 35633 12597 35667 12631
rect 37473 12597 37507 12631
rect 6653 12393 6687 12427
rect 31125 12393 31159 12427
rect 32321 12393 32355 12427
rect 36185 12393 36219 12427
rect 1685 12325 1719 12359
rect 4813 12325 4847 12359
rect 5457 12325 5491 12359
rect 8493 12325 8527 12359
rect 11989 12325 12023 12359
rect 17785 12325 17819 12359
rect 21465 12325 21499 12359
rect 24961 12325 24995 12359
rect 33793 12325 33827 12359
rect 34069 12325 34103 12359
rect 1409 12257 1443 12291
rect 2513 12257 2547 12291
rect 2697 12257 2731 12291
rect 6469 12257 6503 12291
rect 8309 12257 8343 12291
rect 30941 12257 30975 12291
rect 32137 12257 32171 12291
rect 33609 12257 33643 12291
rect 5365 12189 5399 12223
rect 5549 12189 5583 12223
rect 8585 12189 8619 12223
rect 11897 12189 11931 12223
rect 12081 12189 12115 12223
rect 17785 12189 17819 12223
rect 17877 12189 17911 12223
rect 21465 12189 21499 12223
rect 21557 12189 21591 12223
rect 24961 12189 24995 12223
rect 25053 12189 25087 12223
rect 33885 12189 33919 12223
rect 23673 12121 23707 12155
rect 24501 12121 24535 12155
rect 33333 12121 33367 12155
rect 34621 12257 34655 12291
rect 35061 12257 35095 12291
rect 34805 12189 34839 12223
rect 2237 12053 2271 12087
rect 2881 12053 2915 12087
rect 3617 12053 3651 12087
rect 4353 12053 4387 12087
rect 4997 12053 5031 12087
rect 5917 12053 5951 12087
rect 7757 12053 7791 12087
rect 8033 12053 8067 12087
rect 8953 12053 8987 12087
rect 11161 12053 11195 12087
rect 11529 12053 11563 12087
rect 13001 12053 13035 12087
rect 16405 12053 16439 12087
rect 16957 12053 16991 12087
rect 17325 12053 17359 12087
rect 19441 12053 19475 12087
rect 21005 12053 21039 12087
rect 24041 12053 24075 12087
rect 25605 12053 25639 12087
rect 27169 12053 27203 12087
rect 30205 12053 30239 12087
rect 30573 12053 30607 12087
rect 32781 12053 32815 12087
rect 33149 12053 33183 12087
rect 34069 12053 34103 12087
rect 34345 12053 34379 12087
rect 3617 11849 3651 11883
rect 5181 11849 5215 11883
rect 7021 11849 7055 11883
rect 10701 11849 10735 11883
rect 17509 11849 17543 11883
rect 25053 11849 25087 11883
rect 26525 11849 26559 11883
rect 29561 11849 29595 11883
rect 31953 11849 31987 11883
rect 33333 11849 33367 11883
rect 34345 11849 34379 11883
rect 36277 11849 36311 11883
rect 2053 11781 2087 11815
rect 3065 11781 3099 11815
rect 4353 11781 4387 11815
rect 8217 11781 8251 11815
rect 13001 11781 13035 11815
rect 16497 11781 16531 11815
rect 24041 11781 24075 11815
rect 25605 11781 25639 11815
rect 27169 11781 27203 11815
rect 30573 11781 30607 11815
rect 34989 11781 35023 11815
rect 1869 11713 1903 11747
rect 2513 11713 2547 11747
rect 2605 11713 2639 11747
rect 4077 11713 4111 11747
rect 5733 11713 5767 11747
rect 7941 11713 7975 11747
rect 8677 11713 8711 11747
rect 9505 11713 9539 11747
rect 11345 11713 11379 11747
rect 16957 11713 16991 11747
rect 18061 11713 18095 11747
rect 24409 11713 24443 11747
rect 24593 11713 24627 11747
rect 25973 11713 26007 11747
rect 27721 11713 27755 11747
rect 33793 11713 33827 11747
rect 37565 11713 37599 11747
rect 6101 11645 6135 11679
rect 6837 11645 6871 11679
rect 11069 11645 11103 11679
rect 12265 11645 12299 11679
rect 13553 11645 13587 11679
rect 19349 11645 19383 11679
rect 19441 11645 19475 11679
rect 29377 11645 29411 11679
rect 29929 11645 29963 11679
rect 30849 11645 30883 11679
rect 32137 11645 32171 11679
rect 33885 11645 33919 11679
rect 36461 11645 36495 11679
rect 37013 11645 37047 11679
rect 2513 11577 2547 11611
rect 3433 11577 3467 11611
rect 4169 11577 4203 11611
rect 4353 11577 4387 11611
rect 4629 11577 4663 11611
rect 5457 11577 5491 11611
rect 8769 11577 8803 11611
rect 13277 11577 13311 11611
rect 15393 11577 15427 11611
rect 17049 11577 17083 11611
rect 18613 11577 18647 11611
rect 19686 11577 19720 11611
rect 23121 11577 23155 11611
rect 24501 11577 24535 11611
rect 26157 11577 26191 11611
rect 27445 11577 27479 11611
rect 31033 11577 31067 11611
rect 31125 11577 31159 11611
rect 34621 11577 34655 11611
rect 35265 11577 35299 11611
rect 35541 11577 35575 11611
rect 4077 11509 4111 11543
rect 4905 11509 4939 11543
rect 5641 11509 5675 11543
rect 6469 11509 6503 11543
rect 7481 11509 7515 11543
rect 8677 11509 8711 11543
rect 9137 11509 9171 11543
rect 11897 11509 11931 11543
rect 12725 11509 12759 11543
rect 13461 11509 13495 11543
rect 15945 11509 15979 11543
rect 16313 11509 16347 11543
rect 16957 11509 16991 11543
rect 17877 11509 17911 11543
rect 20821 11509 20855 11543
rect 21373 11509 21407 11543
rect 21741 11509 21775 11543
rect 22109 11509 22143 11543
rect 22753 11509 22787 11543
rect 23489 11509 23523 11543
rect 25329 11509 25363 11543
rect 26065 11509 26099 11543
rect 26985 11509 27019 11543
rect 27629 11509 27663 11543
rect 30389 11509 30423 11543
rect 31493 11509 31527 11543
rect 32321 11509 32355 11543
rect 32781 11509 32815 11543
rect 33149 11509 33183 11543
rect 33793 11509 33827 11543
rect 35449 11509 35483 11543
rect 36001 11509 36035 11543
rect 36645 11509 36679 11543
rect 2053 11305 2087 11339
rect 5457 11305 5491 11339
rect 8309 11305 8343 11339
rect 15853 11305 15887 11339
rect 16497 11305 16531 11339
rect 17417 11305 17451 11339
rect 22937 11305 22971 11339
rect 23949 11305 23983 11339
rect 2973 11237 3007 11271
rect 7113 11237 7147 11271
rect 9956 11237 9990 11271
rect 13001 11237 13035 11271
rect 13461 11237 13495 11271
rect 17233 11237 17267 11271
rect 18503 11237 18537 11271
rect 18981 11237 19015 11271
rect 19073 11237 19107 11271
rect 21158 11237 21192 11271
rect 25237 11237 25271 11271
rect 27077 11237 27111 11271
rect 30941 11237 30975 11271
rect 32873 11237 32907 11271
rect 33232 11237 33266 11271
rect 35817 11237 35851 11271
rect 36001 11237 36035 11271
rect 4077 11169 4111 11203
rect 4333 11169 4367 11203
rect 6101 11169 6135 11203
rect 6469 11169 6503 11203
rect 8125 11169 8159 11203
rect 11989 11169 12023 11203
rect 12817 11169 12851 11203
rect 13829 11169 13863 11203
rect 20913 11169 20947 11203
rect 23765 11169 23799 11203
rect 24961 11169 24995 11203
rect 26249 11169 26283 11203
rect 26893 11169 26927 11203
rect 28448 11169 28482 11203
rect 30665 11169 30699 11203
rect 31953 11169 31987 11203
rect 35357 11169 35391 11203
rect 1409 11101 1443 11135
rect 2973 11101 3007 11135
rect 3065 11101 3099 11135
rect 7021 11101 7055 11135
rect 7205 11101 7239 11135
rect 8769 11101 8803 11135
rect 9689 11101 9723 11135
rect 11713 11101 11747 11135
rect 13093 11101 13127 11135
rect 15025 11101 15059 11135
rect 15761 11101 15795 11135
rect 15945 11101 15979 11135
rect 17509 11101 17543 11135
rect 18061 11101 18095 11135
rect 18889 11101 18923 11135
rect 24041 11101 24075 11135
rect 27169 11101 27203 11135
rect 28181 11101 28215 11135
rect 32965 11101 32999 11135
rect 36093 11101 36127 11135
rect 2513 11033 2547 11067
rect 3617 11033 3651 11067
rect 6653 11033 6687 11067
rect 8033 11033 8067 11067
rect 11069 11033 11103 11067
rect 12541 11033 12575 11067
rect 15393 11033 15427 11067
rect 16957 11033 16991 11067
rect 19625 11033 19659 11067
rect 22293 11033 22327 11067
rect 23305 11033 23339 11067
rect 23489 11033 23523 11067
rect 24501 11033 24535 11067
rect 26617 11033 26651 11067
rect 29561 11033 29595 11067
rect 32505 11033 32539 11067
rect 34897 11033 34931 11067
rect 35541 11033 35575 11067
rect 36461 11033 36495 11067
rect 9137 10965 9171 10999
rect 24869 10965 24903 10999
rect 25697 10965 25731 10999
rect 30389 10965 30423 10999
rect 34345 10965 34379 10999
rect 1593 10761 1627 10795
rect 3893 10761 3927 10795
rect 5273 10761 5307 10795
rect 6193 10761 6227 10795
rect 7021 10761 7055 10795
rect 10149 10761 10183 10795
rect 10793 10761 10827 10795
rect 14657 10761 14691 10795
rect 18153 10761 18187 10795
rect 19073 10761 19107 10795
rect 19717 10761 19751 10795
rect 21281 10761 21315 10795
rect 23857 10761 23891 10795
rect 25881 10761 25915 10795
rect 27813 10761 27847 10795
rect 28733 10761 28767 10795
rect 29837 10761 29871 10795
rect 31677 10761 31711 10795
rect 32689 10761 32723 10795
rect 32965 10761 32999 10795
rect 33333 10761 33367 10795
rect 35909 10761 35943 10795
rect 2237 10693 2271 10727
rect 3249 10693 3283 10727
rect 8033 10693 8067 10727
rect 9597 10693 9631 10727
rect 15025 10693 15059 10727
rect 20913 10693 20947 10727
rect 22109 10693 22143 10727
rect 34989 10693 35023 10727
rect 2605 10625 2639 10659
rect 5089 10625 5123 10659
rect 5641 10625 5675 10659
rect 5825 10625 5859 10659
rect 10609 10625 10643 10659
rect 18705 10625 18739 10659
rect 20269 10625 20303 10659
rect 22661 10625 22695 10659
rect 23029 10625 23063 10659
rect 23489 10625 23523 10659
rect 24225 10625 24259 10659
rect 24409 10625 24443 10659
rect 25329 10625 25363 10659
rect 30297 10625 30331 10659
rect 33793 10625 33827 10659
rect 3709 10557 3743 10591
rect 4261 10557 4295 10591
rect 6837 10557 6871 10591
rect 7389 10557 7423 10591
rect 8217 10557 8251 10591
rect 8484 10557 8518 10591
rect 11069 10557 11103 10591
rect 12265 10557 12299 10591
rect 12633 10557 12667 10591
rect 15117 10557 15151 10591
rect 17785 10557 17819 10591
rect 18429 10557 18463 10591
rect 19533 10557 19567 10591
rect 19993 10557 20027 10591
rect 26433 10557 26467 10591
rect 26689 10557 26723 10591
rect 32321 10557 32355 10591
rect 33885 10557 33919 10591
rect 34345 10557 34379 10591
rect 36461 10557 36495 10591
rect 37013 10557 37047 10591
rect 2789 10489 2823 10523
rect 4721 10489 4755 10523
rect 11253 10489 11287 10523
rect 11345 10489 11379 10523
rect 12900 10489 12934 10523
rect 15362 10489 15396 10523
rect 22385 10489 22419 10523
rect 24317 10489 24351 10523
rect 26249 10489 26283 10523
rect 28365 10489 28399 10523
rect 30113 10489 30147 10523
rect 30564 10489 30598 10523
rect 33793 10489 33827 10523
rect 35265 10489 35299 10523
rect 35541 10489 35575 10523
rect 2053 10421 2087 10455
rect 2697 10421 2731 10455
rect 3617 10421 3651 10455
rect 5733 10421 5767 10455
rect 6653 10421 6687 10455
rect 11805 10421 11839 10455
rect 14013 10421 14047 10455
rect 16497 10421 16531 10455
rect 17141 10421 17175 10455
rect 17417 10421 17451 10455
rect 18613 10421 18647 10455
rect 20177 10421 20211 10455
rect 21925 10421 21959 10455
rect 22569 10421 22603 10455
rect 24961 10421 24995 10455
rect 34621 10421 34655 10455
rect 35449 10421 35483 10455
rect 36369 10421 36403 10455
rect 36645 10421 36679 10455
rect 2513 10217 2547 10251
rect 4261 10217 4295 10251
rect 6653 10217 6687 10251
rect 7297 10217 7331 10251
rect 7941 10217 7975 10251
rect 9137 10217 9171 10251
rect 9873 10217 9907 10251
rect 10333 10217 10367 10251
rect 12541 10217 12575 10251
rect 16497 10217 16531 10251
rect 18245 10217 18279 10251
rect 18797 10217 18831 10251
rect 19165 10217 19199 10251
rect 21833 10217 21867 10251
rect 23949 10217 23983 10251
rect 25237 10217 25271 10251
rect 26341 10217 26375 10251
rect 26709 10217 26743 10251
rect 36369 10217 36403 10251
rect 2329 10149 2363 10183
rect 5540 10149 5574 10183
rect 8585 10149 8619 10183
rect 8677 10149 8711 10183
rect 10701 10149 10735 10183
rect 11713 10149 11747 10183
rect 15853 10149 15887 10183
rect 17110 10149 17144 10183
rect 22192 10149 22226 10183
rect 25329 10149 25363 10183
rect 27344 10149 27378 10183
rect 30113 10149 30147 10183
rect 30757 10149 30791 10183
rect 32474 10149 32508 10183
rect 3709 10081 3743 10115
rect 4077 10081 4111 10115
rect 5273 10081 5307 10115
rect 9689 10081 9723 10115
rect 11529 10081 11563 10115
rect 12981 10081 13015 10115
rect 15669 10081 15703 10115
rect 16865 10081 16899 10115
rect 27077 10081 27111 10115
rect 29745 10081 29779 10115
rect 30573 10081 30607 10115
rect 32229 10081 32263 10115
rect 34897 10081 34931 10115
rect 35256 10081 35290 10115
rect 1869 10013 1903 10047
rect 2605 10013 2639 10047
rect 4629 10013 4663 10047
rect 8493 10013 8527 10047
rect 11805 10013 11839 10047
rect 12725 10013 12759 10047
rect 15117 10013 15151 10047
rect 15945 10013 15979 10047
rect 21925 10013 21959 10047
rect 25237 10013 25271 10047
rect 30849 10013 30883 10047
rect 34989 10013 35023 10047
rect 3065 9945 3099 9979
rect 8125 9945 8159 9979
rect 11253 9945 11287 9979
rect 24777 9945 24811 9979
rect 30297 9945 30331 9979
rect 33609 9945 33643 9979
rect 2053 9877 2087 9911
rect 3433 9877 3467 9911
rect 5089 9877 5123 9911
rect 14105 9877 14139 9911
rect 15393 9877 15427 9911
rect 19717 9877 19751 9911
rect 23305 9877 23339 9911
rect 24501 9877 24535 9911
rect 28457 9877 28491 9911
rect 31217 9877 31251 9911
rect 31953 9877 31987 9911
rect 34161 9877 34195 9911
rect 5825 9673 5859 9707
rect 10517 9673 10551 9707
rect 11437 9673 11471 9707
rect 15301 9673 15335 9707
rect 16497 9673 16531 9707
rect 20821 9673 20855 9707
rect 25881 9673 25915 9707
rect 26801 9673 26835 9707
rect 34989 9673 35023 9707
rect 2053 9605 2087 9639
rect 2973 9605 3007 9639
rect 7021 9605 7055 9639
rect 9873 9605 9907 9639
rect 10885 9605 10919 9639
rect 24041 9605 24075 9639
rect 27537 9605 27571 9639
rect 29837 9605 29871 9639
rect 33333 9605 33367 9639
rect 36277 9605 36311 9639
rect 36553 9605 36587 9639
rect 2421 9537 2455 9571
rect 7573 9537 7607 9571
rect 17049 9537 17083 9571
rect 17877 9537 17911 9571
rect 23305 9537 23339 9571
rect 27997 9537 28031 9571
rect 29561 9537 29595 9571
rect 30573 9537 30607 9571
rect 30757 9537 30791 9571
rect 35541 9537 35575 9571
rect 37473 9537 37507 9571
rect 1869 9469 1903 9503
rect 2605 9469 2639 9503
rect 3525 9469 3559 9503
rect 5549 9469 5583 9503
rect 8493 9469 8527 9503
rect 8760 9469 8794 9503
rect 12817 9469 12851 9503
rect 13185 9469 13219 9503
rect 13277 9469 13311 9503
rect 18521 9469 18555 9503
rect 18788 9469 18822 9503
rect 21005 9469 21039 9503
rect 22937 9469 22971 9503
rect 24501 9469 24535 9503
rect 27077 9469 27111 9503
rect 29653 9469 29687 9503
rect 37105 9469 37139 9503
rect 2513 9401 2547 9435
rect 3341 9401 3375 9435
rect 3770 9401 3804 9435
rect 6285 9401 6319 9435
rect 7297 9401 7331 9435
rect 13522 9401 13556 9435
rect 16773 9401 16807 9435
rect 21250 9401 21284 9435
rect 24768 9401 24802 9435
rect 28089 9401 28123 9435
rect 31024 9401 31058 9435
rect 33609 9401 33643 9435
rect 33885 9401 33919 9435
rect 34345 9401 34379 9435
rect 35265 9401 35299 9435
rect 36829 9401 36863 9435
rect 4905 9333 4939 9367
rect 6561 9333 6595 9367
rect 7481 9333 7515 9367
rect 8033 9333 8067 9367
rect 10977 9333 11011 9367
rect 11897 9333 11931 9367
rect 12173 9333 12207 9367
rect 14657 9333 14691 9367
rect 15669 9333 15703 9367
rect 16313 9333 16347 9367
rect 16957 9333 16991 9367
rect 17509 9333 17543 9367
rect 18337 9333 18371 9367
rect 19901 9333 19935 9367
rect 20453 9333 20487 9367
rect 22385 9333 22419 9367
rect 24317 9333 24351 9367
rect 27997 9333 28031 9367
rect 28549 9333 28583 9367
rect 28917 9333 28951 9367
rect 30297 9333 30331 9367
rect 32137 9333 32171 9367
rect 32781 9333 32815 9367
rect 33149 9333 33183 9367
rect 33793 9333 33827 9367
rect 34621 9333 34655 9367
rect 35449 9333 35483 9367
rect 35909 9333 35943 9367
rect 37013 9333 37047 9367
rect 1685 9129 1719 9163
rect 1961 9129 1995 9163
rect 2789 9129 2823 9163
rect 9045 9129 9079 9163
rect 13737 9129 13771 9163
rect 15025 9129 15059 9163
rect 17141 9129 17175 9163
rect 18061 9129 18095 9163
rect 19809 9129 19843 9163
rect 23029 9129 23063 9163
rect 24225 9129 24259 9163
rect 25421 9129 25455 9163
rect 31585 9129 31619 9163
rect 32689 9129 32723 9163
rect 35339 9129 35373 9163
rect 35817 9129 35851 9163
rect 5365 9061 5399 9095
rect 6929 9061 6963 9095
rect 7389 9061 7423 9095
rect 8585 9061 8619 9095
rect 8677 9061 8711 9095
rect 11713 9061 11747 9095
rect 12633 9061 12667 9095
rect 13277 9061 13311 9095
rect 15375 9061 15409 9095
rect 15853 9061 15887 9095
rect 19901 9061 19935 9095
rect 21916 9061 21950 9095
rect 24869 9061 24903 9095
rect 26985 9061 27019 9095
rect 27537 9061 27571 9095
rect 28264 9061 28298 9095
rect 31033 9061 31067 9095
rect 31861 9061 31895 9095
rect 34253 9061 34287 9095
rect 34897 9061 34931 9095
rect 2605 8993 2639 9027
rect 3617 8993 3651 9027
rect 6745 8993 6779 9027
rect 7849 8993 7883 9027
rect 10517 8993 10551 9027
rect 11805 8993 11839 9027
rect 15945 8993 15979 9027
rect 24685 8993 24719 9027
rect 27997 8993 28031 9027
rect 30849 8993 30883 9027
rect 32781 8993 32815 9027
rect 34069 8993 34103 9027
rect 35633 8993 35667 9027
rect 2881 8925 2915 8959
rect 4721 8925 4755 8959
rect 5365 8925 5399 8959
rect 5457 8925 5491 8959
rect 7021 8925 7055 8959
rect 8585 8925 8619 8959
rect 11621 8925 11655 8959
rect 12265 8925 12299 8959
rect 13277 8925 13311 8959
rect 13369 8925 13403 8959
rect 15761 8925 15795 8959
rect 17969 8925 18003 8959
rect 18153 8925 18187 8959
rect 19809 8925 19843 8959
rect 21649 8925 21683 8959
rect 24961 8925 24995 8959
rect 30389 8925 30423 8959
rect 31125 8925 31159 8959
rect 32689 8925 32723 8959
rect 34345 8925 34379 8959
rect 35909 8925 35943 8959
rect 2329 8857 2363 8891
rect 4905 8857 4939 8891
rect 6285 8857 6319 8891
rect 8125 8857 8159 8891
rect 11253 8857 11287 8891
rect 12817 8857 12851 8891
rect 19349 8857 19383 8891
rect 30573 8857 30607 8891
rect 32229 8857 32263 8891
rect 33333 8857 33367 8891
rect 4353 8789 4387 8823
rect 5825 8789 5859 8823
rect 6469 8789 6503 8823
rect 10793 8789 10827 8823
rect 16497 8789 16531 8823
rect 16865 8789 16899 8823
rect 17601 8789 17635 8823
rect 18613 8789 18647 8823
rect 18981 8789 19015 8823
rect 20269 8789 20303 8823
rect 23765 8789 23799 8823
rect 24409 8789 24443 8823
rect 27905 8789 27939 8823
rect 29377 8789 29411 8823
rect 29929 8789 29963 8823
rect 33793 8789 33827 8823
rect 36461 8789 36495 8823
rect 1685 8585 1719 8619
rect 2053 8585 2087 8619
rect 3525 8585 3559 8619
rect 5273 8585 5307 8619
rect 7757 8585 7791 8619
rect 9689 8585 9723 8619
rect 10241 8585 10275 8619
rect 10885 8585 10919 8619
rect 11805 8585 11839 8619
rect 14013 8585 14047 8619
rect 14933 8585 14967 8619
rect 17601 8585 17635 8619
rect 20269 8585 20303 8619
rect 23397 8585 23431 8619
rect 25053 8585 25087 8619
rect 26065 8585 26099 8619
rect 26525 8585 26559 8619
rect 28089 8585 28123 8619
rect 29377 8585 29411 8619
rect 30941 8585 30975 8619
rect 37289 8585 37323 8619
rect 7021 8517 7055 8551
rect 15761 8517 15795 8551
rect 16497 8517 16531 8551
rect 18153 8517 18187 8551
rect 19533 8517 19567 8551
rect 21925 8517 21959 8551
rect 26893 8517 26927 8551
rect 27169 8517 27203 8551
rect 31861 8517 31895 8551
rect 32781 8517 32815 8551
rect 33057 8517 33091 8551
rect 36277 8517 36311 8551
rect 37565 8517 37599 8551
rect 2145 8449 2179 8483
rect 4905 8449 4939 8483
rect 5733 8449 5767 8483
rect 11437 8449 11471 8483
rect 16957 8449 16991 8483
rect 19073 8449 19107 8483
rect 20637 8449 20671 8483
rect 23673 8449 23707 8483
rect 27537 8449 27571 8483
rect 27721 8449 27755 8483
rect 29101 8449 29135 8483
rect 29837 8449 29871 8483
rect 31493 8449 31527 8483
rect 33425 8449 33459 8483
rect 2401 8381 2435 8415
rect 4537 8381 4571 8415
rect 5825 8381 5859 8415
rect 6837 8381 6871 8415
rect 8309 8381 8343 8415
rect 8565 8381 8599 8415
rect 10701 8381 10735 8415
rect 12265 8381 12299 8415
rect 12633 8381 12667 8415
rect 18429 8381 18463 8415
rect 18705 8381 18739 8415
rect 19901 8381 19935 8415
rect 20821 8381 20855 8415
rect 21373 8381 21407 8415
rect 22201 8381 22235 8415
rect 29929 8381 29963 8415
rect 30665 8381 30699 8415
rect 31217 8381 31251 8415
rect 34069 8381 34103 8415
rect 34897 8381 34931 8415
rect 35164 8381 35198 8415
rect 36829 8381 36863 8415
rect 37381 8381 37415 8415
rect 37933 8381 37967 8415
rect 4169 8313 4203 8347
rect 5733 8313 5767 8347
rect 6377 8313 6411 8347
rect 11161 8313 11195 8347
rect 11345 8313 11379 8347
rect 12878 8313 12912 8347
rect 15301 8313 15335 8347
rect 16313 8313 16347 8347
rect 17049 8313 17083 8347
rect 18613 8313 18647 8347
rect 20729 8313 20763 8347
rect 22477 8313 22511 8347
rect 23940 8313 23974 8347
rect 25605 8313 25639 8347
rect 27629 8313 27663 8347
rect 28641 8313 28675 8347
rect 29837 8313 29871 8347
rect 32505 8313 32539 8347
rect 33609 8313 33643 8347
rect 8033 8245 8067 8279
rect 16957 8245 16991 8279
rect 21649 8245 21683 8279
rect 22385 8245 22419 8279
rect 22845 8245 22879 8279
rect 30389 8245 30423 8279
rect 31401 8245 31435 8279
rect 33517 8245 33551 8279
rect 34713 8245 34747 8279
rect 3157 8041 3191 8075
rect 3893 8041 3927 8075
rect 7757 8041 7791 8075
rect 8677 8041 8711 8075
rect 10885 8041 10919 8075
rect 12633 8041 12667 8075
rect 13185 8041 13219 8075
rect 13553 8041 13587 8075
rect 17601 8041 17635 8075
rect 19625 8041 19659 8075
rect 20637 8041 20671 8075
rect 21005 8041 21039 8075
rect 21925 8041 21959 8075
rect 24409 8041 24443 8075
rect 26341 8041 26375 8075
rect 27077 8041 27111 8075
rect 28549 8041 28583 8075
rect 30481 8041 30515 8075
rect 31033 8041 31067 8075
rect 31493 8041 31527 8075
rect 31953 8041 31987 8075
rect 32505 8041 32539 8075
rect 34345 8041 34379 8075
rect 36461 8041 36495 8075
rect 2329 7973 2363 8007
rect 2881 7973 2915 8007
rect 4966 7973 5000 8007
rect 7573 7973 7607 8007
rect 9045 7973 9079 8007
rect 10241 7973 10275 8007
rect 16681 7973 16715 8007
rect 17233 7973 17267 8007
rect 17960 7973 17994 8007
rect 22284 7973 22318 8007
rect 24777 7973 24811 8007
rect 25421 7973 25455 8007
rect 26599 7973 26633 8007
rect 36001 7973 36035 8007
rect 1685 7905 1719 7939
rect 2421 7905 2455 7939
rect 10333 7905 10367 7939
rect 11253 7905 11287 7939
rect 11520 7905 11554 7939
rect 13737 7905 13771 7939
rect 16037 7905 16071 7939
rect 16497 7905 16531 7939
rect 20177 7905 20211 7939
rect 25513 7905 25547 7939
rect 26893 7905 26927 7939
rect 29101 7905 29135 7939
rect 29357 7905 29391 7939
rect 33221 7905 33255 7939
rect 2329 7837 2363 7871
rect 4721 7837 4755 7871
rect 7849 7837 7883 7871
rect 8401 7837 8435 7871
rect 10149 7837 10183 7871
rect 16773 7837 16807 7871
rect 17693 7837 17727 7871
rect 22017 7837 22051 7871
rect 24041 7837 24075 7871
rect 25421 7837 25455 7871
rect 27169 7837 27203 7871
rect 28089 7837 28123 7871
rect 32965 7837 32999 7871
rect 35909 7837 35943 7871
rect 36093 7837 36127 7871
rect 7113 7769 7147 7803
rect 16221 7769 16255 7803
rect 24961 7769 24995 7803
rect 35541 7769 35575 7803
rect 1869 7701 1903 7735
rect 4353 7701 4387 7735
rect 6101 7701 6135 7735
rect 6653 7701 6687 7735
rect 7297 7701 7331 7735
rect 9781 7701 9815 7735
rect 14289 7701 14323 7735
rect 19073 7701 19107 7735
rect 21465 7701 21499 7735
rect 23397 7701 23431 7735
rect 32873 7701 32907 7735
rect 34989 7701 35023 7735
rect 35265 7701 35299 7735
rect 3249 7497 3283 7531
rect 5457 7497 5491 7531
rect 6653 7497 6687 7531
rect 9321 7497 9355 7531
rect 11897 7497 11931 7531
rect 12725 7497 12759 7531
rect 15945 7497 15979 7531
rect 16497 7497 16531 7531
rect 19993 7497 20027 7531
rect 21557 7497 21591 7531
rect 22109 7497 22143 7531
rect 23857 7497 23891 7531
rect 26617 7497 26651 7531
rect 28641 7497 28675 7531
rect 29377 7497 29411 7531
rect 32413 7497 32447 7531
rect 34621 7497 34655 7531
rect 36645 7497 36679 7531
rect 1961 7429 1995 7463
rect 10885 7429 10919 7463
rect 14289 7429 14323 7463
rect 26341 7429 26375 7463
rect 29101 7429 29135 7463
rect 30941 7429 30975 7463
rect 32781 7429 32815 7463
rect 33333 7429 33367 7463
rect 6285 7361 6319 7395
rect 12173 7361 12207 7395
rect 12541 7361 12575 7395
rect 13185 7361 13219 7395
rect 14105 7361 14139 7395
rect 14749 7361 14783 7395
rect 16865 7361 16899 7395
rect 17049 7361 17083 7395
rect 21833 7361 21867 7395
rect 24041 7361 24075 7395
rect 26065 7361 26099 7395
rect 27077 7361 27111 7395
rect 29929 7361 29963 7395
rect 30665 7361 30699 7395
rect 31401 7361 31435 7395
rect 33885 7361 33919 7395
rect 34253 7361 34287 7395
rect 3985 7293 4019 7327
rect 4077 7293 4111 7327
rect 4344 7293 4378 7327
rect 7389 7293 7423 7327
rect 7656 7293 7690 7327
rect 11437 7293 11471 7327
rect 15577 7293 15611 7327
rect 17785 7293 17819 7327
rect 18061 7293 18095 7327
rect 22385 7293 22419 7327
rect 29653 7293 29687 7327
rect 30297 7293 30331 7327
rect 33149 7293 33183 7327
rect 33609 7293 33643 7327
rect 35265 7293 35299 7327
rect 37197 7293 37231 7327
rect 1777 7225 1811 7259
rect 2237 7225 2271 7259
rect 2513 7225 2547 7259
rect 11161 7225 11195 7259
rect 11345 7225 11379 7259
rect 12541 7225 12575 7259
rect 13185 7225 13219 7259
rect 13277 7225 13311 7259
rect 13737 7225 13771 7259
rect 14841 7225 14875 7259
rect 16957 7225 16991 7259
rect 18328 7225 18362 7259
rect 22661 7225 22695 7259
rect 24286 7225 24320 7259
rect 27169 7225 27203 7259
rect 27905 7225 27939 7259
rect 29837 7225 29871 7259
rect 31493 7225 31527 7259
rect 35510 7225 35544 7259
rect 2421 7157 2455 7191
rect 2881 7157 2915 7191
rect 7297 7157 7331 7191
rect 8769 7157 8803 7191
rect 9689 7157 9723 7191
rect 10057 7157 10091 7191
rect 10701 7157 10735 7191
rect 14749 7157 14783 7191
rect 16221 7157 16255 7191
rect 19441 7157 19475 7191
rect 20913 7157 20947 7191
rect 22569 7157 22603 7191
rect 23029 7157 23063 7191
rect 23397 7157 23431 7191
rect 25421 7157 25455 7191
rect 27077 7157 27111 7191
rect 27537 7157 27571 7191
rect 28089 7157 28123 7191
rect 31401 7157 31435 7191
rect 31861 7157 31895 7191
rect 33793 7157 33827 7191
rect 35081 7157 35115 7191
rect 2605 6953 2639 6987
rect 4261 6953 4295 6987
rect 5089 6953 5123 6987
rect 6929 6953 6963 6987
rect 8125 6953 8159 6987
rect 11253 6953 11287 6987
rect 13645 6953 13679 6987
rect 14473 6953 14507 6987
rect 16497 6953 16531 6987
rect 19809 6953 19843 6987
rect 25053 6953 25087 6987
rect 25513 6953 25547 6987
rect 26341 6953 26375 6987
rect 29009 6953 29043 6987
rect 31217 6953 31251 6987
rect 33977 6953 34011 6987
rect 34345 6953 34379 6987
rect 35909 6953 35943 6987
rect 2145 6885 2179 6919
rect 6009 6885 6043 6919
rect 7573 6885 7607 6919
rect 10241 6885 10275 6919
rect 13277 6885 13311 6919
rect 21373 6885 21407 6919
rect 21557 6885 21591 6919
rect 23121 6885 23155 6919
rect 24685 6885 24719 6919
rect 1961 6817 1995 6851
rect 3709 6817 3743 6851
rect 4077 6817 4111 6851
rect 7665 6817 7699 6851
rect 10885 6817 10919 6851
rect 11345 6817 11379 6851
rect 11601 6817 11635 6851
rect 13829 6817 13863 6851
rect 16129 6817 16163 6851
rect 17029 6817 17063 6851
rect 19625 6817 19659 6851
rect 20729 6817 20763 6851
rect 22477 6817 22511 6851
rect 24777 6817 24811 6851
rect 2237 6749 2271 6783
rect 3433 6749 3467 6783
rect 6009 6749 6043 6783
rect 6101 6749 6135 6783
rect 6561 6749 6595 6783
rect 7481 6749 7515 6783
rect 8585 6749 8619 6783
rect 10149 6749 10183 6783
rect 10333 6749 10367 6783
rect 16773 6749 16807 6783
rect 19901 6749 19935 6783
rect 21649 6749 21683 6783
rect 23121 6749 23155 6783
rect 23213 6749 23247 6783
rect 24593 6749 24627 6783
rect 32505 6885 32539 6919
rect 32689 6885 32723 6919
rect 26965 6817 26999 6851
rect 29460 6817 29494 6851
rect 32781 6817 32815 6851
rect 34785 6817 34819 6851
rect 26709 6749 26743 6783
rect 29193 6749 29227 6783
rect 34529 6749 34563 6783
rect 1685 6681 1719 6715
rect 3065 6681 3099 6715
rect 5549 6681 5583 6715
rect 21097 6681 21131 6715
rect 22661 6681 22695 6715
rect 24041 6681 24075 6715
rect 25053 6681 25087 6715
rect 28089 6681 28123 6715
rect 30573 6681 30607 6715
rect 32229 6681 32263 6715
rect 33333 6681 33367 6715
rect 4813 6613 4847 6647
rect 7113 6613 7147 6647
rect 9505 6613 9539 6647
rect 9781 6613 9815 6647
rect 12725 6613 12759 6647
rect 18153 6613 18187 6647
rect 18797 6613 18831 6647
rect 19349 6613 19383 6647
rect 22109 6613 22143 6647
rect 24225 6613 24259 6647
rect 25145 6613 25179 6647
rect 25973 6613 26007 6647
rect 31493 6613 31527 6647
rect 31953 6613 31987 6647
rect 33701 6613 33735 6647
rect 36461 6613 36495 6647
rect 3157 6409 3191 6443
rect 4169 6409 4203 6443
rect 6653 6409 6687 6443
rect 7297 6409 7331 6443
rect 11345 6409 11379 6443
rect 11805 6409 11839 6443
rect 12173 6409 12207 6443
rect 17785 6409 17819 6443
rect 18705 6409 18739 6443
rect 19349 6409 19383 6443
rect 19625 6409 19659 6443
rect 21005 6409 21039 6443
rect 22477 6409 22511 6443
rect 23121 6409 23155 6443
rect 23489 6409 23523 6443
rect 24501 6409 24535 6443
rect 25789 6409 25823 6443
rect 27077 6409 27111 6443
rect 27353 6409 27387 6443
rect 29469 6409 29503 6443
rect 29929 6409 29963 6443
rect 32413 6409 32447 6443
rect 33333 6409 33367 6443
rect 36277 6409 36311 6443
rect 37565 6409 37599 6443
rect 9965 6341 9999 6375
rect 12541 6341 12575 6375
rect 16865 6341 16899 6375
rect 26065 6341 26099 6375
rect 27629 6341 27663 6375
rect 30297 6341 30331 6375
rect 31861 6341 31895 6375
rect 7389 6273 7423 6307
rect 19993 6273 20027 6307
rect 20177 6273 20211 6307
rect 24961 6273 24995 6307
rect 25421 6273 25455 6307
rect 26433 6273 26467 6307
rect 27997 6273 28031 6307
rect 30481 6273 30515 6307
rect 33793 6273 33827 6307
rect 33885 6273 33919 6307
rect 1685 6205 1719 6239
rect 1777 6205 1811 6239
rect 3801 6205 3835 6239
rect 4261 6205 4295 6239
rect 9689 6205 9723 6239
rect 10885 6205 10919 6239
rect 12817 6205 12851 6239
rect 13093 6205 13127 6239
rect 13461 6205 13495 6239
rect 14289 6205 14323 6239
rect 14381 6205 14415 6239
rect 18981 6205 19015 6239
rect 21097 6205 21131 6239
rect 21364 6205 21398 6239
rect 30748 6205 30782 6239
rect 34621 6205 34655 6239
rect 34897 6205 34931 6239
rect 37381 6205 37415 6239
rect 37933 6205 37967 6239
rect 2044 6137 2078 6171
rect 4528 6137 4562 6171
rect 7656 6137 7690 6171
rect 10241 6137 10275 6171
rect 10517 6137 10551 6171
rect 14648 6137 14682 6171
rect 25053 6137 25087 6171
rect 26617 6137 26651 6171
rect 28181 6137 28215 6171
rect 28549 6137 28583 6171
rect 33149 6137 33183 6171
rect 33793 6137 33827 6171
rect 35164 6137 35198 6171
rect 5641 6069 5675 6103
rect 6193 6069 6227 6103
rect 8769 6069 8803 6103
rect 9321 6069 9355 6103
rect 10425 6069 10459 6103
rect 13001 6069 13035 6103
rect 15761 6069 15795 6103
rect 17141 6069 17175 6103
rect 18337 6069 18371 6103
rect 20085 6069 20119 6103
rect 20545 6069 20579 6103
rect 24133 6069 24167 6103
rect 24961 6069 24995 6103
rect 26525 6069 26559 6103
rect 28089 6069 28123 6103
rect 2881 5865 2915 5899
rect 4629 5865 4663 5899
rect 5181 5865 5215 5899
rect 6653 5865 6687 5899
rect 7297 5865 7331 5899
rect 7665 5865 7699 5899
rect 9505 5865 9539 5899
rect 10701 5865 10735 5899
rect 11437 5865 11471 5899
rect 18521 5865 18555 5899
rect 19533 5865 19567 5899
rect 19993 5865 20027 5899
rect 20729 5865 20763 5899
rect 23397 5865 23431 5899
rect 23857 5865 23891 5899
rect 27711 5865 27745 5899
rect 29745 5865 29779 5899
rect 30573 5865 30607 5899
rect 31861 5865 31895 5899
rect 32413 5865 32447 5899
rect 34161 5865 34195 5899
rect 35725 5865 35759 5899
rect 36093 5865 36127 5899
rect 3801 5797 3835 5831
rect 8309 5797 8343 5831
rect 8401 5797 8435 5831
rect 10057 5797 10091 5831
rect 10241 5797 10275 5831
rect 12633 5797 12667 5831
rect 13093 5797 13127 5831
rect 14197 5797 14231 5831
rect 18337 5797 18371 5831
rect 18613 5797 18647 5831
rect 20269 5797 20303 5831
rect 21732 5797 21766 5831
rect 28181 5797 28215 5831
rect 29561 5797 29595 5831
rect 33333 5797 33367 5831
rect 34897 5797 34931 5831
rect 34989 5797 35023 5831
rect 1501 5729 1535 5763
rect 1768 5729 1802 5763
rect 3525 5729 3559 5763
rect 4077 5729 4111 5763
rect 5273 5729 5307 5763
rect 5540 5729 5574 5763
rect 12449 5729 12483 5763
rect 15741 5729 15775 5763
rect 24216 5729 24250 5763
rect 27997 5729 28031 5763
rect 34713 5729 34747 5763
rect 35909 5729 35943 5763
rect 8217 5661 8251 5695
rect 10333 5661 10367 5695
rect 12725 5661 12759 5695
rect 14105 5661 14139 5695
rect 14289 5661 14323 5695
rect 15485 5661 15519 5695
rect 21465 5661 21499 5695
rect 23949 5661 23983 5695
rect 28273 5661 28307 5695
rect 29837 5661 29871 5695
rect 33333 5661 33367 5695
rect 33425 5661 33459 5695
rect 35357 5661 35391 5695
rect 4261 5593 4295 5627
rect 7849 5593 7883 5627
rect 9781 5593 9815 5627
rect 12173 5593 12207 5627
rect 13461 5593 13495 5627
rect 18061 5593 18095 5627
rect 26065 5593 26099 5627
rect 32873 5593 32907 5627
rect 34437 5593 34471 5627
rect 11713 5525 11747 5559
rect 13737 5525 13771 5559
rect 16865 5525 16899 5559
rect 21097 5525 21131 5559
rect 22845 5525 22879 5559
rect 25329 5525 25363 5559
rect 26709 5525 26743 5559
rect 27169 5525 27203 5559
rect 29285 5525 29319 5559
rect 1961 5321 1995 5355
rect 3065 5321 3099 5355
rect 3709 5321 3743 5355
rect 5365 5321 5399 5355
rect 7021 5321 7055 5355
rect 7389 5321 7423 5355
rect 8309 5321 8343 5355
rect 10701 5321 10735 5355
rect 11437 5321 11471 5355
rect 13829 5321 13863 5355
rect 15577 5321 15611 5355
rect 17141 5321 17175 5355
rect 17877 5321 17911 5355
rect 19073 5321 19107 5355
rect 19441 5321 19475 5355
rect 20269 5321 20303 5355
rect 22201 5321 22235 5355
rect 23949 5321 23983 5355
rect 24777 5321 24811 5355
rect 26985 5321 27019 5355
rect 27721 5321 27755 5355
rect 28089 5321 28123 5355
rect 29377 5321 29411 5355
rect 30389 5321 30423 5355
rect 31769 5321 31803 5355
rect 34253 5321 34287 5355
rect 34713 5321 34747 5355
rect 36645 5321 36679 5355
rect 2145 5253 2179 5287
rect 16037 5253 16071 5287
rect 18153 5253 18187 5287
rect 21281 5253 21315 5287
rect 25421 5253 25455 5287
rect 29101 5253 29135 5287
rect 32689 5253 32723 5287
rect 33977 5253 34011 5287
rect 34989 5253 35023 5287
rect 2605 5185 2639 5219
rect 2697 5185 2731 5219
rect 4261 5185 4295 5219
rect 5641 5185 5675 5219
rect 8401 5185 8435 5219
rect 16405 5185 16439 5219
rect 16589 5185 16623 5219
rect 21097 5185 21131 5219
rect 21833 5185 21867 5219
rect 25605 5185 25639 5219
rect 29929 5185 29963 5219
rect 32505 5185 32539 5219
rect 33057 5185 33091 5219
rect 33241 5185 33275 5219
rect 35541 5185 35575 5219
rect 11805 5117 11839 5151
rect 12449 5117 12483 5151
rect 20729 5117 20763 5151
rect 25861 5117 25895 5151
rect 28365 5117 28399 5151
rect 29653 5117 29687 5151
rect 30665 5117 30699 5151
rect 32137 5117 32171 5151
rect 35265 5117 35299 5151
rect 36461 5117 36495 5151
rect 37013 5117 37047 5151
rect 2605 5049 2639 5083
rect 3525 5049 3559 5083
rect 3985 5049 4019 5083
rect 4169 5049 4203 5083
rect 7849 5049 7883 5083
rect 8646 5049 8680 5083
rect 12694 5049 12728 5083
rect 15117 5049 15151 5083
rect 18429 5049 18463 5083
rect 18705 5049 18739 5083
rect 21557 5049 21591 5083
rect 21741 5049 21775 5083
rect 24317 5049 24351 5083
rect 29837 5049 29871 5083
rect 33149 5049 33183 5083
rect 4721 4981 4755 5015
rect 9781 4981 9815 5015
rect 10425 4981 10459 5015
rect 12081 4981 12115 5015
rect 14381 4981 14415 5015
rect 14749 4981 14783 5015
rect 16497 4981 16531 5015
rect 17509 4981 17543 5015
rect 18613 4981 18647 5015
rect 35449 4981 35483 5015
rect 35909 4981 35943 5015
rect 1593 4777 1627 4811
rect 2697 4777 2731 4811
rect 3433 4777 3467 4811
rect 3893 4777 3927 4811
rect 4261 4777 4295 4811
rect 7481 4777 7515 4811
rect 8585 4777 8619 4811
rect 9873 4777 9907 4811
rect 11897 4777 11931 4811
rect 13001 4777 13035 4811
rect 14105 4777 14139 4811
rect 14657 4777 14691 4811
rect 16129 4777 16163 4811
rect 16405 4777 16439 4811
rect 18061 4777 18095 4811
rect 18981 4777 19015 4811
rect 21557 4777 21591 4811
rect 22569 4777 22603 4811
rect 25697 4777 25731 4811
rect 29653 4777 29687 4811
rect 30021 4777 30055 4811
rect 32781 4777 32815 4811
rect 32965 4777 32999 4811
rect 33425 4777 33459 4811
rect 34529 4777 34563 4811
rect 35357 4777 35391 4811
rect 35725 4777 35759 4811
rect 3065 4709 3099 4743
rect 8125 4709 8159 4743
rect 10977 4709 11011 4743
rect 11529 4709 11563 4743
rect 12541 4709 12575 4743
rect 13627 4709 13661 4743
rect 13921 4709 13955 4743
rect 15853 4709 15887 4743
rect 16939 4709 16973 4743
rect 17417 4709 17451 4743
rect 18797 4709 18831 4743
rect 22385 4709 22419 4743
rect 28089 4709 28123 4743
rect 28181 4709 28215 4743
rect 29377 4709 29411 4743
rect 32505 4709 32539 4743
rect 34345 4709 34379 4743
rect 34621 4709 34655 4743
rect 1409 4641 1443 4675
rect 2145 4641 2179 4675
rect 2513 4641 2547 4675
rect 8217 4641 8251 4675
rect 13369 4641 13403 4675
rect 15669 4641 15703 4675
rect 15945 4641 15979 4675
rect 16129 4641 16163 4675
rect 17233 4641 17267 4675
rect 27905 4641 27939 4675
rect 34989 4641 35023 4675
rect 35541 4641 35575 4675
rect 8033 4573 8067 4607
rect 10885 4573 10919 4607
rect 11069 4573 11103 4607
rect 12449 4573 12483 4607
rect 12633 4573 12667 4607
rect 14197 4573 14231 4607
rect 17509 4573 17543 4607
rect 19073 4573 19107 4607
rect 22661 4573 22695 4607
rect 7665 4505 7699 4539
rect 10517 4505 10551 4539
rect 16773 4505 16807 4539
rect 18521 4505 18555 4539
rect 27629 4505 27663 4539
rect 34069 4505 34103 4539
rect 12081 4437 12115 4471
rect 15393 4437 15427 4471
rect 22109 4437 22143 4471
rect 2329 4233 2363 4267
rect 2973 4233 3007 4267
rect 8033 4233 8067 4267
rect 11805 4233 11839 4267
rect 12541 4233 12575 4267
rect 14105 4233 14139 4267
rect 16129 4233 16163 4267
rect 17325 4233 17359 4267
rect 17693 4233 17727 4267
rect 19165 4233 19199 4267
rect 22385 4233 22419 4267
rect 27721 4233 27755 4267
rect 27997 4233 28031 4267
rect 28365 4233 28399 4267
rect 33701 4233 33735 4267
rect 34437 4233 34471 4267
rect 10885 4165 10919 4199
rect 15761 4165 15795 4199
rect 18521 4165 18555 4199
rect 8309 4097 8343 4131
rect 9597 4097 9631 4131
rect 13093 4097 13127 4131
rect 13645 4097 13679 4131
rect 14565 4097 14599 4131
rect 18797 4097 18831 4131
rect 22109 4097 22143 4131
rect 22753 4097 22787 4131
rect 26157 4097 26191 4131
rect 27169 4097 27203 4131
rect 34069 4097 34103 4131
rect 36369 4097 36403 4131
rect 1409 4029 1443 4063
rect 2513 4029 2547 4063
rect 11161 4029 11195 4063
rect 11437 4029 11471 4063
rect 16865 4029 16899 4063
rect 26691 4029 26725 4063
rect 35449 4029 35483 4063
rect 36001 4029 36035 4063
rect 2053 3961 2087 3995
rect 9965 3961 9999 3995
rect 12817 3961 12851 3995
rect 14565 3961 14599 3995
rect 14657 3961 14691 3995
rect 27261 3961 27295 3995
rect 1593 3893 1627 3927
rect 7573 3893 7607 3927
rect 10333 3893 10367 3927
rect 10609 3893 10643 3927
rect 11345 3893 11379 3927
rect 12173 3893 12207 3927
rect 13001 3893 13035 3927
rect 15301 3893 15335 3927
rect 26525 3893 26559 3927
rect 27169 3893 27203 3927
rect 35633 3893 35667 3927
rect 1593 3689 1627 3723
rect 10793 3689 10827 3723
rect 13369 3689 13403 3723
rect 13921 3689 13955 3723
rect 14197 3689 14231 3723
rect 14657 3689 14691 3723
rect 15577 3689 15611 3723
rect 26801 3689 26835 3723
rect 10517 3621 10551 3655
rect 11621 3621 11655 3655
rect 11805 3621 11839 3655
rect 1409 3553 1443 3587
rect 11897 3553 11931 3587
rect 13369 3485 13403 3519
rect 13461 3485 13495 3519
rect 11345 3417 11379 3451
rect 12909 3417 12943 3451
rect 12541 3349 12575 3383
rect 1593 3145 1627 3179
rect 10977 3145 11011 3179
rect 11621 3145 11655 3179
rect 13461 3145 13495 3179
rect 13829 3145 13863 3179
rect 14197 3145 14231 3179
rect 11253 3077 11287 3111
rect 12541 3077 12575 3111
rect 12265 3009 12299 3043
rect 13093 3009 13127 3043
rect 12817 2941 12851 2975
rect 13001 2873 13035 2907
rect 12909 2601 12943 2635
rect 13553 2601 13587 2635
rect 13185 2533 13219 2567
<< metal1 >>
rect 3602 14084 3608 14136
rect 3660 14124 3666 14136
rect 7466 14124 7472 14136
rect 3660 14096 7472 14124
rect 3660 14084 3666 14096
rect 7466 14084 7472 14096
rect 7524 14084 7530 14136
rect 3418 14016 3424 14068
rect 3476 14056 3482 14068
rect 6914 14056 6920 14068
rect 3476 14028 6920 14056
rect 3476 14016 3482 14028
rect 6914 14016 6920 14028
rect 6972 14016 6978 14068
rect 3510 13948 3516 14000
rect 3568 13988 3574 14000
rect 8386 13988 8392 14000
rect 3568 13960 8392 13988
rect 3568 13948 3574 13960
rect 8386 13948 8392 13960
rect 8444 13948 8450 14000
rect 3142 13880 3148 13932
rect 3200 13920 3206 13932
rect 7098 13920 7104 13932
rect 3200 13892 7104 13920
rect 3200 13880 3206 13892
rect 7098 13880 7104 13892
rect 7156 13880 7162 13932
rect 33134 13880 33140 13932
rect 33192 13920 33198 13932
rect 34790 13920 34796 13932
rect 33192 13892 34796 13920
rect 33192 13880 33198 13892
rect 34790 13880 34796 13892
rect 34848 13880 34854 13932
rect 3234 13812 3240 13864
rect 3292 13852 3298 13864
rect 9858 13852 9864 13864
rect 3292 13824 9864 13852
rect 3292 13812 3298 13824
rect 9858 13812 9864 13824
rect 9916 13812 9922 13864
rect 9950 13812 9956 13864
rect 10008 13852 10014 13864
rect 34514 13852 34520 13864
rect 10008 13824 34520 13852
rect 10008 13812 10014 13824
rect 34514 13812 34520 13824
rect 34572 13812 34578 13864
rect 31202 13676 31208 13728
rect 31260 13716 31266 13728
rect 36170 13716 36176 13728
rect 31260 13688 36176 13716
rect 31260 13676 31266 13688
rect 36170 13676 36176 13688
rect 36228 13676 36234 13728
rect 1104 13626 38824 13648
rect 1104 13574 14315 13626
rect 14367 13574 14379 13626
rect 14431 13574 14443 13626
rect 14495 13574 14507 13626
rect 14559 13574 27648 13626
rect 27700 13574 27712 13626
rect 27764 13574 27776 13626
rect 27828 13574 27840 13626
rect 27892 13574 38824 13626
rect 1104 13552 38824 13574
rect 2774 13472 2780 13524
rect 2832 13512 2838 13524
rect 5353 13515 5411 13521
rect 5353 13512 5365 13515
rect 2832 13484 5365 13512
rect 2832 13472 2838 13484
rect 5353 13481 5365 13484
rect 5399 13481 5411 13515
rect 7098 13512 7104 13524
rect 7059 13484 7104 13512
rect 5353 13475 5411 13481
rect 7098 13472 7104 13484
rect 7156 13472 7162 13524
rect 34425 13515 34483 13521
rect 34425 13481 34437 13515
rect 34471 13512 34483 13515
rect 34606 13512 34612 13524
rect 34471 13484 34612 13512
rect 34471 13481 34483 13484
rect 34425 13475 34483 13481
rect 34606 13472 34612 13484
rect 34664 13472 34670 13524
rect 2961 13447 3019 13453
rect 2961 13413 2973 13447
rect 3007 13444 3019 13447
rect 5810 13444 5816 13456
rect 3007 13416 5816 13444
rect 3007 13413 3019 13416
rect 2961 13407 3019 13413
rect 5810 13404 5816 13416
rect 5868 13404 5874 13456
rect 17218 13404 17224 13456
rect 17276 13444 17282 13456
rect 17276 13416 36584 13444
rect 17276 13404 17282 13416
rect 1397 13379 1455 13385
rect 1397 13345 1409 13379
rect 1443 13376 1455 13379
rect 1578 13376 1584 13388
rect 1443 13348 1584 13376
rect 1443 13345 1455 13348
rect 1397 13339 1455 13345
rect 1578 13336 1584 13348
rect 1636 13336 1642 13388
rect 2314 13336 2320 13388
rect 2372 13376 2378 13388
rect 2685 13379 2743 13385
rect 2685 13376 2697 13379
rect 2372 13348 2697 13376
rect 2372 13336 2378 13348
rect 2685 13345 2697 13348
rect 2731 13376 2743 13379
rect 3421 13379 3479 13385
rect 3421 13376 3433 13379
rect 2731 13348 3433 13376
rect 2731 13345 2743 13348
rect 2685 13339 2743 13345
rect 3421 13345 3433 13348
rect 3467 13345 3479 13379
rect 3421 13339 3479 13345
rect 4065 13379 4123 13385
rect 4065 13345 4077 13379
rect 4111 13376 4123 13379
rect 4154 13376 4160 13388
rect 4111 13348 4160 13376
rect 4111 13345 4123 13348
rect 4065 13339 4123 13345
rect 4154 13336 4160 13348
rect 4212 13336 4218 13388
rect 5166 13376 5172 13388
rect 5127 13348 5172 13376
rect 5166 13336 5172 13348
rect 5224 13336 5230 13388
rect 6917 13379 6975 13385
rect 6917 13345 6929 13379
rect 6963 13376 6975 13379
rect 7098 13376 7104 13388
rect 6963 13348 7104 13376
rect 6963 13345 6975 13348
rect 6917 13339 6975 13345
rect 7098 13336 7104 13348
rect 7156 13336 7162 13388
rect 23382 13336 23388 13388
rect 23440 13376 23446 13388
rect 24029 13379 24087 13385
rect 24029 13376 24041 13379
rect 23440 13348 24041 13376
rect 23440 13336 23446 13348
rect 24029 13345 24041 13348
rect 24075 13345 24087 13379
rect 24029 13339 24087 13345
rect 24305 13379 24363 13385
rect 24305 13345 24317 13379
rect 24351 13376 24363 13379
rect 26970 13376 26976 13388
rect 24351 13348 26976 13376
rect 24351 13345 24363 13348
rect 24305 13339 24363 13345
rect 26970 13336 26976 13348
rect 27028 13336 27034 13388
rect 33137 13379 33195 13385
rect 33137 13345 33149 13379
rect 33183 13376 33195 13379
rect 33410 13376 33416 13388
rect 33183 13348 33416 13376
rect 33183 13345 33195 13348
rect 33137 13339 33195 13345
rect 33410 13336 33416 13348
rect 33468 13376 33474 13388
rect 33689 13379 33747 13385
rect 33689 13376 33701 13379
rect 33468 13348 33701 13376
rect 33468 13336 33474 13348
rect 33689 13345 33701 13348
rect 33735 13345 33747 13379
rect 33689 13339 33747 13345
rect 34146 13336 34152 13388
rect 34204 13376 34210 13388
rect 34241 13379 34299 13385
rect 34241 13376 34253 13379
rect 34204 13348 34253 13376
rect 34204 13336 34210 13348
rect 34241 13345 34253 13348
rect 34287 13345 34299 13379
rect 34241 13339 34299 13345
rect 35250 13336 35256 13388
rect 35308 13376 35314 13388
rect 36556 13385 36584 13416
rect 35437 13379 35495 13385
rect 35437 13376 35449 13379
rect 35308 13348 35449 13376
rect 35308 13336 35314 13348
rect 35437 13345 35449 13348
rect 35483 13345 35495 13379
rect 35437 13339 35495 13345
rect 36547 13379 36605 13385
rect 36547 13345 36559 13379
rect 36593 13345 36605 13379
rect 36547 13339 36605 13345
rect 1596 13308 1624 13336
rect 6086 13308 6092 13320
rect 1596 13280 6092 13308
rect 6086 13268 6092 13280
rect 6144 13268 6150 13320
rect 32306 13268 32312 13320
rect 32364 13308 32370 13320
rect 34790 13308 34796 13320
rect 32364 13280 34796 13308
rect 32364 13268 32370 13280
rect 34790 13268 34796 13280
rect 34848 13268 34854 13320
rect 36556 13308 36584 13339
rect 37090 13308 37096 13320
rect 36556 13280 37096 13308
rect 37090 13268 37096 13280
rect 37148 13268 37154 13320
rect 4522 13200 4528 13252
rect 4580 13240 4586 13252
rect 11698 13240 11704 13252
rect 4580 13212 11704 13240
rect 4580 13200 4586 13212
rect 11698 13200 11704 13212
rect 11756 13200 11762 13252
rect 33321 13243 33379 13249
rect 33321 13209 33333 13243
rect 33367 13240 33379 13243
rect 34698 13240 34704 13252
rect 33367 13212 34704 13240
rect 33367 13209 33379 13212
rect 33321 13203 33379 13209
rect 34698 13200 34704 13212
rect 34756 13200 34762 13252
rect 1581 13175 1639 13181
rect 1581 13141 1593 13175
rect 1627 13172 1639 13175
rect 2774 13172 2780 13184
rect 1627 13144 2780 13172
rect 1627 13141 1639 13144
rect 1581 13135 1639 13141
rect 2774 13132 2780 13144
rect 2832 13132 2838 13184
rect 3510 13132 3516 13184
rect 3568 13172 3574 13184
rect 4249 13175 4307 13181
rect 4249 13172 4261 13175
rect 3568 13144 4261 13172
rect 3568 13132 3574 13144
rect 4249 13141 4261 13144
rect 4295 13141 4307 13175
rect 24854 13172 24860 13184
rect 24815 13144 24860 13172
rect 4249 13135 4307 13141
rect 24854 13132 24860 13144
rect 24912 13132 24918 13184
rect 33962 13132 33968 13184
rect 34020 13172 34026 13184
rect 34057 13175 34115 13181
rect 34057 13172 34069 13175
rect 34020 13144 34069 13172
rect 34020 13132 34026 13144
rect 34057 13141 34069 13144
rect 34103 13141 34115 13175
rect 34882 13172 34888 13184
rect 34843 13144 34888 13172
rect 34057 13135 34115 13141
rect 34882 13132 34888 13144
rect 34940 13132 34946 13184
rect 35434 13132 35440 13184
rect 35492 13172 35498 13184
rect 35621 13175 35679 13181
rect 35621 13172 35633 13175
rect 35492 13144 35633 13172
rect 35492 13132 35498 13144
rect 35621 13141 35633 13144
rect 35667 13141 35679 13175
rect 35621 13135 35679 13141
rect 35802 13132 35808 13184
rect 35860 13172 35866 13184
rect 36725 13175 36783 13181
rect 36725 13172 36737 13175
rect 35860 13144 36737 13172
rect 35860 13132 35866 13144
rect 36725 13141 36737 13144
rect 36771 13141 36783 13175
rect 36725 13135 36783 13141
rect 1104 13082 38824 13104
rect 1104 13030 7648 13082
rect 7700 13030 7712 13082
rect 7764 13030 7776 13082
rect 7828 13030 7840 13082
rect 7892 13030 20982 13082
rect 21034 13030 21046 13082
rect 21098 13030 21110 13082
rect 21162 13030 21174 13082
rect 21226 13030 34315 13082
rect 34367 13030 34379 13082
rect 34431 13030 34443 13082
rect 34495 13030 34507 13082
rect 34559 13030 38824 13082
rect 1104 13008 38824 13030
rect 1578 12968 1584 12980
rect 1539 12940 1584 12968
rect 1578 12928 1584 12940
rect 1636 12928 1642 12980
rect 4062 12928 4068 12980
rect 4120 12968 4126 12980
rect 6638 12968 6644 12980
rect 4120 12940 6644 12968
rect 4120 12928 4126 12940
rect 6638 12928 6644 12940
rect 6696 12928 6702 12980
rect 7466 12928 7472 12980
rect 7524 12968 7530 12980
rect 8297 12971 8355 12977
rect 8297 12968 8309 12971
rect 7524 12940 8309 12968
rect 7524 12928 7530 12940
rect 8297 12937 8309 12940
rect 8343 12937 8355 12971
rect 25498 12968 25504 12980
rect 8297 12931 8355 12937
rect 8404 12940 25504 12968
rect 2958 12860 2964 12912
rect 3016 12900 3022 12912
rect 4249 12903 4307 12909
rect 4249 12900 4261 12903
rect 3016 12872 4261 12900
rect 3016 12860 3022 12872
rect 4249 12869 4261 12872
rect 4295 12869 4307 12903
rect 8110 12900 8116 12912
rect 4249 12863 4307 12869
rect 7116 12872 8116 12900
rect 2133 12835 2191 12841
rect 2133 12801 2145 12835
rect 2179 12832 2191 12835
rect 3326 12832 3332 12844
rect 2179 12804 3332 12832
rect 2179 12801 2191 12804
rect 2133 12795 2191 12801
rect 3326 12792 3332 12804
rect 3384 12792 3390 12844
rect 3418 12792 3424 12844
rect 3476 12832 3482 12844
rect 7006 12832 7012 12844
rect 3476 12804 7012 12832
rect 3476 12792 3482 12804
rect 7006 12792 7012 12804
rect 7064 12792 7070 12844
rect 7116 12841 7144 12872
rect 8110 12860 8116 12872
rect 8168 12860 8174 12912
rect 7101 12835 7159 12841
rect 7101 12801 7113 12835
rect 7147 12801 7159 12835
rect 8404 12832 8432 12940
rect 25498 12928 25504 12940
rect 25556 12928 25562 12980
rect 31110 12928 31116 12980
rect 31168 12968 31174 12980
rect 34606 12968 34612 12980
rect 31168 12940 34612 12968
rect 31168 12928 31174 12940
rect 34606 12928 34612 12940
rect 34664 12928 34670 12980
rect 36357 12971 36415 12977
rect 36357 12937 36369 12971
rect 36403 12968 36415 12971
rect 36446 12968 36452 12980
rect 36403 12940 36452 12968
rect 36403 12937 36415 12940
rect 36357 12931 36415 12937
rect 36446 12928 36452 12940
rect 36504 12928 36510 12980
rect 37090 12968 37096 12980
rect 37051 12940 37096 12968
rect 37090 12928 37096 12940
rect 37148 12928 37154 12980
rect 11698 12860 11704 12912
rect 11756 12900 11762 12912
rect 19978 12900 19984 12912
rect 11756 12872 19984 12900
rect 11756 12860 11762 12872
rect 19978 12860 19984 12872
rect 20036 12860 20042 12912
rect 22922 12860 22928 12912
rect 22980 12900 22986 12912
rect 24581 12903 24639 12909
rect 24581 12900 24593 12903
rect 22980 12872 24593 12900
rect 22980 12860 22986 12872
rect 24581 12869 24593 12872
rect 24627 12869 24639 12903
rect 24581 12863 24639 12869
rect 25222 12860 25228 12912
rect 25280 12900 25286 12912
rect 32309 12903 32367 12909
rect 25280 12872 32168 12900
rect 25280 12860 25286 12872
rect 7101 12795 7159 12801
rect 8036 12804 8432 12832
rect 13265 12835 13323 12841
rect 1857 12767 1915 12773
rect 1857 12733 1869 12767
rect 1903 12764 1915 12767
rect 2038 12764 2044 12776
rect 1903 12736 2044 12764
rect 1903 12733 1915 12736
rect 1857 12727 1915 12733
rect 2038 12724 2044 12736
rect 2096 12764 2102 12776
rect 2593 12767 2651 12773
rect 2593 12764 2605 12767
rect 2096 12736 2605 12764
rect 2096 12724 2102 12736
rect 2593 12733 2605 12736
rect 2639 12733 2651 12767
rect 2593 12727 2651 12733
rect 3697 12767 3755 12773
rect 3697 12733 3709 12767
rect 3743 12764 3755 12767
rect 4154 12764 4160 12776
rect 3743 12736 4160 12764
rect 3743 12733 3755 12736
rect 3697 12727 3755 12733
rect 4154 12724 4160 12736
rect 4212 12764 4218 12776
rect 4614 12764 4620 12776
rect 4212 12736 4620 12764
rect 4212 12724 4218 12736
rect 4614 12724 4620 12736
rect 4672 12724 4678 12776
rect 6641 12767 6699 12773
rect 6641 12733 6653 12767
rect 6687 12764 6699 12767
rect 6825 12767 6883 12773
rect 6825 12764 6837 12767
rect 6687 12736 6837 12764
rect 6687 12733 6699 12736
rect 6641 12727 6699 12733
rect 6825 12733 6837 12736
rect 6871 12764 6883 12767
rect 7190 12764 7196 12776
rect 6871 12736 7196 12764
rect 6871 12733 6883 12736
rect 6825 12727 6883 12733
rect 7190 12724 7196 12736
rect 7248 12724 7254 12776
rect 3329 12699 3387 12705
rect 3329 12665 3341 12699
rect 3375 12696 3387 12699
rect 4062 12696 4068 12708
rect 3375 12668 4068 12696
rect 3375 12665 3387 12668
rect 3329 12659 3387 12665
rect 4062 12656 4068 12668
rect 4120 12656 4126 12708
rect 4522 12696 4528 12708
rect 4483 12668 4528 12696
rect 4522 12656 4528 12668
rect 4580 12656 4586 12708
rect 4798 12696 4804 12708
rect 4759 12668 4804 12696
rect 4798 12656 4804 12668
rect 4856 12656 4862 12708
rect 5166 12656 5172 12708
rect 5224 12696 5230 12708
rect 5261 12699 5319 12705
rect 5261 12696 5273 12699
rect 5224 12668 5273 12696
rect 5224 12656 5230 12668
rect 5261 12665 5273 12668
rect 5307 12696 5319 12699
rect 8036 12696 8064 12804
rect 13265 12801 13277 12835
rect 13311 12832 13323 12835
rect 15194 12832 15200 12844
rect 13311 12804 15200 12832
rect 13311 12801 13323 12804
rect 13265 12795 13323 12801
rect 15194 12792 15200 12804
rect 15252 12792 15258 12844
rect 16485 12835 16543 12841
rect 16485 12801 16497 12835
rect 16531 12832 16543 12835
rect 17586 12832 17592 12844
rect 16531 12804 17592 12832
rect 16531 12801 16543 12804
rect 16485 12795 16543 12801
rect 17586 12792 17592 12804
rect 17644 12792 17650 12844
rect 19061 12835 19119 12841
rect 19061 12801 19073 12835
rect 19107 12832 19119 12835
rect 19886 12832 19892 12844
rect 19107 12804 19892 12832
rect 19107 12801 19119 12804
rect 19061 12795 19119 12801
rect 19886 12792 19892 12804
rect 19944 12792 19950 12844
rect 22097 12835 22155 12841
rect 22097 12801 22109 12835
rect 22143 12832 22155 12835
rect 22278 12832 22284 12844
rect 22143 12804 22284 12832
rect 22143 12801 22155 12804
rect 22097 12795 22155 12801
rect 22278 12792 22284 12804
rect 22336 12792 22342 12844
rect 24854 12792 24860 12844
rect 24912 12832 24918 12844
rect 25133 12835 25191 12841
rect 25133 12832 25145 12835
rect 24912 12804 25145 12832
rect 24912 12792 24918 12804
rect 25133 12801 25145 12804
rect 25179 12832 25191 12835
rect 26510 12832 26516 12844
rect 25179 12804 26516 12832
rect 25179 12801 25191 12804
rect 25133 12795 25191 12801
rect 26510 12792 26516 12804
rect 26568 12792 26574 12844
rect 27617 12835 27675 12841
rect 27617 12801 27629 12835
rect 27663 12832 27675 12835
rect 29362 12832 29368 12844
rect 27663 12804 29368 12832
rect 27663 12801 27675 12804
rect 27617 12795 27675 12801
rect 29362 12792 29368 12804
rect 29420 12792 29426 12844
rect 31113 12835 31171 12841
rect 31113 12801 31125 12835
rect 31159 12832 31171 12835
rect 31662 12832 31668 12844
rect 31159 12804 31668 12832
rect 31159 12801 31171 12804
rect 31113 12795 31171 12801
rect 31662 12792 31668 12804
rect 31720 12792 31726 12844
rect 8113 12767 8171 12773
rect 8113 12733 8125 12767
rect 8159 12764 8171 12767
rect 8665 12767 8723 12773
rect 8665 12764 8677 12767
rect 8159 12736 8677 12764
rect 8159 12733 8171 12736
rect 8113 12727 8171 12733
rect 8665 12733 8677 12736
rect 8711 12733 8723 12767
rect 8665 12727 8723 12733
rect 10321 12767 10379 12773
rect 10321 12733 10333 12767
rect 10367 12764 10379 12767
rect 10367 12736 11192 12764
rect 10367 12733 10379 12736
rect 10321 12727 10379 12733
rect 5307 12668 8064 12696
rect 5307 12665 5319 12668
rect 5261 12659 5319 12665
rect 3973 12631 4031 12637
rect 3973 12597 3985 12631
rect 4019 12628 4031 12631
rect 4540 12628 4568 12656
rect 4706 12628 4712 12640
rect 4019 12600 4568 12628
rect 4667 12600 4712 12628
rect 4019 12597 4031 12600
rect 3973 12591 4031 12597
rect 4706 12588 4712 12600
rect 4764 12588 4770 12640
rect 5350 12588 5356 12640
rect 5408 12628 5414 12640
rect 5537 12631 5595 12637
rect 5537 12628 5549 12631
rect 5408 12600 5549 12628
rect 5408 12588 5414 12600
rect 5537 12597 5549 12600
rect 5583 12597 5595 12631
rect 5718 12628 5724 12640
rect 5679 12600 5724 12628
rect 5537 12591 5595 12597
rect 5718 12588 5724 12600
rect 5776 12588 5782 12640
rect 7098 12588 7104 12640
rect 7156 12628 7162 12640
rect 7561 12631 7619 12637
rect 7561 12628 7573 12631
rect 7156 12600 7573 12628
rect 7156 12588 7162 12600
rect 7561 12597 7573 12600
rect 7607 12597 7619 12631
rect 8680 12628 8708 12727
rect 10502 12656 10508 12708
rect 10560 12696 10566 12708
rect 11164 12705 11192 12736
rect 12526 12724 12532 12776
rect 12584 12764 12590 12776
rect 12989 12767 13047 12773
rect 12989 12764 13001 12767
rect 12584 12736 13001 12764
rect 12584 12724 12590 12736
rect 12989 12733 13001 12736
rect 13035 12764 13047 12767
rect 13725 12767 13783 12773
rect 13725 12764 13737 12767
rect 13035 12736 13737 12764
rect 13035 12733 13047 12736
rect 12989 12727 13047 12733
rect 13725 12733 13737 12736
rect 13771 12733 13783 12767
rect 13725 12727 13783 12733
rect 16209 12767 16267 12773
rect 16209 12733 16221 12767
rect 16255 12764 16267 12767
rect 16850 12764 16856 12776
rect 16255 12736 16856 12764
rect 16255 12733 16267 12736
rect 16209 12727 16267 12733
rect 16850 12724 16856 12736
rect 16908 12764 16914 12776
rect 16945 12767 17003 12773
rect 16945 12764 16957 12767
rect 16908 12736 16957 12764
rect 16908 12724 16914 12736
rect 16945 12733 16957 12736
rect 16991 12733 17003 12767
rect 16945 12727 17003 12733
rect 18785 12767 18843 12773
rect 18785 12733 18797 12767
rect 18831 12764 18843 12767
rect 19334 12764 19340 12776
rect 18831 12736 19340 12764
rect 18831 12733 18843 12736
rect 18785 12727 18843 12733
rect 19334 12724 19340 12736
rect 19392 12764 19398 12776
rect 19521 12767 19579 12773
rect 19521 12764 19533 12767
rect 19392 12736 19533 12764
rect 19392 12724 19398 12736
rect 19521 12733 19533 12736
rect 19567 12733 19579 12767
rect 19521 12727 19579 12733
rect 21821 12767 21879 12773
rect 21821 12733 21833 12767
rect 21867 12764 21879 12767
rect 22649 12767 22707 12773
rect 22649 12764 22661 12767
rect 21867 12736 22661 12764
rect 21867 12733 21879 12736
rect 21821 12727 21879 12733
rect 22649 12733 22661 12736
rect 22695 12764 22707 12767
rect 23474 12764 23480 12776
rect 22695 12736 23480 12764
rect 22695 12733 22707 12736
rect 22649 12727 22707 12733
rect 23474 12724 23480 12736
rect 23532 12724 23538 12776
rect 32140 12773 32168 12872
rect 32309 12869 32321 12903
rect 32355 12900 32367 12903
rect 33134 12900 33140 12912
rect 32355 12872 33140 12900
rect 32355 12869 32367 12872
rect 32309 12863 32367 12869
rect 33134 12860 33140 12872
rect 33192 12860 33198 12912
rect 33321 12903 33379 12909
rect 33321 12869 33333 12903
rect 33367 12900 33379 12903
rect 33367 12872 33456 12900
rect 33367 12869 33379 12872
rect 33321 12863 33379 12869
rect 33428 12832 33456 12872
rect 33502 12860 33508 12912
rect 33560 12900 33566 12912
rect 34790 12900 34796 12912
rect 33560 12872 34796 12900
rect 33560 12860 33566 12872
rect 34790 12860 34796 12872
rect 34848 12860 34854 12912
rect 33778 12832 33784 12844
rect 33428 12804 33640 12832
rect 33691 12804 33784 12832
rect 27341 12767 27399 12773
rect 27341 12733 27353 12767
rect 27387 12733 27399 12767
rect 27341 12727 27399 12733
rect 30837 12767 30895 12773
rect 30837 12733 30849 12767
rect 30883 12764 30895 12767
rect 31481 12767 31539 12773
rect 31481 12764 31493 12767
rect 30883 12736 31493 12764
rect 30883 12733 30895 12736
rect 30837 12727 30895 12733
rect 31481 12733 31493 12736
rect 31527 12764 31539 12767
rect 31573 12767 31631 12773
rect 31573 12764 31585 12767
rect 31527 12736 31585 12764
rect 31527 12733 31539 12736
rect 31481 12727 31539 12733
rect 31573 12733 31585 12736
rect 31619 12733 31631 12767
rect 31573 12727 31631 12733
rect 32125 12767 32183 12773
rect 32125 12733 32137 12767
rect 32171 12764 32183 12767
rect 32677 12767 32735 12773
rect 32677 12764 32689 12767
rect 32171 12736 32689 12764
rect 32171 12733 32183 12736
rect 32125 12727 32183 12733
rect 32677 12733 32689 12736
rect 32723 12733 32735 12767
rect 33612 12764 33640 12804
rect 33778 12792 33784 12804
rect 33836 12832 33842 12844
rect 34609 12835 34667 12841
rect 34609 12832 34621 12835
rect 33836 12804 34621 12832
rect 33836 12792 33842 12804
rect 34609 12801 34621 12804
rect 34655 12801 34667 12835
rect 34609 12795 34667 12801
rect 35161 12835 35219 12841
rect 35161 12801 35173 12835
rect 35207 12832 35219 12835
rect 36354 12832 36360 12844
rect 35207 12804 36360 12832
rect 35207 12801 35219 12804
rect 35161 12795 35219 12801
rect 36354 12792 36360 12804
rect 36412 12792 36418 12844
rect 34882 12764 34888 12776
rect 33612 12736 34888 12764
rect 32677 12727 32735 12733
rect 10597 12699 10655 12705
rect 10597 12696 10609 12699
rect 10560 12668 10609 12696
rect 10560 12656 10566 12668
rect 10597 12665 10609 12668
rect 10643 12665 10655 12699
rect 10597 12659 10655 12665
rect 11149 12699 11207 12705
rect 11149 12665 11161 12699
rect 11195 12696 11207 12699
rect 12894 12696 12900 12708
rect 11195 12668 12900 12696
rect 11195 12665 11207 12668
rect 11149 12659 11207 12665
rect 12894 12656 12900 12668
rect 12952 12656 12958 12708
rect 24029 12699 24087 12705
rect 24029 12665 24041 12699
rect 24075 12696 24087 12699
rect 24762 12696 24768 12708
rect 24075 12668 24768 12696
rect 24075 12665 24087 12668
rect 24029 12659 24087 12665
rect 24762 12656 24768 12668
rect 24820 12696 24826 12708
rect 24857 12699 24915 12705
rect 24857 12696 24869 12699
rect 24820 12668 24869 12696
rect 24820 12656 24826 12668
rect 24857 12665 24869 12668
rect 24903 12665 24915 12699
rect 27356 12696 27384 12727
rect 34882 12724 34888 12736
rect 34940 12724 34946 12776
rect 36170 12764 36176 12776
rect 36131 12736 36176 12764
rect 36170 12724 36176 12736
rect 36228 12764 36234 12776
rect 36725 12767 36783 12773
rect 36725 12764 36737 12767
rect 36228 12736 36737 12764
rect 36228 12724 36234 12736
rect 36725 12733 36737 12736
rect 36771 12733 36783 12767
rect 37274 12764 37280 12776
rect 37235 12736 37280 12764
rect 36725 12727 36783 12733
rect 37274 12724 37280 12736
rect 37332 12764 37338 12776
rect 37829 12767 37887 12773
rect 37829 12764 37841 12767
rect 37332 12736 37841 12764
rect 37332 12724 37338 12736
rect 37829 12733 37841 12736
rect 37875 12733 37887 12767
rect 37829 12727 37887 12733
rect 28169 12699 28227 12705
rect 28169 12696 28181 12699
rect 27356 12668 28181 12696
rect 24857 12659 24915 12665
rect 28169 12665 28181 12668
rect 28215 12696 28227 12699
rect 32030 12696 32036 12708
rect 28215 12668 32036 12696
rect 28215 12665 28227 12668
rect 28169 12659 28227 12665
rect 32030 12656 32036 12668
rect 32088 12656 32094 12708
rect 33502 12696 33508 12708
rect 32692 12668 33508 12696
rect 16206 12628 16212 12640
rect 8680 12600 16212 12628
rect 7561 12591 7619 12597
rect 16206 12588 16212 12600
rect 16264 12588 16270 12640
rect 22646 12588 22652 12640
rect 22704 12628 22710 12640
rect 23382 12628 23388 12640
rect 22704 12600 23388 12628
rect 22704 12588 22710 12600
rect 23382 12588 23388 12600
rect 23440 12628 23446 12640
rect 23477 12631 23535 12637
rect 23477 12628 23489 12631
rect 23440 12600 23489 12628
rect 23440 12588 23446 12600
rect 23477 12597 23489 12600
rect 23523 12597 23535 12631
rect 23477 12591 23535 12597
rect 24397 12631 24455 12637
rect 24397 12597 24409 12631
rect 24443 12628 24455 12631
rect 25041 12631 25099 12637
rect 25041 12628 25053 12631
rect 24443 12600 25053 12628
rect 24443 12597 24455 12600
rect 24397 12591 24455 12597
rect 25041 12597 25053 12600
rect 25087 12628 25099 12631
rect 25130 12628 25136 12640
rect 25087 12600 25136 12628
rect 25087 12597 25099 12600
rect 25041 12591 25099 12597
rect 25130 12588 25136 12600
rect 25188 12588 25194 12640
rect 31481 12631 31539 12637
rect 31481 12597 31493 12631
rect 31527 12628 31539 12631
rect 32692 12628 32720 12668
rect 33502 12656 33508 12668
rect 33560 12656 33566 12708
rect 33873 12699 33931 12705
rect 33873 12696 33885 12699
rect 33704 12668 33885 12696
rect 31527 12600 32720 12628
rect 33137 12631 33195 12637
rect 31527 12597 31539 12600
rect 31481 12591 31539 12597
rect 33137 12597 33149 12631
rect 33183 12628 33195 12631
rect 33704 12628 33732 12668
rect 33873 12665 33885 12668
rect 33919 12696 33931 12699
rect 36262 12696 36268 12708
rect 33919 12668 36268 12696
rect 33919 12665 33931 12668
rect 33873 12659 33931 12665
rect 36262 12656 36268 12668
rect 36320 12696 36326 12708
rect 38746 12696 38752 12708
rect 36320 12668 38752 12696
rect 36320 12656 36326 12668
rect 38746 12656 38752 12668
rect 38804 12656 38810 12708
rect 33183 12600 33732 12628
rect 33781 12631 33839 12637
rect 33183 12597 33195 12600
rect 33137 12591 33195 12597
rect 33781 12597 33793 12631
rect 33827 12628 33839 12631
rect 33962 12628 33968 12640
rect 33827 12600 33968 12628
rect 33827 12597 33839 12600
rect 33781 12591 33839 12597
rect 33962 12588 33968 12600
rect 34020 12588 34026 12640
rect 34330 12628 34336 12640
rect 34291 12600 34336 12628
rect 34330 12588 34336 12600
rect 34388 12588 34394 12640
rect 35250 12588 35256 12640
rect 35308 12628 35314 12640
rect 35621 12631 35679 12637
rect 35621 12628 35633 12631
rect 35308 12600 35633 12628
rect 35308 12588 35314 12600
rect 35621 12597 35633 12600
rect 35667 12597 35679 12631
rect 37458 12628 37464 12640
rect 37419 12600 37464 12628
rect 35621 12591 35679 12597
rect 37458 12588 37464 12600
rect 37516 12588 37522 12640
rect 1104 12538 38824 12560
rect 1104 12486 14315 12538
rect 14367 12486 14379 12538
rect 14431 12486 14443 12538
rect 14495 12486 14507 12538
rect 14559 12486 27648 12538
rect 27700 12486 27712 12538
rect 27764 12486 27776 12538
rect 27828 12486 27840 12538
rect 27892 12486 38824 12538
rect 1104 12464 38824 12486
rect 4154 12384 4160 12436
rect 4212 12424 4218 12436
rect 4706 12424 4712 12436
rect 4212 12396 4712 12424
rect 4212 12384 4218 12396
rect 4706 12384 4712 12396
rect 4764 12384 4770 12436
rect 6638 12424 6644 12436
rect 6599 12396 6644 12424
rect 6638 12384 6644 12396
rect 6696 12384 6702 12436
rect 31110 12424 31116 12436
rect 31071 12396 31116 12424
rect 31110 12384 31116 12396
rect 31168 12384 31174 12436
rect 32306 12424 32312 12436
rect 32267 12396 32312 12424
rect 32306 12384 32312 12396
rect 32364 12384 32370 12436
rect 36173 12427 36231 12433
rect 36173 12393 36185 12427
rect 36219 12424 36231 12427
rect 36262 12424 36268 12436
rect 36219 12396 36268 12424
rect 36219 12393 36231 12396
rect 36173 12387 36231 12393
rect 36262 12384 36268 12396
rect 36320 12384 36326 12436
rect 1118 12316 1124 12368
rect 1176 12356 1182 12368
rect 1673 12359 1731 12365
rect 1673 12356 1685 12359
rect 1176 12328 1685 12356
rect 1176 12316 1182 12328
rect 1673 12325 1685 12328
rect 1719 12325 1731 12359
rect 1673 12319 1731 12325
rect 4801 12359 4859 12365
rect 4801 12325 4813 12359
rect 4847 12356 4859 12359
rect 5258 12356 5264 12368
rect 4847 12328 5264 12356
rect 4847 12325 4859 12328
rect 4801 12319 4859 12325
rect 5258 12316 5264 12328
rect 5316 12356 5322 12368
rect 5445 12359 5503 12365
rect 5445 12356 5457 12359
rect 5316 12328 5457 12356
rect 5316 12316 5322 12328
rect 5445 12325 5457 12328
rect 5491 12325 5503 12359
rect 8481 12359 8539 12365
rect 8481 12356 8493 12359
rect 5445 12319 5503 12325
rect 7760 12328 8493 12356
rect 1397 12291 1455 12297
rect 1397 12257 1409 12291
rect 1443 12288 1455 12291
rect 2498 12288 2504 12300
rect 1443 12260 2504 12288
rect 1443 12257 1455 12260
rect 1397 12251 1455 12257
rect 2498 12248 2504 12260
rect 2556 12248 2562 12300
rect 2682 12288 2688 12300
rect 2643 12260 2688 12288
rect 2682 12248 2688 12260
rect 2740 12248 2746 12300
rect 6270 12248 6276 12300
rect 6328 12288 6334 12300
rect 6457 12291 6515 12297
rect 6457 12288 6469 12291
rect 6328 12260 6469 12288
rect 6328 12248 6334 12260
rect 6457 12257 6469 12260
rect 6503 12257 6515 12291
rect 6457 12251 6515 12257
rect 5350 12220 5356 12232
rect 5311 12192 5356 12220
rect 5350 12180 5356 12192
rect 5408 12180 5414 12232
rect 5537 12223 5595 12229
rect 5537 12189 5549 12223
rect 5583 12220 5595 12223
rect 5626 12220 5632 12232
rect 5583 12192 5632 12220
rect 5583 12189 5595 12192
rect 5537 12183 5595 12189
rect 5626 12180 5632 12192
rect 5684 12180 5690 12232
rect 2225 12087 2283 12093
rect 2225 12053 2237 12087
rect 2271 12084 2283 12087
rect 2590 12084 2596 12096
rect 2271 12056 2596 12084
rect 2271 12053 2283 12056
rect 2225 12047 2283 12053
rect 2590 12044 2596 12056
rect 2648 12044 2654 12096
rect 2866 12084 2872 12096
rect 2827 12056 2872 12084
rect 2866 12044 2872 12056
rect 2924 12044 2930 12096
rect 3602 12084 3608 12096
rect 3563 12056 3608 12084
rect 3602 12044 3608 12056
rect 3660 12044 3666 12096
rect 4338 12084 4344 12096
rect 4299 12056 4344 12084
rect 4338 12044 4344 12056
rect 4396 12084 4402 12096
rect 4798 12084 4804 12096
rect 4396 12056 4804 12084
rect 4396 12044 4402 12056
rect 4798 12044 4804 12056
rect 4856 12044 4862 12096
rect 4982 12084 4988 12096
rect 4943 12056 4988 12084
rect 4982 12044 4988 12056
rect 5040 12044 5046 12096
rect 5902 12084 5908 12096
rect 5863 12056 5908 12084
rect 5902 12044 5908 12056
rect 5960 12044 5966 12096
rect 7466 12044 7472 12096
rect 7524 12084 7530 12096
rect 7760 12093 7788 12328
rect 8481 12325 8493 12328
rect 8527 12325 8539 12359
rect 8481 12319 8539 12325
rect 11698 12316 11704 12368
rect 11756 12356 11762 12368
rect 11977 12359 12035 12365
rect 11977 12356 11989 12359
rect 11756 12328 11989 12356
rect 11756 12316 11762 12328
rect 11977 12325 11989 12328
rect 12023 12325 12035 12359
rect 11977 12319 12035 12325
rect 17773 12359 17831 12365
rect 17773 12325 17785 12359
rect 17819 12356 17831 12359
rect 17862 12356 17868 12368
rect 17819 12328 17868 12356
rect 17819 12325 17831 12328
rect 17773 12319 17831 12325
rect 17862 12316 17868 12328
rect 17920 12316 17926 12368
rect 21358 12316 21364 12368
rect 21416 12356 21422 12368
rect 21453 12359 21511 12365
rect 21453 12356 21465 12359
rect 21416 12328 21465 12356
rect 21416 12316 21422 12328
rect 21453 12325 21465 12328
rect 21499 12325 21511 12359
rect 21453 12319 21511 12325
rect 24949 12359 25007 12365
rect 24949 12325 24961 12359
rect 24995 12356 25007 12359
rect 25038 12356 25044 12368
rect 24995 12328 25044 12356
rect 24995 12325 25007 12328
rect 24949 12319 25007 12325
rect 25038 12316 25044 12328
rect 25096 12316 25102 12368
rect 33781 12359 33839 12365
rect 33781 12325 33793 12359
rect 33827 12356 33839 12359
rect 34057 12359 34115 12365
rect 34057 12356 34069 12359
rect 33827 12328 34069 12356
rect 33827 12325 33839 12328
rect 33781 12319 33839 12325
rect 34057 12325 34069 12328
rect 34103 12325 34115 12359
rect 34057 12319 34115 12325
rect 8294 12288 8300 12300
rect 8255 12260 8300 12288
rect 8294 12248 8300 12260
rect 8352 12248 8358 12300
rect 30929 12291 30987 12297
rect 30929 12257 30941 12291
rect 30975 12288 30987 12291
rect 31294 12288 31300 12300
rect 30975 12260 31300 12288
rect 30975 12257 30987 12260
rect 30929 12251 30987 12257
rect 31294 12248 31300 12260
rect 31352 12248 31358 12300
rect 32125 12291 32183 12297
rect 32125 12257 32137 12291
rect 32171 12288 32183 12291
rect 32950 12288 32956 12300
rect 32171 12260 32956 12288
rect 32171 12257 32183 12260
rect 32125 12251 32183 12257
rect 32950 12248 32956 12260
rect 33008 12248 33014 12300
rect 33318 12248 33324 12300
rect 33376 12288 33382 12300
rect 33597 12291 33655 12297
rect 33597 12288 33609 12291
rect 33376 12260 33609 12288
rect 33376 12248 33382 12260
rect 33597 12257 33609 12260
rect 33643 12288 33655 12291
rect 34609 12291 34667 12297
rect 34609 12288 34621 12291
rect 33643 12260 34621 12288
rect 33643 12257 33655 12260
rect 33597 12251 33655 12257
rect 34609 12257 34621 12260
rect 34655 12257 34667 12291
rect 35049 12291 35107 12297
rect 35049 12288 35061 12291
rect 34609 12251 34667 12257
rect 34716 12260 35061 12288
rect 8570 12220 8576 12232
rect 8531 12192 8576 12220
rect 8570 12180 8576 12192
rect 8628 12180 8634 12232
rect 11882 12220 11888 12232
rect 11843 12192 11888 12220
rect 11882 12180 11888 12192
rect 11940 12180 11946 12232
rect 12069 12223 12127 12229
rect 12069 12189 12081 12223
rect 12115 12220 12127 12223
rect 12250 12220 12256 12232
rect 12115 12192 12256 12220
rect 12115 12189 12127 12192
rect 12069 12183 12127 12189
rect 12250 12180 12256 12192
rect 12308 12180 12314 12232
rect 17770 12220 17776 12232
rect 17731 12192 17776 12220
rect 17770 12180 17776 12192
rect 17828 12180 17834 12232
rect 17865 12223 17923 12229
rect 17865 12189 17877 12223
rect 17911 12189 17923 12223
rect 17865 12183 17923 12189
rect 21453 12223 21511 12229
rect 21453 12189 21465 12223
rect 21499 12189 21511 12223
rect 21453 12183 21511 12189
rect 21545 12223 21603 12229
rect 21545 12189 21557 12223
rect 21591 12220 21603 12223
rect 21818 12220 21824 12232
rect 21591 12192 21824 12220
rect 21591 12189 21603 12192
rect 21545 12183 21603 12189
rect 17494 12112 17500 12164
rect 17552 12152 17558 12164
rect 17880 12152 17908 12183
rect 17552 12124 17908 12152
rect 21468 12152 21496 12183
rect 21818 12180 21824 12192
rect 21876 12180 21882 12232
rect 24946 12220 24952 12232
rect 24907 12192 24952 12220
rect 24946 12180 24952 12192
rect 25004 12180 25010 12232
rect 25041 12223 25099 12229
rect 25041 12189 25053 12223
rect 25087 12220 25099 12223
rect 25866 12220 25872 12232
rect 25087 12192 25872 12220
rect 25087 12189 25099 12192
rect 25041 12183 25099 12189
rect 25866 12180 25872 12192
rect 25924 12180 25930 12232
rect 33873 12223 33931 12229
rect 33873 12220 33885 12223
rect 32784 12192 33885 12220
rect 21726 12152 21732 12164
rect 21468 12124 21732 12152
rect 17552 12112 17558 12124
rect 21726 12112 21732 12124
rect 21784 12112 21790 12164
rect 23661 12155 23719 12161
rect 23661 12121 23673 12155
rect 23707 12152 23719 12155
rect 24394 12152 24400 12164
rect 23707 12124 24400 12152
rect 23707 12121 23719 12124
rect 23661 12115 23719 12121
rect 24394 12112 24400 12124
rect 24452 12152 24458 12164
rect 24489 12155 24547 12161
rect 24489 12152 24501 12155
rect 24452 12124 24501 12152
rect 24452 12112 24458 12124
rect 24489 12121 24501 12124
rect 24535 12121 24547 12155
rect 24489 12115 24547 12121
rect 32784 12096 32812 12192
rect 33873 12189 33885 12192
rect 33919 12220 33931 12223
rect 34716 12220 34744 12260
rect 35049 12257 35061 12260
rect 35095 12288 35107 12291
rect 36262 12288 36268 12300
rect 35095 12260 36268 12288
rect 35095 12257 35107 12260
rect 35049 12251 35107 12257
rect 36262 12248 36268 12260
rect 36320 12248 36326 12300
rect 33919 12192 34744 12220
rect 34793 12223 34851 12229
rect 33919 12189 33931 12192
rect 33873 12183 33931 12189
rect 34793 12189 34805 12223
rect 34839 12189 34851 12223
rect 34793 12183 34851 12189
rect 33321 12155 33379 12161
rect 33321 12121 33333 12155
rect 33367 12152 33379 12155
rect 33778 12152 33784 12164
rect 33367 12124 33784 12152
rect 33367 12121 33379 12124
rect 33321 12115 33379 12121
rect 33778 12112 33784 12124
rect 33836 12112 33842 12164
rect 34606 12112 34612 12164
rect 34664 12152 34670 12164
rect 34808 12152 34836 12183
rect 34664 12124 34836 12152
rect 34664 12112 34670 12124
rect 7745 12087 7803 12093
rect 7745 12084 7757 12087
rect 7524 12056 7757 12084
rect 7524 12044 7530 12056
rect 7745 12053 7757 12056
rect 7791 12053 7803 12087
rect 8018 12084 8024 12096
rect 7979 12056 8024 12084
rect 7745 12047 7803 12053
rect 8018 12044 8024 12056
rect 8076 12044 8082 12096
rect 8938 12084 8944 12096
rect 8899 12056 8944 12084
rect 8938 12044 8944 12056
rect 8996 12044 9002 12096
rect 11054 12044 11060 12096
rect 11112 12084 11118 12096
rect 11149 12087 11207 12093
rect 11149 12084 11161 12087
rect 11112 12056 11161 12084
rect 11112 12044 11118 12056
rect 11149 12053 11161 12056
rect 11195 12084 11207 12087
rect 11517 12087 11575 12093
rect 11517 12084 11529 12087
rect 11195 12056 11529 12084
rect 11195 12053 11207 12056
rect 11149 12047 11207 12053
rect 11517 12053 11529 12056
rect 11563 12053 11575 12087
rect 12986 12084 12992 12096
rect 12947 12056 12992 12084
rect 11517 12047 11575 12053
rect 12986 12044 12992 12056
rect 13044 12044 13050 12096
rect 15838 12044 15844 12096
rect 15896 12084 15902 12096
rect 16393 12087 16451 12093
rect 16393 12084 16405 12087
rect 15896 12056 16405 12084
rect 15896 12044 15902 12056
rect 16393 12053 16405 12056
rect 16439 12053 16451 12087
rect 16393 12047 16451 12053
rect 16945 12087 17003 12093
rect 16945 12053 16957 12087
rect 16991 12084 17003 12087
rect 17313 12087 17371 12093
rect 17313 12084 17325 12087
rect 16991 12056 17325 12084
rect 16991 12053 17003 12056
rect 16945 12047 17003 12053
rect 17313 12053 17325 12056
rect 17359 12084 17371 12087
rect 17402 12084 17408 12096
rect 17359 12056 17408 12084
rect 17359 12053 17371 12056
rect 17313 12047 17371 12053
rect 17402 12044 17408 12056
rect 17460 12044 17466 12096
rect 18230 12044 18236 12096
rect 18288 12084 18294 12096
rect 19429 12087 19487 12093
rect 19429 12084 19441 12087
rect 18288 12056 19441 12084
rect 18288 12044 18294 12056
rect 19429 12053 19441 12056
rect 19475 12053 19487 12087
rect 19429 12047 19487 12053
rect 20622 12044 20628 12096
rect 20680 12084 20686 12096
rect 20993 12087 21051 12093
rect 20993 12084 21005 12087
rect 20680 12056 21005 12084
rect 20680 12044 20686 12056
rect 20993 12053 21005 12056
rect 21039 12053 21051 12087
rect 20993 12047 21051 12053
rect 24029 12087 24087 12093
rect 24029 12053 24041 12087
rect 24075 12084 24087 12087
rect 24670 12084 24676 12096
rect 24075 12056 24676 12084
rect 24075 12053 24087 12056
rect 24029 12047 24087 12053
rect 24670 12044 24676 12056
rect 24728 12044 24734 12096
rect 25498 12044 25504 12096
rect 25556 12084 25562 12096
rect 25593 12087 25651 12093
rect 25593 12084 25605 12087
rect 25556 12056 25605 12084
rect 25556 12044 25562 12056
rect 25593 12053 25605 12056
rect 25639 12084 25651 12087
rect 25958 12084 25964 12096
rect 25639 12056 25964 12084
rect 25639 12053 25651 12056
rect 25593 12047 25651 12053
rect 25958 12044 25964 12056
rect 26016 12044 26022 12096
rect 27157 12087 27215 12093
rect 27157 12053 27169 12087
rect 27203 12084 27215 12087
rect 27430 12084 27436 12096
rect 27203 12056 27436 12084
rect 27203 12053 27215 12056
rect 27157 12047 27215 12053
rect 27430 12044 27436 12056
rect 27488 12044 27494 12096
rect 30190 12084 30196 12096
rect 30151 12056 30196 12084
rect 30190 12044 30196 12056
rect 30248 12044 30254 12096
rect 30561 12087 30619 12093
rect 30561 12053 30573 12087
rect 30607 12084 30619 12087
rect 31018 12084 31024 12096
rect 30607 12056 31024 12084
rect 30607 12053 30619 12056
rect 30561 12047 30619 12053
rect 31018 12044 31024 12056
rect 31076 12044 31082 12096
rect 32766 12084 32772 12096
rect 32727 12056 32772 12084
rect 32766 12044 32772 12056
rect 32824 12044 32830 12096
rect 33137 12087 33195 12093
rect 33137 12053 33149 12087
rect 33183 12084 33195 12087
rect 33686 12084 33692 12096
rect 33183 12056 33692 12084
rect 33183 12053 33195 12056
rect 33137 12047 33195 12053
rect 33686 12044 33692 12056
rect 33744 12044 33750 12096
rect 34057 12087 34115 12093
rect 34057 12053 34069 12087
rect 34103 12084 34115 12087
rect 34333 12087 34391 12093
rect 34333 12084 34345 12087
rect 34103 12056 34345 12084
rect 34103 12053 34115 12056
rect 34057 12047 34115 12053
rect 34333 12053 34345 12056
rect 34379 12084 34391 12087
rect 35526 12084 35532 12096
rect 34379 12056 35532 12084
rect 34379 12053 34391 12056
rect 34333 12047 34391 12053
rect 35526 12044 35532 12056
rect 35584 12044 35590 12096
rect 1104 11994 38824 12016
rect 1104 11942 7648 11994
rect 7700 11942 7712 11994
rect 7764 11942 7776 11994
rect 7828 11942 7840 11994
rect 7892 11942 20982 11994
rect 21034 11942 21046 11994
rect 21098 11942 21110 11994
rect 21162 11942 21174 11994
rect 21226 11942 34315 11994
rect 34367 11942 34379 11994
rect 34431 11942 34443 11994
rect 34495 11942 34507 11994
rect 34559 11942 38824 11994
rect 1104 11920 38824 11942
rect 2498 11840 2504 11892
rect 2556 11880 2562 11892
rect 3605 11883 3663 11889
rect 3605 11880 3617 11883
rect 2556 11852 3617 11880
rect 2556 11840 2562 11852
rect 3605 11849 3617 11852
rect 3651 11849 3663 11883
rect 3605 11843 3663 11849
rect 4706 11840 4712 11892
rect 4764 11880 4770 11892
rect 5169 11883 5227 11889
rect 5169 11880 5181 11883
rect 4764 11852 5181 11880
rect 4764 11840 4770 11852
rect 5169 11849 5181 11852
rect 5215 11849 5227 11883
rect 7006 11880 7012 11892
rect 6967 11852 7012 11880
rect 5169 11843 5227 11849
rect 7006 11840 7012 11852
rect 7064 11840 7070 11892
rect 8294 11880 8300 11892
rect 7944 11852 8300 11880
rect 1670 11772 1676 11824
rect 1728 11812 1734 11824
rect 2041 11815 2099 11821
rect 2041 11812 2053 11815
rect 1728 11784 2053 11812
rect 1728 11772 1734 11784
rect 2041 11781 2053 11784
rect 2087 11781 2099 11815
rect 2041 11775 2099 11781
rect 2682 11772 2688 11824
rect 2740 11812 2746 11824
rect 3053 11815 3111 11821
rect 3053 11812 3065 11815
rect 2740 11784 3065 11812
rect 2740 11772 2746 11784
rect 3053 11781 3065 11784
rect 3099 11812 3111 11815
rect 4341 11815 4399 11821
rect 4341 11812 4353 11815
rect 3099 11784 4353 11812
rect 3099 11781 3111 11784
rect 3053 11775 3111 11781
rect 4341 11781 4353 11784
rect 4387 11781 4399 11815
rect 4341 11775 4399 11781
rect 1857 11747 1915 11753
rect 1857 11713 1869 11747
rect 1903 11744 1915 11747
rect 2498 11744 2504 11756
rect 1903 11716 2504 11744
rect 1903 11713 1915 11716
rect 1857 11707 1915 11713
rect 2498 11704 2504 11716
rect 2556 11704 2562 11756
rect 2590 11704 2596 11756
rect 2648 11744 2654 11756
rect 2648 11716 2693 11744
rect 2648 11704 2654 11716
rect 3602 11704 3608 11756
rect 3660 11744 3666 11756
rect 4065 11747 4123 11753
rect 4065 11744 4077 11747
rect 3660 11716 4077 11744
rect 3660 11704 3666 11716
rect 4065 11713 4077 11716
rect 4111 11744 4123 11747
rect 4982 11744 4988 11756
rect 4111 11716 4988 11744
rect 4111 11713 4123 11716
rect 4065 11707 4123 11713
rect 4982 11704 4988 11716
rect 5040 11704 5046 11756
rect 5721 11747 5779 11753
rect 5721 11713 5733 11747
rect 5767 11744 5779 11747
rect 5902 11744 5908 11756
rect 5767 11716 5908 11744
rect 5767 11713 5779 11716
rect 5721 11707 5779 11713
rect 5902 11704 5908 11716
rect 5960 11704 5966 11756
rect 7374 11704 7380 11756
rect 7432 11744 7438 11756
rect 7944 11753 7972 11852
rect 8294 11840 8300 11852
rect 8352 11840 8358 11892
rect 10686 11880 10692 11892
rect 10647 11852 10692 11880
rect 10686 11840 10692 11852
rect 10744 11880 10750 11892
rect 10962 11880 10968 11892
rect 10744 11852 10968 11880
rect 10744 11840 10750 11852
rect 10962 11840 10968 11852
rect 11020 11840 11026 11892
rect 17494 11880 17500 11892
rect 17455 11852 17500 11880
rect 17494 11840 17500 11852
rect 17552 11840 17558 11892
rect 25038 11880 25044 11892
rect 24999 11852 25044 11880
rect 25038 11840 25044 11852
rect 25096 11840 25102 11892
rect 26510 11880 26516 11892
rect 26471 11852 26516 11880
rect 26510 11840 26516 11852
rect 26568 11880 26574 11892
rect 29546 11880 29552 11892
rect 26568 11852 27752 11880
rect 29507 11852 29552 11880
rect 26568 11840 26574 11852
rect 8018 11772 8024 11824
rect 8076 11812 8082 11824
rect 8205 11815 8263 11821
rect 8205 11812 8217 11815
rect 8076 11784 8217 11812
rect 8076 11772 8082 11784
rect 8205 11781 8217 11784
rect 8251 11781 8263 11815
rect 8205 11775 8263 11781
rect 12989 11815 13047 11821
rect 12989 11781 13001 11815
rect 13035 11812 13047 11815
rect 13170 11812 13176 11824
rect 13035 11784 13176 11812
rect 13035 11781 13047 11784
rect 12989 11775 13047 11781
rect 13170 11772 13176 11784
rect 13228 11772 13234 11824
rect 16482 11812 16488 11824
rect 16443 11784 16488 11812
rect 16482 11772 16488 11784
rect 16540 11772 16546 11824
rect 23750 11772 23756 11824
rect 23808 11812 23814 11824
rect 24029 11815 24087 11821
rect 24029 11812 24041 11815
rect 23808 11784 24041 11812
rect 23808 11772 23814 11784
rect 24029 11781 24041 11784
rect 24075 11781 24087 11815
rect 25593 11815 25651 11821
rect 25593 11812 25605 11815
rect 24029 11775 24087 11781
rect 24504 11784 25605 11812
rect 7929 11747 7987 11753
rect 7929 11744 7941 11747
rect 7432 11716 7941 11744
rect 7432 11704 7438 11716
rect 7929 11713 7941 11716
rect 7975 11713 7987 11747
rect 7929 11707 7987 11713
rect 8110 11704 8116 11756
rect 8168 11744 8174 11756
rect 8665 11747 8723 11753
rect 8665 11744 8677 11747
rect 8168 11716 8677 11744
rect 8168 11704 8174 11716
rect 8665 11713 8677 11716
rect 8711 11744 8723 11747
rect 9493 11747 9551 11753
rect 9493 11744 9505 11747
rect 8711 11716 9505 11744
rect 8711 11713 8723 11716
rect 8665 11707 8723 11713
rect 9493 11713 9505 11716
rect 9539 11713 9551 11747
rect 9493 11707 9551 11713
rect 11333 11747 11391 11753
rect 11333 11713 11345 11747
rect 11379 11744 11391 11747
rect 12802 11744 12808 11756
rect 11379 11716 12808 11744
rect 11379 11713 11391 11716
rect 11333 11707 11391 11713
rect 12802 11704 12808 11716
rect 12860 11704 12866 11756
rect 16942 11744 16948 11756
rect 16855 11716 16948 11744
rect 16942 11704 16948 11716
rect 17000 11744 17006 11756
rect 18049 11747 18107 11753
rect 18049 11744 18061 11747
rect 17000 11716 18061 11744
rect 17000 11704 17006 11716
rect 18049 11713 18061 11716
rect 18095 11713 18107 11747
rect 24394 11744 24400 11756
rect 24355 11716 24400 11744
rect 18049 11707 18107 11713
rect 24394 11704 24400 11716
rect 24452 11704 24458 11756
rect 5626 11636 5632 11688
rect 5684 11676 5690 11688
rect 6089 11679 6147 11685
rect 6089 11676 6101 11679
rect 5684 11648 6101 11676
rect 5684 11636 5690 11648
rect 6089 11645 6101 11648
rect 6135 11645 6147 11679
rect 6822 11676 6828 11688
rect 6735 11648 6828 11676
rect 6089 11639 6147 11645
rect 6822 11636 6828 11648
rect 6880 11676 6886 11688
rect 11054 11676 11060 11688
rect 6880 11648 7512 11676
rect 11015 11648 11060 11676
rect 6880 11636 6886 11648
rect 2406 11568 2412 11620
rect 2464 11608 2470 11620
rect 2501 11611 2559 11617
rect 2501 11608 2513 11611
rect 2464 11580 2513 11608
rect 2464 11568 2470 11580
rect 2501 11577 2513 11580
rect 2547 11577 2559 11611
rect 2501 11571 2559 11577
rect 3421 11611 3479 11617
rect 3421 11577 3433 11611
rect 3467 11608 3479 11611
rect 4154 11608 4160 11620
rect 3467 11580 4160 11608
rect 3467 11577 3479 11580
rect 3421 11571 3479 11577
rect 4154 11568 4160 11580
rect 4212 11568 4218 11620
rect 4341 11611 4399 11617
rect 4341 11577 4353 11611
rect 4387 11608 4399 11611
rect 4617 11611 4675 11617
rect 4617 11608 4629 11611
rect 4387 11580 4629 11608
rect 4387 11577 4399 11580
rect 4341 11571 4399 11577
rect 4617 11577 4629 11580
rect 4663 11608 4675 11611
rect 5445 11611 5503 11617
rect 5445 11608 5457 11611
rect 4663 11580 5457 11608
rect 4663 11577 4675 11580
rect 4617 11571 4675 11577
rect 5445 11577 5457 11580
rect 5491 11608 5503 11611
rect 5994 11608 6000 11620
rect 5491 11580 6000 11608
rect 5491 11577 5503 11580
rect 5445 11571 5503 11577
rect 5994 11568 6000 11580
rect 6052 11568 6058 11620
rect 3602 11500 3608 11552
rect 3660 11540 3666 11552
rect 4065 11543 4123 11549
rect 4065 11540 4077 11543
rect 3660 11512 4077 11540
rect 3660 11500 3666 11512
rect 4065 11509 4077 11512
rect 4111 11509 4123 11543
rect 4890 11540 4896 11552
rect 4851 11512 4896 11540
rect 4065 11503 4123 11509
rect 4890 11500 4896 11512
rect 4948 11540 4954 11552
rect 5629 11543 5687 11549
rect 5629 11540 5641 11543
rect 4948 11512 5641 11540
rect 4948 11500 4954 11512
rect 5629 11509 5641 11512
rect 5675 11509 5687 11543
rect 5629 11503 5687 11509
rect 6270 11500 6276 11552
rect 6328 11540 6334 11552
rect 7484 11549 7512 11648
rect 11054 11636 11060 11648
rect 11112 11636 11118 11688
rect 12253 11679 12311 11685
rect 12253 11645 12265 11679
rect 12299 11676 12311 11679
rect 13446 11676 13452 11688
rect 12299 11648 13452 11676
rect 12299 11645 12311 11648
rect 12253 11639 12311 11645
rect 13446 11636 13452 11648
rect 13504 11676 13510 11688
rect 13541 11679 13599 11685
rect 13541 11676 13553 11679
rect 13504 11648 13553 11676
rect 13504 11636 13510 11648
rect 13541 11645 13553 11648
rect 13587 11645 13599 11679
rect 13541 11639 13599 11645
rect 19337 11679 19395 11685
rect 19337 11645 19349 11679
rect 19383 11676 19395 11679
rect 19429 11679 19487 11685
rect 19429 11676 19441 11679
rect 19383 11648 19441 11676
rect 19383 11645 19395 11648
rect 19337 11639 19395 11645
rect 19429 11645 19441 11648
rect 19475 11676 19487 11679
rect 20898 11676 20904 11688
rect 19475 11648 20904 11676
rect 19475 11645 19487 11648
rect 19429 11639 19487 11645
rect 20898 11636 20904 11648
rect 20956 11636 20962 11688
rect 8570 11568 8576 11620
rect 8628 11608 8634 11620
rect 8757 11611 8815 11617
rect 8757 11608 8769 11611
rect 8628 11580 8769 11608
rect 8628 11568 8634 11580
rect 8757 11577 8769 11580
rect 8803 11608 8815 11611
rect 8803 11580 9168 11608
rect 8803 11577 8815 11580
rect 8757 11571 8815 11577
rect 9140 11552 9168 11580
rect 12986 11568 12992 11620
rect 13044 11608 13050 11620
rect 13265 11611 13323 11617
rect 13265 11608 13277 11611
rect 13044 11580 13277 11608
rect 13044 11568 13050 11580
rect 13265 11577 13277 11580
rect 13311 11577 13323 11611
rect 13265 11571 13323 11577
rect 15381 11611 15439 11617
rect 15381 11577 15393 11611
rect 15427 11608 15439 11611
rect 15838 11608 15844 11620
rect 15427 11580 15844 11608
rect 15427 11577 15439 11580
rect 15381 11571 15439 11577
rect 15838 11568 15844 11580
rect 15896 11608 15902 11620
rect 17037 11611 17095 11617
rect 17037 11608 17049 11611
rect 15896 11580 17049 11608
rect 15896 11568 15902 11580
rect 17037 11577 17049 11580
rect 17083 11608 17095 11611
rect 17678 11608 17684 11620
rect 17083 11580 17684 11608
rect 17083 11577 17095 11580
rect 17037 11571 17095 11577
rect 17678 11568 17684 11580
rect 17736 11568 17742 11620
rect 17770 11568 17776 11620
rect 17828 11608 17834 11620
rect 18601 11611 18659 11617
rect 18601 11608 18613 11611
rect 17828 11580 18613 11608
rect 17828 11568 17834 11580
rect 18601 11577 18613 11580
rect 18647 11608 18659 11611
rect 19518 11608 19524 11620
rect 18647 11580 19524 11608
rect 18647 11577 18659 11580
rect 18601 11571 18659 11577
rect 19518 11568 19524 11580
rect 19576 11568 19582 11620
rect 19610 11568 19616 11620
rect 19668 11617 19674 11620
rect 24504 11617 24532 11784
rect 25593 11781 25605 11784
rect 25639 11781 25651 11815
rect 27154 11812 27160 11824
rect 27115 11784 27160 11812
rect 25593 11775 25651 11781
rect 27154 11772 27160 11784
rect 27212 11772 27218 11824
rect 24581 11747 24639 11753
rect 24581 11713 24593 11747
rect 24627 11744 24639 11747
rect 24670 11744 24676 11756
rect 24627 11716 24676 11744
rect 24627 11713 24639 11716
rect 24581 11707 24639 11713
rect 24670 11704 24676 11716
rect 24728 11704 24734 11756
rect 25961 11747 26019 11753
rect 25961 11744 25973 11747
rect 25332 11716 25973 11744
rect 19668 11611 19732 11617
rect 19668 11577 19686 11611
rect 19720 11577 19732 11611
rect 19668 11571 19732 11577
rect 23109 11611 23167 11617
rect 23109 11577 23121 11611
rect 23155 11608 23167 11611
rect 24489 11611 24547 11617
rect 24489 11608 24501 11611
rect 23155 11580 24501 11608
rect 23155 11577 23167 11580
rect 23109 11571 23167 11577
rect 24489 11577 24501 11580
rect 24535 11577 24547 11611
rect 24489 11571 24547 11577
rect 19668 11568 19674 11571
rect 6457 11543 6515 11549
rect 6457 11540 6469 11543
rect 6328 11512 6469 11540
rect 6328 11500 6334 11512
rect 6457 11509 6469 11512
rect 6503 11509 6515 11543
rect 6457 11503 6515 11509
rect 7469 11543 7527 11549
rect 7469 11509 7481 11543
rect 7515 11540 7527 11543
rect 7558 11540 7564 11552
rect 7515 11512 7564 11540
rect 7515 11509 7527 11512
rect 7469 11503 7527 11509
rect 7558 11500 7564 11512
rect 7616 11500 7622 11552
rect 8294 11500 8300 11552
rect 8352 11540 8358 11552
rect 8665 11543 8723 11549
rect 8665 11540 8677 11543
rect 8352 11512 8677 11540
rect 8352 11500 8358 11512
rect 8665 11509 8677 11512
rect 8711 11540 8723 11543
rect 8938 11540 8944 11552
rect 8711 11512 8944 11540
rect 8711 11509 8723 11512
rect 8665 11503 8723 11509
rect 8938 11500 8944 11512
rect 8996 11500 9002 11552
rect 9122 11540 9128 11552
rect 9083 11512 9128 11540
rect 9122 11500 9128 11512
rect 9180 11500 9186 11552
rect 11885 11543 11943 11549
rect 11885 11509 11897 11543
rect 11931 11540 11943 11543
rect 12250 11540 12256 11552
rect 11931 11512 12256 11540
rect 11931 11509 11943 11512
rect 11885 11503 11943 11509
rect 12250 11500 12256 11512
rect 12308 11500 12314 11552
rect 12618 11500 12624 11552
rect 12676 11540 12682 11552
rect 12713 11543 12771 11549
rect 12713 11540 12725 11543
rect 12676 11512 12725 11540
rect 12676 11500 12682 11512
rect 12713 11509 12725 11512
rect 12759 11540 12771 11543
rect 13449 11543 13507 11549
rect 13449 11540 13461 11543
rect 12759 11512 13461 11540
rect 12759 11509 12771 11512
rect 12713 11503 12771 11509
rect 13449 11509 13461 11512
rect 13495 11509 13507 11543
rect 15930 11540 15936 11552
rect 15891 11512 15936 11540
rect 13449 11503 13507 11509
rect 15930 11500 15936 11512
rect 15988 11500 15994 11552
rect 16206 11500 16212 11552
rect 16264 11540 16270 11552
rect 16301 11543 16359 11549
rect 16301 11540 16313 11543
rect 16264 11512 16313 11540
rect 16264 11500 16270 11512
rect 16301 11509 16313 11512
rect 16347 11540 16359 11543
rect 16945 11543 17003 11549
rect 16945 11540 16957 11543
rect 16347 11512 16957 11540
rect 16347 11509 16359 11512
rect 16301 11503 16359 11509
rect 16945 11509 16957 11512
rect 16991 11540 17003 11543
rect 17126 11540 17132 11552
rect 16991 11512 17132 11540
rect 16991 11509 17003 11512
rect 16945 11503 17003 11509
rect 17126 11500 17132 11512
rect 17184 11500 17190 11552
rect 17862 11540 17868 11552
rect 17823 11512 17868 11540
rect 17862 11500 17868 11512
rect 17920 11500 17926 11552
rect 20806 11540 20812 11552
rect 20767 11512 20812 11540
rect 20806 11500 20812 11512
rect 20864 11500 20870 11552
rect 21358 11540 21364 11552
rect 21319 11512 21364 11540
rect 21358 11500 21364 11512
rect 21416 11500 21422 11552
rect 21726 11540 21732 11552
rect 21687 11512 21732 11540
rect 21726 11500 21732 11512
rect 21784 11500 21790 11552
rect 21818 11500 21824 11552
rect 21876 11540 21882 11552
rect 22097 11543 22155 11549
rect 22097 11540 22109 11543
rect 21876 11512 22109 11540
rect 21876 11500 21882 11512
rect 22097 11509 22109 11512
rect 22143 11509 22155 11543
rect 22097 11503 22155 11509
rect 22741 11543 22799 11549
rect 22741 11509 22753 11543
rect 22787 11540 22799 11543
rect 23290 11540 23296 11552
rect 22787 11512 23296 11540
rect 22787 11509 22799 11512
rect 22741 11503 22799 11509
rect 23290 11500 23296 11512
rect 23348 11500 23354 11552
rect 23477 11543 23535 11549
rect 23477 11509 23489 11543
rect 23523 11540 23535 11543
rect 23566 11540 23572 11552
rect 23523 11512 23572 11540
rect 23523 11509 23535 11512
rect 23477 11503 23535 11509
rect 23566 11500 23572 11512
rect 23624 11500 23630 11552
rect 24394 11500 24400 11552
rect 24452 11540 24458 11552
rect 25332 11549 25360 11716
rect 25961 11713 25973 11716
rect 26007 11744 26019 11747
rect 27246 11744 27252 11756
rect 26007 11716 27252 11744
rect 26007 11713 26019 11716
rect 25961 11707 26019 11713
rect 27246 11704 27252 11716
rect 27304 11704 27310 11756
rect 27724 11753 27752 11852
rect 29546 11840 29552 11852
rect 29604 11840 29610 11892
rect 31938 11880 31944 11892
rect 31899 11852 31944 11880
rect 31938 11840 31944 11852
rect 31996 11840 32002 11892
rect 33318 11880 33324 11892
rect 33279 11852 33324 11880
rect 33318 11840 33324 11852
rect 33376 11840 33382 11892
rect 34333 11883 34391 11889
rect 34333 11880 34345 11883
rect 33428 11852 34345 11880
rect 30374 11772 30380 11824
rect 30432 11812 30438 11824
rect 30561 11815 30619 11821
rect 30561 11812 30573 11815
rect 30432 11784 30573 11812
rect 30432 11772 30438 11784
rect 30561 11781 30573 11784
rect 30607 11781 30619 11815
rect 30561 11775 30619 11781
rect 32858 11772 32864 11824
rect 32916 11812 32922 11824
rect 33428 11812 33456 11852
rect 34333 11849 34345 11852
rect 34379 11880 34391 11883
rect 34606 11880 34612 11892
rect 34379 11852 34612 11880
rect 34379 11849 34391 11852
rect 34333 11843 34391 11849
rect 34606 11840 34612 11852
rect 34664 11840 34670 11892
rect 36262 11880 36268 11892
rect 36223 11852 36268 11880
rect 36262 11840 36268 11852
rect 36320 11840 36326 11892
rect 32916 11784 33456 11812
rect 32916 11772 32922 11784
rect 34146 11772 34152 11824
rect 34204 11812 34210 11824
rect 34977 11815 35035 11821
rect 34977 11812 34989 11815
rect 34204 11784 34989 11812
rect 34204 11772 34210 11784
rect 34977 11781 34989 11784
rect 35023 11781 35035 11815
rect 34977 11775 35035 11781
rect 27709 11747 27767 11753
rect 27709 11713 27721 11747
rect 27755 11713 27767 11747
rect 33778 11744 33784 11756
rect 33739 11716 33784 11744
rect 27709 11707 27767 11713
rect 33778 11704 33784 11716
rect 33836 11704 33842 11756
rect 37550 11744 37556 11756
rect 37511 11716 37556 11744
rect 37550 11704 37556 11716
rect 37608 11704 37614 11756
rect 29362 11676 29368 11688
rect 29323 11648 29368 11676
rect 29362 11636 29368 11648
rect 29420 11676 29426 11688
rect 29914 11676 29920 11688
rect 29420 11648 29920 11676
rect 29420 11636 29426 11648
rect 29914 11636 29920 11648
rect 29972 11636 29978 11688
rect 30190 11636 30196 11688
rect 30248 11676 30254 11688
rect 30837 11679 30895 11685
rect 30837 11676 30849 11679
rect 30248 11648 30849 11676
rect 30248 11636 30254 11648
rect 30837 11645 30849 11648
rect 30883 11645 30895 11679
rect 31662 11676 31668 11688
rect 30837 11639 30895 11645
rect 31036 11648 31668 11676
rect 31036 11620 31064 11648
rect 31662 11636 31668 11648
rect 31720 11636 31726 11688
rect 31938 11636 31944 11688
rect 31996 11676 32002 11688
rect 32125 11679 32183 11685
rect 32125 11676 32137 11679
rect 31996 11648 32137 11676
rect 31996 11636 32002 11648
rect 32125 11645 32137 11648
rect 32171 11645 32183 11679
rect 33870 11676 33876 11688
rect 33783 11648 33876 11676
rect 32125 11639 32183 11645
rect 33870 11636 33876 11648
rect 33928 11676 33934 11688
rect 33928 11648 35572 11676
rect 33928 11636 33934 11648
rect 25866 11568 25872 11620
rect 25924 11608 25930 11620
rect 26145 11611 26203 11617
rect 26145 11608 26157 11611
rect 25924 11580 26157 11608
rect 25924 11568 25930 11580
rect 26145 11577 26157 11580
rect 26191 11577 26203 11611
rect 27430 11608 27436 11620
rect 27391 11580 27436 11608
rect 26145 11571 26203 11577
rect 27430 11568 27436 11580
rect 27488 11568 27494 11620
rect 31018 11608 31024 11620
rect 30979 11580 31024 11608
rect 31018 11568 31024 11580
rect 31076 11568 31082 11620
rect 31113 11611 31171 11617
rect 31113 11577 31125 11611
rect 31159 11577 31171 11611
rect 34606 11608 34612 11620
rect 34567 11580 34612 11608
rect 31113 11571 31171 11577
rect 25317 11543 25375 11549
rect 25317 11540 25329 11543
rect 24452 11512 25329 11540
rect 24452 11500 24458 11512
rect 25317 11509 25329 11512
rect 25363 11509 25375 11543
rect 25317 11503 25375 11509
rect 25958 11500 25964 11552
rect 26016 11540 26022 11552
rect 26053 11543 26111 11549
rect 26053 11540 26065 11543
rect 26016 11512 26065 11540
rect 26016 11500 26022 11512
rect 26053 11509 26065 11512
rect 26099 11509 26111 11543
rect 26053 11503 26111 11509
rect 26973 11543 27031 11549
rect 26973 11509 26985 11543
rect 27019 11540 27031 11543
rect 27617 11543 27675 11549
rect 27617 11540 27629 11543
rect 27019 11512 27629 11540
rect 27019 11509 27031 11512
rect 26973 11503 27031 11509
rect 27617 11509 27629 11512
rect 27663 11540 27675 11543
rect 28258 11540 28264 11552
rect 27663 11512 28264 11540
rect 27663 11509 27675 11512
rect 27617 11503 27675 11509
rect 28258 11500 28264 11512
rect 28316 11500 28322 11552
rect 30377 11543 30435 11549
rect 30377 11509 30389 11543
rect 30423 11540 30435 11543
rect 31128 11540 31156 11571
rect 34606 11568 34612 11580
rect 34664 11608 34670 11620
rect 35544 11617 35572 11648
rect 35986 11636 35992 11688
rect 36044 11676 36050 11688
rect 36449 11679 36507 11685
rect 36449 11676 36461 11679
rect 36044 11648 36461 11676
rect 36044 11636 36050 11648
rect 36449 11645 36461 11648
rect 36495 11676 36507 11679
rect 37001 11679 37059 11685
rect 37001 11676 37013 11679
rect 36495 11648 37013 11676
rect 36495 11645 36507 11648
rect 36449 11639 36507 11645
rect 37001 11645 37013 11648
rect 37047 11645 37059 11679
rect 37001 11639 37059 11645
rect 35253 11611 35311 11617
rect 35253 11608 35265 11611
rect 34664 11580 35265 11608
rect 34664 11568 34670 11580
rect 35253 11577 35265 11580
rect 35299 11577 35311 11611
rect 35253 11571 35311 11577
rect 35529 11611 35587 11617
rect 35529 11577 35541 11611
rect 35575 11577 35587 11611
rect 35529 11571 35587 11577
rect 31202 11540 31208 11552
rect 30423 11512 31208 11540
rect 30423 11509 30435 11512
rect 30377 11503 30435 11509
rect 31202 11500 31208 11512
rect 31260 11500 31266 11552
rect 31294 11500 31300 11552
rect 31352 11540 31358 11552
rect 31481 11543 31539 11549
rect 31481 11540 31493 11543
rect 31352 11512 31493 11540
rect 31352 11500 31358 11512
rect 31481 11509 31493 11512
rect 31527 11509 31539 11543
rect 32306 11540 32312 11552
rect 32267 11512 32312 11540
rect 31481 11503 31539 11509
rect 32306 11500 32312 11512
rect 32364 11500 32370 11552
rect 32769 11543 32827 11549
rect 32769 11509 32781 11543
rect 32815 11540 32827 11543
rect 32950 11540 32956 11552
rect 32815 11512 32956 11540
rect 32815 11509 32827 11512
rect 32769 11503 32827 11509
rect 32950 11500 32956 11512
rect 33008 11500 33014 11552
rect 33134 11540 33140 11552
rect 33047 11512 33140 11540
rect 33134 11500 33140 11512
rect 33192 11540 33198 11552
rect 33778 11540 33784 11552
rect 33192 11512 33784 11540
rect 33192 11500 33198 11512
rect 33778 11500 33784 11512
rect 33836 11500 33842 11552
rect 34882 11500 34888 11552
rect 34940 11540 34946 11552
rect 35437 11543 35495 11549
rect 35437 11540 35449 11543
rect 34940 11512 35449 11540
rect 34940 11500 34946 11512
rect 35437 11509 35449 11512
rect 35483 11509 35495 11543
rect 35544 11540 35572 11571
rect 35989 11543 36047 11549
rect 35989 11540 36001 11543
rect 35544 11512 36001 11540
rect 35437 11503 35495 11509
rect 35989 11509 36001 11512
rect 36035 11540 36047 11543
rect 36078 11540 36084 11552
rect 36035 11512 36084 11540
rect 36035 11509 36047 11512
rect 35989 11503 36047 11509
rect 36078 11500 36084 11512
rect 36136 11500 36142 11552
rect 36633 11543 36691 11549
rect 36633 11509 36645 11543
rect 36679 11540 36691 11543
rect 36814 11540 36820 11552
rect 36679 11512 36820 11540
rect 36679 11509 36691 11512
rect 36633 11503 36691 11509
rect 36814 11500 36820 11512
rect 36872 11500 36878 11552
rect 1104 11450 38824 11472
rect 1104 11398 14315 11450
rect 14367 11398 14379 11450
rect 14431 11398 14443 11450
rect 14495 11398 14507 11450
rect 14559 11398 27648 11450
rect 27700 11398 27712 11450
rect 27764 11398 27776 11450
rect 27828 11398 27840 11450
rect 27892 11398 38824 11450
rect 1104 11376 38824 11398
rect 2041 11339 2099 11345
rect 2041 11305 2053 11339
rect 2087 11336 2099 11339
rect 2406 11336 2412 11348
rect 2087 11308 2412 11336
rect 2087 11305 2099 11308
rect 2041 11299 2099 11305
rect 2406 11296 2412 11308
rect 2464 11296 2470 11348
rect 4154 11296 4160 11348
rect 4212 11336 4218 11348
rect 5445 11339 5503 11345
rect 5445 11336 5457 11339
rect 4212 11308 5457 11336
rect 4212 11296 4218 11308
rect 5445 11305 5457 11308
rect 5491 11336 5503 11339
rect 5534 11336 5540 11348
rect 5491 11308 5540 11336
rect 5491 11305 5503 11308
rect 5445 11299 5503 11305
rect 5534 11296 5540 11308
rect 5592 11296 5598 11348
rect 8297 11339 8355 11345
rect 8297 11305 8309 11339
rect 8343 11336 8355 11339
rect 8386 11336 8392 11348
rect 8343 11308 8392 11336
rect 8343 11305 8355 11308
rect 8297 11299 8355 11305
rect 8386 11296 8392 11308
rect 8444 11296 8450 11348
rect 15102 11296 15108 11348
rect 15160 11336 15166 11348
rect 15841 11339 15899 11345
rect 15841 11336 15853 11339
rect 15160 11308 15853 11336
rect 15160 11296 15166 11308
rect 15841 11305 15853 11308
rect 15887 11336 15899 11339
rect 16022 11336 16028 11348
rect 15887 11308 16028 11336
rect 15887 11305 15899 11308
rect 15841 11299 15899 11305
rect 16022 11296 16028 11308
rect 16080 11296 16086 11348
rect 16485 11339 16543 11345
rect 16485 11305 16497 11339
rect 16531 11336 16543 11339
rect 16942 11336 16948 11348
rect 16531 11308 16948 11336
rect 16531 11305 16543 11308
rect 16485 11299 16543 11305
rect 16942 11296 16948 11308
rect 17000 11296 17006 11348
rect 17402 11336 17408 11348
rect 17363 11308 17408 11336
rect 17402 11296 17408 11308
rect 17460 11296 17466 11348
rect 17494 11296 17500 11348
rect 17552 11336 17558 11348
rect 22922 11336 22928 11348
rect 17552 11308 19104 11336
rect 22883 11308 22928 11336
rect 17552 11296 17558 11308
rect 19076 11280 19104 11308
rect 22922 11296 22928 11308
rect 22980 11296 22986 11348
rect 23290 11296 23296 11348
rect 23348 11336 23354 11348
rect 23842 11336 23848 11348
rect 23348 11308 23848 11336
rect 23348 11296 23354 11308
rect 23842 11296 23848 11308
rect 23900 11336 23906 11348
rect 23937 11339 23995 11345
rect 23937 11336 23949 11339
rect 23900 11308 23949 11336
rect 23900 11296 23906 11308
rect 23937 11305 23949 11308
rect 23983 11305 23995 11339
rect 23937 11299 23995 11305
rect 2961 11271 3019 11277
rect 2961 11237 2973 11271
rect 3007 11268 3019 11271
rect 3418 11268 3424 11280
rect 3007 11240 3424 11268
rect 3007 11237 3019 11240
rect 2961 11231 3019 11237
rect 3418 11228 3424 11240
rect 3476 11228 3482 11280
rect 7098 11268 7104 11280
rect 7059 11240 7104 11268
rect 7098 11228 7104 11240
rect 7156 11228 7162 11280
rect 9950 11277 9956 11280
rect 9944 11268 9956 11277
rect 9911 11240 9956 11268
rect 9944 11231 9956 11240
rect 9950 11228 9956 11231
rect 10008 11228 10014 11280
rect 12434 11228 12440 11280
rect 12492 11268 12498 11280
rect 12989 11271 13047 11277
rect 12989 11268 13001 11271
rect 12492 11240 13001 11268
rect 12492 11228 12498 11240
rect 12989 11237 13001 11240
rect 13035 11268 13047 11271
rect 13449 11271 13507 11277
rect 13449 11268 13461 11271
rect 13035 11240 13461 11268
rect 13035 11237 13047 11240
rect 12989 11231 13047 11237
rect 13449 11237 13461 11240
rect 13495 11237 13507 11271
rect 13449 11231 13507 11237
rect 15930 11228 15936 11280
rect 15988 11268 15994 11280
rect 17221 11271 17279 11277
rect 17221 11268 17233 11271
rect 15988 11240 17233 11268
rect 15988 11228 15994 11240
rect 17221 11237 17233 11240
rect 17267 11268 17279 11271
rect 18491 11271 18549 11277
rect 18491 11268 18503 11271
rect 17267 11240 18503 11268
rect 17267 11237 17279 11240
rect 17221 11231 17279 11237
rect 18491 11237 18503 11240
rect 18537 11237 18549 11271
rect 18491 11231 18549 11237
rect 18969 11271 19027 11277
rect 18969 11237 18981 11271
rect 19015 11237 19027 11271
rect 18969 11231 19027 11237
rect 3694 11160 3700 11212
rect 3752 11200 3758 11212
rect 4065 11203 4123 11209
rect 4065 11200 4077 11203
rect 3752 11172 4077 11200
rect 3752 11160 3758 11172
rect 4065 11169 4077 11172
rect 4111 11169 4123 11203
rect 4065 11163 4123 11169
rect 4154 11160 4160 11212
rect 4212 11200 4218 11212
rect 4321 11203 4379 11209
rect 4321 11200 4333 11203
rect 4212 11172 4333 11200
rect 4212 11160 4218 11172
rect 4321 11169 4333 11172
rect 4367 11200 4379 11203
rect 5626 11200 5632 11212
rect 4367 11172 5632 11200
rect 4367 11169 4379 11172
rect 4321 11163 4379 11169
rect 5626 11160 5632 11172
rect 5684 11160 5690 11212
rect 5810 11160 5816 11212
rect 5868 11200 5874 11212
rect 6089 11203 6147 11209
rect 6089 11200 6101 11203
rect 5868 11172 6101 11200
rect 5868 11160 5874 11172
rect 6089 11169 6101 11172
rect 6135 11200 6147 11203
rect 6457 11203 6515 11209
rect 6457 11200 6469 11203
rect 6135 11172 6469 11200
rect 6135 11169 6147 11172
rect 6089 11163 6147 11169
rect 6457 11169 6469 11172
rect 6503 11200 6515 11203
rect 8113 11203 8171 11209
rect 6503 11172 7236 11200
rect 6503 11169 6515 11172
rect 6457 11163 6515 11169
rect 1394 11132 1400 11144
rect 1355 11104 1400 11132
rect 1394 11092 1400 11104
rect 1452 11092 1458 11144
rect 2958 11132 2964 11144
rect 2919 11104 2964 11132
rect 2958 11092 2964 11104
rect 3016 11092 3022 11144
rect 3053 11135 3111 11141
rect 3053 11101 3065 11135
rect 3099 11132 3111 11135
rect 3970 11132 3976 11144
rect 3099 11104 3976 11132
rect 3099 11101 3111 11104
rect 3053 11095 3111 11101
rect 3970 11092 3976 11104
rect 4028 11092 4034 11144
rect 7208 11141 7236 11172
rect 8113 11169 8125 11203
rect 8159 11200 8171 11203
rect 8386 11200 8392 11212
rect 8159 11172 8392 11200
rect 8159 11169 8171 11172
rect 8113 11163 8171 11169
rect 8386 11160 8392 11172
rect 8444 11160 8450 11212
rect 10686 11160 10692 11212
rect 10744 11200 10750 11212
rect 11882 11200 11888 11212
rect 10744 11172 11888 11200
rect 10744 11160 10750 11172
rect 11882 11160 11888 11172
rect 11940 11200 11946 11212
rect 11977 11203 12035 11209
rect 11977 11200 11989 11203
rect 11940 11172 11989 11200
rect 11940 11160 11946 11172
rect 11977 11169 11989 11172
rect 12023 11169 12035 11203
rect 12802 11200 12808 11212
rect 12763 11172 12808 11200
rect 11977 11163 12035 11169
rect 12802 11160 12808 11172
rect 12860 11200 12866 11212
rect 13817 11203 13875 11209
rect 13817 11200 13829 11203
rect 12860 11172 13829 11200
rect 12860 11160 12866 11172
rect 13817 11169 13829 11172
rect 13863 11169 13875 11203
rect 18782 11200 18788 11212
rect 13817 11163 13875 11169
rect 15396 11172 18788 11200
rect 7009 11135 7067 11141
rect 7009 11132 7021 11135
rect 6932 11104 7021 11132
rect 2498 11064 2504 11076
rect 2459 11036 2504 11064
rect 2498 11024 2504 11036
rect 2556 11024 2562 11076
rect 2682 11024 2688 11076
rect 2740 11024 2746 11076
rect 3602 11064 3608 11076
rect 3563 11036 3608 11064
rect 3602 11024 3608 11036
rect 3660 11024 3666 11076
rect 5350 11024 5356 11076
rect 5408 11064 5414 11076
rect 6641 11067 6699 11073
rect 6641 11064 6653 11067
rect 5408 11036 6653 11064
rect 5408 11024 5414 11036
rect 6641 11033 6653 11036
rect 6687 11033 6699 11067
rect 6641 11027 6699 11033
rect 2700 10996 2728 11024
rect 3142 10996 3148 11008
rect 2700 10968 3148 10996
rect 3142 10956 3148 10968
rect 3200 10996 3206 11008
rect 4338 10996 4344 11008
rect 3200 10968 4344 10996
rect 3200 10956 3206 10968
rect 4338 10956 4344 10968
rect 4396 10956 4402 11008
rect 6822 10956 6828 11008
rect 6880 10996 6886 11008
rect 6932 10996 6960 11104
rect 7009 11101 7021 11104
rect 7055 11101 7067 11135
rect 7009 11095 7067 11101
rect 7193 11135 7251 11141
rect 7193 11101 7205 11135
rect 7239 11101 7251 11135
rect 7193 11095 7251 11101
rect 7208 11064 7236 11095
rect 8294 11092 8300 11144
rect 8352 11132 8358 11144
rect 8662 11132 8668 11144
rect 8352 11104 8668 11132
rect 8352 11092 8358 11104
rect 8662 11092 8668 11104
rect 8720 11132 8726 11144
rect 8757 11135 8815 11141
rect 8757 11132 8769 11135
rect 8720 11104 8769 11132
rect 8720 11092 8726 11104
rect 8757 11101 8769 11104
rect 8803 11132 8815 11135
rect 9674 11132 9680 11144
rect 8803 11104 9680 11132
rect 8803 11101 8815 11104
rect 8757 11095 8815 11101
rect 9674 11092 9680 11104
rect 9732 11092 9738 11144
rect 11698 11132 11704 11144
rect 11659 11104 11704 11132
rect 11698 11092 11704 11104
rect 11756 11092 11762 11144
rect 13078 11132 13084 11144
rect 13039 11104 13084 11132
rect 13078 11092 13084 11104
rect 13136 11132 13142 11144
rect 15013 11135 15071 11141
rect 15013 11132 15025 11135
rect 13136 11104 15025 11132
rect 13136 11092 13142 11104
rect 15013 11101 15025 11104
rect 15059 11101 15071 11135
rect 15013 11095 15071 11101
rect 8021 11067 8079 11073
rect 8021 11064 8033 11067
rect 7208 11036 8033 11064
rect 8021 11033 8033 11036
rect 8067 11064 8079 11067
rect 11057 11067 11115 11073
rect 8067 11036 9168 11064
rect 8067 11033 8079 11036
rect 8021 11027 8079 11033
rect 9140 11008 9168 11036
rect 11057 11033 11069 11067
rect 11103 11064 11115 11067
rect 11146 11064 11152 11076
rect 11103 11036 11152 11064
rect 11103 11033 11115 11036
rect 11057 11027 11115 11033
rect 11146 11024 11152 11036
rect 11204 11024 11210 11076
rect 12526 11064 12532 11076
rect 12487 11036 12532 11064
rect 12526 11024 12532 11036
rect 12584 11024 12590 11076
rect 15396 11073 15424 11172
rect 18782 11160 18788 11172
rect 18840 11200 18846 11212
rect 18984 11200 19012 11231
rect 19058 11228 19064 11280
rect 19116 11268 19122 11280
rect 19116 11240 19209 11268
rect 19116 11228 19122 11240
rect 20806 11228 20812 11280
rect 20864 11268 20870 11280
rect 21146 11271 21204 11277
rect 21146 11268 21158 11271
rect 20864 11240 21158 11268
rect 20864 11228 20870 11240
rect 21146 11237 21158 11240
rect 21192 11237 21204 11271
rect 21146 11231 21204 11237
rect 21634 11228 21640 11280
rect 21692 11268 21698 11280
rect 24394 11268 24400 11280
rect 21692 11240 24400 11268
rect 21692 11228 21698 11240
rect 24394 11228 24400 11240
rect 24452 11228 24458 11280
rect 24578 11228 24584 11280
rect 24636 11268 24642 11280
rect 25225 11271 25283 11277
rect 25225 11268 25237 11271
rect 24636 11240 25237 11268
rect 24636 11228 24642 11240
rect 25225 11237 25237 11240
rect 25271 11237 25283 11271
rect 25225 11231 25283 11237
rect 26326 11228 26332 11280
rect 26384 11268 26390 11280
rect 27065 11271 27123 11277
rect 27065 11268 27077 11271
rect 26384 11240 27077 11268
rect 26384 11228 26390 11240
rect 27065 11237 27077 11240
rect 27111 11268 27123 11271
rect 27154 11268 27160 11280
rect 27111 11240 27160 11268
rect 27111 11237 27123 11240
rect 27065 11231 27123 11237
rect 27154 11228 27160 11240
rect 27212 11228 27218 11280
rect 30926 11268 30932 11280
rect 30887 11240 30932 11268
rect 30926 11228 30932 11240
rect 30984 11228 30990 11280
rect 32674 11228 32680 11280
rect 32732 11268 32738 11280
rect 32861 11271 32919 11277
rect 32861 11268 32873 11271
rect 32732 11240 32873 11268
rect 32732 11228 32738 11240
rect 32861 11237 32873 11240
rect 32907 11268 32919 11271
rect 33220 11271 33278 11277
rect 33220 11268 33232 11271
rect 32907 11240 33232 11268
rect 32907 11237 32919 11240
rect 32861 11231 32919 11237
rect 33220 11237 33232 11240
rect 33266 11268 33278 11271
rect 33870 11268 33876 11280
rect 33266 11240 33876 11268
rect 33266 11237 33278 11240
rect 33220 11231 33278 11237
rect 33870 11228 33876 11240
rect 33928 11228 33934 11280
rect 35710 11228 35716 11280
rect 35768 11268 35774 11280
rect 35805 11271 35863 11277
rect 35805 11268 35817 11271
rect 35768 11240 35817 11268
rect 35768 11228 35774 11240
rect 35805 11237 35817 11240
rect 35851 11237 35863 11271
rect 35805 11231 35863 11237
rect 35989 11271 36047 11277
rect 35989 11237 36001 11271
rect 36035 11268 36047 11271
rect 36354 11268 36360 11280
rect 36035 11240 36360 11268
rect 36035 11237 36047 11240
rect 35989 11231 36047 11237
rect 36354 11228 36360 11240
rect 36412 11228 36418 11280
rect 18840 11172 19012 11200
rect 18840 11160 18846 11172
rect 20714 11160 20720 11212
rect 20772 11200 20778 11212
rect 20898 11200 20904 11212
rect 20772 11172 20904 11200
rect 20772 11160 20778 11172
rect 20898 11160 20904 11172
rect 20956 11160 20962 11212
rect 23750 11200 23756 11212
rect 23711 11172 23756 11200
rect 23750 11160 23756 11172
rect 23808 11160 23814 11212
rect 24854 11160 24860 11212
rect 24912 11200 24918 11212
rect 24949 11203 25007 11209
rect 24949 11200 24961 11203
rect 24912 11172 24961 11200
rect 24912 11160 24918 11172
rect 24949 11169 24961 11172
rect 24995 11169 25007 11203
rect 26234 11200 26240 11212
rect 26195 11172 26240 11200
rect 24949 11163 25007 11169
rect 26234 11160 26240 11172
rect 26292 11200 26298 11212
rect 28442 11209 28448 11212
rect 26881 11203 26939 11209
rect 26881 11200 26893 11203
rect 26292 11172 26893 11200
rect 26292 11160 26298 11172
rect 26881 11169 26893 11172
rect 26927 11169 26939 11203
rect 28436 11200 28448 11209
rect 28403 11172 28448 11200
rect 26881 11163 26939 11169
rect 28436 11163 28448 11172
rect 28442 11160 28448 11163
rect 28500 11160 28506 11212
rect 30374 11160 30380 11212
rect 30432 11200 30438 11212
rect 30653 11203 30711 11209
rect 30653 11200 30665 11203
rect 30432 11172 30665 11200
rect 30432 11160 30438 11172
rect 30653 11169 30665 11172
rect 30699 11169 30711 11203
rect 30653 11163 30711 11169
rect 31941 11203 31999 11209
rect 31941 11169 31953 11203
rect 31987 11200 31999 11203
rect 33042 11200 33048 11212
rect 31987 11172 33048 11200
rect 31987 11169 31999 11172
rect 31941 11163 31999 11169
rect 33042 11160 33048 11172
rect 33100 11160 33106 11212
rect 35345 11203 35403 11209
rect 35345 11169 35357 11203
rect 35391 11200 35403 11203
rect 35391 11172 36124 11200
rect 35391 11169 35403 11172
rect 35345 11163 35403 11169
rect 36096 11144 36124 11172
rect 15746 11132 15752 11144
rect 15488 11104 15752 11132
rect 15381 11067 15439 11073
rect 15381 11033 15393 11067
rect 15427 11033 15439 11067
rect 15381 11027 15439 11033
rect 9122 10996 9128 11008
rect 6880 10968 6960 10996
rect 9035 10968 9128 10996
rect 6880 10956 6886 10968
rect 9122 10956 9128 10968
rect 9180 10996 9186 11008
rect 9582 10996 9588 11008
rect 9180 10968 9588 10996
rect 9180 10956 9186 10968
rect 9582 10956 9588 10968
rect 9640 10956 9646 11008
rect 15010 10956 15016 11008
rect 15068 10996 15074 11008
rect 15488 10996 15516 11104
rect 15746 11092 15752 11104
rect 15804 11092 15810 11144
rect 15838 11092 15844 11144
rect 15896 11132 15902 11144
rect 15933 11135 15991 11141
rect 15933 11132 15945 11135
rect 15896 11104 15945 11132
rect 15896 11092 15902 11104
rect 15933 11101 15945 11104
rect 15979 11101 15991 11135
rect 15933 11095 15991 11101
rect 17126 11092 17132 11144
rect 17184 11132 17190 11144
rect 17497 11135 17555 11141
rect 17497 11132 17509 11135
rect 17184 11104 17509 11132
rect 17184 11092 17190 11104
rect 17497 11101 17509 11104
rect 17543 11101 17555 11135
rect 17497 11095 17555 11101
rect 17678 11092 17684 11144
rect 17736 11132 17742 11144
rect 18049 11135 18107 11141
rect 18049 11132 18061 11135
rect 17736 11104 18061 11132
rect 17736 11092 17742 11104
rect 18049 11101 18061 11104
rect 18095 11132 18107 11135
rect 18230 11132 18236 11144
rect 18095 11104 18236 11132
rect 18095 11101 18107 11104
rect 18049 11095 18107 11101
rect 18230 11092 18236 11104
rect 18288 11092 18294 11144
rect 18874 11132 18880 11144
rect 18835 11104 18880 11132
rect 18874 11092 18880 11104
rect 18932 11092 18938 11144
rect 24026 11132 24032 11144
rect 23987 11104 24032 11132
rect 24026 11092 24032 11104
rect 24084 11092 24090 11144
rect 26694 11092 26700 11144
rect 26752 11132 26758 11144
rect 27157 11135 27215 11141
rect 27157 11132 27169 11135
rect 26752 11104 27169 11132
rect 26752 11092 26758 11104
rect 27157 11101 27169 11104
rect 27203 11101 27215 11135
rect 28166 11132 28172 11144
rect 28127 11104 28172 11132
rect 27157 11095 27215 11101
rect 28166 11092 28172 11104
rect 28224 11092 28230 11144
rect 32858 11092 32864 11144
rect 32916 11132 32922 11144
rect 32953 11135 33011 11141
rect 32953 11132 32965 11135
rect 32916 11104 32965 11132
rect 32916 11092 32922 11104
rect 32953 11101 32965 11104
rect 32999 11101 33011 11135
rect 36078 11132 36084 11144
rect 36039 11104 36084 11132
rect 32953 11095 33011 11101
rect 36078 11092 36084 11104
rect 36136 11092 36142 11144
rect 16850 11024 16856 11076
rect 16908 11064 16914 11076
rect 16945 11067 17003 11073
rect 16945 11064 16957 11067
rect 16908 11036 16957 11064
rect 16908 11024 16914 11036
rect 16945 11033 16957 11036
rect 16991 11033 17003 11067
rect 18248 11064 18276 11092
rect 19610 11064 19616 11076
rect 18248 11036 19616 11064
rect 16945 11027 17003 11033
rect 19610 11024 19616 11036
rect 19668 11024 19674 11076
rect 22278 11064 22284 11076
rect 22239 11036 22284 11064
rect 22278 11024 22284 11036
rect 22336 11024 22342 11076
rect 23293 11067 23351 11073
rect 23293 11033 23305 11067
rect 23339 11033 23351 11067
rect 23474 11064 23480 11076
rect 23435 11036 23480 11064
rect 23293 11027 23351 11033
rect 15068 10968 15516 10996
rect 23308 10996 23336 11027
rect 23474 11024 23480 11036
rect 23532 11024 23538 11076
rect 24489 11067 24547 11073
rect 24489 11033 24501 11067
rect 24535 11064 24547 11067
rect 24946 11064 24952 11076
rect 24535 11036 24952 11064
rect 24535 11033 24547 11036
rect 24489 11027 24547 11033
rect 24946 11024 24952 11036
rect 25004 11064 25010 11076
rect 25314 11064 25320 11076
rect 25004 11036 25320 11064
rect 25004 11024 25010 11036
rect 25314 11024 25320 11036
rect 25372 11024 25378 11076
rect 26602 11064 26608 11076
rect 26563 11036 26608 11064
rect 26602 11024 26608 11036
rect 26660 11024 26666 11076
rect 29546 11064 29552 11076
rect 29507 11036 29552 11064
rect 29546 11024 29552 11036
rect 29604 11024 29610 11076
rect 32493 11067 32551 11073
rect 32493 11033 32505 11067
rect 32539 11064 32551 11067
rect 32539 11036 32996 11064
rect 32539 11033 32551 11036
rect 32493 11027 32551 11033
rect 24302 10996 24308 11008
rect 23308 10968 24308 10996
rect 15068 10956 15074 10968
rect 24302 10956 24308 10968
rect 24360 10956 24366 11008
rect 24857 10999 24915 11005
rect 24857 10965 24869 10999
rect 24903 10996 24915 10999
rect 25038 10996 25044 11008
rect 24903 10968 25044 10996
rect 24903 10965 24915 10968
rect 24857 10959 24915 10965
rect 25038 10956 25044 10968
rect 25096 10996 25102 11008
rect 25685 10999 25743 11005
rect 25685 10996 25697 10999
rect 25096 10968 25697 10996
rect 25096 10956 25102 10968
rect 25685 10965 25697 10968
rect 25731 10996 25743 10999
rect 25866 10996 25872 11008
rect 25731 10968 25872 10996
rect 25731 10965 25743 10968
rect 25685 10959 25743 10965
rect 25866 10956 25872 10968
rect 25924 10956 25930 11008
rect 30377 10999 30435 11005
rect 30377 10965 30389 10999
rect 30423 10996 30435 10999
rect 30834 10996 30840 11008
rect 30423 10968 30840 10996
rect 30423 10965 30435 10968
rect 30377 10959 30435 10965
rect 30834 10956 30840 10968
rect 30892 10956 30898 11008
rect 32968 10996 32996 11036
rect 34514 11024 34520 11076
rect 34572 11064 34578 11076
rect 34882 11064 34888 11076
rect 34572 11036 34888 11064
rect 34572 11024 34578 11036
rect 34882 11024 34888 11036
rect 34940 11024 34946 11076
rect 35526 11064 35532 11076
rect 35487 11036 35532 11064
rect 35526 11024 35532 11036
rect 35584 11024 35590 11076
rect 36449 11067 36507 11073
rect 36449 11064 36461 11067
rect 35820 11036 36461 11064
rect 33686 10996 33692 11008
rect 32968 10968 33692 10996
rect 33686 10956 33692 10968
rect 33744 10956 33750 11008
rect 33870 10956 33876 11008
rect 33928 10996 33934 11008
rect 34333 10999 34391 11005
rect 34333 10996 34345 10999
rect 33928 10968 34345 10996
rect 33928 10956 33934 10968
rect 34333 10965 34345 10968
rect 34379 10965 34391 10999
rect 34333 10959 34391 10965
rect 35618 10956 35624 11008
rect 35676 10996 35682 11008
rect 35820 10996 35848 11036
rect 36449 11033 36461 11036
rect 36495 11033 36507 11067
rect 36449 11027 36507 11033
rect 35676 10968 35848 10996
rect 35676 10956 35682 10968
rect 1104 10906 38824 10928
rect 1104 10854 7648 10906
rect 7700 10854 7712 10906
rect 7764 10854 7776 10906
rect 7828 10854 7840 10906
rect 7892 10854 20982 10906
rect 21034 10854 21046 10906
rect 21098 10854 21110 10906
rect 21162 10854 21174 10906
rect 21226 10854 34315 10906
rect 34367 10854 34379 10906
rect 34431 10854 34443 10906
rect 34495 10854 34507 10906
rect 34559 10854 38824 10906
rect 1104 10832 38824 10854
rect 1394 10752 1400 10804
rect 1452 10792 1458 10804
rect 1581 10795 1639 10801
rect 1581 10792 1593 10795
rect 1452 10764 1593 10792
rect 1452 10752 1458 10764
rect 1581 10761 1593 10764
rect 1627 10761 1639 10795
rect 3878 10792 3884 10804
rect 3839 10764 3884 10792
rect 1581 10755 1639 10761
rect 1596 10656 1624 10755
rect 3878 10752 3884 10764
rect 3936 10752 3942 10804
rect 5258 10792 5264 10804
rect 5219 10764 5264 10792
rect 5258 10752 5264 10764
rect 5316 10752 5322 10804
rect 5718 10752 5724 10804
rect 5776 10792 5782 10804
rect 6181 10795 6239 10801
rect 6181 10792 6193 10795
rect 5776 10764 6193 10792
rect 5776 10752 5782 10764
rect 6181 10761 6193 10764
rect 6227 10792 6239 10795
rect 6822 10792 6828 10804
rect 6227 10764 6828 10792
rect 6227 10761 6239 10764
rect 6181 10755 6239 10761
rect 6822 10752 6828 10764
rect 6880 10752 6886 10804
rect 6914 10752 6920 10804
rect 6972 10792 6978 10804
rect 7009 10795 7067 10801
rect 7009 10792 7021 10795
rect 6972 10764 7021 10792
rect 6972 10752 6978 10764
rect 7009 10761 7021 10764
rect 7055 10761 7067 10795
rect 8386 10792 8392 10804
rect 7009 10755 7067 10761
rect 8220 10764 8392 10792
rect 2222 10724 2228 10736
rect 2183 10696 2228 10724
rect 2222 10684 2228 10696
rect 2280 10684 2286 10736
rect 3237 10727 3295 10733
rect 3237 10693 3249 10727
rect 3283 10724 3295 10727
rect 4154 10724 4160 10736
rect 3283 10696 4160 10724
rect 3283 10693 3295 10696
rect 3237 10687 3295 10693
rect 4154 10684 4160 10696
rect 4212 10684 4218 10736
rect 7926 10724 7932 10736
rect 4908 10696 7932 10724
rect 2593 10659 2651 10665
rect 2593 10656 2605 10659
rect 1596 10628 2605 10656
rect 2593 10625 2605 10628
rect 2639 10625 2651 10659
rect 4908 10656 4936 10696
rect 7926 10684 7932 10696
rect 7984 10724 7990 10736
rect 8021 10727 8079 10733
rect 8021 10724 8033 10727
rect 7984 10696 8033 10724
rect 7984 10684 7990 10696
rect 8021 10693 8033 10696
rect 8067 10724 8079 10727
rect 8220 10724 8248 10764
rect 8386 10752 8392 10764
rect 8444 10752 8450 10804
rect 9950 10752 9956 10804
rect 10008 10792 10014 10804
rect 10137 10795 10195 10801
rect 10137 10792 10149 10795
rect 10008 10764 10149 10792
rect 10008 10752 10014 10764
rect 10137 10761 10149 10764
rect 10183 10761 10195 10795
rect 10778 10792 10784 10804
rect 10739 10764 10784 10792
rect 10137 10755 10195 10761
rect 10778 10752 10784 10764
rect 10836 10752 10842 10804
rect 14645 10795 14703 10801
rect 14645 10761 14657 10795
rect 14691 10792 14703 10795
rect 15102 10792 15108 10804
rect 14691 10764 15108 10792
rect 14691 10761 14703 10764
rect 14645 10755 14703 10761
rect 15102 10752 15108 10764
rect 15160 10752 15166 10804
rect 17862 10752 17868 10804
rect 17920 10792 17926 10804
rect 18141 10795 18199 10801
rect 18141 10792 18153 10795
rect 17920 10764 18153 10792
rect 17920 10752 17926 10764
rect 18141 10761 18153 10764
rect 18187 10761 18199 10795
rect 19058 10792 19064 10804
rect 19019 10764 19064 10792
rect 18141 10755 18199 10761
rect 19058 10752 19064 10764
rect 19116 10752 19122 10804
rect 19518 10752 19524 10804
rect 19576 10792 19582 10804
rect 19705 10795 19763 10801
rect 19705 10792 19717 10795
rect 19576 10764 19717 10792
rect 19576 10752 19582 10764
rect 19705 10761 19717 10764
rect 19751 10761 19763 10795
rect 19705 10755 19763 10761
rect 20806 10752 20812 10804
rect 20864 10792 20870 10804
rect 21269 10795 21327 10801
rect 21269 10792 21281 10795
rect 20864 10764 21281 10792
rect 20864 10752 20870 10764
rect 21269 10761 21281 10764
rect 21315 10761 21327 10795
rect 23842 10792 23848 10804
rect 23803 10764 23848 10792
rect 21269 10755 21327 10761
rect 23842 10752 23848 10764
rect 23900 10752 23906 10804
rect 25866 10792 25872 10804
rect 25827 10764 25872 10792
rect 25866 10752 25872 10764
rect 25924 10752 25930 10804
rect 27798 10792 27804 10804
rect 27759 10764 27804 10792
rect 27798 10752 27804 10764
rect 27856 10792 27862 10804
rect 28442 10792 28448 10804
rect 27856 10764 28448 10792
rect 27856 10752 27862 10764
rect 28442 10752 28448 10764
rect 28500 10792 28506 10804
rect 28721 10795 28779 10801
rect 28721 10792 28733 10795
rect 28500 10764 28733 10792
rect 28500 10752 28506 10764
rect 28721 10761 28733 10764
rect 28767 10761 28779 10795
rect 28721 10755 28779 10761
rect 29825 10795 29883 10801
rect 29825 10761 29837 10795
rect 29871 10792 29883 10795
rect 30282 10792 30288 10804
rect 29871 10764 30288 10792
rect 29871 10761 29883 10764
rect 29825 10755 29883 10761
rect 30282 10752 30288 10764
rect 30340 10752 30346 10804
rect 31202 10752 31208 10804
rect 31260 10792 31266 10804
rect 31662 10792 31668 10804
rect 31260 10764 31668 10792
rect 31260 10752 31266 10764
rect 31662 10752 31668 10764
rect 31720 10752 31726 10804
rect 32674 10792 32680 10804
rect 32635 10764 32680 10792
rect 32674 10752 32680 10764
rect 32732 10752 32738 10804
rect 32858 10752 32864 10804
rect 32916 10792 32922 10804
rect 32953 10795 33011 10801
rect 32953 10792 32965 10795
rect 32916 10764 32965 10792
rect 32916 10752 32922 10764
rect 32953 10761 32965 10764
rect 32999 10761 33011 10795
rect 32953 10755 33011 10761
rect 33321 10795 33379 10801
rect 33321 10761 33333 10795
rect 33367 10792 33379 10795
rect 33962 10792 33968 10804
rect 33367 10764 33968 10792
rect 33367 10761 33379 10764
rect 33321 10755 33379 10761
rect 33962 10752 33968 10764
rect 34020 10752 34026 10804
rect 35710 10752 35716 10804
rect 35768 10792 35774 10804
rect 35897 10795 35955 10801
rect 35897 10792 35909 10795
rect 35768 10764 35909 10792
rect 35768 10752 35774 10764
rect 35897 10761 35909 10764
rect 35943 10761 35955 10795
rect 35897 10755 35955 10761
rect 8067 10696 8248 10724
rect 8067 10693 8079 10696
rect 8021 10687 8079 10693
rect 9490 10684 9496 10736
rect 9548 10724 9554 10736
rect 9585 10727 9643 10733
rect 9585 10724 9597 10727
rect 9548 10696 9597 10724
rect 9548 10684 9554 10696
rect 9585 10693 9597 10696
rect 9631 10693 9643 10727
rect 9585 10687 9643 10693
rect 14090 10684 14096 10736
rect 14148 10724 14154 10736
rect 15010 10724 15016 10736
rect 14148 10696 15016 10724
rect 14148 10684 14154 10696
rect 15010 10684 15016 10696
rect 15068 10684 15074 10736
rect 20714 10684 20720 10736
rect 20772 10724 20778 10736
rect 20901 10727 20959 10733
rect 20901 10724 20913 10727
rect 20772 10696 20913 10724
rect 20772 10684 20778 10696
rect 20901 10693 20913 10696
rect 20947 10693 20959 10727
rect 20901 10687 20959 10693
rect 22097 10727 22155 10733
rect 22097 10693 22109 10727
rect 22143 10724 22155 10727
rect 23566 10724 23572 10736
rect 22143 10696 23572 10724
rect 22143 10693 22155 10696
rect 22097 10687 22155 10693
rect 23566 10684 23572 10696
rect 23624 10724 23630 10736
rect 23624 10696 24256 10724
rect 23624 10684 23630 10696
rect 2593 10619 2651 10625
rect 2700 10628 4936 10656
rect 2700 10461 2728 10628
rect 4982 10616 4988 10668
rect 5040 10656 5046 10668
rect 5077 10659 5135 10665
rect 5077 10656 5089 10659
rect 5040 10628 5089 10656
rect 5040 10616 5046 10628
rect 5077 10625 5089 10628
rect 5123 10656 5135 10659
rect 5626 10656 5632 10668
rect 5123 10628 5632 10656
rect 5123 10625 5135 10628
rect 5077 10619 5135 10625
rect 5626 10616 5632 10628
rect 5684 10616 5690 10668
rect 5810 10656 5816 10668
rect 5771 10628 5816 10656
rect 5810 10616 5816 10628
rect 5868 10616 5874 10668
rect 9674 10616 9680 10668
rect 9732 10656 9738 10668
rect 10597 10659 10655 10665
rect 10597 10656 10609 10659
rect 9732 10628 10609 10656
rect 9732 10616 9738 10628
rect 10597 10625 10609 10628
rect 10643 10656 10655 10659
rect 10643 10628 12296 10656
rect 10643 10625 10655 10628
rect 10597 10619 10655 10625
rect 3697 10591 3755 10597
rect 3697 10557 3709 10591
rect 3743 10588 3755 10591
rect 4249 10591 4307 10597
rect 4249 10588 4261 10591
rect 3743 10560 4261 10588
rect 3743 10557 3755 10560
rect 3697 10551 3755 10557
rect 4249 10557 4261 10560
rect 4295 10588 4307 10591
rect 4798 10588 4804 10600
rect 4295 10560 4804 10588
rect 4295 10557 4307 10560
rect 4249 10551 4307 10557
rect 4798 10548 4804 10560
rect 4856 10548 4862 10600
rect 6546 10548 6552 10600
rect 6604 10588 6610 10600
rect 6825 10591 6883 10597
rect 6825 10588 6837 10591
rect 6604 10560 6837 10588
rect 6604 10548 6610 10560
rect 6825 10557 6837 10560
rect 6871 10588 6883 10591
rect 7377 10591 7435 10597
rect 7377 10588 7389 10591
rect 6871 10560 7389 10588
rect 6871 10557 6883 10560
rect 6825 10551 6883 10557
rect 7377 10557 7389 10560
rect 7423 10557 7435 10591
rect 7377 10551 7435 10557
rect 8205 10591 8263 10597
rect 8205 10557 8217 10591
rect 8251 10588 8263 10591
rect 8294 10588 8300 10600
rect 8251 10560 8300 10588
rect 8251 10557 8263 10560
rect 8205 10551 8263 10557
rect 8294 10548 8300 10560
rect 8352 10548 8358 10600
rect 8472 10591 8530 10597
rect 8472 10557 8484 10591
rect 8518 10588 8530 10591
rect 9582 10588 9588 10600
rect 8518 10560 9588 10588
rect 8518 10557 8530 10560
rect 8472 10551 8530 10557
rect 9582 10548 9588 10560
rect 9640 10548 9646 10600
rect 11054 10588 11060 10600
rect 11015 10560 11060 10588
rect 11054 10548 11060 10560
rect 11112 10548 11118 10600
rect 12268 10597 12296 10628
rect 18230 10616 18236 10668
rect 18288 10656 18294 10668
rect 18693 10659 18751 10665
rect 18693 10656 18705 10659
rect 18288 10628 18705 10656
rect 18288 10616 18294 10628
rect 18693 10625 18705 10628
rect 18739 10625 18751 10659
rect 18693 10619 18751 10625
rect 19610 10616 19616 10668
rect 19668 10656 19674 10668
rect 20257 10659 20315 10665
rect 20257 10656 20269 10659
rect 19668 10628 20269 10656
rect 19668 10616 19674 10628
rect 20257 10625 20269 10628
rect 20303 10625 20315 10659
rect 20257 10619 20315 10625
rect 22649 10659 22707 10665
rect 22649 10625 22661 10659
rect 22695 10656 22707 10659
rect 23014 10656 23020 10668
rect 22695 10628 23020 10656
rect 22695 10625 22707 10628
rect 22649 10619 22707 10625
rect 23014 10616 23020 10628
rect 23072 10616 23078 10668
rect 23477 10659 23535 10665
rect 23477 10625 23489 10659
rect 23523 10656 23535 10659
rect 24026 10656 24032 10668
rect 23523 10628 24032 10656
rect 23523 10625 23535 10628
rect 23477 10619 23535 10625
rect 24026 10616 24032 10628
rect 24084 10616 24090 10668
rect 24228 10665 24256 10696
rect 24213 10659 24271 10665
rect 24213 10625 24225 10659
rect 24259 10625 24271 10659
rect 24394 10656 24400 10668
rect 24307 10628 24400 10656
rect 24213 10619 24271 10625
rect 24394 10616 24400 10628
rect 24452 10656 24458 10668
rect 24762 10656 24768 10668
rect 24452 10628 24768 10656
rect 24452 10616 24458 10628
rect 24762 10616 24768 10628
rect 24820 10616 24826 10668
rect 25314 10656 25320 10668
rect 25275 10628 25320 10656
rect 25314 10616 25320 10628
rect 25372 10616 25378 10668
rect 25884 10656 25912 10752
rect 33686 10684 33692 10736
rect 33744 10724 33750 10736
rect 34977 10727 35035 10733
rect 34977 10724 34989 10727
rect 33744 10696 34989 10724
rect 33744 10684 33750 10696
rect 34977 10693 34989 10696
rect 35023 10693 35035 10727
rect 34977 10687 35035 10693
rect 35158 10684 35164 10736
rect 35216 10724 35222 10736
rect 35986 10724 35992 10736
rect 35216 10696 35992 10724
rect 35216 10684 35222 10696
rect 35986 10684 35992 10696
rect 36044 10684 36050 10736
rect 30285 10659 30343 10665
rect 30285 10656 30297 10659
rect 25884 10628 26556 10656
rect 12253 10591 12311 10597
rect 12253 10557 12265 10591
rect 12299 10588 12311 10591
rect 12621 10591 12679 10597
rect 12621 10588 12633 10591
rect 12299 10560 12633 10588
rect 12299 10557 12311 10560
rect 12253 10551 12311 10557
rect 12621 10557 12633 10560
rect 12667 10588 12679 10591
rect 12710 10588 12716 10600
rect 12667 10560 12716 10588
rect 12667 10557 12679 10560
rect 12621 10551 12679 10557
rect 12710 10548 12716 10560
rect 12768 10548 12774 10600
rect 15102 10588 15108 10600
rect 15063 10560 15108 10588
rect 15102 10548 15108 10560
rect 15160 10548 15166 10600
rect 16942 10548 16948 10600
rect 17000 10588 17006 10600
rect 17773 10591 17831 10597
rect 17773 10588 17785 10591
rect 17000 10560 17785 10588
rect 17000 10548 17006 10560
rect 17773 10557 17785 10560
rect 17819 10588 17831 10591
rect 18322 10588 18328 10600
rect 17819 10560 18328 10588
rect 17819 10557 17831 10560
rect 17773 10551 17831 10557
rect 18322 10548 18328 10560
rect 18380 10588 18386 10600
rect 18417 10591 18475 10597
rect 18417 10588 18429 10591
rect 18380 10560 18429 10588
rect 18380 10548 18386 10560
rect 18417 10557 18429 10560
rect 18463 10557 18475 10591
rect 18417 10551 18475 10557
rect 19521 10591 19579 10597
rect 19521 10557 19533 10591
rect 19567 10588 19579 10591
rect 19978 10588 19984 10600
rect 19567 10560 19984 10588
rect 19567 10557 19579 10560
rect 19521 10551 19579 10557
rect 19978 10548 19984 10560
rect 20036 10548 20042 10600
rect 26421 10591 26479 10597
rect 26421 10557 26433 10591
rect 26467 10557 26479 10591
rect 26528 10588 26556 10628
rect 30116 10628 30297 10656
rect 26694 10597 26700 10600
rect 26677 10591 26700 10597
rect 26677 10588 26689 10591
rect 26528 10560 26689 10588
rect 26421 10551 26479 10557
rect 26677 10557 26689 10560
rect 26752 10588 26758 10600
rect 26752 10560 26825 10588
rect 26677 10551 26700 10557
rect 2777 10523 2835 10529
rect 2777 10489 2789 10523
rect 2823 10520 2835 10523
rect 3142 10520 3148 10532
rect 2823 10492 3148 10520
rect 2823 10489 2835 10492
rect 2777 10483 2835 10489
rect 3142 10480 3148 10492
rect 3200 10480 3206 10532
rect 4614 10480 4620 10532
rect 4672 10520 4678 10532
rect 4709 10523 4767 10529
rect 4709 10520 4721 10523
rect 4672 10492 4721 10520
rect 4672 10480 4678 10492
rect 4709 10489 4721 10492
rect 4755 10520 4767 10523
rect 4755 10492 5488 10520
rect 4755 10489 4767 10492
rect 4709 10483 4767 10489
rect 2041 10455 2099 10461
rect 2041 10421 2053 10455
rect 2087 10452 2099 10455
rect 2685 10455 2743 10461
rect 2685 10452 2697 10455
rect 2087 10424 2697 10452
rect 2087 10421 2099 10424
rect 2041 10415 2099 10421
rect 2685 10421 2697 10424
rect 2731 10421 2743 10455
rect 2685 10415 2743 10421
rect 3605 10455 3663 10461
rect 3605 10421 3617 10455
rect 3651 10452 3663 10455
rect 3694 10452 3700 10464
rect 3651 10424 3700 10452
rect 3651 10421 3663 10424
rect 3605 10415 3663 10421
rect 3694 10412 3700 10424
rect 3752 10452 3758 10464
rect 5350 10452 5356 10464
rect 3752 10424 5356 10452
rect 3752 10412 3758 10424
rect 5350 10412 5356 10424
rect 5408 10412 5414 10464
rect 5460 10452 5488 10492
rect 10318 10480 10324 10532
rect 10376 10520 10382 10532
rect 11241 10523 11299 10529
rect 11241 10520 11253 10523
rect 10376 10492 11253 10520
rect 10376 10480 10382 10492
rect 11241 10489 11253 10492
rect 11287 10489 11299 10523
rect 11241 10483 11299 10489
rect 11330 10480 11336 10532
rect 11388 10520 11394 10532
rect 12888 10523 12946 10529
rect 12888 10520 12900 10523
rect 11388 10492 11433 10520
rect 11808 10492 12900 10520
rect 11388 10480 11394 10492
rect 11808 10464 11836 10492
rect 12888 10489 12900 10492
rect 12934 10520 12946 10523
rect 13538 10520 13544 10532
rect 12934 10492 13544 10520
rect 12934 10489 12946 10492
rect 12888 10483 12946 10489
rect 13538 10480 13544 10492
rect 13596 10480 13602 10532
rect 15350 10523 15408 10529
rect 15350 10520 15362 10523
rect 14016 10492 15362 10520
rect 5721 10455 5779 10461
rect 5721 10452 5733 10455
rect 5460 10424 5733 10452
rect 5721 10421 5733 10424
rect 5767 10452 5779 10455
rect 5810 10452 5816 10464
rect 5767 10424 5816 10452
rect 5767 10421 5779 10424
rect 5721 10415 5779 10421
rect 5810 10412 5816 10424
rect 5868 10412 5874 10464
rect 6641 10455 6699 10461
rect 6641 10421 6653 10455
rect 6687 10452 6699 10455
rect 6822 10452 6828 10464
rect 6687 10424 6828 10452
rect 6687 10421 6699 10424
rect 6641 10415 6699 10421
rect 6822 10412 6828 10424
rect 6880 10412 6886 10464
rect 11790 10452 11796 10464
rect 11751 10424 11796 10452
rect 11790 10412 11796 10424
rect 11848 10412 11854 10464
rect 13078 10412 13084 10464
rect 13136 10452 13142 10464
rect 14016 10461 14044 10492
rect 15350 10489 15362 10492
rect 15396 10489 15408 10523
rect 22373 10523 22431 10529
rect 15350 10483 15408 10489
rect 17420 10492 17908 10520
rect 17420 10464 17448 10492
rect 14001 10455 14059 10461
rect 14001 10452 14013 10455
rect 13136 10424 14013 10452
rect 13136 10412 13142 10424
rect 14001 10421 14013 10424
rect 14047 10421 14059 10455
rect 16482 10452 16488 10464
rect 16443 10424 16488 10452
rect 14001 10415 14059 10421
rect 16482 10412 16488 10424
rect 16540 10412 16546 10464
rect 17126 10452 17132 10464
rect 17087 10424 17132 10452
rect 17126 10412 17132 10424
rect 17184 10412 17190 10464
rect 17402 10452 17408 10464
rect 17363 10424 17408 10452
rect 17402 10412 17408 10424
rect 17460 10412 17466 10464
rect 17880 10452 17908 10492
rect 22373 10489 22385 10523
rect 22419 10489 22431 10523
rect 24302 10520 24308 10532
rect 24263 10492 24308 10520
rect 22373 10483 22431 10489
rect 18601 10455 18659 10461
rect 18601 10452 18613 10455
rect 17880 10424 18613 10452
rect 18601 10421 18613 10424
rect 18647 10421 18659 10455
rect 20162 10452 20168 10464
rect 20123 10424 20168 10452
rect 18601 10415 18659 10421
rect 20162 10412 20168 10424
rect 20220 10412 20226 10464
rect 21913 10455 21971 10461
rect 21913 10421 21925 10455
rect 21959 10452 21971 10455
rect 22002 10452 22008 10464
rect 21959 10424 22008 10452
rect 21959 10421 21971 10424
rect 21913 10415 21971 10421
rect 22002 10412 22008 10424
rect 22060 10452 22066 10464
rect 22388 10452 22416 10483
rect 24302 10480 24308 10492
rect 24360 10480 24366 10532
rect 24486 10480 24492 10532
rect 24544 10520 24550 10532
rect 26237 10523 26295 10529
rect 26237 10520 26249 10523
rect 24544 10492 26249 10520
rect 24544 10480 24550 10492
rect 26237 10489 26249 10492
rect 26283 10520 26295 10523
rect 26436 10520 26464 10551
rect 26694 10548 26700 10551
rect 26752 10548 26758 10560
rect 27062 10520 27068 10532
rect 26283 10492 27068 10520
rect 26283 10489 26295 10492
rect 26237 10483 26295 10489
rect 27062 10480 27068 10492
rect 27120 10520 27126 10532
rect 28166 10520 28172 10532
rect 27120 10492 28172 10520
rect 27120 10480 27126 10492
rect 28166 10480 28172 10492
rect 28224 10520 28230 10532
rect 28353 10523 28411 10529
rect 28353 10520 28365 10523
rect 28224 10492 28365 10520
rect 28224 10480 28230 10492
rect 28353 10489 28365 10492
rect 28399 10520 28411 10523
rect 29086 10520 29092 10532
rect 28399 10492 29092 10520
rect 28399 10489 28411 10492
rect 28353 10483 28411 10489
rect 29086 10480 29092 10492
rect 29144 10520 29150 10532
rect 30116 10529 30144 10628
rect 30285 10625 30297 10628
rect 30331 10625 30343 10659
rect 30285 10619 30343 10625
rect 33134 10616 33140 10668
rect 33192 10656 33198 10668
rect 33781 10659 33839 10665
rect 33781 10656 33793 10659
rect 33192 10628 33793 10656
rect 33192 10616 33198 10628
rect 33781 10625 33793 10628
rect 33827 10656 33839 10659
rect 34146 10656 34152 10668
rect 33827 10628 34152 10656
rect 33827 10625 33839 10628
rect 33781 10619 33839 10625
rect 34146 10616 34152 10628
rect 34204 10616 34210 10668
rect 36262 10656 36268 10668
rect 34256 10628 36268 10656
rect 32309 10591 32367 10597
rect 32309 10557 32321 10591
rect 32355 10588 32367 10591
rect 32766 10588 32772 10600
rect 32355 10560 32772 10588
rect 32355 10557 32367 10560
rect 32309 10551 32367 10557
rect 32766 10548 32772 10560
rect 32824 10588 32830 10600
rect 33870 10588 33876 10600
rect 32824 10560 33876 10588
rect 32824 10548 32830 10560
rect 33870 10548 33876 10560
rect 33928 10548 33934 10600
rect 30101 10523 30159 10529
rect 30101 10520 30113 10523
rect 29144 10492 30113 10520
rect 29144 10480 29150 10492
rect 30101 10489 30113 10492
rect 30147 10489 30159 10523
rect 30101 10483 30159 10489
rect 30552 10523 30610 10529
rect 30552 10489 30564 10523
rect 30598 10520 30610 10523
rect 30834 10520 30840 10532
rect 30598 10492 30840 10520
rect 30598 10489 30610 10492
rect 30552 10483 30610 10489
rect 30834 10480 30840 10492
rect 30892 10480 30898 10532
rect 33686 10480 33692 10532
rect 33744 10520 33750 10532
rect 33781 10523 33839 10529
rect 33781 10520 33793 10523
rect 33744 10492 33793 10520
rect 33744 10480 33750 10492
rect 33781 10489 33793 10492
rect 33827 10489 33839 10523
rect 33781 10483 33839 10489
rect 22060 10424 22416 10452
rect 22557 10455 22615 10461
rect 22060 10412 22066 10424
rect 22557 10421 22569 10455
rect 22603 10452 22615 10455
rect 22922 10452 22928 10464
rect 22603 10424 22928 10452
rect 22603 10421 22615 10424
rect 22557 10415 22615 10421
rect 22922 10412 22928 10424
rect 22980 10412 22986 10464
rect 24854 10412 24860 10464
rect 24912 10452 24918 10464
rect 24949 10455 25007 10461
rect 24949 10452 24961 10455
rect 24912 10424 24961 10452
rect 24912 10412 24918 10424
rect 24949 10421 24961 10424
rect 24995 10421 25007 10455
rect 24949 10415 25007 10421
rect 30006 10412 30012 10464
rect 30064 10452 30070 10464
rect 34256 10452 34284 10628
rect 36262 10616 36268 10628
rect 36320 10656 36326 10668
rect 37274 10656 37280 10668
rect 36320 10628 37280 10656
rect 36320 10616 36326 10628
rect 37274 10616 37280 10628
rect 37332 10616 37338 10668
rect 34333 10591 34391 10597
rect 34333 10557 34345 10591
rect 34379 10588 34391 10591
rect 34379 10560 35572 10588
rect 34379 10557 34391 10560
rect 34333 10551 34391 10557
rect 35544 10532 35572 10560
rect 35986 10548 35992 10600
rect 36044 10588 36050 10600
rect 36449 10591 36507 10597
rect 36449 10588 36461 10591
rect 36044 10560 36461 10588
rect 36044 10548 36050 10560
rect 36449 10557 36461 10560
rect 36495 10588 36507 10591
rect 37001 10591 37059 10597
rect 37001 10588 37013 10591
rect 36495 10560 37013 10588
rect 36495 10557 36507 10560
rect 36449 10551 36507 10557
rect 37001 10557 37013 10560
rect 37047 10557 37059 10591
rect 37001 10551 37059 10557
rect 35253 10523 35311 10529
rect 35253 10489 35265 10523
rect 35299 10489 35311 10523
rect 35526 10520 35532 10532
rect 35487 10492 35532 10520
rect 35253 10483 35311 10489
rect 34606 10452 34612 10464
rect 30064 10424 34284 10452
rect 34567 10424 34612 10452
rect 30064 10412 30070 10424
rect 34606 10412 34612 10424
rect 34664 10452 34670 10464
rect 35158 10452 35164 10464
rect 34664 10424 35164 10452
rect 34664 10412 34670 10424
rect 35158 10412 35164 10424
rect 35216 10452 35222 10464
rect 35268 10452 35296 10483
rect 35526 10480 35532 10492
rect 35584 10480 35590 10532
rect 35216 10424 35296 10452
rect 35437 10455 35495 10461
rect 35216 10412 35222 10424
rect 35437 10421 35449 10455
rect 35483 10452 35495 10455
rect 35618 10452 35624 10464
rect 35483 10424 35624 10452
rect 35483 10421 35495 10424
rect 35437 10415 35495 10421
rect 35618 10412 35624 10424
rect 35676 10412 35682 10464
rect 36354 10452 36360 10464
rect 36315 10424 36360 10452
rect 36354 10412 36360 10424
rect 36412 10412 36418 10464
rect 36633 10455 36691 10461
rect 36633 10421 36645 10455
rect 36679 10452 36691 10455
rect 36906 10452 36912 10464
rect 36679 10424 36912 10452
rect 36679 10421 36691 10424
rect 36633 10415 36691 10421
rect 36906 10412 36912 10424
rect 36964 10412 36970 10464
rect 1104 10362 38824 10384
rect 1104 10310 14315 10362
rect 14367 10310 14379 10362
rect 14431 10310 14443 10362
rect 14495 10310 14507 10362
rect 14559 10310 27648 10362
rect 27700 10310 27712 10362
rect 27764 10310 27776 10362
rect 27828 10310 27840 10362
rect 27892 10310 38824 10362
rect 1104 10288 38824 10310
rect 1670 10208 1676 10260
rect 1728 10248 1734 10260
rect 2501 10251 2559 10257
rect 2501 10248 2513 10251
rect 1728 10220 2513 10248
rect 1728 10208 1734 10220
rect 2501 10217 2513 10220
rect 2547 10217 2559 10251
rect 2501 10211 2559 10217
rect 4062 10208 4068 10260
rect 4120 10248 4126 10260
rect 4249 10251 4307 10257
rect 4249 10248 4261 10251
rect 4120 10220 4261 10248
rect 4120 10208 4126 10220
rect 4249 10217 4261 10220
rect 4295 10217 4307 10251
rect 4249 10211 4307 10217
rect 5902 10208 5908 10260
rect 5960 10248 5966 10260
rect 6638 10248 6644 10260
rect 5960 10220 6644 10248
rect 5960 10208 5966 10220
rect 6638 10208 6644 10220
rect 6696 10208 6702 10260
rect 7285 10251 7343 10257
rect 7285 10217 7297 10251
rect 7331 10248 7343 10251
rect 7929 10251 7987 10257
rect 7929 10248 7941 10251
rect 7331 10220 7941 10248
rect 7331 10217 7343 10220
rect 7285 10211 7343 10217
rect 7929 10217 7941 10220
rect 7975 10248 7987 10251
rect 9122 10248 9128 10260
rect 7975 10220 9128 10248
rect 7975 10217 7987 10220
rect 7929 10211 7987 10217
rect 2222 10140 2228 10192
rect 2280 10180 2286 10192
rect 5534 10189 5540 10192
rect 2317 10183 2375 10189
rect 2317 10180 2329 10183
rect 2280 10152 2329 10180
rect 2280 10140 2286 10152
rect 2317 10149 2329 10152
rect 2363 10149 2375 10183
rect 5528 10180 5540 10189
rect 5495 10152 5540 10180
rect 2317 10143 2375 10149
rect 5528 10143 5540 10152
rect 2332 10112 2360 10143
rect 5534 10140 5540 10143
rect 5592 10140 5598 10192
rect 8294 10140 8300 10192
rect 8352 10180 8358 10192
rect 8680 10189 8708 10220
rect 9122 10208 9128 10220
rect 9180 10208 9186 10260
rect 9858 10248 9864 10260
rect 9819 10220 9864 10248
rect 9858 10208 9864 10220
rect 9916 10208 9922 10260
rect 10318 10248 10324 10260
rect 10279 10220 10324 10248
rect 10318 10208 10324 10220
rect 10376 10208 10382 10260
rect 12529 10251 12587 10257
rect 12529 10217 12541 10251
rect 12575 10248 12587 10251
rect 13078 10248 13084 10260
rect 12575 10220 13084 10248
rect 12575 10217 12587 10220
rect 12529 10211 12587 10217
rect 13078 10208 13084 10220
rect 13136 10208 13142 10260
rect 16482 10248 16488 10260
rect 16443 10220 16488 10248
rect 16482 10208 16488 10220
rect 16540 10208 16546 10260
rect 18230 10248 18236 10260
rect 18191 10220 18236 10248
rect 18230 10208 18236 10220
rect 18288 10208 18294 10260
rect 18782 10248 18788 10260
rect 18743 10220 18788 10248
rect 18782 10208 18788 10220
rect 18840 10208 18846 10260
rect 18874 10208 18880 10260
rect 18932 10248 18938 10260
rect 19153 10251 19211 10257
rect 19153 10248 19165 10251
rect 18932 10220 19165 10248
rect 18932 10208 18938 10220
rect 19153 10217 19165 10220
rect 19199 10217 19211 10251
rect 21818 10248 21824 10260
rect 21779 10220 21824 10248
rect 19153 10211 19211 10217
rect 21818 10208 21824 10220
rect 21876 10208 21882 10260
rect 23937 10251 23995 10257
rect 23937 10217 23949 10251
rect 23983 10248 23995 10251
rect 24394 10248 24400 10260
rect 23983 10220 24400 10248
rect 23983 10217 23995 10220
rect 23937 10211 23995 10217
rect 24394 10208 24400 10220
rect 24452 10208 24458 10260
rect 25225 10251 25283 10257
rect 25225 10217 25237 10251
rect 25271 10248 25283 10251
rect 26142 10248 26148 10260
rect 25271 10220 26148 10248
rect 25271 10217 25283 10220
rect 25225 10211 25283 10217
rect 8573 10183 8631 10189
rect 8573 10180 8585 10183
rect 8352 10152 8585 10180
rect 8352 10140 8358 10152
rect 8573 10149 8585 10152
rect 8619 10149 8631 10183
rect 8573 10143 8631 10149
rect 8665 10183 8723 10189
rect 8665 10149 8677 10183
rect 8711 10149 8723 10183
rect 8665 10143 8723 10149
rect 9490 10140 9496 10192
rect 9548 10180 9554 10192
rect 10689 10183 10747 10189
rect 10689 10180 10701 10183
rect 9548 10152 10701 10180
rect 9548 10140 9554 10152
rect 10689 10149 10701 10152
rect 10735 10180 10747 10183
rect 11330 10180 11336 10192
rect 10735 10152 11336 10180
rect 10735 10149 10747 10152
rect 10689 10143 10747 10149
rect 11330 10140 11336 10152
rect 11388 10140 11394 10192
rect 11698 10180 11704 10192
rect 11659 10152 11704 10180
rect 11698 10140 11704 10152
rect 11756 10140 11762 10192
rect 15286 10140 15292 10192
rect 15344 10180 15350 10192
rect 15841 10183 15899 10189
rect 15841 10180 15853 10183
rect 15344 10152 15853 10180
rect 15344 10140 15350 10152
rect 15841 10149 15853 10152
rect 15887 10149 15899 10183
rect 16500 10180 16528 10208
rect 17034 10180 17040 10192
rect 16500 10152 17040 10180
rect 15841 10143 15899 10149
rect 17034 10140 17040 10152
rect 17092 10189 17098 10192
rect 17092 10183 17156 10189
rect 17092 10149 17110 10183
rect 17144 10149 17156 10183
rect 17092 10143 17156 10149
rect 22180 10183 22238 10189
rect 22180 10149 22192 10183
rect 22226 10180 22238 10183
rect 22370 10180 22376 10192
rect 22226 10152 22376 10180
rect 22226 10149 22238 10152
rect 22180 10143 22238 10149
rect 17092 10140 17098 10143
rect 22370 10140 22376 10152
rect 22428 10140 22434 10192
rect 3697 10115 3755 10121
rect 3697 10112 3709 10115
rect 2332 10084 3709 10112
rect 3697 10081 3709 10084
rect 3743 10081 3755 10115
rect 3697 10075 3755 10081
rect 4065 10115 4123 10121
rect 4065 10081 4077 10115
rect 4111 10112 4123 10115
rect 4338 10112 4344 10124
rect 4111 10084 4344 10112
rect 4111 10081 4123 10084
rect 4065 10075 4123 10081
rect 4338 10072 4344 10084
rect 4396 10072 4402 10124
rect 5261 10115 5319 10121
rect 5261 10081 5273 10115
rect 5307 10112 5319 10115
rect 5350 10112 5356 10124
rect 5307 10084 5356 10112
rect 5307 10081 5319 10084
rect 5261 10075 5319 10081
rect 5350 10072 5356 10084
rect 5408 10072 5414 10124
rect 9677 10115 9735 10121
rect 9677 10081 9689 10115
rect 9723 10112 9735 10115
rect 10502 10112 10508 10124
rect 9723 10084 10508 10112
rect 9723 10081 9735 10084
rect 9677 10075 9735 10081
rect 10502 10072 10508 10084
rect 10560 10072 10566 10124
rect 11514 10112 11520 10124
rect 11475 10084 11520 10112
rect 11514 10072 11520 10084
rect 11572 10072 11578 10124
rect 12158 10072 12164 10124
rect 12216 10112 12222 10124
rect 12969 10115 13027 10121
rect 12969 10112 12981 10115
rect 12216 10084 12981 10112
rect 12216 10072 12222 10084
rect 12969 10081 12981 10084
rect 13015 10081 13027 10115
rect 15654 10112 15660 10124
rect 15615 10084 15660 10112
rect 12969 10075 13027 10081
rect 15654 10072 15660 10084
rect 15712 10072 15718 10124
rect 16853 10115 16911 10121
rect 16853 10112 16865 10115
rect 15764 10084 16865 10112
rect 1857 10047 1915 10053
rect 1857 10013 1869 10047
rect 1903 10044 1915 10047
rect 1946 10044 1952 10056
rect 1903 10016 1952 10044
rect 1903 10013 1915 10016
rect 1857 10007 1915 10013
rect 1946 10004 1952 10016
rect 2004 10044 2010 10056
rect 2590 10044 2596 10056
rect 2004 10016 2596 10044
rect 2004 10004 2010 10016
rect 2590 10004 2596 10016
rect 2648 10004 2654 10056
rect 4614 10044 4620 10056
rect 4575 10016 4620 10044
rect 4614 10004 4620 10016
rect 4672 10004 4678 10056
rect 8478 10044 8484 10056
rect 8439 10016 8484 10044
rect 8478 10004 8484 10016
rect 8536 10004 8542 10056
rect 11790 10044 11796 10056
rect 11751 10016 11796 10044
rect 11790 10004 11796 10016
rect 11848 10004 11854 10056
rect 12710 10044 12716 10056
rect 12671 10016 12716 10044
rect 12710 10004 12716 10016
rect 12768 10004 12774 10056
rect 13722 10004 13728 10056
rect 13780 10044 13786 10056
rect 15102 10044 15108 10056
rect 13780 10016 15108 10044
rect 13780 10004 13786 10016
rect 15102 10004 15108 10016
rect 15160 10044 15166 10056
rect 15764 10044 15792 10084
rect 16853 10081 16865 10084
rect 16899 10112 16911 10115
rect 17678 10112 17684 10124
rect 16899 10084 17684 10112
rect 16899 10081 16911 10084
rect 16853 10075 16911 10081
rect 17678 10072 17684 10084
rect 17736 10072 17742 10124
rect 24394 10072 24400 10124
rect 24452 10112 24458 10124
rect 25240 10112 25268 10211
rect 26142 10208 26148 10220
rect 26200 10208 26206 10260
rect 26326 10248 26332 10260
rect 26287 10220 26332 10248
rect 26326 10208 26332 10220
rect 26384 10208 26390 10260
rect 26694 10248 26700 10260
rect 26655 10220 26700 10248
rect 26694 10208 26700 10220
rect 26752 10208 26758 10260
rect 35526 10208 35532 10260
rect 35584 10248 35590 10260
rect 36078 10248 36084 10260
rect 35584 10220 36084 10248
rect 35584 10208 35590 10220
rect 36078 10208 36084 10220
rect 36136 10248 36142 10260
rect 36357 10251 36415 10257
rect 36357 10248 36369 10251
rect 36136 10220 36369 10248
rect 36136 10208 36142 10220
rect 36357 10217 36369 10220
rect 36403 10217 36415 10251
rect 36357 10211 36415 10217
rect 25317 10183 25375 10189
rect 25317 10149 25329 10183
rect 25363 10180 25375 10183
rect 25406 10180 25412 10192
rect 25363 10152 25412 10180
rect 25363 10149 25375 10152
rect 25317 10143 25375 10149
rect 25406 10140 25412 10152
rect 25464 10180 25470 10192
rect 26510 10180 26516 10192
rect 25464 10152 26516 10180
rect 25464 10140 25470 10152
rect 26510 10140 26516 10152
rect 26568 10140 26574 10192
rect 27338 10189 27344 10192
rect 27332 10180 27344 10189
rect 27299 10152 27344 10180
rect 27332 10143 27344 10152
rect 27338 10140 27344 10143
rect 27396 10140 27402 10192
rect 28902 10140 28908 10192
rect 28960 10140 28966 10192
rect 28994 10140 29000 10192
rect 29052 10180 29058 10192
rect 30006 10180 30012 10192
rect 29052 10152 30012 10180
rect 29052 10140 29058 10152
rect 30006 10140 30012 10152
rect 30064 10140 30070 10192
rect 30101 10183 30159 10189
rect 30101 10149 30113 10183
rect 30147 10180 30159 10183
rect 30745 10183 30803 10189
rect 30745 10180 30757 10183
rect 30147 10152 30757 10180
rect 30147 10149 30159 10152
rect 30101 10143 30159 10149
rect 30745 10149 30757 10152
rect 30791 10180 30803 10183
rect 30926 10180 30932 10192
rect 30791 10152 30932 10180
rect 30791 10149 30803 10152
rect 30745 10143 30803 10149
rect 30926 10140 30932 10152
rect 30984 10140 30990 10192
rect 31662 10140 31668 10192
rect 31720 10180 31726 10192
rect 31846 10180 31852 10192
rect 31720 10152 31852 10180
rect 31720 10140 31726 10152
rect 31846 10140 31852 10152
rect 31904 10180 31910 10192
rect 32462 10183 32520 10189
rect 32462 10180 32474 10183
rect 31904 10152 32474 10180
rect 31904 10140 31910 10152
rect 32462 10149 32474 10152
rect 32508 10149 32520 10183
rect 32462 10143 32520 10149
rect 27062 10112 27068 10124
rect 24452 10084 25268 10112
rect 27023 10084 27068 10112
rect 24452 10072 24458 10084
rect 27062 10072 27068 10084
rect 27120 10072 27126 10124
rect 28920 10112 28948 10140
rect 27172 10084 28948 10112
rect 29733 10115 29791 10121
rect 15930 10044 15936 10056
rect 15160 10016 15792 10044
rect 15891 10016 15936 10044
rect 15160 10004 15166 10016
rect 15930 10004 15936 10016
rect 15988 10004 15994 10056
rect 20714 10004 20720 10056
rect 20772 10044 20778 10056
rect 21913 10047 21971 10053
rect 21913 10044 21925 10047
rect 20772 10016 21925 10044
rect 20772 10004 20778 10016
rect 21913 10013 21925 10016
rect 21959 10013 21971 10047
rect 25222 10044 25228 10056
rect 25183 10016 25228 10044
rect 21913 10007 21971 10013
rect 25222 10004 25228 10016
rect 25280 10004 25286 10056
rect 25314 10004 25320 10056
rect 25372 10044 25378 10056
rect 27172 10044 27200 10084
rect 29733 10081 29745 10115
rect 29779 10112 29791 10115
rect 30558 10112 30564 10124
rect 29779 10084 30564 10112
rect 29779 10081 29791 10084
rect 29733 10075 29791 10081
rect 30558 10072 30564 10084
rect 30616 10072 30622 10124
rect 32217 10115 32275 10121
rect 32217 10081 32229 10115
rect 32263 10112 32275 10115
rect 32858 10112 32864 10124
rect 32263 10084 32864 10112
rect 32263 10081 32275 10084
rect 32217 10075 32275 10081
rect 32858 10072 32864 10084
rect 32916 10072 32922 10124
rect 34885 10115 34943 10121
rect 34885 10081 34897 10115
rect 34931 10112 34943 10115
rect 35244 10115 35302 10121
rect 35244 10112 35256 10115
rect 34931 10084 35256 10112
rect 34931 10081 34943 10084
rect 34885 10075 34943 10081
rect 35244 10081 35256 10084
rect 35290 10112 35302 10115
rect 35526 10112 35532 10124
rect 35290 10084 35532 10112
rect 35290 10081 35302 10084
rect 35244 10075 35302 10081
rect 30834 10044 30840 10056
rect 25372 10016 27200 10044
rect 30747 10016 30840 10044
rect 25372 10004 25378 10016
rect 30834 10004 30840 10016
rect 30892 10044 30898 10056
rect 31662 10044 31668 10056
rect 30892 10016 31668 10044
rect 30892 10004 30898 10016
rect 31662 10004 31668 10016
rect 31720 10004 31726 10056
rect 3053 9979 3111 9985
rect 3053 9945 3065 9979
rect 3099 9976 3111 9979
rect 3142 9976 3148 9988
rect 3099 9948 3148 9976
rect 3099 9945 3111 9948
rect 3053 9939 3111 9945
rect 3142 9936 3148 9948
rect 3200 9976 3206 9988
rect 3694 9976 3700 9988
rect 3200 9948 3700 9976
rect 3200 9936 3206 9948
rect 3694 9936 3700 9948
rect 3752 9936 3758 9988
rect 8110 9976 8116 9988
rect 8071 9948 8116 9976
rect 8110 9936 8116 9948
rect 8168 9936 8174 9988
rect 11241 9979 11299 9985
rect 11241 9945 11253 9979
rect 11287 9976 11299 9979
rect 12342 9976 12348 9988
rect 11287 9948 12348 9976
rect 11287 9945 11299 9948
rect 11241 9939 11299 9945
rect 12342 9936 12348 9948
rect 12400 9936 12406 9988
rect 24670 9936 24676 9988
rect 24728 9976 24734 9988
rect 24765 9979 24823 9985
rect 24765 9976 24777 9979
rect 24728 9948 24777 9976
rect 24728 9936 24734 9948
rect 24765 9945 24777 9948
rect 24811 9945 24823 9979
rect 24765 9939 24823 9945
rect 30190 9936 30196 9988
rect 30248 9976 30254 9988
rect 30285 9979 30343 9985
rect 30285 9976 30297 9979
rect 30248 9948 30297 9976
rect 30248 9936 30254 9948
rect 30285 9945 30297 9948
rect 30331 9945 30343 9979
rect 30285 9939 30343 9945
rect 33597 9979 33655 9985
rect 33597 9945 33609 9979
rect 33643 9976 33655 9979
rect 34900 9976 34928 10075
rect 35526 10072 35532 10084
rect 35584 10072 35590 10124
rect 34977 10047 35035 10053
rect 34977 10013 34989 10047
rect 35023 10013 35035 10047
rect 34977 10007 35035 10013
rect 33643 9948 34928 9976
rect 33643 9945 33655 9948
rect 33597 9939 33655 9945
rect 2041 9911 2099 9917
rect 2041 9877 2053 9911
rect 2087 9908 2099 9911
rect 2406 9908 2412 9920
rect 2087 9880 2412 9908
rect 2087 9877 2099 9880
rect 2041 9871 2099 9877
rect 2406 9868 2412 9880
rect 2464 9868 2470 9920
rect 3418 9908 3424 9920
rect 3331 9880 3424 9908
rect 3418 9868 3424 9880
rect 3476 9908 3482 9920
rect 4062 9908 4068 9920
rect 3476 9880 4068 9908
rect 3476 9868 3482 9880
rect 4062 9868 4068 9880
rect 4120 9868 4126 9920
rect 5074 9908 5080 9920
rect 5035 9880 5080 9908
rect 5074 9868 5080 9880
rect 5132 9868 5138 9920
rect 13630 9868 13636 9920
rect 13688 9908 13694 9920
rect 14093 9911 14151 9917
rect 14093 9908 14105 9911
rect 13688 9880 14105 9908
rect 13688 9868 13694 9880
rect 14093 9877 14105 9880
rect 14139 9877 14151 9911
rect 15378 9908 15384 9920
rect 15339 9880 15384 9908
rect 14093 9871 14151 9877
rect 15378 9868 15384 9880
rect 15436 9868 15442 9920
rect 19705 9911 19763 9917
rect 19705 9877 19717 9911
rect 19751 9908 19763 9911
rect 20162 9908 20168 9920
rect 19751 9880 20168 9908
rect 19751 9877 19763 9880
rect 19705 9871 19763 9877
rect 20162 9868 20168 9880
rect 20220 9908 20226 9920
rect 20530 9908 20536 9920
rect 20220 9880 20536 9908
rect 20220 9868 20226 9880
rect 20530 9868 20536 9880
rect 20588 9868 20594 9920
rect 23293 9911 23351 9917
rect 23293 9877 23305 9911
rect 23339 9908 23351 9911
rect 23474 9908 23480 9920
rect 23339 9880 23480 9908
rect 23339 9877 23351 9880
rect 23293 9871 23351 9877
rect 23474 9868 23480 9880
rect 23532 9868 23538 9920
rect 24486 9908 24492 9920
rect 24447 9880 24492 9908
rect 24486 9868 24492 9880
rect 24544 9868 24550 9920
rect 28442 9908 28448 9920
rect 28403 9880 28448 9908
rect 28442 9868 28448 9880
rect 28500 9868 28506 9920
rect 31018 9868 31024 9920
rect 31076 9908 31082 9920
rect 31205 9911 31263 9917
rect 31205 9908 31217 9911
rect 31076 9880 31217 9908
rect 31076 9868 31082 9880
rect 31205 9877 31217 9880
rect 31251 9877 31263 9911
rect 31205 9871 31263 9877
rect 31941 9911 31999 9917
rect 31941 9877 31953 9911
rect 31987 9908 31999 9911
rect 32582 9908 32588 9920
rect 31987 9880 32588 9908
rect 31987 9877 31999 9880
rect 31941 9871 31999 9877
rect 32582 9868 32588 9880
rect 32640 9868 32646 9920
rect 33870 9868 33876 9920
rect 33928 9908 33934 9920
rect 34149 9911 34207 9917
rect 34149 9908 34161 9911
rect 33928 9880 34161 9908
rect 33928 9868 33934 9880
rect 34149 9877 34161 9880
rect 34195 9877 34207 9911
rect 34149 9871 34207 9877
rect 34698 9868 34704 9920
rect 34756 9908 34762 9920
rect 34992 9908 35020 10007
rect 34756 9880 35020 9908
rect 34756 9868 34762 9880
rect 1104 9818 38824 9840
rect 1104 9766 7648 9818
rect 7700 9766 7712 9818
rect 7764 9766 7776 9818
rect 7828 9766 7840 9818
rect 7892 9766 20982 9818
rect 21034 9766 21046 9818
rect 21098 9766 21110 9818
rect 21162 9766 21174 9818
rect 21226 9766 34315 9818
rect 34367 9766 34379 9818
rect 34431 9766 34443 9818
rect 34495 9766 34507 9818
rect 34559 9766 38824 9818
rect 1104 9744 38824 9766
rect 3786 9664 3792 9716
rect 3844 9704 3850 9716
rect 4522 9704 4528 9716
rect 3844 9676 4528 9704
rect 3844 9664 3850 9676
rect 4522 9664 4528 9676
rect 4580 9664 4586 9716
rect 5534 9664 5540 9716
rect 5592 9704 5598 9716
rect 5813 9707 5871 9713
rect 5813 9704 5825 9707
rect 5592 9676 5825 9704
rect 5592 9664 5598 9676
rect 5813 9673 5825 9676
rect 5859 9673 5871 9707
rect 10502 9704 10508 9716
rect 10463 9676 10508 9704
rect 5813 9667 5871 9673
rect 10502 9664 10508 9676
rect 10560 9664 10566 9716
rect 11425 9707 11483 9713
rect 11425 9673 11437 9707
rect 11471 9704 11483 9707
rect 11790 9704 11796 9716
rect 11471 9676 11796 9704
rect 11471 9673 11483 9676
rect 11425 9667 11483 9673
rect 11790 9664 11796 9676
rect 11848 9664 11854 9716
rect 15286 9704 15292 9716
rect 15247 9676 15292 9704
rect 15286 9664 15292 9676
rect 15344 9664 15350 9716
rect 16485 9707 16543 9713
rect 16485 9673 16497 9707
rect 16531 9704 16543 9707
rect 17402 9704 17408 9716
rect 16531 9676 17408 9704
rect 16531 9673 16543 9676
rect 16485 9667 16543 9673
rect 17402 9664 17408 9676
rect 17460 9664 17466 9716
rect 20714 9664 20720 9716
rect 20772 9704 20778 9716
rect 20809 9707 20867 9713
rect 20809 9704 20821 9707
rect 20772 9676 20821 9704
rect 20772 9664 20778 9676
rect 20809 9673 20821 9676
rect 20855 9673 20867 9707
rect 25222 9704 25228 9716
rect 20809 9667 20867 9673
rect 24504 9676 25228 9704
rect 2038 9636 2044 9648
rect 1999 9608 2044 9636
rect 2038 9596 2044 9608
rect 2096 9596 2102 9648
rect 2958 9636 2964 9648
rect 2919 9608 2964 9636
rect 2958 9596 2964 9608
rect 3016 9596 3022 9648
rect 7009 9639 7067 9645
rect 7009 9605 7021 9639
rect 7055 9636 7067 9639
rect 7466 9636 7472 9648
rect 7055 9608 7472 9636
rect 7055 9605 7067 9608
rect 7009 9599 7067 9605
rect 7466 9596 7472 9608
rect 7524 9596 7530 9648
rect 9582 9596 9588 9648
rect 9640 9636 9646 9648
rect 9861 9639 9919 9645
rect 9861 9636 9873 9639
rect 9640 9608 9873 9636
rect 9640 9596 9646 9608
rect 9861 9605 9873 9608
rect 9907 9605 9919 9639
rect 9861 9599 9919 9605
rect 10873 9639 10931 9645
rect 10873 9605 10885 9639
rect 10919 9636 10931 9639
rect 11514 9636 11520 9648
rect 10919 9608 11520 9636
rect 10919 9605 10931 9608
rect 10873 9599 10931 9605
rect 11514 9596 11520 9608
rect 11572 9596 11578 9648
rect 2406 9568 2412 9580
rect 2367 9540 2412 9568
rect 2406 9528 2412 9540
rect 2464 9568 2470 9580
rect 2682 9568 2688 9580
rect 2464 9540 2688 9568
rect 2464 9528 2470 9540
rect 2682 9528 2688 9540
rect 2740 9528 2746 9580
rect 4522 9528 4528 9580
rect 4580 9568 4586 9580
rect 7374 9568 7380 9580
rect 4580 9540 7380 9568
rect 4580 9528 4586 9540
rect 7374 9528 7380 9540
rect 7432 9528 7438 9580
rect 7561 9571 7619 9577
rect 7561 9537 7573 9571
rect 7607 9568 7619 9571
rect 17034 9568 17040 9580
rect 7607 9540 8616 9568
rect 16995 9540 17040 9568
rect 7607 9537 7619 9540
rect 7561 9531 7619 9537
rect 1857 9503 1915 9509
rect 1857 9469 1869 9503
rect 1903 9500 1915 9503
rect 2593 9503 2651 9509
rect 2593 9500 2605 9503
rect 1903 9472 2605 9500
rect 1903 9469 1915 9472
rect 1857 9463 1915 9469
rect 2593 9469 2605 9472
rect 2639 9500 2651 9503
rect 3418 9500 3424 9512
rect 2639 9472 3424 9500
rect 2639 9469 2651 9472
rect 2593 9463 2651 9469
rect 3418 9460 3424 9472
rect 3476 9460 3482 9512
rect 3513 9503 3571 9509
rect 3513 9469 3525 9503
rect 3559 9500 3571 9503
rect 3602 9500 3608 9512
rect 3559 9472 3608 9500
rect 3559 9469 3571 9472
rect 3513 9463 3571 9469
rect 2498 9432 2504 9444
rect 2459 9404 2504 9432
rect 2498 9392 2504 9404
rect 2556 9392 2562 9444
rect 3329 9435 3387 9441
rect 3329 9401 3341 9435
rect 3375 9432 3387 9435
rect 3528 9432 3556 9463
rect 3602 9460 3608 9472
rect 3660 9460 3666 9512
rect 5350 9460 5356 9512
rect 5408 9500 5414 9512
rect 5537 9503 5595 9509
rect 5537 9500 5549 9503
rect 5408 9472 5549 9500
rect 5408 9460 5414 9472
rect 5537 9469 5549 9472
rect 5583 9500 5595 9503
rect 8481 9503 8539 9509
rect 8481 9500 8493 9503
rect 5583 9472 8493 9500
rect 5583 9469 5595 9472
rect 5537 9463 5595 9469
rect 8481 9469 8493 9472
rect 8527 9469 8539 9503
rect 8588 9500 8616 9540
rect 17034 9528 17040 9540
rect 17092 9528 17098 9580
rect 17126 9528 17132 9580
rect 17184 9568 17190 9580
rect 17865 9571 17923 9577
rect 17865 9568 17877 9571
rect 17184 9540 17877 9568
rect 17184 9528 17190 9540
rect 17865 9537 17877 9540
rect 17911 9568 17923 9571
rect 17911 9540 18644 9568
rect 17911 9537 17923 9540
rect 17865 9531 17923 9537
rect 8748 9503 8806 9509
rect 8748 9500 8760 9503
rect 8588 9472 8760 9500
rect 8481 9463 8539 9469
rect 8748 9469 8760 9472
rect 8794 9500 8806 9503
rect 9122 9500 9128 9512
rect 8794 9472 9128 9500
rect 8794 9469 8806 9472
rect 8748 9463 8806 9469
rect 3375 9404 3556 9432
rect 3375 9401 3387 9404
rect 3329 9395 3387 9401
rect 2590 9324 2596 9376
rect 2648 9364 2654 9376
rect 3344 9364 3372 9395
rect 3694 9392 3700 9444
rect 3752 9441 3758 9444
rect 3752 9435 3816 9441
rect 3752 9401 3770 9435
rect 3804 9401 3816 9435
rect 3752 9395 3816 9401
rect 3752 9392 3758 9395
rect 6086 9392 6092 9444
rect 6144 9432 6150 9444
rect 6273 9435 6331 9441
rect 6273 9432 6285 9435
rect 6144 9404 6285 9432
rect 6144 9392 6150 9404
rect 6273 9401 6285 9404
rect 6319 9432 6331 9435
rect 7282 9432 7288 9444
rect 6319 9404 7288 9432
rect 6319 9401 6331 9404
rect 6273 9395 6331 9401
rect 7282 9392 7288 9404
rect 7340 9392 7346 9444
rect 8496 9432 8524 9463
rect 9122 9460 9128 9472
rect 9180 9460 9186 9512
rect 12710 9460 12716 9512
rect 12768 9500 12774 9512
rect 12805 9503 12863 9509
rect 12805 9500 12817 9503
rect 12768 9472 12817 9500
rect 12768 9460 12774 9472
rect 12805 9469 12817 9472
rect 12851 9500 12863 9503
rect 13173 9503 13231 9509
rect 13173 9500 13185 9503
rect 12851 9472 13185 9500
rect 12851 9469 12863 9472
rect 12805 9463 12863 9469
rect 13173 9469 13185 9472
rect 13219 9500 13231 9503
rect 13265 9503 13323 9509
rect 13265 9500 13277 9503
rect 13219 9472 13277 9500
rect 13219 9469 13231 9472
rect 13173 9463 13231 9469
rect 13265 9469 13277 9472
rect 13311 9500 13323 9503
rect 18509 9503 18567 9509
rect 18509 9500 18521 9503
rect 13311 9472 13768 9500
rect 13311 9469 13323 9472
rect 13265 9463 13323 9469
rect 13740 9444 13768 9472
rect 18340 9472 18521 9500
rect 8662 9432 8668 9444
rect 8496 9404 8668 9432
rect 8662 9392 8668 9404
rect 8720 9392 8726 9444
rect 13446 9392 13452 9444
rect 13504 9441 13510 9444
rect 13504 9435 13568 9441
rect 13504 9401 13522 9435
rect 13556 9401 13568 9435
rect 13504 9395 13568 9401
rect 13504 9392 13510 9395
rect 13722 9392 13728 9444
rect 13780 9392 13786 9444
rect 16574 9392 16580 9444
rect 16632 9432 16638 9444
rect 16761 9435 16819 9441
rect 16761 9432 16773 9435
rect 16632 9404 16773 9432
rect 16632 9392 16638 9404
rect 16761 9401 16773 9404
rect 16807 9401 16819 9435
rect 16761 9395 16819 9401
rect 2648 9336 3372 9364
rect 2648 9324 2654 9336
rect 4246 9324 4252 9376
rect 4304 9364 4310 9376
rect 4893 9367 4951 9373
rect 4893 9364 4905 9367
rect 4304 9336 4905 9364
rect 4304 9324 4310 9336
rect 4893 9333 4905 9336
rect 4939 9333 4951 9367
rect 4893 9327 4951 9333
rect 5902 9324 5908 9376
rect 5960 9364 5966 9376
rect 6549 9367 6607 9373
rect 6549 9364 6561 9367
rect 5960 9336 6561 9364
rect 5960 9324 5966 9336
rect 6549 9333 6561 9336
rect 6595 9364 6607 9367
rect 7469 9367 7527 9373
rect 7469 9364 7481 9367
rect 6595 9336 7481 9364
rect 6595 9333 6607 9336
rect 6549 9327 6607 9333
rect 7469 9333 7481 9336
rect 7515 9333 7527 9367
rect 7469 9327 7527 9333
rect 7926 9324 7932 9376
rect 7984 9364 7990 9376
rect 8021 9367 8079 9373
rect 8021 9364 8033 9367
rect 7984 9336 8033 9364
rect 7984 9324 7990 9336
rect 8021 9333 8033 9336
rect 8067 9364 8079 9367
rect 8294 9364 8300 9376
rect 8067 9336 8300 9364
rect 8067 9333 8079 9336
rect 8021 9327 8079 9333
rect 8294 9324 8300 9336
rect 8352 9324 8358 9376
rect 10778 9324 10784 9376
rect 10836 9364 10842 9376
rect 10965 9367 11023 9373
rect 10965 9364 10977 9367
rect 10836 9336 10977 9364
rect 10836 9324 10842 9336
rect 10965 9333 10977 9336
rect 11011 9333 11023 9367
rect 10965 9327 11023 9333
rect 11698 9324 11704 9376
rect 11756 9364 11762 9376
rect 11885 9367 11943 9373
rect 11885 9364 11897 9367
rect 11756 9336 11897 9364
rect 11756 9324 11762 9336
rect 11885 9333 11897 9336
rect 11931 9364 11943 9367
rect 11974 9364 11980 9376
rect 11931 9336 11980 9364
rect 11931 9333 11943 9336
rect 11885 9327 11943 9333
rect 11974 9324 11980 9336
rect 12032 9324 12038 9376
rect 12158 9364 12164 9376
rect 12119 9336 12164 9364
rect 12158 9324 12164 9336
rect 12216 9324 12222 9376
rect 13354 9324 13360 9376
rect 13412 9364 13418 9376
rect 14645 9367 14703 9373
rect 14645 9364 14657 9367
rect 13412 9336 14657 9364
rect 13412 9324 13418 9336
rect 14645 9333 14657 9336
rect 14691 9364 14703 9367
rect 14918 9364 14924 9376
rect 14691 9336 14924 9364
rect 14691 9333 14703 9336
rect 14645 9327 14703 9333
rect 14918 9324 14924 9336
rect 14976 9324 14982 9376
rect 15654 9364 15660 9376
rect 15615 9336 15660 9364
rect 15654 9324 15660 9336
rect 15712 9324 15718 9376
rect 16301 9367 16359 9373
rect 16301 9333 16313 9367
rect 16347 9364 16359 9367
rect 16945 9367 17003 9373
rect 16945 9364 16957 9367
rect 16347 9336 16957 9364
rect 16347 9333 16359 9336
rect 16301 9327 16359 9333
rect 16945 9333 16957 9336
rect 16991 9364 17003 9367
rect 17310 9364 17316 9376
rect 16991 9336 17316 9364
rect 16991 9333 17003 9336
rect 16945 9327 17003 9333
rect 17310 9324 17316 9336
rect 17368 9324 17374 9376
rect 17497 9367 17555 9373
rect 17497 9333 17509 9367
rect 17543 9364 17555 9367
rect 17678 9364 17684 9376
rect 17543 9336 17684 9364
rect 17543 9333 17555 9336
rect 17497 9327 17555 9333
rect 17678 9324 17684 9336
rect 17736 9364 17742 9376
rect 18340 9373 18368 9472
rect 18509 9469 18521 9472
rect 18555 9469 18567 9503
rect 18616 9500 18644 9540
rect 18776 9503 18834 9509
rect 18776 9500 18788 9503
rect 18616 9472 18788 9500
rect 18509 9463 18567 9469
rect 18776 9469 18788 9472
rect 18822 9500 18834 9503
rect 19058 9500 19064 9512
rect 18822 9472 19064 9500
rect 18822 9469 18834 9472
rect 18776 9463 18834 9469
rect 19058 9460 19064 9472
rect 19116 9460 19122 9512
rect 20824 9500 20852 9667
rect 24026 9636 24032 9648
rect 23939 9608 24032 9636
rect 24026 9596 24032 9608
rect 24084 9636 24090 9648
rect 24504 9636 24532 9676
rect 25222 9664 25228 9676
rect 25280 9664 25286 9716
rect 25866 9704 25872 9716
rect 25827 9676 25872 9704
rect 25866 9664 25872 9676
rect 25924 9664 25930 9716
rect 26789 9707 26847 9713
rect 26789 9673 26801 9707
rect 26835 9704 26847 9707
rect 27338 9704 27344 9716
rect 26835 9676 27344 9704
rect 26835 9673 26847 9676
rect 26789 9667 26847 9673
rect 27338 9664 27344 9676
rect 27396 9664 27402 9716
rect 29086 9664 29092 9716
rect 29144 9704 29150 9716
rect 30282 9704 30288 9716
rect 29144 9676 30288 9704
rect 29144 9664 29150 9676
rect 30282 9664 30288 9676
rect 30340 9664 30346 9716
rect 30742 9704 30748 9716
rect 30392 9676 30748 9704
rect 24084 9608 24532 9636
rect 24084 9596 24090 9608
rect 26050 9596 26056 9648
rect 26108 9636 26114 9648
rect 27525 9639 27583 9645
rect 27525 9636 27537 9639
rect 26108 9608 27537 9636
rect 26108 9596 26114 9608
rect 27525 9605 27537 9608
rect 27571 9605 27583 9639
rect 29822 9636 29828 9648
rect 29783 9608 29828 9636
rect 27525 9599 27583 9605
rect 29822 9596 29828 9608
rect 29880 9596 29886 9648
rect 30392 9636 30420 9676
rect 30742 9664 30748 9676
rect 30800 9664 30806 9716
rect 34977 9707 35035 9713
rect 34977 9673 34989 9707
rect 35023 9704 35035 9707
rect 35618 9704 35624 9716
rect 35023 9676 35624 9704
rect 35023 9673 35035 9676
rect 34977 9667 35035 9673
rect 35618 9664 35624 9676
rect 35676 9664 35682 9716
rect 30300 9608 30420 9636
rect 33321 9639 33379 9645
rect 22370 9528 22376 9580
rect 22428 9568 22434 9580
rect 23293 9571 23351 9577
rect 23293 9568 23305 9571
rect 22428 9540 23305 9568
rect 22428 9528 22434 9540
rect 23293 9537 23305 9540
rect 23339 9537 23351 9571
rect 23293 9531 23351 9537
rect 27985 9571 28043 9577
rect 27985 9537 27997 9571
rect 28031 9568 28043 9571
rect 28902 9568 28908 9580
rect 28031 9540 28908 9568
rect 28031 9537 28043 9540
rect 27985 9531 28043 9537
rect 28902 9528 28908 9540
rect 28960 9528 28966 9580
rect 29549 9571 29607 9577
rect 29549 9537 29561 9571
rect 29595 9568 29607 9571
rect 30300 9568 30328 9608
rect 33321 9605 33333 9639
rect 33367 9636 33379 9639
rect 35802 9636 35808 9648
rect 33367 9608 35808 9636
rect 33367 9605 33379 9608
rect 33321 9599 33379 9605
rect 35802 9596 35808 9608
rect 35860 9596 35866 9648
rect 36262 9636 36268 9648
rect 36223 9608 36268 9636
rect 36262 9596 36268 9608
rect 36320 9596 36326 9648
rect 36538 9636 36544 9648
rect 36499 9608 36544 9636
rect 36538 9596 36544 9608
rect 36596 9596 36602 9648
rect 29595 9540 30328 9568
rect 29595 9537 29607 9540
rect 29549 9531 29607 9537
rect 30374 9528 30380 9580
rect 30432 9568 30438 9580
rect 30561 9571 30619 9577
rect 30561 9568 30573 9571
rect 30432 9540 30573 9568
rect 30432 9528 30438 9540
rect 30561 9537 30573 9540
rect 30607 9568 30619 9571
rect 30745 9571 30803 9577
rect 30745 9568 30757 9571
rect 30607 9540 30757 9568
rect 30607 9537 30619 9540
rect 30561 9531 30619 9537
rect 30745 9537 30757 9540
rect 30791 9537 30803 9571
rect 35526 9568 35532 9580
rect 35439 9540 35532 9568
rect 30745 9531 30803 9537
rect 20993 9503 21051 9509
rect 20993 9500 21005 9503
rect 20824 9472 21005 9500
rect 20993 9469 21005 9472
rect 21039 9500 21051 9503
rect 21634 9500 21640 9512
rect 21039 9472 21640 9500
rect 21039 9469 21051 9472
rect 20993 9463 21051 9469
rect 21634 9460 21640 9472
rect 21692 9500 21698 9512
rect 22925 9503 22983 9509
rect 22925 9500 22937 9503
rect 21692 9472 22937 9500
rect 21692 9460 21698 9472
rect 22925 9469 22937 9472
rect 22971 9500 22983 9503
rect 23382 9500 23388 9512
rect 22971 9472 23388 9500
rect 22971 9469 22983 9472
rect 22925 9463 22983 9469
rect 23382 9460 23388 9472
rect 23440 9500 23446 9512
rect 24486 9500 24492 9512
rect 23440 9472 24492 9500
rect 23440 9460 23446 9472
rect 24486 9460 24492 9472
rect 24544 9500 24550 9512
rect 27062 9500 27068 9512
rect 24544 9472 27068 9500
rect 24544 9460 24550 9472
rect 27062 9460 27068 9472
rect 27120 9460 27126 9512
rect 29641 9503 29699 9509
rect 29641 9469 29653 9503
rect 29687 9500 29699 9503
rect 30760 9500 30788 9531
rect 35526 9528 35532 9540
rect 35584 9568 35590 9580
rect 37461 9571 37519 9577
rect 37461 9568 37473 9571
rect 35584 9540 37473 9568
rect 35584 9528 35590 9540
rect 37461 9537 37473 9540
rect 37507 9537 37519 9571
rect 37461 9531 37519 9537
rect 37093 9503 37151 9509
rect 37093 9500 37105 9503
rect 29687 9472 30328 9500
rect 30760 9472 32812 9500
rect 29687 9469 29699 9472
rect 29641 9463 29699 9469
rect 21238 9435 21296 9441
rect 21238 9432 21250 9435
rect 20456 9404 21250 9432
rect 18325 9367 18383 9373
rect 18325 9364 18337 9367
rect 17736 9336 18337 9364
rect 17736 9324 17742 9336
rect 18325 9333 18337 9336
rect 18371 9333 18383 9367
rect 18325 9327 18383 9333
rect 19889 9367 19947 9373
rect 19889 9333 19901 9367
rect 19935 9364 19947 9367
rect 19978 9364 19984 9376
rect 19935 9336 19984 9364
rect 19935 9333 19947 9336
rect 19889 9327 19947 9333
rect 19978 9324 19984 9336
rect 20036 9324 20042 9376
rect 20162 9324 20168 9376
rect 20220 9364 20226 9376
rect 20456 9373 20484 9404
rect 21238 9401 21250 9404
rect 21284 9432 21296 9435
rect 23014 9432 23020 9444
rect 21284 9404 23020 9432
rect 21284 9401 21296 9404
rect 21238 9395 21296 9401
rect 23014 9392 23020 9404
rect 23072 9392 23078 9444
rect 24756 9435 24814 9441
rect 24756 9401 24768 9435
rect 24802 9432 24814 9435
rect 25406 9432 25412 9444
rect 24802 9404 25412 9432
rect 24802 9401 24814 9404
rect 24756 9395 24814 9401
rect 25406 9392 25412 9404
rect 25464 9392 25470 9444
rect 28077 9435 28135 9441
rect 28077 9401 28089 9435
rect 28123 9432 28135 9435
rect 28166 9432 28172 9444
rect 28123 9404 28172 9432
rect 28123 9401 28135 9404
rect 28077 9395 28135 9401
rect 28166 9392 28172 9404
rect 28224 9392 28230 9444
rect 30300 9376 30328 9472
rect 31018 9441 31024 9444
rect 31012 9432 31024 9441
rect 30979 9404 31024 9432
rect 31012 9395 31024 9404
rect 31018 9392 31024 9395
rect 31076 9392 31082 9444
rect 20441 9367 20499 9373
rect 20441 9364 20453 9367
rect 20220 9336 20453 9364
rect 20220 9324 20226 9336
rect 20441 9333 20453 9336
rect 20487 9333 20499 9367
rect 22370 9364 22376 9376
rect 22331 9336 22376 9364
rect 20441 9327 20499 9333
rect 22370 9324 22376 9336
rect 22428 9324 22434 9376
rect 24118 9324 24124 9376
rect 24176 9364 24182 9376
rect 24305 9367 24363 9373
rect 24305 9364 24317 9367
rect 24176 9336 24317 9364
rect 24176 9324 24182 9336
rect 24305 9333 24317 9336
rect 24351 9364 24363 9367
rect 24394 9364 24400 9376
rect 24351 9336 24400 9364
rect 24351 9333 24363 9336
rect 24305 9327 24363 9333
rect 24394 9324 24400 9336
rect 24452 9324 24458 9376
rect 27985 9367 28043 9373
rect 27985 9333 27997 9367
rect 28031 9364 28043 9367
rect 28534 9364 28540 9376
rect 28031 9336 28540 9364
rect 28031 9333 28043 9336
rect 27985 9327 28043 9333
rect 28534 9324 28540 9336
rect 28592 9324 28598 9376
rect 28902 9364 28908 9376
rect 28863 9336 28908 9364
rect 28902 9324 28908 9336
rect 28960 9324 28966 9376
rect 30282 9364 30288 9376
rect 30243 9336 30288 9364
rect 30282 9324 30288 9336
rect 30340 9324 30346 9376
rect 31662 9324 31668 9376
rect 31720 9364 31726 9376
rect 31938 9364 31944 9376
rect 31720 9336 31944 9364
rect 31720 9324 31726 9336
rect 31938 9324 31944 9336
rect 31996 9364 32002 9376
rect 32784 9373 32812 9472
rect 35912 9472 37105 9500
rect 33597 9435 33655 9441
rect 33597 9401 33609 9435
rect 33643 9432 33655 9435
rect 33686 9432 33692 9444
rect 33643 9404 33692 9432
rect 33643 9401 33655 9404
rect 33597 9395 33655 9401
rect 33686 9392 33692 9404
rect 33744 9392 33750 9444
rect 33870 9432 33876 9444
rect 33831 9404 33876 9432
rect 33870 9392 33876 9404
rect 33928 9392 33934 9444
rect 34333 9435 34391 9441
rect 34333 9401 34345 9435
rect 34379 9432 34391 9435
rect 34698 9432 34704 9444
rect 34379 9404 34704 9432
rect 34379 9401 34391 9404
rect 34333 9395 34391 9401
rect 34698 9392 34704 9404
rect 34756 9392 34762 9444
rect 34882 9392 34888 9444
rect 34940 9432 34946 9444
rect 35253 9435 35311 9441
rect 35253 9432 35265 9435
rect 34940 9404 35265 9432
rect 34940 9392 34946 9404
rect 35253 9401 35265 9404
rect 35299 9401 35311 9435
rect 35253 9395 35311 9401
rect 35912 9376 35940 9472
rect 37093 9469 37105 9472
rect 37139 9469 37151 9503
rect 37093 9463 37151 9469
rect 36262 9392 36268 9444
rect 36320 9432 36326 9444
rect 36817 9435 36875 9441
rect 36817 9432 36829 9435
rect 36320 9404 36829 9432
rect 36320 9392 36326 9404
rect 36817 9401 36829 9404
rect 36863 9401 36875 9435
rect 36817 9395 36875 9401
rect 32125 9367 32183 9373
rect 32125 9364 32137 9367
rect 31996 9336 32137 9364
rect 31996 9324 32002 9336
rect 32125 9333 32137 9336
rect 32171 9333 32183 9367
rect 32125 9327 32183 9333
rect 32769 9367 32827 9373
rect 32769 9333 32781 9367
rect 32815 9364 32827 9367
rect 32950 9364 32956 9376
rect 32815 9336 32956 9364
rect 32815 9333 32827 9336
rect 32769 9327 32827 9333
rect 32950 9324 32956 9336
rect 33008 9324 33014 9376
rect 33134 9364 33140 9376
rect 33095 9336 33140 9364
rect 33134 9324 33140 9336
rect 33192 9364 33198 9376
rect 33781 9367 33839 9373
rect 33781 9364 33793 9367
rect 33192 9336 33793 9364
rect 33192 9324 33198 9336
rect 33781 9333 33793 9336
rect 33827 9333 33839 9367
rect 34606 9364 34612 9376
rect 34567 9336 34612 9364
rect 33781 9327 33839 9333
rect 34606 9324 34612 9336
rect 34664 9364 34670 9376
rect 35437 9367 35495 9373
rect 35437 9364 35449 9367
rect 34664 9336 35449 9364
rect 34664 9324 34670 9336
rect 35437 9333 35449 9336
rect 35483 9333 35495 9367
rect 35894 9364 35900 9376
rect 35855 9336 35900 9364
rect 35437 9327 35495 9333
rect 35894 9324 35900 9336
rect 35952 9324 35958 9376
rect 36998 9364 37004 9376
rect 36959 9336 37004 9364
rect 36998 9324 37004 9336
rect 37056 9324 37062 9376
rect 1104 9274 38824 9296
rect 1104 9222 14315 9274
rect 14367 9222 14379 9274
rect 14431 9222 14443 9274
rect 14495 9222 14507 9274
rect 14559 9222 27648 9274
rect 27700 9222 27712 9274
rect 27764 9222 27776 9274
rect 27828 9222 27840 9274
rect 27892 9222 38824 9274
rect 1104 9200 38824 9222
rect 1670 9160 1676 9172
rect 1631 9132 1676 9160
rect 1670 9120 1676 9132
rect 1728 9120 1734 9172
rect 1946 9160 1952 9172
rect 1907 9132 1952 9160
rect 1946 9120 1952 9132
rect 2004 9120 2010 9172
rect 2777 9163 2835 9169
rect 2777 9129 2789 9163
rect 2823 9160 2835 9163
rect 5074 9160 5080 9172
rect 2823 9132 5080 9160
rect 2823 9129 2835 9132
rect 2777 9123 2835 9129
rect 5074 9120 5080 9132
rect 5132 9120 5138 9172
rect 7282 9120 7288 9172
rect 7340 9160 7346 9172
rect 7926 9160 7932 9172
rect 7340 9132 7932 9160
rect 7340 9120 7346 9132
rect 7926 9120 7932 9132
rect 7984 9120 7990 9172
rect 8754 9120 8760 9172
rect 8812 9160 8818 9172
rect 9033 9163 9091 9169
rect 9033 9160 9045 9163
rect 8812 9132 9045 9160
rect 8812 9120 8818 9132
rect 9033 9129 9045 9132
rect 9079 9129 9091 9163
rect 9033 9123 9091 9129
rect 13446 9120 13452 9172
rect 13504 9160 13510 9172
rect 13725 9163 13783 9169
rect 13725 9160 13737 9163
rect 13504 9132 13737 9160
rect 13504 9120 13510 9132
rect 13725 9129 13737 9132
rect 13771 9160 13783 9163
rect 13998 9160 14004 9172
rect 13771 9132 14004 9160
rect 13771 9129 13783 9132
rect 13725 9123 13783 9129
rect 13998 9120 14004 9132
rect 14056 9120 14062 9172
rect 14918 9120 14924 9172
rect 14976 9160 14982 9172
rect 15013 9163 15071 9169
rect 15013 9160 15025 9163
rect 14976 9132 15025 9160
rect 14976 9120 14982 9132
rect 15013 9129 15025 9132
rect 15059 9160 15071 9163
rect 15059 9132 15516 9160
rect 15059 9129 15071 9132
rect 15013 9123 15071 9129
rect 5353 9095 5411 9101
rect 5353 9061 5365 9095
rect 5399 9092 5411 9095
rect 5442 9092 5448 9104
rect 5399 9064 5448 9092
rect 5399 9061 5411 9064
rect 5353 9055 5411 9061
rect 5442 9052 5448 9064
rect 5500 9052 5506 9104
rect 6638 9052 6644 9104
rect 6696 9092 6702 9104
rect 6917 9095 6975 9101
rect 6917 9092 6929 9095
rect 6696 9064 6929 9092
rect 6696 9052 6702 9064
rect 6917 9061 6929 9064
rect 6963 9061 6975 9095
rect 7374 9092 7380 9104
rect 7335 9064 7380 9092
rect 6917 9055 6975 9061
rect 1670 8984 1676 9036
rect 1728 9024 1734 9036
rect 2593 9027 2651 9033
rect 2593 9024 2605 9027
rect 1728 8996 2605 9024
rect 1728 8984 1734 8996
rect 2593 8993 2605 8996
rect 2639 9024 2651 9027
rect 2682 9024 2688 9036
rect 2639 8996 2688 9024
rect 2639 8993 2651 8996
rect 2593 8987 2651 8993
rect 2682 8984 2688 8996
rect 2740 8984 2746 9036
rect 3605 9027 3663 9033
rect 3605 8993 3617 9027
rect 3651 9024 3663 9027
rect 3694 9024 3700 9036
rect 3651 8996 3700 9024
rect 3651 8993 3663 8996
rect 3605 8987 3663 8993
rect 3694 8984 3700 8996
rect 3752 9024 3758 9036
rect 5258 9024 5264 9036
rect 3752 8996 5264 9024
rect 3752 8984 3758 8996
rect 5258 8984 5264 8996
rect 5316 9024 5322 9036
rect 5316 8996 5488 9024
rect 5316 8984 5322 8996
rect 2866 8956 2872 8968
rect 2827 8928 2872 8956
rect 2866 8916 2872 8928
rect 2924 8916 2930 8968
rect 4709 8959 4767 8965
rect 4709 8925 4721 8959
rect 4755 8956 4767 8959
rect 5350 8956 5356 8968
rect 4755 8928 5356 8956
rect 4755 8925 4767 8928
rect 4709 8919 4767 8925
rect 5350 8916 5356 8928
rect 5408 8916 5414 8968
rect 5460 8965 5488 8996
rect 6362 8984 6368 9036
rect 6420 9024 6426 9036
rect 6733 9027 6791 9033
rect 6733 9024 6745 9027
rect 6420 8996 6745 9024
rect 6420 8984 6426 8996
rect 6733 8993 6745 8996
rect 6779 8993 6791 9027
rect 6932 9024 6960 9055
rect 7374 9052 7380 9064
rect 7432 9052 7438 9104
rect 8110 9052 8116 9104
rect 8168 9092 8174 9104
rect 8573 9095 8631 9101
rect 8573 9092 8585 9095
rect 8168 9064 8585 9092
rect 8168 9052 8174 9064
rect 8573 9061 8585 9064
rect 8619 9061 8631 9095
rect 8573 9055 8631 9061
rect 8662 9052 8668 9104
rect 8720 9092 8726 9104
rect 9122 9092 9128 9104
rect 8720 9064 9128 9092
rect 8720 9052 8726 9064
rect 9122 9052 9128 9064
rect 9180 9052 9186 9104
rect 10226 9052 10232 9104
rect 10284 9092 10290 9104
rect 11698 9092 11704 9104
rect 10284 9064 11704 9092
rect 10284 9052 10290 9064
rect 11698 9052 11704 9064
rect 11756 9052 11762 9104
rect 12621 9095 12679 9101
rect 12621 9061 12633 9095
rect 12667 9092 12679 9095
rect 13265 9095 13323 9101
rect 13265 9092 13277 9095
rect 12667 9064 13277 9092
rect 12667 9061 12679 9064
rect 12621 9055 12679 9061
rect 13265 9061 13277 9064
rect 13311 9092 13323 9095
rect 15363 9095 15421 9101
rect 15363 9092 15375 9095
rect 13311 9064 15375 9092
rect 13311 9061 13323 9064
rect 13265 9055 13323 9061
rect 15363 9061 15375 9064
rect 15409 9061 15421 9095
rect 15363 9055 15421 9061
rect 7837 9027 7895 9033
rect 7837 9024 7849 9027
rect 6932 8996 7849 9024
rect 6733 8987 6791 8993
rect 7837 8993 7849 8996
rect 7883 9024 7895 9027
rect 8478 9024 8484 9036
rect 7883 8996 8484 9024
rect 7883 8993 7895 8996
rect 7837 8987 7895 8993
rect 8478 8984 8484 8996
rect 8536 8984 8542 9036
rect 10505 9027 10563 9033
rect 10505 8993 10517 9027
rect 10551 9024 10563 9027
rect 11793 9027 11851 9033
rect 11793 9024 11805 9027
rect 10551 8996 11805 9024
rect 10551 8993 10563 8996
rect 10505 8987 10563 8993
rect 11793 8993 11805 8996
rect 11839 9024 11851 9027
rect 12158 9024 12164 9036
rect 11839 8996 12164 9024
rect 11839 8993 11851 8996
rect 11793 8987 11851 8993
rect 12158 8984 12164 8996
rect 12216 8984 12222 9036
rect 15488 9024 15516 9132
rect 17034 9120 17040 9172
rect 17092 9160 17098 9172
rect 17129 9163 17187 9169
rect 17129 9160 17141 9163
rect 17092 9132 17141 9160
rect 17092 9120 17098 9132
rect 17129 9129 17141 9132
rect 17175 9129 17187 9163
rect 18046 9160 18052 9172
rect 18007 9132 18052 9160
rect 17129 9123 17187 9129
rect 18046 9120 18052 9132
rect 18104 9120 18110 9172
rect 19518 9120 19524 9172
rect 19576 9160 19582 9172
rect 19797 9163 19855 9169
rect 19797 9160 19809 9163
rect 19576 9132 19809 9160
rect 19576 9120 19582 9132
rect 19797 9129 19809 9132
rect 19843 9129 19855 9163
rect 23014 9160 23020 9172
rect 22975 9132 23020 9160
rect 19797 9123 19855 9129
rect 23014 9120 23020 9132
rect 23072 9120 23078 9172
rect 23474 9120 23480 9172
rect 23532 9160 23538 9172
rect 24213 9163 24271 9169
rect 24213 9160 24225 9163
rect 23532 9132 24225 9160
rect 23532 9120 23538 9132
rect 24213 9129 24225 9132
rect 24259 9160 24271 9163
rect 25406 9160 25412 9172
rect 24259 9132 25412 9160
rect 24259 9129 24271 9132
rect 24213 9123 24271 9129
rect 25406 9120 25412 9132
rect 25464 9120 25470 9172
rect 31573 9163 31631 9169
rect 31573 9129 31585 9163
rect 31619 9160 31631 9163
rect 32677 9163 32735 9169
rect 32677 9160 32689 9163
rect 31619 9132 32689 9160
rect 31619 9129 31631 9132
rect 31573 9123 31631 9129
rect 32677 9129 32689 9132
rect 32723 9160 32735 9163
rect 35327 9163 35385 9169
rect 35327 9160 35339 9163
rect 32723 9132 35339 9160
rect 32723 9129 32735 9132
rect 32677 9123 32735 9129
rect 35327 9129 35339 9132
rect 35373 9129 35385 9163
rect 35802 9160 35808 9172
rect 35763 9132 35808 9160
rect 35327 9123 35385 9129
rect 35802 9120 35808 9132
rect 35860 9120 35866 9172
rect 15746 9052 15752 9104
rect 15804 9092 15810 9104
rect 15841 9095 15899 9101
rect 15841 9092 15853 9095
rect 15804 9064 15853 9092
rect 15804 9052 15810 9064
rect 15841 9061 15853 9064
rect 15887 9061 15899 9095
rect 19886 9092 19892 9104
rect 19847 9064 19892 9092
rect 15841 9055 15899 9061
rect 19886 9052 19892 9064
rect 19944 9052 19950 9104
rect 21910 9101 21916 9104
rect 21904 9092 21916 9101
rect 21871 9064 21916 9092
rect 21904 9055 21916 9064
rect 21910 9052 21916 9055
rect 21968 9052 21974 9104
rect 24857 9095 24915 9101
rect 24857 9061 24869 9095
rect 24903 9092 24915 9095
rect 24946 9092 24952 9104
rect 24903 9064 24952 9092
rect 24903 9061 24915 9064
rect 24857 9055 24915 9061
rect 24946 9052 24952 9064
rect 25004 9052 25010 9104
rect 26970 9092 26976 9104
rect 26931 9064 26976 9092
rect 26970 9052 26976 9064
rect 27028 9052 27034 9104
rect 27525 9095 27583 9101
rect 27525 9061 27537 9095
rect 27571 9092 27583 9095
rect 27706 9092 27712 9104
rect 27571 9064 27712 9092
rect 27571 9061 27583 9064
rect 27525 9055 27583 9061
rect 27706 9052 27712 9064
rect 27764 9092 27770 9104
rect 28252 9095 28310 9101
rect 28252 9092 28264 9095
rect 27764 9064 28264 9092
rect 27764 9052 27770 9064
rect 28252 9061 28264 9064
rect 28298 9092 28310 9095
rect 28442 9092 28448 9104
rect 28298 9064 28448 9092
rect 28298 9061 28310 9064
rect 28252 9055 28310 9061
rect 28442 9052 28448 9064
rect 28500 9052 28506 9104
rect 30742 9052 30748 9104
rect 30800 9092 30806 9104
rect 31021 9095 31079 9101
rect 31021 9092 31033 9095
rect 30800 9064 31033 9092
rect 30800 9052 30806 9064
rect 31021 9061 31033 9064
rect 31067 9061 31079 9095
rect 31846 9092 31852 9104
rect 31807 9064 31852 9092
rect 31021 9055 31079 9061
rect 31846 9052 31852 9064
rect 31904 9052 31910 9104
rect 34146 9052 34152 9104
rect 34204 9092 34210 9104
rect 34241 9095 34299 9101
rect 34241 9092 34253 9095
rect 34204 9064 34253 9092
rect 34204 9052 34210 9064
rect 34241 9061 34253 9064
rect 34287 9061 34299 9095
rect 34882 9092 34888 9104
rect 34843 9064 34888 9092
rect 34241 9055 34299 9061
rect 34882 9052 34888 9064
rect 34940 9052 34946 9104
rect 15930 9024 15936 9036
rect 15488 8996 15936 9024
rect 15930 8984 15936 8996
rect 15988 8984 15994 9036
rect 24673 9027 24731 9033
rect 24673 8993 24685 9027
rect 24719 9024 24731 9027
rect 26050 9024 26056 9036
rect 24719 8996 26056 9024
rect 24719 8993 24731 8996
rect 24673 8987 24731 8993
rect 26050 8984 26056 8996
rect 26108 8984 26114 9036
rect 27062 8984 27068 9036
rect 27120 9024 27126 9036
rect 27985 9027 28043 9033
rect 27985 9024 27997 9027
rect 27120 8996 27997 9024
rect 27120 8984 27126 8996
rect 27985 8993 27997 8996
rect 28031 9024 28043 9027
rect 28074 9024 28080 9036
rect 28031 8996 28080 9024
rect 28031 8993 28043 8996
rect 27985 8987 28043 8993
rect 28074 8984 28080 8996
rect 28132 8984 28138 9036
rect 30834 9024 30840 9036
rect 30795 8996 30840 9024
rect 30834 8984 30840 8996
rect 30892 8984 30898 9036
rect 31938 8984 31944 9036
rect 31996 9024 32002 9036
rect 32769 9027 32827 9033
rect 32769 9024 32781 9027
rect 31996 8996 32781 9024
rect 31996 8984 32002 8996
rect 32769 8993 32781 8996
rect 32815 8993 32827 9027
rect 32769 8987 32827 8993
rect 33134 8984 33140 9036
rect 33192 9024 33198 9036
rect 34057 9027 34115 9033
rect 34057 9024 34069 9027
rect 33192 8996 34069 9024
rect 33192 8984 33198 8996
rect 34057 8993 34069 8996
rect 34103 8993 34115 9027
rect 35618 9024 35624 9036
rect 35579 8996 35624 9024
rect 34057 8987 34115 8993
rect 35618 8984 35624 8996
rect 35676 9024 35682 9036
rect 35986 9024 35992 9036
rect 35676 8996 35992 9024
rect 35676 8984 35682 8996
rect 35986 8984 35992 8996
rect 36044 8984 36050 9036
rect 5445 8959 5503 8965
rect 5445 8925 5457 8959
rect 5491 8925 5503 8959
rect 5445 8919 5503 8925
rect 7009 8959 7067 8965
rect 7009 8925 7021 8959
rect 7055 8925 7067 8959
rect 8570 8956 8576 8968
rect 8531 8928 8576 8956
rect 7009 8919 7067 8925
rect 2314 8888 2320 8900
rect 2275 8860 2320 8888
rect 2314 8848 2320 8860
rect 2372 8848 2378 8900
rect 4154 8848 4160 8900
rect 4212 8888 4218 8900
rect 4893 8891 4951 8897
rect 4893 8888 4905 8891
rect 4212 8860 4905 8888
rect 4212 8848 4218 8860
rect 4893 8857 4905 8860
rect 4939 8857 4951 8891
rect 4893 8851 4951 8857
rect 6273 8891 6331 8897
rect 6273 8857 6285 8891
rect 6319 8888 6331 8891
rect 6730 8888 6736 8900
rect 6319 8860 6736 8888
rect 6319 8857 6331 8860
rect 6273 8851 6331 8857
rect 6730 8848 6736 8860
rect 6788 8888 6794 8900
rect 7024 8888 7052 8919
rect 8570 8916 8576 8928
rect 8628 8916 8634 8968
rect 11606 8956 11612 8968
rect 11567 8928 11612 8956
rect 11606 8916 11612 8928
rect 11664 8916 11670 8968
rect 12253 8959 12311 8965
rect 12253 8925 12265 8959
rect 12299 8956 12311 8959
rect 13262 8956 13268 8968
rect 12299 8928 13268 8956
rect 12299 8925 12311 8928
rect 12253 8919 12311 8925
rect 13262 8916 13268 8928
rect 13320 8916 13326 8968
rect 13357 8959 13415 8965
rect 13357 8925 13369 8959
rect 13403 8956 13415 8959
rect 13538 8956 13544 8968
rect 13403 8928 13544 8956
rect 13403 8925 13415 8928
rect 13357 8919 13415 8925
rect 13538 8916 13544 8928
rect 13596 8916 13602 8968
rect 15286 8916 15292 8968
rect 15344 8956 15350 8968
rect 15749 8959 15807 8965
rect 15749 8956 15761 8959
rect 15344 8928 15761 8956
rect 15344 8916 15350 8928
rect 15749 8925 15761 8928
rect 15795 8925 15807 8959
rect 15749 8919 15807 8925
rect 17957 8959 18015 8965
rect 17957 8925 17969 8959
rect 18003 8925 18015 8959
rect 17957 8919 18015 8925
rect 6788 8860 7052 8888
rect 8113 8891 8171 8897
rect 6788 8848 6794 8860
rect 8113 8857 8125 8891
rect 8159 8888 8171 8891
rect 8202 8888 8208 8900
rect 8159 8860 8208 8888
rect 8159 8857 8171 8860
rect 8113 8851 8171 8857
rect 8202 8848 8208 8860
rect 8260 8848 8266 8900
rect 11241 8891 11299 8897
rect 11241 8857 11253 8891
rect 11287 8888 11299 8891
rect 11514 8888 11520 8900
rect 11287 8860 11520 8888
rect 11287 8857 11299 8860
rect 11241 8851 11299 8857
rect 11514 8848 11520 8860
rect 11572 8848 11578 8900
rect 12802 8888 12808 8900
rect 12763 8860 12808 8888
rect 12802 8848 12808 8860
rect 12860 8848 12866 8900
rect 17972 8888 18000 8919
rect 18046 8916 18052 8968
rect 18104 8956 18110 8968
rect 18141 8959 18199 8965
rect 18141 8956 18153 8959
rect 18104 8928 18153 8956
rect 18104 8916 18110 8928
rect 18141 8925 18153 8928
rect 18187 8956 18199 8959
rect 19794 8956 19800 8968
rect 18187 8928 19012 8956
rect 19755 8928 19800 8956
rect 18187 8925 18199 8928
rect 18141 8919 18199 8925
rect 18230 8888 18236 8900
rect 17972 8860 18236 8888
rect 18230 8848 18236 8860
rect 18288 8848 18294 8900
rect 4338 8820 4344 8832
rect 4299 8792 4344 8820
rect 4338 8780 4344 8792
rect 4396 8780 4402 8832
rect 5718 8780 5724 8832
rect 5776 8820 5782 8832
rect 5813 8823 5871 8829
rect 5813 8820 5825 8823
rect 5776 8792 5825 8820
rect 5776 8780 5782 8792
rect 5813 8789 5825 8792
rect 5859 8789 5871 8823
rect 6454 8820 6460 8832
rect 6415 8792 6460 8820
rect 5813 8783 5871 8789
rect 6454 8780 6460 8792
rect 6512 8780 6518 8832
rect 10318 8780 10324 8832
rect 10376 8820 10382 8832
rect 10781 8823 10839 8829
rect 10781 8820 10793 8823
rect 10376 8792 10793 8820
rect 10376 8780 10382 8792
rect 10781 8789 10793 8792
rect 10827 8789 10839 8823
rect 10781 8783 10839 8789
rect 12158 8780 12164 8832
rect 12216 8820 12222 8832
rect 13262 8820 13268 8832
rect 12216 8792 13268 8820
rect 12216 8780 12222 8792
rect 13262 8780 13268 8792
rect 13320 8780 13326 8832
rect 16485 8823 16543 8829
rect 16485 8789 16497 8823
rect 16531 8820 16543 8823
rect 16574 8820 16580 8832
rect 16531 8792 16580 8820
rect 16531 8789 16543 8792
rect 16485 8783 16543 8789
rect 16574 8780 16580 8792
rect 16632 8780 16638 8832
rect 16853 8823 16911 8829
rect 16853 8789 16865 8823
rect 16899 8820 16911 8823
rect 16942 8820 16948 8832
rect 16899 8792 16948 8820
rect 16899 8789 16911 8792
rect 16853 8783 16911 8789
rect 16942 8780 16948 8792
rect 17000 8780 17006 8832
rect 17589 8823 17647 8829
rect 17589 8789 17601 8823
rect 17635 8820 17647 8823
rect 17862 8820 17868 8832
rect 17635 8792 17868 8820
rect 17635 8789 17647 8792
rect 17589 8783 17647 8789
rect 17862 8780 17868 8792
rect 17920 8780 17926 8832
rect 18598 8820 18604 8832
rect 18559 8792 18604 8820
rect 18598 8780 18604 8792
rect 18656 8780 18662 8832
rect 18984 8829 19012 8928
rect 19794 8916 19800 8928
rect 19852 8916 19858 8968
rect 21634 8956 21640 8968
rect 21595 8928 21640 8956
rect 21634 8916 21640 8928
rect 21692 8916 21698 8968
rect 24949 8959 25007 8965
rect 24949 8925 24961 8959
rect 24995 8956 25007 8959
rect 25038 8956 25044 8968
rect 24995 8928 25044 8956
rect 24995 8925 25007 8928
rect 24949 8919 25007 8925
rect 25038 8916 25044 8928
rect 25096 8916 25102 8968
rect 30377 8959 30435 8965
rect 30377 8925 30389 8959
rect 30423 8956 30435 8959
rect 31018 8956 31024 8968
rect 30423 8928 31024 8956
rect 30423 8925 30435 8928
rect 30377 8919 30435 8925
rect 31018 8916 31024 8928
rect 31076 8956 31082 8968
rect 31113 8959 31171 8965
rect 31113 8956 31125 8959
rect 31076 8928 31125 8956
rect 31076 8916 31082 8928
rect 31113 8925 31125 8928
rect 31159 8956 31171 8959
rect 31478 8956 31484 8968
rect 31159 8928 31484 8956
rect 31159 8925 31171 8928
rect 31113 8919 31171 8925
rect 31478 8916 31484 8928
rect 31536 8916 31542 8968
rect 32674 8956 32680 8968
rect 32635 8928 32680 8956
rect 32674 8916 32680 8928
rect 32732 8916 32738 8968
rect 33594 8916 33600 8968
rect 33652 8956 33658 8968
rect 34333 8959 34391 8965
rect 34333 8956 34345 8959
rect 33652 8928 34345 8956
rect 33652 8916 33658 8928
rect 34333 8925 34345 8928
rect 34379 8925 34391 8959
rect 35894 8956 35900 8968
rect 35807 8928 35900 8956
rect 34333 8919 34391 8925
rect 35894 8916 35900 8928
rect 35952 8956 35958 8968
rect 36262 8956 36268 8968
rect 35952 8928 36268 8956
rect 35952 8916 35958 8928
rect 36262 8916 36268 8928
rect 36320 8916 36326 8968
rect 19334 8888 19340 8900
rect 19295 8860 19340 8888
rect 19334 8848 19340 8860
rect 19392 8848 19398 8900
rect 30558 8888 30564 8900
rect 30519 8860 30564 8888
rect 30558 8848 30564 8860
rect 30616 8848 30622 8900
rect 31754 8848 31760 8900
rect 31812 8888 31818 8900
rect 32217 8891 32275 8897
rect 32217 8888 32229 8891
rect 31812 8860 32229 8888
rect 31812 8848 31818 8860
rect 32217 8857 32229 8860
rect 32263 8857 32275 8891
rect 32217 8851 32275 8857
rect 33321 8891 33379 8897
rect 33321 8857 33333 8891
rect 33367 8888 33379 8891
rect 33686 8888 33692 8900
rect 33367 8860 33692 8888
rect 33367 8857 33379 8860
rect 33321 8851 33379 8857
rect 33686 8848 33692 8860
rect 33744 8848 33750 8900
rect 33962 8848 33968 8900
rect 34020 8888 34026 8900
rect 34514 8888 34520 8900
rect 34020 8860 34520 8888
rect 34020 8848 34026 8860
rect 34514 8848 34520 8860
rect 34572 8848 34578 8900
rect 18969 8823 19027 8829
rect 18969 8789 18981 8823
rect 19015 8820 19027 8823
rect 19978 8820 19984 8832
rect 19015 8792 19984 8820
rect 19015 8789 19027 8792
rect 18969 8783 19027 8789
rect 19978 8780 19984 8792
rect 20036 8780 20042 8832
rect 20254 8820 20260 8832
rect 20215 8792 20260 8820
rect 20254 8780 20260 8792
rect 20312 8780 20318 8832
rect 23750 8820 23756 8832
rect 23711 8792 23756 8820
rect 23750 8780 23756 8792
rect 23808 8780 23814 8832
rect 24397 8823 24455 8829
rect 24397 8789 24409 8823
rect 24443 8820 24455 8823
rect 24762 8820 24768 8832
rect 24443 8792 24768 8820
rect 24443 8789 24455 8792
rect 24397 8783 24455 8789
rect 24762 8780 24768 8792
rect 24820 8780 24826 8832
rect 27893 8823 27951 8829
rect 27893 8789 27905 8823
rect 27939 8820 27951 8823
rect 28166 8820 28172 8832
rect 27939 8792 28172 8820
rect 27939 8789 27951 8792
rect 27893 8783 27951 8789
rect 28166 8780 28172 8792
rect 28224 8780 28230 8832
rect 29178 8780 29184 8832
rect 29236 8820 29242 8832
rect 29365 8823 29423 8829
rect 29365 8820 29377 8823
rect 29236 8792 29377 8820
rect 29236 8780 29242 8792
rect 29365 8789 29377 8792
rect 29411 8820 29423 8823
rect 29917 8823 29975 8829
rect 29917 8820 29929 8823
rect 29411 8792 29929 8820
rect 29411 8789 29423 8792
rect 29365 8783 29423 8789
rect 29917 8789 29929 8792
rect 29963 8789 29975 8823
rect 33778 8820 33784 8832
rect 33739 8792 33784 8820
rect 29917 8783 29975 8789
rect 33778 8780 33784 8792
rect 33836 8780 33842 8832
rect 35894 8780 35900 8832
rect 35952 8820 35958 8832
rect 36449 8823 36507 8829
rect 36449 8820 36461 8823
rect 35952 8792 36461 8820
rect 35952 8780 35958 8792
rect 36449 8789 36461 8792
rect 36495 8820 36507 8823
rect 36998 8820 37004 8832
rect 36495 8792 37004 8820
rect 36495 8789 36507 8792
rect 36449 8783 36507 8789
rect 36998 8780 37004 8792
rect 37056 8780 37062 8832
rect 1104 8730 38824 8752
rect 1104 8678 7648 8730
rect 7700 8678 7712 8730
rect 7764 8678 7776 8730
rect 7828 8678 7840 8730
rect 7892 8678 20982 8730
rect 21034 8678 21046 8730
rect 21098 8678 21110 8730
rect 21162 8678 21174 8730
rect 21226 8678 34315 8730
rect 34367 8678 34379 8730
rect 34431 8678 34443 8730
rect 34495 8678 34507 8730
rect 34559 8678 38824 8730
rect 1104 8656 38824 8678
rect 1673 8619 1731 8625
rect 1673 8585 1685 8619
rect 1719 8616 1731 8619
rect 1946 8616 1952 8628
rect 1719 8588 1952 8616
rect 1719 8585 1731 8588
rect 1673 8579 1731 8585
rect 1946 8576 1952 8588
rect 2004 8576 2010 8628
rect 2041 8619 2099 8625
rect 2041 8585 2053 8619
rect 2087 8616 2099 8619
rect 2498 8616 2504 8628
rect 2087 8588 2504 8616
rect 2087 8585 2099 8588
rect 2041 8579 2099 8585
rect 2148 8489 2176 8588
rect 2498 8576 2504 8588
rect 2556 8576 2562 8628
rect 3418 8576 3424 8628
rect 3476 8616 3482 8628
rect 3513 8619 3571 8625
rect 3513 8616 3525 8619
rect 3476 8588 3525 8616
rect 3476 8576 3482 8588
rect 3513 8585 3525 8588
rect 3559 8616 3571 8619
rect 4154 8616 4160 8628
rect 3559 8588 4160 8616
rect 3559 8585 3571 8588
rect 3513 8579 3571 8585
rect 4154 8576 4160 8588
rect 4212 8576 4218 8628
rect 5074 8576 5080 8628
rect 5132 8616 5138 8628
rect 5261 8619 5319 8625
rect 5261 8616 5273 8619
rect 5132 8588 5273 8616
rect 5132 8576 5138 8588
rect 5261 8585 5273 8588
rect 5307 8585 5319 8619
rect 5261 8579 5319 8585
rect 7745 8619 7803 8625
rect 7745 8585 7757 8619
rect 7791 8616 7803 8619
rect 8570 8616 8576 8628
rect 7791 8588 8576 8616
rect 7791 8585 7803 8588
rect 7745 8579 7803 8585
rect 7852 8560 7880 8588
rect 8570 8576 8576 8588
rect 8628 8576 8634 8628
rect 9674 8616 9680 8628
rect 9635 8588 9680 8616
rect 9674 8576 9680 8588
rect 9732 8576 9738 8628
rect 10226 8616 10232 8628
rect 10187 8588 10232 8616
rect 10226 8576 10232 8588
rect 10284 8576 10290 8628
rect 10870 8616 10876 8628
rect 10831 8588 10876 8616
rect 10870 8576 10876 8588
rect 10928 8576 10934 8628
rect 11606 8576 11612 8628
rect 11664 8616 11670 8628
rect 11793 8619 11851 8625
rect 11793 8616 11805 8619
rect 11664 8588 11805 8616
rect 11664 8576 11670 8588
rect 11793 8585 11805 8588
rect 11839 8585 11851 8619
rect 13998 8616 14004 8628
rect 13959 8588 14004 8616
rect 11793 8579 11851 8585
rect 13998 8576 14004 8588
rect 14056 8576 14062 8628
rect 14918 8616 14924 8628
rect 14879 8588 14924 8616
rect 14918 8576 14924 8588
rect 14976 8576 14982 8628
rect 17589 8619 17647 8625
rect 17589 8585 17601 8619
rect 17635 8616 17647 8619
rect 17954 8616 17960 8628
rect 17635 8588 17960 8616
rect 17635 8585 17647 8588
rect 17589 8579 17647 8585
rect 17954 8576 17960 8588
rect 18012 8576 18018 8628
rect 19794 8576 19800 8628
rect 19852 8616 19858 8628
rect 20257 8619 20315 8625
rect 20257 8616 20269 8619
rect 19852 8588 20269 8616
rect 19852 8576 19858 8588
rect 20257 8585 20269 8588
rect 20303 8585 20315 8619
rect 23382 8616 23388 8628
rect 23343 8588 23388 8616
rect 20257 8579 20315 8585
rect 23382 8576 23388 8588
rect 23440 8576 23446 8628
rect 25038 8616 25044 8628
rect 24999 8588 25044 8616
rect 25038 8576 25044 8588
rect 25096 8576 25102 8628
rect 26050 8616 26056 8628
rect 26011 8588 26056 8616
rect 26050 8576 26056 8588
rect 26108 8576 26114 8628
rect 26510 8616 26516 8628
rect 26471 8588 26516 8616
rect 26510 8576 26516 8588
rect 26568 8616 26574 8628
rect 28074 8616 28080 8628
rect 26568 8588 27568 8616
rect 28035 8588 28080 8616
rect 26568 8576 26574 8588
rect 3970 8508 3976 8560
rect 4028 8548 4034 8560
rect 7009 8551 7067 8557
rect 7009 8548 7021 8551
rect 4028 8520 7021 8548
rect 4028 8508 4034 8520
rect 7009 8517 7021 8520
rect 7055 8517 7067 8551
rect 7009 8511 7067 8517
rect 7834 8508 7840 8560
rect 7892 8508 7898 8560
rect 15746 8548 15752 8560
rect 15707 8520 15752 8548
rect 15746 8508 15752 8520
rect 15804 8508 15810 8560
rect 16390 8508 16396 8560
rect 16448 8548 16454 8560
rect 16485 8551 16543 8557
rect 16485 8548 16497 8551
rect 16448 8520 16497 8548
rect 16448 8508 16454 8520
rect 16485 8517 16497 8520
rect 16531 8517 16543 8551
rect 18138 8548 18144 8560
rect 18099 8520 18144 8548
rect 16485 8511 16543 8517
rect 18138 8508 18144 8520
rect 18196 8508 18202 8560
rect 19521 8551 19579 8557
rect 19521 8517 19533 8551
rect 19567 8548 19579 8551
rect 19886 8548 19892 8560
rect 19567 8520 19892 8548
rect 19567 8517 19579 8520
rect 19521 8511 19579 8517
rect 19886 8508 19892 8520
rect 19944 8508 19950 8560
rect 21913 8551 21971 8557
rect 21913 8517 21925 8551
rect 21959 8548 21971 8551
rect 22002 8548 22008 8560
rect 21959 8520 22008 8548
rect 21959 8517 21971 8520
rect 21913 8511 21971 8517
rect 22002 8508 22008 8520
rect 22060 8508 22066 8560
rect 2133 8483 2191 8489
rect 2133 8449 2145 8483
rect 2179 8449 2191 8483
rect 2133 8443 2191 8449
rect 4893 8483 4951 8489
rect 4893 8449 4905 8483
rect 4939 8480 4951 8483
rect 5258 8480 5264 8492
rect 4939 8452 5264 8480
rect 4939 8449 4951 8452
rect 4893 8443 4951 8449
rect 5258 8440 5264 8452
rect 5316 8440 5322 8492
rect 5534 8440 5540 8492
rect 5592 8480 5598 8492
rect 5721 8483 5779 8489
rect 5721 8480 5733 8483
rect 5592 8452 5733 8480
rect 5592 8440 5598 8452
rect 5721 8449 5733 8452
rect 5767 8480 5779 8483
rect 6454 8480 6460 8492
rect 5767 8452 6460 8480
rect 5767 8449 5779 8452
rect 5721 8443 5779 8449
rect 6454 8440 6460 8452
rect 6512 8440 6518 8492
rect 10318 8440 10324 8492
rect 10376 8480 10382 8492
rect 11425 8483 11483 8489
rect 11425 8480 11437 8483
rect 10376 8452 11437 8480
rect 10376 8440 10382 8452
rect 11425 8449 11437 8452
rect 11471 8449 11483 8483
rect 16942 8480 16948 8492
rect 16903 8452 16948 8480
rect 11425 8443 11483 8449
rect 16942 8440 16948 8452
rect 17000 8440 17006 8492
rect 19058 8480 19064 8492
rect 18432 8452 19064 8480
rect 18432 8424 18460 8452
rect 19058 8440 19064 8452
rect 19116 8440 19122 8492
rect 20622 8480 20628 8492
rect 20583 8452 20628 8480
rect 20622 8440 20628 8452
rect 20680 8440 20686 8492
rect 23400 8480 23428 8576
rect 26878 8548 26884 8560
rect 26839 8520 26884 8548
rect 26878 8508 26884 8520
rect 26936 8508 26942 8560
rect 27154 8548 27160 8560
rect 27115 8520 27160 8548
rect 27154 8508 27160 8520
rect 27212 8508 27218 8560
rect 27540 8548 27568 8588
rect 28074 8576 28080 8588
rect 28132 8576 28138 8628
rect 28534 8576 28540 8628
rect 28592 8616 28598 8628
rect 29365 8619 29423 8625
rect 29365 8616 29377 8619
rect 28592 8588 29377 8616
rect 28592 8576 28598 8588
rect 29365 8585 29377 8588
rect 29411 8585 29423 8619
rect 30926 8616 30932 8628
rect 30887 8588 30932 8616
rect 29365 8579 29423 8585
rect 30926 8576 30932 8588
rect 30984 8576 30990 8628
rect 37274 8616 37280 8628
rect 37235 8588 37280 8616
rect 37274 8576 37280 8588
rect 37332 8576 37338 8628
rect 28350 8548 28356 8560
rect 27540 8520 28356 8548
rect 23658 8480 23664 8492
rect 23400 8452 23664 8480
rect 23658 8440 23664 8452
rect 23716 8440 23722 8492
rect 27540 8489 27568 8520
rect 28350 8508 28356 8520
rect 28408 8508 28414 8560
rect 30834 8508 30840 8560
rect 30892 8548 30898 8560
rect 31849 8551 31907 8557
rect 31849 8548 31861 8551
rect 30892 8520 31861 8548
rect 30892 8508 30898 8520
rect 31849 8517 31861 8520
rect 31895 8517 31907 8551
rect 32766 8548 32772 8560
rect 32727 8520 32772 8548
rect 31849 8511 31907 8517
rect 32766 8508 32772 8520
rect 32824 8508 32830 8560
rect 33042 8548 33048 8560
rect 33003 8520 33048 8548
rect 33042 8508 33048 8520
rect 33100 8508 33106 8560
rect 36262 8548 36268 8560
rect 36223 8520 36268 8548
rect 36262 8508 36268 8520
rect 36320 8508 36326 8560
rect 37550 8548 37556 8560
rect 37511 8520 37556 8548
rect 37550 8508 37556 8520
rect 37608 8508 37614 8560
rect 27525 8483 27583 8489
rect 27525 8449 27537 8483
rect 27571 8449 27583 8483
rect 27706 8480 27712 8492
rect 27667 8452 27712 8480
rect 27525 8443 27583 8449
rect 27706 8440 27712 8452
rect 27764 8440 27770 8492
rect 29089 8483 29147 8489
rect 29089 8449 29101 8483
rect 29135 8480 29147 8483
rect 29825 8483 29883 8489
rect 29825 8480 29837 8483
rect 29135 8452 29837 8480
rect 29135 8449 29147 8452
rect 29089 8443 29147 8449
rect 29825 8449 29837 8452
rect 29871 8480 29883 8483
rect 30006 8480 30012 8492
rect 29871 8452 30012 8480
rect 29871 8449 29883 8452
rect 29825 8443 29883 8449
rect 30006 8440 30012 8452
rect 30064 8440 30070 8492
rect 31478 8480 31484 8492
rect 31439 8452 31484 8480
rect 31478 8440 31484 8452
rect 31536 8440 31542 8492
rect 32784 8480 32812 8508
rect 33410 8480 33416 8492
rect 32784 8452 33416 8480
rect 33410 8440 33416 8452
rect 33468 8440 33474 8492
rect 33520 8452 34744 8480
rect 1946 8372 1952 8424
rect 2004 8412 2010 8424
rect 2389 8415 2447 8421
rect 2389 8412 2401 8415
rect 2004 8384 2401 8412
rect 2004 8372 2010 8384
rect 2389 8381 2401 8384
rect 2435 8381 2447 8415
rect 2389 8375 2447 8381
rect 4525 8415 4583 8421
rect 4525 8381 4537 8415
rect 4571 8412 4583 8415
rect 5350 8412 5356 8424
rect 4571 8384 5356 8412
rect 4571 8381 4583 8384
rect 4525 8375 4583 8381
rect 5350 8372 5356 8384
rect 5408 8412 5414 8424
rect 5813 8415 5871 8421
rect 5813 8412 5825 8415
rect 5408 8384 5825 8412
rect 5408 8372 5414 8384
rect 5813 8381 5825 8384
rect 5859 8381 5871 8415
rect 6822 8412 6828 8424
rect 6783 8384 6828 8412
rect 5813 8375 5871 8381
rect 6822 8372 6828 8384
rect 6880 8372 6886 8424
rect 8297 8415 8355 8421
rect 8297 8381 8309 8415
rect 8343 8381 8355 8415
rect 8297 8375 8355 8381
rect 4157 8347 4215 8353
rect 4157 8313 4169 8347
rect 4203 8344 4215 8347
rect 5442 8344 5448 8356
rect 4203 8316 5448 8344
rect 4203 8313 4215 8316
rect 4157 8307 4215 8313
rect 5442 8304 5448 8316
rect 5500 8304 5506 8356
rect 5718 8344 5724 8356
rect 5679 8316 5724 8344
rect 5718 8304 5724 8316
rect 5776 8304 5782 8356
rect 6362 8344 6368 8356
rect 6323 8316 6368 8344
rect 6362 8304 6368 8316
rect 6420 8304 6426 8356
rect 8312 8344 8340 8375
rect 8386 8372 8392 8424
rect 8444 8412 8450 8424
rect 8553 8415 8611 8421
rect 8553 8412 8565 8415
rect 8444 8384 8565 8412
rect 8444 8372 8450 8384
rect 8553 8381 8565 8384
rect 8599 8381 8611 8415
rect 8553 8375 8611 8381
rect 10410 8372 10416 8424
rect 10468 8412 10474 8424
rect 10689 8415 10747 8421
rect 10689 8412 10701 8415
rect 10468 8384 10701 8412
rect 10468 8372 10474 8384
rect 10689 8381 10701 8384
rect 10735 8412 10747 8415
rect 10735 8384 11376 8412
rect 10735 8381 10747 8384
rect 10689 8375 10747 8381
rect 11348 8356 11376 8384
rect 11882 8372 11888 8424
rect 11940 8412 11946 8424
rect 12253 8415 12311 8421
rect 12253 8412 12265 8415
rect 11940 8384 12265 8412
rect 11940 8372 11946 8384
rect 12253 8381 12265 8384
rect 12299 8412 12311 8415
rect 12621 8415 12679 8421
rect 12621 8412 12633 8415
rect 12299 8384 12633 8412
rect 12299 8381 12311 8384
rect 12253 8375 12311 8381
rect 12621 8381 12633 8384
rect 12667 8381 12679 8415
rect 18414 8412 18420 8424
rect 18375 8384 18420 8412
rect 12621 8375 12679 8381
rect 18414 8372 18420 8384
rect 18472 8372 18478 8424
rect 18693 8415 18751 8421
rect 18693 8381 18705 8415
rect 18739 8412 18751 8415
rect 19889 8415 19947 8421
rect 19889 8412 19901 8415
rect 18739 8384 19901 8412
rect 18739 8381 18751 8384
rect 18693 8375 18751 8381
rect 19889 8381 19901 8384
rect 19935 8412 19947 8415
rect 19978 8412 19984 8424
rect 19935 8384 19984 8412
rect 19935 8381 19947 8384
rect 19889 8375 19947 8381
rect 19978 8372 19984 8384
rect 20036 8372 20042 8424
rect 20162 8372 20168 8424
rect 20220 8412 20226 8424
rect 20809 8415 20867 8421
rect 20809 8412 20821 8415
rect 20220 8384 20821 8412
rect 20220 8372 20226 8384
rect 20809 8381 20821 8384
rect 20855 8381 20867 8415
rect 20809 8375 20867 8381
rect 20898 8372 20904 8424
rect 20956 8412 20962 8424
rect 21361 8415 21419 8421
rect 21361 8412 21373 8415
rect 20956 8384 21373 8412
rect 20956 8372 20962 8384
rect 21361 8381 21373 8384
rect 21407 8412 21419 8415
rect 21910 8412 21916 8424
rect 21407 8384 21916 8412
rect 21407 8381 21419 8384
rect 21361 8375 21419 8381
rect 21910 8372 21916 8384
rect 21968 8372 21974 8424
rect 22094 8372 22100 8424
rect 22152 8412 22158 8424
rect 22189 8415 22247 8421
rect 22189 8412 22201 8415
rect 22152 8384 22201 8412
rect 22152 8372 22158 8384
rect 22189 8381 22201 8384
rect 22235 8381 22247 8415
rect 28534 8412 28540 8424
rect 22189 8375 22247 8381
rect 27632 8384 28540 8412
rect 8754 8344 8760 8356
rect 8312 8316 8760 8344
rect 8754 8304 8760 8316
rect 8812 8304 8818 8356
rect 10962 8304 10968 8356
rect 11020 8344 11026 8356
rect 11149 8347 11207 8353
rect 11149 8344 11161 8347
rect 11020 8316 11161 8344
rect 11020 8304 11026 8316
rect 11149 8313 11161 8316
rect 11195 8313 11207 8347
rect 11330 8344 11336 8356
rect 11291 8316 11336 8344
rect 11149 8307 11207 8313
rect 11330 8304 11336 8316
rect 11388 8304 11394 8356
rect 12526 8304 12532 8356
rect 12584 8344 12590 8356
rect 12866 8347 12924 8353
rect 12866 8344 12878 8347
rect 12584 8316 12878 8344
rect 12584 8304 12590 8316
rect 12866 8313 12878 8316
rect 12912 8313 12924 8347
rect 15286 8344 15292 8356
rect 15247 8316 15292 8344
rect 12866 8307 12924 8313
rect 15286 8304 15292 8316
rect 15344 8304 15350 8356
rect 16298 8344 16304 8356
rect 16211 8316 16304 8344
rect 16298 8304 16304 8316
rect 16356 8344 16362 8356
rect 17034 8344 17040 8356
rect 16356 8316 16896 8344
rect 16995 8316 17040 8344
rect 16356 8304 16362 8316
rect 6454 8236 6460 8288
rect 6512 8276 6518 8288
rect 6638 8276 6644 8288
rect 6512 8248 6644 8276
rect 6512 8236 6518 8248
rect 6638 8236 6644 8248
rect 6696 8236 6702 8288
rect 7006 8236 7012 8288
rect 7064 8276 7070 8288
rect 7190 8276 7196 8288
rect 7064 8248 7196 8276
rect 7064 8236 7070 8248
rect 7190 8236 7196 8248
rect 7248 8236 7254 8288
rect 7466 8236 7472 8288
rect 7524 8276 7530 8288
rect 8021 8279 8079 8285
rect 8021 8276 8033 8279
rect 7524 8248 8033 8276
rect 7524 8236 7530 8248
rect 8021 8245 8033 8248
rect 8067 8276 8079 8279
rect 8110 8276 8116 8288
rect 8067 8248 8116 8276
rect 8067 8245 8079 8248
rect 8021 8239 8079 8245
rect 8110 8236 8116 8248
rect 8168 8236 8174 8288
rect 16868 8276 16896 8316
rect 17034 8304 17040 8316
rect 17092 8304 17098 8356
rect 17218 8344 17224 8356
rect 17144 8316 17224 8344
rect 16945 8279 17003 8285
rect 16945 8276 16957 8279
rect 16868 8248 16957 8276
rect 16945 8245 16957 8248
rect 16991 8276 17003 8279
rect 17144 8276 17172 8316
rect 17218 8304 17224 8316
rect 17276 8304 17282 8356
rect 18598 8344 18604 8356
rect 18559 8316 18604 8344
rect 18598 8304 18604 8316
rect 18656 8304 18662 8356
rect 19610 8304 19616 8356
rect 19668 8344 19674 8356
rect 20254 8344 20260 8356
rect 19668 8316 20260 8344
rect 19668 8304 19674 8316
rect 20254 8304 20260 8316
rect 20312 8344 20318 8356
rect 20717 8347 20775 8353
rect 20717 8344 20729 8347
rect 20312 8316 20729 8344
rect 20312 8304 20318 8316
rect 20717 8313 20729 8316
rect 20763 8313 20775 8347
rect 22462 8344 22468 8356
rect 20717 8307 20775 8313
rect 22020 8316 22468 8344
rect 21634 8276 21640 8288
rect 16991 8248 17172 8276
rect 21595 8248 21640 8276
rect 16991 8245 17003 8248
rect 16945 8239 17003 8245
rect 21634 8236 21640 8248
rect 21692 8236 21698 8288
rect 21910 8236 21916 8288
rect 21968 8276 21974 8288
rect 22020 8276 22048 8316
rect 22462 8304 22468 8316
rect 22520 8304 22526 8356
rect 23750 8304 23756 8356
rect 23808 8344 23814 8356
rect 23928 8347 23986 8353
rect 23928 8344 23940 8347
rect 23808 8316 23940 8344
rect 23808 8304 23814 8316
rect 23928 8313 23940 8316
rect 23974 8344 23986 8347
rect 23974 8316 24808 8344
rect 23974 8313 23986 8316
rect 23928 8307 23986 8313
rect 22370 8276 22376 8288
rect 21968 8248 22048 8276
rect 22331 8248 22376 8276
rect 21968 8236 21974 8248
rect 22370 8236 22376 8248
rect 22428 8276 22434 8288
rect 22833 8279 22891 8285
rect 22833 8276 22845 8279
rect 22428 8248 22845 8276
rect 22428 8236 22434 8248
rect 22833 8245 22845 8248
rect 22879 8245 22891 8279
rect 24780 8276 24808 8316
rect 24946 8304 24952 8356
rect 25004 8344 25010 8356
rect 25593 8347 25651 8353
rect 25593 8344 25605 8347
rect 25004 8316 25605 8344
rect 25004 8304 25010 8316
rect 25593 8313 25605 8316
rect 25639 8313 25651 8347
rect 25593 8307 25651 8313
rect 26878 8304 26884 8356
rect 26936 8344 26942 8356
rect 27632 8353 27660 8384
rect 28534 8372 28540 8384
rect 28592 8372 28598 8424
rect 29178 8372 29184 8424
rect 29236 8412 29242 8424
rect 29917 8415 29975 8421
rect 29917 8412 29929 8415
rect 29236 8384 29929 8412
rect 29236 8372 29242 8384
rect 29917 8381 29929 8384
rect 29963 8381 29975 8415
rect 30650 8412 30656 8424
rect 30611 8384 30656 8412
rect 29917 8375 29975 8381
rect 30650 8372 30656 8384
rect 30708 8412 30714 8424
rect 31110 8412 31116 8424
rect 30708 8384 31116 8412
rect 30708 8372 30714 8384
rect 31110 8372 31116 8384
rect 31168 8412 31174 8424
rect 31205 8415 31263 8421
rect 31205 8412 31217 8415
rect 31168 8384 31217 8412
rect 31168 8372 31174 8384
rect 31205 8381 31217 8384
rect 31251 8381 31263 8415
rect 31205 8375 31263 8381
rect 32950 8372 32956 8424
rect 33008 8412 33014 8424
rect 33520 8412 33548 8452
rect 34716 8424 34744 8452
rect 34054 8412 34060 8424
rect 33008 8384 33548 8412
rect 34015 8384 34060 8412
rect 33008 8372 33014 8384
rect 34054 8372 34060 8384
rect 34112 8372 34118 8424
rect 34698 8372 34704 8424
rect 34756 8412 34762 8424
rect 34885 8415 34943 8421
rect 34885 8412 34897 8415
rect 34756 8384 34897 8412
rect 34756 8372 34762 8384
rect 34885 8381 34897 8384
rect 34931 8381 34943 8415
rect 35152 8415 35210 8421
rect 35152 8412 35164 8415
rect 34885 8375 34943 8381
rect 34992 8384 35164 8412
rect 27617 8347 27675 8353
rect 27617 8344 27629 8347
rect 26936 8316 27629 8344
rect 26936 8304 26942 8316
rect 27617 8313 27629 8316
rect 27663 8313 27675 8347
rect 27617 8307 27675 8313
rect 27706 8304 27712 8356
rect 27764 8344 27770 8356
rect 28629 8347 28687 8353
rect 28629 8344 28641 8347
rect 27764 8316 28641 8344
rect 27764 8304 27770 8316
rect 28629 8313 28641 8316
rect 28675 8344 28687 8347
rect 29825 8347 29883 8353
rect 29825 8344 29837 8347
rect 28675 8316 29837 8344
rect 28675 8313 28687 8316
rect 28629 8307 28687 8313
rect 29825 8313 29837 8316
rect 29871 8313 29883 8347
rect 32490 8344 32496 8356
rect 32403 8316 32496 8344
rect 29825 8307 29883 8313
rect 32490 8304 32496 8316
rect 32548 8344 32554 8356
rect 33594 8344 33600 8356
rect 32548 8316 33456 8344
rect 33555 8316 33600 8344
rect 32548 8304 32554 8316
rect 25498 8276 25504 8288
rect 24780 8248 25504 8276
rect 22833 8239 22891 8245
rect 25498 8236 25504 8248
rect 25556 8236 25562 8288
rect 30374 8276 30380 8288
rect 30287 8248 30380 8276
rect 30374 8236 30380 8248
rect 30432 8276 30438 8288
rect 31389 8279 31447 8285
rect 31389 8276 31401 8279
rect 30432 8248 31401 8276
rect 30432 8236 30438 8248
rect 31389 8245 31401 8248
rect 31435 8276 31447 8279
rect 32214 8276 32220 8288
rect 31435 8248 32220 8276
rect 31435 8245 31447 8248
rect 31389 8239 31447 8245
rect 32214 8236 32220 8248
rect 32272 8236 32278 8288
rect 33428 8276 33456 8316
rect 33594 8304 33600 8316
rect 33652 8304 33658 8356
rect 33870 8304 33876 8356
rect 33928 8344 33934 8356
rect 34330 8344 34336 8356
rect 33928 8316 34336 8344
rect 33928 8304 33934 8316
rect 34330 8304 34336 8316
rect 34388 8344 34394 8356
rect 34992 8344 35020 8384
rect 35152 8381 35164 8384
rect 35198 8412 35210 8415
rect 36817 8415 36875 8421
rect 36817 8412 36829 8415
rect 35198 8384 36829 8412
rect 35198 8381 35210 8384
rect 35152 8375 35210 8381
rect 36817 8381 36829 8384
rect 36863 8381 36875 8415
rect 37366 8412 37372 8424
rect 37327 8384 37372 8412
rect 36817 8375 36875 8381
rect 37366 8372 37372 8384
rect 37424 8412 37430 8424
rect 37921 8415 37979 8421
rect 37921 8412 37933 8415
rect 37424 8384 37933 8412
rect 37424 8372 37430 8384
rect 37921 8381 37933 8384
rect 37967 8381 37979 8415
rect 37921 8375 37979 8381
rect 34388 8316 35020 8344
rect 34388 8304 34394 8316
rect 33502 8276 33508 8288
rect 33428 8248 33508 8276
rect 33502 8236 33508 8248
rect 33560 8236 33566 8288
rect 34698 8276 34704 8288
rect 34611 8248 34704 8276
rect 34698 8236 34704 8248
rect 34756 8276 34762 8288
rect 35158 8276 35164 8288
rect 34756 8248 35164 8276
rect 34756 8236 34762 8248
rect 35158 8236 35164 8248
rect 35216 8236 35222 8288
rect 1104 8186 38824 8208
rect 1104 8134 14315 8186
rect 14367 8134 14379 8186
rect 14431 8134 14443 8186
rect 14495 8134 14507 8186
rect 14559 8134 27648 8186
rect 27700 8134 27712 8186
rect 27764 8134 27776 8186
rect 27828 8134 27840 8186
rect 27892 8134 38824 8186
rect 1104 8112 38824 8134
rect 2774 8032 2780 8084
rect 2832 8072 2838 8084
rect 3145 8075 3203 8081
rect 3145 8072 3157 8075
rect 2832 8044 3157 8072
rect 2832 8032 2838 8044
rect 3145 8041 3157 8044
rect 3191 8041 3203 8075
rect 3878 8072 3884 8084
rect 3839 8044 3884 8072
rect 3145 8035 3203 8041
rect 3878 8032 3884 8044
rect 3936 8032 3942 8084
rect 7466 8032 7472 8084
rect 7524 8072 7530 8084
rect 7745 8075 7803 8081
rect 7745 8072 7757 8075
rect 7524 8044 7757 8072
rect 7524 8032 7530 8044
rect 7745 8041 7757 8044
rect 7791 8041 7803 8075
rect 8662 8072 8668 8084
rect 8623 8044 8668 8072
rect 7745 8035 7803 8041
rect 8662 8032 8668 8044
rect 8720 8032 8726 8084
rect 10873 8075 10931 8081
rect 10873 8041 10885 8075
rect 10919 8072 10931 8075
rect 10962 8072 10968 8084
rect 10919 8044 10968 8072
rect 10919 8041 10931 8044
rect 10873 8035 10931 8041
rect 10962 8032 10968 8044
rect 11020 8032 11026 8084
rect 12526 8032 12532 8084
rect 12584 8072 12590 8084
rect 12621 8075 12679 8081
rect 12621 8072 12633 8075
rect 12584 8044 12633 8072
rect 12584 8032 12590 8044
rect 12621 8041 12633 8044
rect 12667 8072 12679 8075
rect 13173 8075 13231 8081
rect 13173 8072 13185 8075
rect 12667 8044 13185 8072
rect 12667 8041 12679 8044
rect 12621 8035 12679 8041
rect 13173 8041 13185 8044
rect 13219 8041 13231 8075
rect 13538 8072 13544 8084
rect 13499 8044 13544 8072
rect 13173 8035 13231 8041
rect 13538 8032 13544 8044
rect 13596 8032 13602 8084
rect 17586 8072 17592 8084
rect 17547 8044 17592 8072
rect 17586 8032 17592 8044
rect 17644 8032 17650 8084
rect 19518 8032 19524 8084
rect 19576 8072 19582 8084
rect 19613 8075 19671 8081
rect 19613 8072 19625 8075
rect 19576 8044 19625 8072
rect 19576 8032 19582 8044
rect 19613 8041 19625 8044
rect 19659 8041 19671 8075
rect 20622 8072 20628 8084
rect 20583 8044 20628 8072
rect 19613 8035 19671 8041
rect 20622 8032 20628 8044
rect 20680 8032 20686 8084
rect 20993 8075 21051 8081
rect 20993 8041 21005 8075
rect 21039 8072 21051 8075
rect 21726 8072 21732 8084
rect 21039 8044 21732 8072
rect 21039 8041 21051 8044
rect 20993 8035 21051 8041
rect 21726 8032 21732 8044
rect 21784 8032 21790 8084
rect 21910 8072 21916 8084
rect 21871 8044 21916 8072
rect 21910 8032 21916 8044
rect 21968 8032 21974 8084
rect 24397 8075 24455 8081
rect 24397 8041 24409 8075
rect 24443 8072 24455 8075
rect 25038 8072 25044 8084
rect 24443 8044 25044 8072
rect 24443 8041 24455 8044
rect 24397 8035 24455 8041
rect 2314 8004 2320 8016
rect 2275 7976 2320 8004
rect 2314 7964 2320 7976
rect 2372 7964 2378 8016
rect 2866 8004 2872 8016
rect 2827 7976 2872 8004
rect 2866 7964 2872 7976
rect 2924 7964 2930 8016
rect 4154 7964 4160 8016
rect 4212 8004 4218 8016
rect 4954 8007 5012 8013
rect 4954 8004 4966 8007
rect 4212 7976 4966 8004
rect 4212 7964 4218 7976
rect 4954 7973 4966 7976
rect 5000 8004 5012 8007
rect 5074 8004 5080 8016
rect 5000 7976 5080 8004
rect 5000 7973 5012 7976
rect 4954 7967 5012 7973
rect 5074 7964 5080 7976
rect 5132 7964 5138 8016
rect 6638 7964 6644 8016
rect 6696 8004 6702 8016
rect 7561 8007 7619 8013
rect 7561 8004 7573 8007
rect 6696 7976 7573 8004
rect 6696 7964 6702 7976
rect 7561 7973 7573 7976
rect 7607 8004 7619 8007
rect 7834 8004 7840 8016
rect 7607 7976 7840 8004
rect 7607 7973 7619 7976
rect 7561 7967 7619 7973
rect 7834 7964 7840 7976
rect 7892 7964 7898 8016
rect 8386 7964 8392 8016
rect 8444 8004 8450 8016
rect 9033 8007 9091 8013
rect 9033 8004 9045 8007
rect 8444 7976 9045 8004
rect 8444 7964 8450 7976
rect 9033 7973 9045 7976
rect 9079 8004 9091 8007
rect 9306 8004 9312 8016
rect 9079 7976 9312 8004
rect 9079 7973 9091 7976
rect 9033 7967 9091 7973
rect 9306 7964 9312 7976
rect 9364 7964 9370 8016
rect 9674 7964 9680 8016
rect 9732 8004 9738 8016
rect 10229 8007 10287 8013
rect 10229 8004 10241 8007
rect 9732 7976 10241 8004
rect 9732 7964 9738 7976
rect 10229 7973 10241 7976
rect 10275 7973 10287 8007
rect 11882 8004 11888 8016
rect 10229 7967 10287 7973
rect 11256 7976 11888 8004
rect 1673 7939 1731 7945
rect 1673 7905 1685 7939
rect 1719 7936 1731 7939
rect 2409 7939 2467 7945
rect 2409 7936 2421 7939
rect 1719 7908 2421 7936
rect 1719 7905 1731 7908
rect 1673 7899 1731 7905
rect 2409 7905 2421 7908
rect 2455 7936 2467 7939
rect 2498 7936 2504 7948
rect 2455 7908 2504 7936
rect 2455 7905 2467 7908
rect 2409 7899 2467 7905
rect 2498 7896 2504 7908
rect 2556 7896 2562 7948
rect 9324 7936 9352 7964
rect 10318 7936 10324 7948
rect 9324 7908 10324 7936
rect 10318 7896 10324 7908
rect 10376 7896 10382 7948
rect 11256 7945 11284 7976
rect 11882 7964 11888 7976
rect 11940 7964 11946 8016
rect 16666 8004 16672 8016
rect 16627 7976 16672 8004
rect 16666 7964 16672 7976
rect 16724 7964 16730 8016
rect 17034 7964 17040 8016
rect 17092 8004 17098 8016
rect 17221 8007 17279 8013
rect 17221 8004 17233 8007
rect 17092 7976 17233 8004
rect 17092 7964 17098 7976
rect 17221 7973 17233 7976
rect 17267 8004 17279 8007
rect 17770 8004 17776 8016
rect 17267 7976 17776 8004
rect 17267 7973 17279 7976
rect 17221 7967 17279 7973
rect 17770 7964 17776 7976
rect 17828 8004 17834 8016
rect 17948 8007 18006 8013
rect 17948 8004 17960 8007
rect 17828 7976 17960 8004
rect 17828 7964 17834 7976
rect 17948 7973 17960 7976
rect 17994 8004 18006 8007
rect 18046 8004 18052 8016
rect 17994 7976 18052 8004
rect 17994 7973 18006 7976
rect 17948 7967 18006 7973
rect 18046 7964 18052 7976
rect 18104 7964 18110 8016
rect 21358 7964 21364 8016
rect 21416 8004 21422 8016
rect 22094 8004 22100 8016
rect 21416 7976 22100 8004
rect 21416 7964 21422 7976
rect 22094 7964 22100 7976
rect 22152 7964 22158 8016
rect 22272 8007 22330 8013
rect 22272 8004 22284 8007
rect 22204 7976 22284 8004
rect 11514 7945 11520 7948
rect 11241 7939 11299 7945
rect 11241 7905 11253 7939
rect 11287 7905 11299 7939
rect 11508 7936 11520 7945
rect 11475 7908 11520 7936
rect 11241 7899 11299 7905
rect 11508 7899 11520 7908
rect 11514 7896 11520 7899
rect 11572 7896 11578 7948
rect 13722 7936 13728 7948
rect 13683 7908 13728 7936
rect 13722 7896 13728 7908
rect 13780 7896 13786 7948
rect 16025 7939 16083 7945
rect 16025 7905 16037 7939
rect 16071 7936 16083 7939
rect 16482 7936 16488 7948
rect 16071 7908 16488 7936
rect 16071 7905 16083 7908
rect 16025 7899 16083 7905
rect 16482 7896 16488 7908
rect 16540 7896 16546 7948
rect 20162 7936 20168 7948
rect 16776 7908 20168 7936
rect 2317 7871 2375 7877
rect 2317 7837 2329 7871
rect 2363 7868 2375 7871
rect 2682 7868 2688 7880
rect 2363 7840 2688 7868
rect 2363 7837 2375 7840
rect 2317 7831 2375 7837
rect 2682 7828 2688 7840
rect 2740 7828 2746 7880
rect 4706 7868 4712 7880
rect 4667 7840 4712 7868
rect 4706 7828 4712 7840
rect 4764 7828 4770 7880
rect 7837 7871 7895 7877
rect 7837 7837 7849 7871
rect 7883 7868 7895 7871
rect 8018 7868 8024 7880
rect 7883 7840 8024 7868
rect 7883 7837 7895 7840
rect 7837 7831 7895 7837
rect 8018 7828 8024 7840
rect 8076 7828 8082 7880
rect 8110 7828 8116 7880
rect 8168 7868 8174 7880
rect 8389 7871 8447 7877
rect 8389 7868 8401 7871
rect 8168 7840 8401 7868
rect 8168 7828 8174 7840
rect 8389 7837 8401 7840
rect 8435 7868 8447 7871
rect 8754 7868 8760 7880
rect 8435 7840 8760 7868
rect 8435 7837 8447 7840
rect 8389 7831 8447 7837
rect 8754 7828 8760 7840
rect 8812 7828 8818 7880
rect 10042 7828 10048 7880
rect 10100 7868 10106 7880
rect 10137 7871 10195 7877
rect 10137 7868 10149 7871
rect 10100 7840 10149 7868
rect 10100 7828 10106 7840
rect 10137 7837 10149 7840
rect 10183 7837 10195 7871
rect 10137 7831 10195 7837
rect 15930 7828 15936 7880
rect 15988 7868 15994 7880
rect 16776 7877 16804 7908
rect 20162 7896 20168 7908
rect 20220 7896 20226 7948
rect 21542 7896 21548 7948
rect 21600 7936 21606 7948
rect 22204 7936 22232 7976
rect 22272 7973 22284 7976
rect 22318 8004 22330 8007
rect 24412 8004 24440 8035
rect 25038 8032 25044 8044
rect 25096 8032 25102 8084
rect 26329 8075 26387 8081
rect 26329 8041 26341 8075
rect 26375 8072 26387 8075
rect 27065 8075 27123 8081
rect 27065 8072 27077 8075
rect 26375 8044 27077 8072
rect 26375 8041 26387 8044
rect 26329 8035 26387 8041
rect 27065 8041 27077 8044
rect 27111 8072 27123 8075
rect 27154 8072 27160 8084
rect 27111 8044 27160 8072
rect 27111 8041 27123 8044
rect 27065 8035 27123 8041
rect 27154 8032 27160 8044
rect 27212 8032 27218 8084
rect 28442 8032 28448 8084
rect 28500 8072 28506 8084
rect 28537 8075 28595 8081
rect 28537 8072 28549 8075
rect 28500 8044 28549 8072
rect 28500 8032 28506 8044
rect 28537 8041 28549 8044
rect 28583 8041 28595 8075
rect 30466 8072 30472 8084
rect 30427 8044 30472 8072
rect 28537 8035 28595 8041
rect 30466 8032 30472 8044
rect 30524 8032 30530 8084
rect 30742 8032 30748 8084
rect 30800 8072 30806 8084
rect 31021 8075 31079 8081
rect 31021 8072 31033 8075
rect 30800 8044 31033 8072
rect 30800 8032 30806 8044
rect 31021 8041 31033 8044
rect 31067 8041 31079 8075
rect 31478 8072 31484 8084
rect 31439 8044 31484 8072
rect 31021 8035 31079 8041
rect 31478 8032 31484 8044
rect 31536 8032 31542 8084
rect 31938 8072 31944 8084
rect 31899 8044 31944 8072
rect 31938 8032 31944 8044
rect 31996 8032 32002 8084
rect 32493 8075 32551 8081
rect 32493 8041 32505 8075
rect 32539 8072 32551 8075
rect 33594 8072 33600 8084
rect 32539 8044 33600 8072
rect 32539 8041 32551 8044
rect 32493 8035 32551 8041
rect 33594 8032 33600 8044
rect 33652 8032 33658 8084
rect 34330 8072 34336 8084
rect 34291 8044 34336 8072
rect 34330 8032 34336 8044
rect 34388 8032 34394 8084
rect 36262 8032 36268 8084
rect 36320 8072 36326 8084
rect 36449 8075 36507 8081
rect 36449 8072 36461 8075
rect 36320 8044 36461 8072
rect 36320 8032 36326 8044
rect 36449 8041 36461 8044
rect 36495 8041 36507 8075
rect 36449 8035 36507 8041
rect 22318 7976 24440 8004
rect 24765 8007 24823 8013
rect 22318 7973 22330 7976
rect 22272 7967 22330 7973
rect 24765 7973 24777 8007
rect 24811 8004 24823 8007
rect 25409 8007 25467 8013
rect 25409 8004 25421 8007
rect 24811 7976 25421 8004
rect 24811 7973 24823 7976
rect 24765 7967 24823 7973
rect 25409 7973 25421 7976
rect 25455 8004 25467 8007
rect 26587 8007 26645 8013
rect 26587 8004 26599 8007
rect 25455 7976 26599 8004
rect 25455 7973 25467 7976
rect 25409 7967 25467 7973
rect 26587 7973 26599 7976
rect 26633 7973 26645 8007
rect 35986 8004 35992 8016
rect 35947 7976 35992 8004
rect 26587 7967 26645 7973
rect 35986 7964 35992 7976
rect 36044 7964 36050 8016
rect 25498 7936 25504 7948
rect 21600 7908 22232 7936
rect 25459 7908 25504 7936
rect 21600 7896 21606 7908
rect 25498 7896 25504 7908
rect 25556 7896 25562 7948
rect 26326 7896 26332 7948
rect 26384 7936 26390 7948
rect 26881 7939 26939 7945
rect 26881 7936 26893 7939
rect 26384 7908 26893 7936
rect 26384 7896 26390 7908
rect 26881 7905 26893 7908
rect 26927 7936 26939 7939
rect 27338 7936 27344 7948
rect 26927 7908 27344 7936
rect 26927 7905 26939 7908
rect 26881 7899 26939 7905
rect 27338 7896 27344 7908
rect 27396 7896 27402 7948
rect 28902 7896 28908 7948
rect 28960 7936 28966 7948
rect 29086 7936 29092 7948
rect 28960 7908 29092 7936
rect 28960 7896 28966 7908
rect 29086 7896 29092 7908
rect 29144 7896 29150 7948
rect 29178 7896 29184 7948
rect 29236 7936 29242 7948
rect 29345 7939 29403 7945
rect 29345 7936 29357 7939
rect 29236 7908 29357 7936
rect 29236 7896 29242 7908
rect 29345 7905 29357 7908
rect 29391 7905 29403 7939
rect 29345 7899 29403 7905
rect 32398 7896 32404 7948
rect 32456 7936 32462 7948
rect 33209 7939 33267 7945
rect 33209 7936 33221 7939
rect 32456 7908 33221 7936
rect 32456 7896 32462 7908
rect 33209 7905 33221 7908
rect 33255 7905 33267 7939
rect 33209 7899 33267 7905
rect 34974 7896 34980 7948
rect 35032 7936 35038 7948
rect 35526 7936 35532 7948
rect 35032 7908 35532 7936
rect 35032 7896 35038 7908
rect 35526 7896 35532 7908
rect 35584 7896 35590 7948
rect 36446 7936 36452 7948
rect 35912 7908 36452 7936
rect 16761 7871 16819 7877
rect 16761 7868 16773 7871
rect 15988 7840 16773 7868
rect 15988 7828 15994 7840
rect 16761 7837 16773 7840
rect 16807 7837 16819 7871
rect 17678 7868 17684 7880
rect 17639 7840 17684 7868
rect 16761 7831 16819 7837
rect 17678 7828 17684 7840
rect 17736 7828 17742 7880
rect 21634 7828 21640 7880
rect 21692 7868 21698 7880
rect 21910 7868 21916 7880
rect 21692 7840 21916 7868
rect 21692 7828 21698 7840
rect 21910 7828 21916 7840
rect 21968 7868 21974 7880
rect 22005 7871 22063 7877
rect 22005 7868 22017 7871
rect 21968 7840 22017 7868
rect 21968 7828 21974 7840
rect 22005 7837 22017 7840
rect 22051 7837 22063 7871
rect 22005 7831 22063 7837
rect 24029 7871 24087 7877
rect 24029 7837 24041 7871
rect 24075 7868 24087 7871
rect 25406 7868 25412 7880
rect 24075 7840 25412 7868
rect 24075 7837 24087 7840
rect 24029 7831 24087 7837
rect 25406 7828 25412 7840
rect 25464 7828 25470 7880
rect 27154 7868 27160 7880
rect 27115 7840 27160 7868
rect 27154 7828 27160 7840
rect 27212 7828 27218 7880
rect 28074 7868 28080 7880
rect 28035 7840 28080 7868
rect 28074 7828 28080 7840
rect 28132 7828 28138 7880
rect 32950 7868 32956 7880
rect 32911 7840 32956 7868
rect 32950 7828 32956 7840
rect 33008 7828 33014 7880
rect 35912 7877 35940 7908
rect 36446 7896 36452 7908
rect 36504 7896 36510 7948
rect 35897 7871 35955 7877
rect 35897 7837 35909 7871
rect 35943 7837 35955 7871
rect 35897 7831 35955 7837
rect 35986 7828 35992 7880
rect 36044 7868 36050 7880
rect 36081 7871 36139 7877
rect 36081 7868 36093 7871
rect 36044 7840 36093 7868
rect 36044 7828 36050 7840
rect 36081 7837 36093 7840
rect 36127 7837 36139 7871
rect 36081 7831 36139 7837
rect 6822 7760 6828 7812
rect 6880 7800 6886 7812
rect 7101 7803 7159 7809
rect 7101 7800 7113 7803
rect 6880 7772 7113 7800
rect 6880 7760 6886 7772
rect 7101 7769 7113 7772
rect 7147 7800 7159 7803
rect 8202 7800 8208 7812
rect 7147 7772 8208 7800
rect 7147 7769 7159 7772
rect 7101 7763 7159 7769
rect 8202 7760 8208 7772
rect 8260 7760 8266 7812
rect 16206 7800 16212 7812
rect 16167 7772 16212 7800
rect 16206 7760 16212 7772
rect 16264 7760 16270 7812
rect 24946 7800 24952 7812
rect 24907 7772 24952 7800
rect 24946 7760 24952 7772
rect 25004 7760 25010 7812
rect 34790 7760 34796 7812
rect 34848 7800 34854 7812
rect 35529 7803 35587 7809
rect 35529 7800 35541 7803
rect 34848 7772 35541 7800
rect 34848 7760 34854 7772
rect 35529 7769 35541 7772
rect 35575 7769 35587 7803
rect 35529 7763 35587 7769
rect 1854 7732 1860 7744
rect 1815 7704 1860 7732
rect 1854 7692 1860 7704
rect 1912 7692 1918 7744
rect 4338 7732 4344 7744
rect 4299 7704 4344 7732
rect 4338 7692 4344 7704
rect 4396 7692 4402 7744
rect 6086 7732 6092 7744
rect 6047 7704 6092 7732
rect 6086 7692 6092 7704
rect 6144 7692 6150 7744
rect 6454 7692 6460 7744
rect 6512 7732 6518 7744
rect 6641 7735 6699 7741
rect 6641 7732 6653 7735
rect 6512 7704 6653 7732
rect 6512 7692 6518 7704
rect 6641 7701 6653 7704
rect 6687 7701 6699 7735
rect 6641 7695 6699 7701
rect 7006 7692 7012 7744
rect 7064 7732 7070 7744
rect 7285 7735 7343 7741
rect 7285 7732 7297 7735
rect 7064 7704 7297 7732
rect 7064 7692 7070 7704
rect 7285 7701 7297 7704
rect 7331 7701 7343 7735
rect 9766 7732 9772 7744
rect 9727 7704 9772 7732
rect 7285 7695 7343 7701
rect 9766 7692 9772 7704
rect 9824 7692 9830 7744
rect 14090 7692 14096 7744
rect 14148 7732 14154 7744
rect 14277 7735 14335 7741
rect 14277 7732 14289 7735
rect 14148 7704 14289 7732
rect 14148 7692 14154 7704
rect 14277 7701 14289 7704
rect 14323 7732 14335 7735
rect 14642 7732 14648 7744
rect 14323 7704 14648 7732
rect 14323 7701 14335 7704
rect 14277 7695 14335 7701
rect 14642 7692 14648 7704
rect 14700 7692 14706 7744
rect 17586 7692 17592 7744
rect 17644 7732 17650 7744
rect 19061 7735 19119 7741
rect 19061 7732 19073 7735
rect 17644 7704 19073 7732
rect 17644 7692 17650 7704
rect 19061 7701 19073 7704
rect 19107 7732 19119 7735
rect 19242 7732 19248 7744
rect 19107 7704 19248 7732
rect 19107 7701 19119 7704
rect 19061 7695 19119 7701
rect 19242 7692 19248 7704
rect 19300 7692 19306 7744
rect 21358 7692 21364 7744
rect 21416 7732 21422 7744
rect 21453 7735 21511 7741
rect 21453 7732 21465 7735
rect 21416 7704 21465 7732
rect 21416 7692 21422 7704
rect 21453 7701 21465 7704
rect 21499 7701 21511 7735
rect 23382 7732 23388 7744
rect 23343 7704 23388 7732
rect 21453 7695 21511 7701
rect 23382 7692 23388 7704
rect 23440 7692 23446 7744
rect 32861 7735 32919 7741
rect 32861 7701 32873 7735
rect 32907 7732 32919 7735
rect 32950 7732 32956 7744
rect 32907 7704 32956 7732
rect 32907 7701 32919 7704
rect 32861 7695 32919 7701
rect 32950 7692 32956 7704
rect 33008 7732 33014 7744
rect 33134 7732 33140 7744
rect 33008 7704 33140 7732
rect 33008 7692 33014 7704
rect 33134 7692 33140 7704
rect 33192 7692 33198 7744
rect 34974 7732 34980 7744
rect 34935 7704 34980 7732
rect 34974 7692 34980 7704
rect 35032 7692 35038 7744
rect 35250 7732 35256 7744
rect 35211 7704 35256 7732
rect 35250 7692 35256 7704
rect 35308 7732 35314 7744
rect 35618 7732 35624 7744
rect 35308 7704 35624 7732
rect 35308 7692 35314 7704
rect 35618 7692 35624 7704
rect 35676 7692 35682 7744
rect 1104 7642 38824 7664
rect 1104 7590 7648 7642
rect 7700 7590 7712 7642
rect 7764 7590 7776 7642
rect 7828 7590 7840 7642
rect 7892 7590 20982 7642
rect 21034 7590 21046 7642
rect 21098 7590 21110 7642
rect 21162 7590 21174 7642
rect 21226 7590 34315 7642
rect 34367 7590 34379 7642
rect 34431 7590 34443 7642
rect 34495 7590 34507 7642
rect 34559 7590 38824 7642
rect 1104 7568 38824 7590
rect 2682 7488 2688 7540
rect 2740 7528 2746 7540
rect 3237 7531 3295 7537
rect 3237 7528 3249 7531
rect 2740 7500 3249 7528
rect 2740 7488 2746 7500
rect 3237 7497 3249 7500
rect 3283 7497 3295 7531
rect 3237 7491 3295 7497
rect 5350 7488 5356 7540
rect 5408 7528 5414 7540
rect 5445 7531 5503 7537
rect 5445 7528 5457 7531
rect 5408 7500 5457 7528
rect 5408 7488 5414 7500
rect 5445 7497 5457 7500
rect 5491 7497 5503 7531
rect 5445 7491 5503 7497
rect 5534 7488 5540 7540
rect 5592 7528 5598 7540
rect 6638 7528 6644 7540
rect 5592 7500 6644 7528
rect 5592 7488 5598 7500
rect 6638 7488 6644 7500
rect 6696 7488 6702 7540
rect 7374 7488 7380 7540
rect 7432 7528 7438 7540
rect 8110 7528 8116 7540
rect 7432 7500 8116 7528
rect 7432 7488 7438 7500
rect 8110 7488 8116 7500
rect 8168 7488 8174 7540
rect 9306 7528 9312 7540
rect 9267 7500 9312 7528
rect 9306 7488 9312 7500
rect 9364 7488 9370 7540
rect 11882 7528 11888 7540
rect 11843 7500 11888 7528
rect 11882 7488 11888 7500
rect 11940 7488 11946 7540
rect 11974 7488 11980 7540
rect 12032 7528 12038 7540
rect 12713 7531 12771 7537
rect 12713 7528 12725 7531
rect 12032 7500 12725 7528
rect 12032 7488 12038 7500
rect 12713 7497 12725 7500
rect 12759 7497 12771 7531
rect 15930 7528 15936 7540
rect 15891 7500 15936 7528
rect 12713 7491 12771 7497
rect 15930 7488 15936 7500
rect 15988 7488 15994 7540
rect 16482 7528 16488 7540
rect 16443 7500 16488 7528
rect 16482 7488 16488 7500
rect 16540 7488 16546 7540
rect 19794 7488 19800 7540
rect 19852 7528 19858 7540
rect 19981 7531 20039 7537
rect 19981 7528 19993 7531
rect 19852 7500 19993 7528
rect 19852 7488 19858 7500
rect 19981 7497 19993 7500
rect 20027 7497 20039 7531
rect 21542 7528 21548 7540
rect 21503 7500 21548 7528
rect 19981 7491 20039 7497
rect 21542 7488 21548 7500
rect 21600 7488 21606 7540
rect 22097 7531 22155 7537
rect 22097 7497 22109 7531
rect 22143 7528 22155 7531
rect 22370 7528 22376 7540
rect 22143 7500 22376 7528
rect 22143 7497 22155 7500
rect 22097 7491 22155 7497
rect 22370 7488 22376 7500
rect 22428 7488 22434 7540
rect 23658 7488 23664 7540
rect 23716 7528 23722 7540
rect 23845 7531 23903 7537
rect 23845 7528 23857 7531
rect 23716 7500 23857 7528
rect 23716 7488 23722 7500
rect 23845 7497 23857 7500
rect 23891 7497 23903 7531
rect 23845 7491 23903 7497
rect 1949 7463 2007 7469
rect 1949 7429 1961 7463
rect 1995 7460 2007 7463
rect 2130 7460 2136 7472
rect 1995 7432 2136 7460
rect 1995 7429 2007 7432
rect 1949 7423 2007 7429
rect 2130 7420 2136 7432
rect 2188 7420 2194 7472
rect 2314 7420 2320 7472
rect 2372 7460 2378 7472
rect 3142 7460 3148 7472
rect 2372 7432 3148 7460
rect 2372 7420 2378 7432
rect 3142 7420 3148 7432
rect 3200 7420 3206 7472
rect 10873 7463 10931 7469
rect 10873 7429 10885 7463
rect 10919 7460 10931 7463
rect 10962 7460 10968 7472
rect 10919 7432 10968 7460
rect 10919 7429 10931 7432
rect 10873 7423 10931 7429
rect 10962 7420 10968 7432
rect 11020 7420 11026 7472
rect 13630 7420 13636 7472
rect 13688 7460 13694 7472
rect 14277 7463 14335 7469
rect 14277 7460 14289 7463
rect 13688 7432 14289 7460
rect 13688 7420 13694 7432
rect 14277 7429 14289 7432
rect 14323 7429 14335 7463
rect 14277 7423 14335 7429
rect 2774 7392 2780 7404
rect 2240 7364 2780 7392
rect 2240 7265 2268 7364
rect 2774 7352 2780 7364
rect 2832 7352 2838 7404
rect 6086 7352 6092 7404
rect 6144 7392 6150 7404
rect 6273 7395 6331 7401
rect 6273 7392 6285 7395
rect 6144 7364 6285 7392
rect 6144 7352 6150 7364
rect 6273 7361 6285 7364
rect 6319 7392 6331 7395
rect 12158 7392 12164 7404
rect 6319 7364 7512 7392
rect 12119 7364 12164 7392
rect 6319 7361 6331 7364
rect 6273 7355 6331 7361
rect 7484 7336 7512 7364
rect 12158 7352 12164 7364
rect 12216 7352 12222 7404
rect 12529 7395 12587 7401
rect 12529 7361 12541 7395
rect 12575 7392 12587 7395
rect 13173 7395 13231 7401
rect 13173 7392 13185 7395
rect 12575 7364 13185 7392
rect 12575 7361 12587 7364
rect 12529 7355 12587 7361
rect 13173 7361 13185 7364
rect 13219 7392 13231 7395
rect 13354 7392 13360 7404
rect 13219 7364 13360 7392
rect 13219 7361 13231 7364
rect 13173 7355 13231 7361
rect 13354 7352 13360 7364
rect 13412 7352 13418 7404
rect 14090 7392 14096 7404
rect 14003 7364 14096 7392
rect 14090 7352 14096 7364
rect 14148 7392 14154 7404
rect 14734 7392 14740 7404
rect 14148 7364 14740 7392
rect 14148 7352 14154 7364
rect 14734 7352 14740 7364
rect 14792 7352 14798 7404
rect 16206 7352 16212 7404
rect 16264 7392 16270 7404
rect 16853 7395 16911 7401
rect 16853 7392 16865 7395
rect 16264 7364 16865 7392
rect 16264 7352 16270 7364
rect 16853 7361 16865 7364
rect 16899 7361 16911 7395
rect 16853 7355 16911 7361
rect 17037 7395 17095 7401
rect 17037 7361 17049 7395
rect 17083 7392 17095 7395
rect 17126 7392 17132 7404
rect 17083 7364 17132 7392
rect 17083 7361 17095 7364
rect 17037 7355 17095 7361
rect 17126 7352 17132 7364
rect 17184 7392 17190 7404
rect 17586 7392 17592 7404
rect 17184 7364 17592 7392
rect 17184 7352 17190 7364
rect 17586 7352 17592 7364
rect 17644 7352 17650 7404
rect 20806 7352 20812 7404
rect 20864 7392 20870 7404
rect 21821 7395 21879 7401
rect 21821 7392 21833 7395
rect 20864 7364 21833 7392
rect 20864 7352 20870 7364
rect 21821 7361 21833 7364
rect 21867 7361 21879 7395
rect 23860 7392 23888 7491
rect 25406 7488 25412 7540
rect 25464 7528 25470 7540
rect 26605 7531 26663 7537
rect 26605 7528 26617 7531
rect 25464 7500 26617 7528
rect 25464 7488 25470 7500
rect 26605 7497 26617 7500
rect 26651 7497 26663 7531
rect 26605 7491 26663 7497
rect 27982 7488 27988 7540
rect 28040 7528 28046 7540
rect 28629 7531 28687 7537
rect 28629 7528 28641 7531
rect 28040 7500 28641 7528
rect 28040 7488 28046 7500
rect 28629 7497 28641 7500
rect 28675 7497 28687 7531
rect 28629 7491 28687 7497
rect 28994 7488 29000 7540
rect 29052 7528 29058 7540
rect 29365 7531 29423 7537
rect 29365 7528 29377 7531
rect 29052 7500 29377 7528
rect 29052 7488 29058 7500
rect 29365 7497 29377 7500
rect 29411 7497 29423 7531
rect 32398 7528 32404 7540
rect 32359 7500 32404 7528
rect 29365 7491 29423 7497
rect 32398 7488 32404 7500
rect 32456 7528 32462 7540
rect 34609 7531 34667 7537
rect 34609 7528 34621 7531
rect 32456 7500 34621 7528
rect 32456 7488 32462 7500
rect 34609 7497 34621 7500
rect 34655 7528 34667 7531
rect 35986 7528 35992 7540
rect 34655 7500 35992 7528
rect 34655 7497 34667 7500
rect 34609 7491 34667 7497
rect 35986 7488 35992 7500
rect 36044 7528 36050 7540
rect 36633 7531 36691 7537
rect 36633 7528 36645 7531
rect 36044 7500 36645 7528
rect 36044 7488 36050 7500
rect 36633 7497 36645 7500
rect 36679 7497 36691 7531
rect 36633 7491 36691 7497
rect 26326 7460 26332 7472
rect 26287 7432 26332 7460
rect 26326 7420 26332 7432
rect 26384 7420 26390 7472
rect 29086 7460 29092 7472
rect 29047 7432 29092 7460
rect 29086 7420 29092 7432
rect 29144 7420 29150 7472
rect 30929 7463 30987 7469
rect 30929 7429 30941 7463
rect 30975 7460 30987 7463
rect 31754 7460 31760 7472
rect 30975 7432 31760 7460
rect 30975 7429 30987 7432
rect 30929 7423 30987 7429
rect 31754 7420 31760 7432
rect 31812 7420 31818 7472
rect 32769 7463 32827 7469
rect 32769 7429 32781 7463
rect 32815 7460 32827 7463
rect 32858 7460 32864 7472
rect 32815 7432 32864 7460
rect 32815 7429 32827 7432
rect 32769 7423 32827 7429
rect 32858 7420 32864 7432
rect 32916 7420 32922 7472
rect 33318 7460 33324 7472
rect 33279 7432 33324 7460
rect 33318 7420 33324 7432
rect 33376 7420 33382 7472
rect 33594 7420 33600 7472
rect 33652 7460 33658 7472
rect 33652 7432 33916 7460
rect 33652 7420 33658 7432
rect 24029 7395 24087 7401
rect 24029 7392 24041 7395
rect 23860 7364 24041 7392
rect 21821 7355 21879 7361
rect 24029 7361 24041 7364
rect 24075 7361 24087 7395
rect 26050 7392 26056 7404
rect 25963 7364 26056 7392
rect 24029 7355 24087 7361
rect 4338 7333 4344 7336
rect 3973 7327 4031 7333
rect 3973 7293 3985 7327
rect 4019 7324 4031 7327
rect 4065 7327 4123 7333
rect 4065 7324 4077 7327
rect 4019 7296 4077 7324
rect 4019 7293 4031 7296
rect 3973 7287 4031 7293
rect 4065 7293 4077 7296
rect 4111 7293 4123 7327
rect 4332 7324 4344 7333
rect 4299 7296 4344 7324
rect 4065 7287 4123 7293
rect 4332 7287 4344 7296
rect 1765 7259 1823 7265
rect 1765 7225 1777 7259
rect 1811 7256 1823 7259
rect 2225 7259 2283 7265
rect 2225 7256 2237 7259
rect 1811 7228 2237 7256
rect 1811 7225 1823 7228
rect 1765 7219 1823 7225
rect 2225 7225 2237 7228
rect 2271 7225 2283 7259
rect 2498 7256 2504 7268
rect 2459 7228 2504 7256
rect 2225 7219 2283 7225
rect 2498 7216 2504 7228
rect 2556 7256 2562 7268
rect 2958 7256 2964 7268
rect 2556 7228 2964 7256
rect 2556 7216 2562 7228
rect 2958 7216 2964 7228
rect 3016 7216 3022 7268
rect 4080 7256 4108 7287
rect 4338 7284 4344 7287
rect 4396 7284 4402 7336
rect 7374 7324 7380 7336
rect 7335 7296 7380 7324
rect 7374 7284 7380 7296
rect 7432 7284 7438 7336
rect 7466 7284 7472 7336
rect 7524 7324 7530 7336
rect 7644 7327 7702 7333
rect 7644 7324 7656 7327
rect 7524 7296 7656 7324
rect 7524 7284 7530 7296
rect 7644 7293 7656 7296
rect 7690 7324 7702 7327
rect 8018 7324 8024 7336
rect 7690 7296 8024 7324
rect 7690 7293 7702 7296
rect 7644 7287 7702 7293
rect 8018 7284 8024 7296
rect 8076 7284 8082 7336
rect 11238 7284 11244 7336
rect 11296 7324 11302 7336
rect 11425 7327 11483 7333
rect 11425 7324 11437 7327
rect 11296 7296 11437 7324
rect 11296 7284 11302 7296
rect 11425 7293 11437 7296
rect 11471 7324 11483 7327
rect 15565 7327 15623 7333
rect 11471 7296 13768 7324
rect 11471 7293 11483 7296
rect 11425 7287 11483 7293
rect 4706 7256 4712 7268
rect 4080 7228 4712 7256
rect 4706 7216 4712 7228
rect 4764 7216 4770 7268
rect 6822 7216 6828 7268
rect 6880 7256 6886 7268
rect 6880 7228 8800 7256
rect 6880 7216 6886 7228
rect 2409 7191 2467 7197
rect 2409 7157 2421 7191
rect 2455 7188 2467 7191
rect 2590 7188 2596 7200
rect 2455 7160 2596 7188
rect 2455 7157 2467 7160
rect 2409 7151 2467 7157
rect 2590 7148 2596 7160
rect 2648 7148 2654 7200
rect 2869 7191 2927 7197
rect 2869 7157 2881 7191
rect 2915 7188 2927 7191
rect 3142 7188 3148 7200
rect 2915 7160 3148 7188
rect 2915 7157 2927 7160
rect 2869 7151 2927 7157
rect 3142 7148 3148 7160
rect 3200 7148 3206 7200
rect 6638 7148 6644 7200
rect 6696 7188 6702 7200
rect 7006 7188 7012 7200
rect 6696 7160 7012 7188
rect 6696 7148 6702 7160
rect 7006 7148 7012 7160
rect 7064 7148 7070 7200
rect 7285 7191 7343 7197
rect 7285 7157 7297 7191
rect 7331 7188 7343 7191
rect 7558 7188 7564 7200
rect 7331 7160 7564 7188
rect 7331 7157 7343 7160
rect 7285 7151 7343 7157
rect 7558 7148 7564 7160
rect 7616 7148 7622 7200
rect 8772 7197 8800 7228
rect 11054 7216 11060 7268
rect 11112 7256 11118 7268
rect 11149 7259 11207 7265
rect 11149 7256 11161 7259
rect 11112 7228 11161 7256
rect 11112 7216 11118 7228
rect 11149 7225 11161 7228
rect 11195 7225 11207 7259
rect 11330 7256 11336 7268
rect 11291 7228 11336 7256
rect 11149 7219 11207 7225
rect 11330 7216 11336 7228
rect 11388 7216 11394 7268
rect 12250 7216 12256 7268
rect 12308 7256 12314 7268
rect 12529 7259 12587 7265
rect 12529 7256 12541 7259
rect 12308 7228 12541 7256
rect 12308 7216 12314 7228
rect 12529 7225 12541 7228
rect 12575 7225 12587 7259
rect 13170 7256 13176 7268
rect 13131 7228 13176 7256
rect 12529 7219 12587 7225
rect 13170 7216 13176 7228
rect 13228 7216 13234 7268
rect 13262 7216 13268 7268
rect 13320 7256 13326 7268
rect 13740 7265 13768 7296
rect 15565 7293 15577 7327
rect 15611 7324 15623 7327
rect 16390 7324 16396 7336
rect 15611 7296 16396 7324
rect 15611 7293 15623 7296
rect 15565 7287 15623 7293
rect 16390 7284 16396 7296
rect 16448 7324 16454 7336
rect 16448 7296 16988 7324
rect 16448 7284 16454 7296
rect 13725 7259 13783 7265
rect 13320 7228 13365 7256
rect 13320 7216 13326 7228
rect 13725 7225 13737 7259
rect 13771 7256 13783 7259
rect 14826 7256 14832 7268
rect 13771 7228 14832 7256
rect 13771 7225 13783 7228
rect 13725 7219 13783 7225
rect 14826 7216 14832 7228
rect 14884 7216 14890 7268
rect 16960 7265 16988 7296
rect 17678 7284 17684 7336
rect 17736 7324 17742 7336
rect 17773 7327 17831 7333
rect 17773 7324 17785 7327
rect 17736 7296 17785 7324
rect 17736 7284 17742 7296
rect 17773 7293 17785 7296
rect 17819 7324 17831 7327
rect 18049 7327 18107 7333
rect 18049 7324 18061 7327
rect 17819 7296 18061 7324
rect 17819 7293 17831 7296
rect 17773 7287 17831 7293
rect 18049 7293 18061 7296
rect 18095 7324 18107 7327
rect 18874 7324 18880 7336
rect 18095 7296 18880 7324
rect 18095 7293 18107 7296
rect 18049 7287 18107 7293
rect 18874 7284 18880 7296
rect 18932 7284 18938 7336
rect 21836 7324 21864 7355
rect 26050 7352 26056 7364
rect 26108 7392 26114 7404
rect 27062 7392 27068 7404
rect 26108 7364 27068 7392
rect 26108 7352 26114 7364
rect 27062 7352 27068 7364
rect 27120 7352 27126 7404
rect 29178 7352 29184 7404
rect 29236 7392 29242 7404
rect 29917 7395 29975 7401
rect 29917 7392 29929 7395
rect 29236 7364 29929 7392
rect 29236 7352 29242 7364
rect 29917 7361 29929 7364
rect 29963 7392 29975 7395
rect 30653 7395 30711 7401
rect 30653 7392 30665 7395
rect 29963 7364 30665 7392
rect 29963 7361 29975 7364
rect 29917 7355 29975 7361
rect 30653 7361 30665 7364
rect 30699 7361 30711 7395
rect 30653 7355 30711 7361
rect 31389 7395 31447 7401
rect 31389 7361 31401 7395
rect 31435 7392 31447 7395
rect 31570 7392 31576 7404
rect 31435 7364 31576 7392
rect 31435 7361 31447 7364
rect 31389 7355 31447 7361
rect 31570 7352 31576 7364
rect 31628 7352 31634 7404
rect 33888 7401 33916 7432
rect 33873 7395 33931 7401
rect 33873 7361 33885 7395
rect 33919 7392 33931 7395
rect 33962 7392 33968 7404
rect 33919 7364 33968 7392
rect 33919 7361 33931 7364
rect 33873 7355 33931 7361
rect 33962 7352 33968 7364
rect 34020 7392 34026 7404
rect 34241 7395 34299 7401
rect 34241 7392 34253 7395
rect 34020 7364 34253 7392
rect 34020 7352 34026 7364
rect 34241 7361 34253 7364
rect 34287 7361 34299 7395
rect 34241 7355 34299 7361
rect 22373 7327 22431 7333
rect 22373 7324 22385 7327
rect 21836 7296 22385 7324
rect 22373 7293 22385 7296
rect 22419 7324 22431 7327
rect 24118 7324 24124 7336
rect 22419 7296 24124 7324
rect 22419 7293 22431 7296
rect 22373 7287 22431 7293
rect 24118 7284 24124 7296
rect 24176 7284 24182 7336
rect 28074 7284 28080 7336
rect 28132 7324 28138 7336
rect 29641 7327 29699 7333
rect 29641 7324 29653 7327
rect 28132 7296 29653 7324
rect 28132 7284 28138 7296
rect 29641 7293 29653 7296
rect 29687 7324 29699 7327
rect 30285 7327 30343 7333
rect 30285 7324 30297 7327
rect 29687 7296 30297 7324
rect 29687 7293 29699 7296
rect 29641 7287 29699 7293
rect 30285 7293 30297 7296
rect 30331 7293 30343 7327
rect 30285 7287 30343 7293
rect 33137 7327 33195 7333
rect 33137 7293 33149 7327
rect 33183 7324 33195 7327
rect 33226 7324 33232 7336
rect 33183 7296 33232 7324
rect 33183 7293 33195 7296
rect 33137 7287 33195 7293
rect 33226 7284 33232 7296
rect 33284 7324 33290 7336
rect 33597 7327 33655 7333
rect 33597 7324 33609 7327
rect 33284 7296 33609 7324
rect 33284 7284 33290 7296
rect 33597 7293 33609 7296
rect 33643 7293 33655 7327
rect 33597 7287 33655 7293
rect 35066 7284 35072 7336
rect 35124 7324 35130 7336
rect 35253 7327 35311 7333
rect 35253 7324 35265 7327
rect 35124 7296 35265 7324
rect 35124 7284 35130 7296
rect 35253 7293 35265 7296
rect 35299 7293 35311 7327
rect 35253 7287 35311 7293
rect 36078 7284 36084 7336
rect 36136 7324 36142 7336
rect 37185 7327 37243 7333
rect 37185 7324 37197 7327
rect 36136 7296 37197 7324
rect 36136 7284 36142 7296
rect 37185 7293 37197 7296
rect 37231 7293 37243 7327
rect 37185 7287 37243 7293
rect 16945 7259 17003 7265
rect 16945 7225 16957 7259
rect 16991 7225 17003 7259
rect 16945 7219 17003 7225
rect 18316 7259 18374 7265
rect 18316 7225 18328 7259
rect 18362 7256 18374 7259
rect 18506 7256 18512 7268
rect 18362 7228 18512 7256
rect 18362 7225 18374 7228
rect 18316 7219 18374 7225
rect 18506 7216 18512 7228
rect 18564 7216 18570 7268
rect 22649 7259 22707 7265
rect 22649 7225 22661 7259
rect 22695 7256 22707 7259
rect 22738 7256 22744 7268
rect 22695 7228 22744 7256
rect 22695 7225 22707 7228
rect 22649 7219 22707 7225
rect 22738 7216 22744 7228
rect 22796 7216 22802 7268
rect 24274 7259 24332 7265
rect 24274 7256 24286 7259
rect 23400 7228 24286 7256
rect 8757 7191 8815 7197
rect 8757 7157 8769 7191
rect 8803 7157 8815 7191
rect 9674 7188 9680 7200
rect 9635 7160 9680 7188
rect 8757 7151 8815 7157
rect 9674 7148 9680 7160
rect 9732 7148 9738 7200
rect 10042 7188 10048 7200
rect 10003 7160 10048 7188
rect 10042 7148 10048 7160
rect 10100 7148 10106 7200
rect 10134 7148 10140 7200
rect 10192 7188 10198 7200
rect 10689 7191 10747 7197
rect 10689 7188 10701 7191
rect 10192 7160 10701 7188
rect 10192 7148 10198 7160
rect 10689 7157 10701 7160
rect 10735 7188 10747 7191
rect 11348 7188 11376 7216
rect 23400 7200 23428 7228
rect 24274 7225 24286 7228
rect 24320 7225 24332 7259
rect 27154 7256 27160 7268
rect 27115 7228 27160 7256
rect 24274 7219 24332 7225
rect 27154 7216 27160 7228
rect 27212 7256 27218 7268
rect 27893 7259 27951 7265
rect 27893 7256 27905 7259
rect 27212 7228 27905 7256
rect 27212 7216 27218 7228
rect 27893 7225 27905 7228
rect 27939 7225 27951 7259
rect 27893 7219 27951 7225
rect 29086 7216 29092 7268
rect 29144 7256 29150 7268
rect 29822 7256 29828 7268
rect 29144 7228 29828 7256
rect 29144 7216 29150 7228
rect 29822 7216 29828 7228
rect 29880 7216 29886 7268
rect 31478 7256 31484 7268
rect 31439 7228 31484 7256
rect 31478 7216 31484 7228
rect 31536 7216 31542 7268
rect 34606 7216 34612 7268
rect 34664 7256 34670 7268
rect 34974 7256 34980 7268
rect 34664 7228 34980 7256
rect 34664 7216 34670 7228
rect 34974 7216 34980 7228
rect 35032 7256 35038 7268
rect 35498 7259 35556 7265
rect 35498 7256 35510 7259
rect 35032 7228 35510 7256
rect 35032 7216 35038 7228
rect 35498 7225 35510 7228
rect 35544 7256 35556 7259
rect 35710 7256 35716 7268
rect 35544 7228 35716 7256
rect 35544 7225 35556 7228
rect 35498 7219 35556 7225
rect 35710 7216 35716 7228
rect 35768 7216 35774 7268
rect 14734 7188 14740 7200
rect 10735 7160 11376 7188
rect 14695 7160 14740 7188
rect 10735 7157 10747 7160
rect 10689 7151 10747 7157
rect 14734 7148 14740 7160
rect 14792 7148 14798 7200
rect 16206 7188 16212 7200
rect 16167 7160 16212 7188
rect 16206 7148 16212 7160
rect 16264 7148 16270 7200
rect 19426 7188 19432 7200
rect 19387 7160 19432 7188
rect 19426 7148 19432 7160
rect 19484 7148 19490 7200
rect 20898 7188 20904 7200
rect 20859 7160 20904 7188
rect 20898 7148 20904 7160
rect 20956 7148 20962 7200
rect 22554 7188 22560 7200
rect 22467 7160 22560 7188
rect 22554 7148 22560 7160
rect 22612 7188 22618 7200
rect 23017 7191 23075 7197
rect 23017 7188 23029 7191
rect 22612 7160 23029 7188
rect 22612 7148 22618 7160
rect 23017 7157 23029 7160
rect 23063 7157 23075 7191
rect 23382 7188 23388 7200
rect 23343 7160 23388 7188
rect 23017 7151 23075 7157
rect 23382 7148 23388 7160
rect 23440 7148 23446 7200
rect 25406 7188 25412 7200
rect 25367 7160 25412 7188
rect 25406 7148 25412 7160
rect 25464 7148 25470 7200
rect 27062 7188 27068 7200
rect 27023 7160 27068 7188
rect 27062 7148 27068 7160
rect 27120 7188 27126 7200
rect 27522 7188 27528 7200
rect 27120 7160 27528 7188
rect 27120 7148 27126 7160
rect 27522 7148 27528 7160
rect 27580 7148 27586 7200
rect 27982 7148 27988 7200
rect 28040 7188 28046 7200
rect 28077 7191 28135 7197
rect 28077 7188 28089 7191
rect 28040 7160 28089 7188
rect 28040 7148 28046 7160
rect 28077 7157 28089 7160
rect 28123 7157 28135 7191
rect 31386 7188 31392 7200
rect 31347 7160 31392 7188
rect 28077 7151 28135 7157
rect 31386 7148 31392 7160
rect 31444 7188 31450 7200
rect 31849 7191 31907 7197
rect 31849 7188 31861 7191
rect 31444 7160 31861 7188
rect 31444 7148 31450 7160
rect 31849 7157 31861 7160
rect 31895 7157 31907 7191
rect 31849 7151 31907 7157
rect 33134 7148 33140 7200
rect 33192 7188 33198 7200
rect 33781 7191 33839 7197
rect 33781 7188 33793 7191
rect 33192 7160 33793 7188
rect 33192 7148 33198 7160
rect 33781 7157 33793 7160
rect 33827 7157 33839 7191
rect 35066 7188 35072 7200
rect 35027 7160 35072 7188
rect 33781 7151 33839 7157
rect 35066 7148 35072 7160
rect 35124 7148 35130 7200
rect 1104 7098 38824 7120
rect 1104 7046 14315 7098
rect 14367 7046 14379 7098
rect 14431 7046 14443 7098
rect 14495 7046 14507 7098
rect 14559 7046 27648 7098
rect 27700 7046 27712 7098
rect 27764 7046 27776 7098
rect 27828 7046 27840 7098
rect 27892 7046 38824 7098
rect 1104 7024 38824 7046
rect 2590 6984 2596 6996
rect 2551 6956 2596 6984
rect 2590 6944 2596 6956
rect 2648 6944 2654 6996
rect 4246 6984 4252 6996
rect 4207 6956 4252 6984
rect 4246 6944 4252 6956
rect 4304 6944 4310 6996
rect 5074 6984 5080 6996
rect 5035 6956 5080 6984
rect 5074 6944 5080 6956
rect 5132 6944 5138 6996
rect 6917 6987 6975 6993
rect 6917 6953 6929 6987
rect 6963 6984 6975 6987
rect 7466 6984 7472 6996
rect 6963 6956 7472 6984
rect 6963 6953 6975 6956
rect 6917 6947 6975 6953
rect 7466 6944 7472 6956
rect 7524 6944 7530 6996
rect 8110 6984 8116 6996
rect 8071 6956 8116 6984
rect 8110 6944 8116 6956
rect 8168 6944 8174 6996
rect 11238 6984 11244 6996
rect 11199 6956 11244 6984
rect 11238 6944 11244 6956
rect 11296 6944 11302 6996
rect 13170 6944 13176 6996
rect 13228 6984 13234 6996
rect 13633 6987 13691 6993
rect 13633 6984 13645 6987
rect 13228 6956 13645 6984
rect 13228 6944 13234 6956
rect 13633 6953 13645 6956
rect 13679 6953 13691 6987
rect 13633 6947 13691 6953
rect 14461 6987 14519 6993
rect 14461 6953 14473 6987
rect 14507 6984 14519 6987
rect 14826 6984 14832 6996
rect 14507 6956 14832 6984
rect 14507 6953 14519 6956
rect 14461 6947 14519 6953
rect 14826 6944 14832 6956
rect 14884 6944 14890 6996
rect 16485 6987 16543 6993
rect 16485 6953 16497 6987
rect 16531 6984 16543 6987
rect 17126 6984 17132 6996
rect 16531 6956 17132 6984
rect 16531 6953 16543 6956
rect 16485 6947 16543 6953
rect 17126 6944 17132 6956
rect 17184 6944 17190 6996
rect 19794 6984 19800 6996
rect 19755 6956 19800 6984
rect 19794 6944 19800 6956
rect 19852 6944 19858 6996
rect 25041 6987 25099 6993
rect 25041 6984 25053 6987
rect 21376 6956 25053 6984
rect 2130 6916 2136 6928
rect 2091 6888 2136 6916
rect 2130 6876 2136 6888
rect 2188 6876 2194 6928
rect 5350 6916 5356 6928
rect 3988 6888 5356 6916
rect 1854 6808 1860 6860
rect 1912 6848 1918 6860
rect 1949 6851 2007 6857
rect 1949 6848 1961 6851
rect 1912 6820 1961 6848
rect 1912 6808 1918 6820
rect 1949 6817 1961 6820
rect 1995 6817 2007 6851
rect 2148 6848 2176 6876
rect 3697 6851 3755 6857
rect 3697 6848 3709 6851
rect 2148 6820 3709 6848
rect 1949 6811 2007 6817
rect 3697 6817 3709 6820
rect 3743 6817 3755 6851
rect 3697 6811 3755 6817
rect 2222 6780 2228 6792
rect 2183 6752 2228 6780
rect 2222 6740 2228 6752
rect 2280 6780 2286 6792
rect 3421 6783 3479 6789
rect 3421 6780 3433 6783
rect 2280 6752 3433 6780
rect 2280 6740 2286 6752
rect 3421 6749 3433 6752
rect 3467 6780 3479 6783
rect 3510 6780 3516 6792
rect 3467 6752 3516 6780
rect 3467 6749 3479 6752
rect 3421 6743 3479 6749
rect 3510 6740 3516 6752
rect 3568 6780 3574 6792
rect 3988 6780 4016 6888
rect 5350 6876 5356 6888
rect 5408 6876 5414 6928
rect 5997 6919 6055 6925
rect 5997 6885 6009 6919
rect 6043 6885 6055 6919
rect 7561 6919 7619 6925
rect 7561 6916 7573 6919
rect 5997 6879 6055 6885
rect 7300 6888 7573 6916
rect 4065 6851 4123 6857
rect 4065 6817 4077 6851
rect 4111 6817 4123 6851
rect 4065 6811 4123 6817
rect 4080 6780 4108 6811
rect 5166 6808 5172 6860
rect 5224 6848 5230 6860
rect 6012 6848 6040 6879
rect 6638 6848 6644 6860
rect 5224 6820 6644 6848
rect 5224 6808 5230 6820
rect 6638 6808 6644 6820
rect 6696 6808 6702 6860
rect 7006 6808 7012 6860
rect 7064 6848 7070 6860
rect 7300 6848 7328 6888
rect 7561 6885 7573 6888
rect 7607 6885 7619 6919
rect 7561 6879 7619 6885
rect 10229 6919 10287 6925
rect 10229 6885 10241 6919
rect 10275 6916 10287 6919
rect 10502 6916 10508 6928
rect 10275 6888 10508 6916
rect 10275 6885 10287 6888
rect 10229 6879 10287 6885
rect 7064 6820 7328 6848
rect 7064 6808 7070 6820
rect 7374 6808 7380 6860
rect 7432 6848 7438 6860
rect 7653 6851 7711 6857
rect 7653 6848 7665 6851
rect 7432 6820 7665 6848
rect 7432 6808 7438 6820
rect 7653 6817 7665 6820
rect 7699 6817 7711 6851
rect 7653 6811 7711 6817
rect 9306 6808 9312 6860
rect 9364 6848 9370 6860
rect 10244 6848 10272 6879
rect 10502 6876 10508 6888
rect 10560 6876 10566 6928
rect 11054 6876 11060 6928
rect 11112 6876 11118 6928
rect 11882 6916 11888 6928
rect 11348 6888 11888 6916
rect 9364 6820 10272 6848
rect 10873 6851 10931 6857
rect 9364 6808 9370 6820
rect 10873 6817 10885 6851
rect 10919 6848 10931 6851
rect 11072 6848 11100 6876
rect 11348 6860 11376 6888
rect 11882 6876 11888 6888
rect 11940 6916 11946 6928
rect 12526 6916 12532 6928
rect 11940 6888 12532 6916
rect 11940 6876 11946 6888
rect 12526 6876 12532 6888
rect 12584 6876 12590 6928
rect 13262 6916 13268 6928
rect 13223 6888 13268 6916
rect 13262 6876 13268 6888
rect 13320 6876 13326 6928
rect 16666 6916 16672 6928
rect 16579 6888 16672 6916
rect 11330 6848 11336 6860
rect 10919 6820 11100 6848
rect 11243 6820 11336 6848
rect 10919 6817 10931 6820
rect 10873 6811 10931 6817
rect 11330 6808 11336 6820
rect 11388 6808 11394 6860
rect 11422 6808 11428 6860
rect 11480 6848 11486 6860
rect 11589 6851 11647 6857
rect 11589 6848 11601 6851
rect 11480 6820 11601 6848
rect 11480 6808 11486 6820
rect 11589 6817 11601 6820
rect 11635 6817 11647 6851
rect 13814 6848 13820 6860
rect 13775 6820 13820 6848
rect 11589 6811 11647 6817
rect 13814 6808 13820 6820
rect 13872 6808 13878 6860
rect 16117 6851 16175 6857
rect 16117 6817 16129 6851
rect 16163 6848 16175 6851
rect 16592 6848 16620 6888
rect 16666 6876 16672 6888
rect 16724 6916 16730 6928
rect 17862 6916 17868 6928
rect 16724 6888 17868 6916
rect 16724 6876 16730 6888
rect 17862 6876 17868 6888
rect 17920 6876 17926 6928
rect 20898 6916 20904 6928
rect 20640 6888 20904 6916
rect 16163 6820 16620 6848
rect 16163 6817 16175 6820
rect 16117 6811 16175 6817
rect 16850 6808 16856 6860
rect 16908 6848 16914 6860
rect 17017 6851 17075 6857
rect 17017 6848 17029 6851
rect 16908 6820 17029 6848
rect 16908 6808 16914 6820
rect 17017 6817 17029 6820
rect 17063 6817 17075 6851
rect 17017 6811 17075 6817
rect 18690 6808 18696 6860
rect 18748 6848 18754 6860
rect 19613 6851 19671 6857
rect 19613 6848 19625 6851
rect 18748 6820 19625 6848
rect 18748 6808 18754 6820
rect 19613 6817 19625 6820
rect 19659 6848 19671 6851
rect 20640 6848 20668 6888
rect 20898 6876 20904 6888
rect 20956 6876 20962 6928
rect 21266 6876 21272 6928
rect 21324 6916 21330 6928
rect 21376 6925 21404 6956
rect 25041 6953 25053 6956
rect 25087 6953 25099 6987
rect 25498 6984 25504 6996
rect 25459 6956 25504 6984
rect 25041 6947 25099 6953
rect 25498 6944 25504 6956
rect 25556 6944 25562 6996
rect 26329 6987 26387 6993
rect 26329 6953 26341 6987
rect 26375 6984 26387 6987
rect 27154 6984 27160 6996
rect 26375 6956 27160 6984
rect 26375 6953 26387 6956
rect 26329 6947 26387 6953
rect 27154 6944 27160 6956
rect 27212 6984 27218 6996
rect 28997 6987 29055 6993
rect 28997 6984 29009 6987
rect 27212 6956 29009 6984
rect 27212 6944 27218 6956
rect 28997 6953 29009 6956
rect 29043 6984 29055 6987
rect 29178 6984 29184 6996
rect 29043 6956 29184 6984
rect 29043 6953 29055 6956
rect 28997 6947 29055 6953
rect 29178 6944 29184 6956
rect 29236 6944 29242 6996
rect 31205 6987 31263 6993
rect 31205 6953 31217 6987
rect 31251 6984 31263 6987
rect 31478 6984 31484 6996
rect 31251 6956 31484 6984
rect 31251 6953 31263 6956
rect 31205 6947 31263 6953
rect 21361 6919 21419 6925
rect 21361 6916 21373 6919
rect 21324 6888 21373 6916
rect 21324 6876 21330 6888
rect 21361 6885 21373 6888
rect 21407 6885 21419 6919
rect 21542 6916 21548 6928
rect 21503 6888 21548 6916
rect 21361 6879 21419 6885
rect 21542 6876 21548 6888
rect 21600 6876 21606 6928
rect 23106 6916 23112 6928
rect 23067 6888 23112 6916
rect 23106 6876 23112 6888
rect 23164 6876 23170 6928
rect 24670 6916 24676 6928
rect 24631 6888 24676 6916
rect 24670 6876 24676 6888
rect 24728 6876 24734 6928
rect 25406 6916 25412 6928
rect 24780 6888 25412 6916
rect 19659 6820 20668 6848
rect 20717 6851 20775 6857
rect 19659 6817 19671 6820
rect 19613 6811 19671 6817
rect 20717 6817 20729 6851
rect 20763 6848 20775 6851
rect 22465 6851 22523 6857
rect 20763 6820 21680 6848
rect 20763 6817 20775 6820
rect 20717 6811 20775 6817
rect 4154 6780 4160 6792
rect 3568 6752 4016 6780
rect 4067 6752 4160 6780
rect 3568 6740 3574 6752
rect 4154 6740 4160 6752
rect 4212 6780 4218 6792
rect 5442 6780 5448 6792
rect 4212 6752 5448 6780
rect 4212 6740 4218 6752
rect 5442 6740 5448 6752
rect 5500 6740 5506 6792
rect 5997 6783 6055 6789
rect 5997 6749 6009 6783
rect 6043 6749 6055 6783
rect 5997 6743 6055 6749
rect 6089 6783 6147 6789
rect 6089 6749 6101 6783
rect 6135 6749 6147 6783
rect 6089 6743 6147 6749
rect 6549 6783 6607 6789
rect 6549 6749 6561 6783
rect 6595 6780 6607 6783
rect 7466 6780 7472 6792
rect 6595 6752 7472 6780
rect 6595 6749 6607 6752
rect 6549 6743 6607 6749
rect 1670 6712 1676 6724
rect 1631 6684 1676 6712
rect 1670 6672 1676 6684
rect 1728 6672 1734 6724
rect 2958 6672 2964 6724
rect 3016 6712 3022 6724
rect 3053 6715 3111 6721
rect 3053 6712 3065 6715
rect 3016 6684 3065 6712
rect 3016 6672 3022 6684
rect 3053 6681 3065 6684
rect 3099 6712 3111 6715
rect 4338 6712 4344 6724
rect 3099 6684 4344 6712
rect 3099 6681 3111 6684
rect 3053 6675 3111 6681
rect 4338 6672 4344 6684
rect 4396 6672 4402 6724
rect 5537 6715 5595 6721
rect 5537 6681 5549 6715
rect 5583 6712 5595 6715
rect 5718 6712 5724 6724
rect 5583 6684 5724 6712
rect 5583 6681 5595 6684
rect 5537 6675 5595 6681
rect 5718 6672 5724 6684
rect 5776 6672 5782 6724
rect 4706 6604 4712 6656
rect 4764 6644 4770 6656
rect 4801 6647 4859 6653
rect 4801 6644 4813 6647
rect 4764 6616 4813 6644
rect 4764 6604 4770 6616
rect 4801 6613 4813 6616
rect 4847 6644 4859 6647
rect 5350 6644 5356 6656
rect 4847 6616 5356 6644
rect 4847 6613 4859 6616
rect 4801 6607 4859 6613
rect 5350 6604 5356 6616
rect 5408 6604 5414 6656
rect 6012 6644 6040 6743
rect 6104 6712 6132 6743
rect 7466 6740 7472 6752
rect 7524 6740 7530 6792
rect 8570 6780 8576 6792
rect 8531 6752 8576 6780
rect 8570 6740 8576 6752
rect 8628 6740 8634 6792
rect 9674 6740 9680 6792
rect 9732 6780 9738 6792
rect 10137 6783 10195 6789
rect 10137 6780 10149 6783
rect 9732 6752 10149 6780
rect 9732 6740 9738 6752
rect 10137 6749 10149 6752
rect 10183 6749 10195 6783
rect 10318 6780 10324 6792
rect 10279 6752 10324 6780
rect 10137 6743 10195 6749
rect 6822 6712 6828 6724
rect 6104 6684 6828 6712
rect 6822 6672 6828 6684
rect 6880 6672 6886 6724
rect 10152 6712 10180 6743
rect 10318 6740 10324 6752
rect 10376 6740 10382 6792
rect 16758 6780 16764 6792
rect 16719 6752 16764 6780
rect 16758 6740 16764 6752
rect 16816 6740 16822 6792
rect 19889 6783 19947 6789
rect 19889 6749 19901 6783
rect 19935 6780 19947 6783
rect 20732 6780 20760 6811
rect 21652 6792 21680 6820
rect 22465 6817 22477 6851
rect 22511 6848 22523 6851
rect 22738 6848 22744 6860
rect 22511 6820 22744 6848
rect 22511 6817 22523 6820
rect 22465 6811 22523 6817
rect 21634 6780 21640 6792
rect 19935 6752 20760 6780
rect 21547 6752 21640 6780
rect 19935 6749 19947 6752
rect 19889 6743 19947 6749
rect 21634 6740 21640 6752
rect 21692 6780 21698 6792
rect 22480 6780 22508 6811
rect 22738 6808 22744 6820
rect 22796 6848 22802 6860
rect 23842 6848 23848 6860
rect 22796 6820 23848 6848
rect 22796 6808 22802 6820
rect 23842 6808 23848 6820
rect 23900 6848 23906 6860
rect 24780 6857 24808 6888
rect 25406 6876 25412 6888
rect 25464 6876 25470 6928
rect 25682 6876 25688 6928
rect 25740 6916 25746 6928
rect 28902 6916 28908 6928
rect 25740 6888 28908 6916
rect 25740 6876 25746 6888
rect 28902 6876 28908 6888
rect 28960 6876 28966 6928
rect 24765 6851 24823 6857
rect 24765 6848 24777 6851
rect 23900 6820 24777 6848
rect 23900 6808 23906 6820
rect 24765 6817 24777 6820
rect 24811 6817 24823 6851
rect 24765 6811 24823 6817
rect 26602 6808 26608 6860
rect 26660 6848 26666 6860
rect 26953 6851 27011 6857
rect 26953 6848 26965 6851
rect 26660 6820 26965 6848
rect 26660 6808 26666 6820
rect 26953 6817 26965 6820
rect 26999 6817 27011 6851
rect 29448 6851 29506 6857
rect 29448 6848 29460 6851
rect 26953 6811 27011 6817
rect 28092 6820 29460 6848
rect 21692 6752 22508 6780
rect 23109 6783 23167 6789
rect 21692 6740 21698 6752
rect 23109 6749 23121 6783
rect 23155 6749 23167 6783
rect 23109 6743 23167 6749
rect 23201 6783 23259 6789
rect 23201 6749 23213 6783
rect 23247 6780 23259 6783
rect 23382 6780 23388 6792
rect 23247 6752 23388 6780
rect 23247 6749 23259 6752
rect 23201 6743 23259 6749
rect 11146 6712 11152 6724
rect 10152 6684 11152 6712
rect 11146 6672 11152 6684
rect 11204 6672 11210 6724
rect 21085 6715 21143 6721
rect 21085 6681 21097 6715
rect 21131 6712 21143 6715
rect 21358 6712 21364 6724
rect 21131 6684 21364 6712
rect 21131 6681 21143 6684
rect 21085 6675 21143 6681
rect 21358 6672 21364 6684
rect 21416 6672 21422 6724
rect 22554 6672 22560 6724
rect 22612 6712 22618 6724
rect 22649 6715 22707 6721
rect 22649 6712 22661 6715
rect 22612 6684 22661 6712
rect 22612 6672 22618 6684
rect 22649 6681 22661 6684
rect 22695 6681 22707 6715
rect 23124 6712 23152 6743
rect 23382 6740 23388 6752
rect 23440 6740 23446 6792
rect 24118 6740 24124 6792
rect 24176 6780 24182 6792
rect 24581 6783 24639 6789
rect 24581 6780 24593 6783
rect 24176 6752 24593 6780
rect 24176 6740 24182 6752
rect 24581 6749 24593 6752
rect 24627 6749 24639 6783
rect 26694 6780 26700 6792
rect 26655 6752 26700 6780
rect 24581 6743 24639 6749
rect 26694 6740 26700 6752
rect 26752 6740 26758 6792
rect 23474 6712 23480 6724
rect 23124 6684 23480 6712
rect 22649 6675 22707 6681
rect 23474 6672 23480 6684
rect 23532 6672 23538 6724
rect 24026 6712 24032 6724
rect 23939 6684 24032 6712
rect 24026 6672 24032 6684
rect 24084 6712 24090 6724
rect 24670 6712 24676 6724
rect 24084 6684 24676 6712
rect 24084 6672 24090 6684
rect 24670 6672 24676 6684
rect 24728 6672 24734 6724
rect 28092 6721 28120 6820
rect 29448 6817 29460 6820
rect 29494 6848 29506 6851
rect 29914 6848 29920 6860
rect 29494 6820 29920 6848
rect 29494 6817 29506 6820
rect 29448 6811 29506 6817
rect 29914 6808 29920 6820
rect 29972 6848 29978 6860
rect 31220 6848 31248 6947
rect 31478 6944 31484 6956
rect 31536 6944 31542 6996
rect 33962 6984 33968 6996
rect 33923 6956 33968 6984
rect 33962 6944 33968 6956
rect 34020 6984 34026 6996
rect 34333 6987 34391 6993
rect 34333 6984 34345 6987
rect 34020 6956 34345 6984
rect 34020 6944 34026 6956
rect 34333 6953 34345 6956
rect 34379 6953 34391 6987
rect 34333 6947 34391 6953
rect 32493 6919 32551 6925
rect 32493 6916 32505 6919
rect 32324 6888 32505 6916
rect 29972 6820 31248 6848
rect 29972 6808 29978 6820
rect 31754 6808 31760 6860
rect 31812 6848 31818 6860
rect 32324 6848 32352 6888
rect 32493 6885 32505 6888
rect 32539 6885 32551 6919
rect 32674 6916 32680 6928
rect 32635 6888 32680 6916
rect 32493 6879 32551 6885
rect 32674 6876 32680 6888
rect 32732 6876 32738 6928
rect 32769 6851 32827 6857
rect 32769 6848 32781 6851
rect 31812 6820 32352 6848
rect 32416 6820 32781 6848
rect 31812 6808 31818 6820
rect 32416 6792 32444 6820
rect 32769 6817 32781 6820
rect 32815 6817 32827 6851
rect 34348 6848 34376 6947
rect 35710 6944 35716 6996
rect 35768 6984 35774 6996
rect 35897 6987 35955 6993
rect 35897 6984 35909 6987
rect 35768 6956 35909 6984
rect 35768 6944 35774 6956
rect 35897 6953 35909 6956
rect 35943 6953 35955 6987
rect 35897 6947 35955 6953
rect 34514 6876 34520 6928
rect 34572 6916 34578 6928
rect 34974 6916 34980 6928
rect 34572 6888 34980 6916
rect 34572 6876 34578 6888
rect 34974 6876 34980 6888
rect 35032 6876 35038 6928
rect 34790 6857 34796 6860
rect 34773 6851 34796 6857
rect 34773 6848 34785 6851
rect 34348 6820 34785 6848
rect 32769 6811 32827 6817
rect 34773 6817 34785 6820
rect 34848 6848 34854 6860
rect 36262 6848 36268 6860
rect 34848 6820 36268 6848
rect 34773 6811 34796 6817
rect 34790 6808 34796 6811
rect 34848 6808 34854 6820
rect 36262 6808 36268 6820
rect 36320 6808 36326 6860
rect 28994 6740 29000 6792
rect 29052 6780 29058 6792
rect 29181 6783 29239 6789
rect 29181 6780 29193 6783
rect 29052 6752 29193 6780
rect 29052 6740 29058 6752
rect 29181 6749 29193 6752
rect 29227 6749 29239 6783
rect 30742 6780 30748 6792
rect 29181 6743 29239 6749
rect 30576 6752 30748 6780
rect 30576 6721 30604 6752
rect 30742 6740 30748 6752
rect 30800 6780 30806 6792
rect 32398 6780 32404 6792
rect 30800 6752 32404 6780
rect 30800 6740 30806 6752
rect 32398 6740 32404 6752
rect 32456 6740 32462 6792
rect 34514 6780 34520 6792
rect 34475 6752 34520 6780
rect 34514 6740 34520 6752
rect 34572 6740 34578 6792
rect 25041 6715 25099 6721
rect 25041 6681 25053 6715
rect 25087 6712 25099 6715
rect 28077 6715 28135 6721
rect 25087 6684 26096 6712
rect 25087 6681 25099 6684
rect 25041 6675 25099 6681
rect 6178 6644 6184 6656
rect 6012 6616 6184 6644
rect 6178 6604 6184 6616
rect 6236 6604 6242 6656
rect 7098 6644 7104 6656
rect 7059 6616 7104 6644
rect 7098 6604 7104 6616
rect 7156 6604 7162 6656
rect 9490 6644 9496 6656
rect 9451 6616 9496 6644
rect 9490 6604 9496 6616
rect 9548 6604 9554 6656
rect 9766 6644 9772 6656
rect 9727 6616 9772 6644
rect 9766 6604 9772 6616
rect 9824 6604 9830 6656
rect 11698 6604 11704 6656
rect 11756 6644 11762 6656
rect 12713 6647 12771 6653
rect 12713 6644 12725 6647
rect 11756 6616 12725 6644
rect 11756 6604 11762 6616
rect 12713 6613 12725 6616
rect 12759 6613 12771 6647
rect 12713 6607 12771 6613
rect 18141 6647 18199 6653
rect 18141 6613 18153 6647
rect 18187 6644 18199 6647
rect 18506 6644 18512 6656
rect 18187 6616 18512 6644
rect 18187 6613 18199 6616
rect 18141 6607 18199 6613
rect 18506 6604 18512 6616
rect 18564 6604 18570 6656
rect 18785 6647 18843 6653
rect 18785 6613 18797 6647
rect 18831 6644 18843 6647
rect 18874 6644 18880 6656
rect 18831 6616 18880 6644
rect 18831 6613 18843 6616
rect 18785 6607 18843 6613
rect 18874 6604 18880 6616
rect 18932 6604 18938 6656
rect 19337 6647 19395 6653
rect 19337 6613 19349 6647
rect 19383 6644 19395 6647
rect 20254 6644 20260 6656
rect 19383 6616 20260 6644
rect 19383 6613 19395 6616
rect 19337 6607 19395 6613
rect 20254 6604 20260 6616
rect 20312 6604 20318 6656
rect 20530 6604 20536 6656
rect 20588 6644 20594 6656
rect 21542 6644 21548 6656
rect 20588 6616 21548 6644
rect 20588 6604 20594 6616
rect 21542 6604 21548 6616
rect 21600 6604 21606 6656
rect 21910 6604 21916 6656
rect 21968 6644 21974 6656
rect 22094 6644 22100 6656
rect 21968 6616 22100 6644
rect 21968 6604 21974 6616
rect 22094 6604 22100 6616
rect 22152 6604 22158 6656
rect 24210 6644 24216 6656
rect 24171 6616 24216 6644
rect 24210 6604 24216 6616
rect 24268 6604 24274 6656
rect 24946 6604 24952 6656
rect 25004 6644 25010 6656
rect 25133 6647 25191 6653
rect 25133 6644 25145 6647
rect 25004 6616 25145 6644
rect 25004 6604 25010 6616
rect 25133 6613 25145 6616
rect 25179 6613 25191 6647
rect 25958 6644 25964 6656
rect 25919 6616 25964 6644
rect 25133 6607 25191 6613
rect 25958 6604 25964 6616
rect 26016 6604 26022 6656
rect 26068 6644 26096 6684
rect 28077 6681 28089 6715
rect 28123 6681 28135 6715
rect 28077 6675 28135 6681
rect 30561 6715 30619 6721
rect 30561 6681 30573 6715
rect 30607 6681 30619 6715
rect 30561 6675 30619 6681
rect 32030 6672 32036 6724
rect 32088 6712 32094 6724
rect 32217 6715 32275 6721
rect 32217 6712 32229 6715
rect 32088 6684 32229 6712
rect 32088 6672 32094 6684
rect 32217 6681 32229 6684
rect 32263 6681 32275 6715
rect 32217 6675 32275 6681
rect 33321 6715 33379 6721
rect 33321 6681 33333 6715
rect 33367 6712 33379 6715
rect 33778 6712 33784 6724
rect 33367 6684 33784 6712
rect 33367 6681 33379 6684
rect 33321 6675 33379 6681
rect 33778 6672 33784 6684
rect 33836 6672 33842 6724
rect 28810 6644 28816 6656
rect 26068 6616 28816 6644
rect 28810 6604 28816 6616
rect 28868 6604 28874 6656
rect 31478 6644 31484 6656
rect 31439 6616 31484 6644
rect 31478 6604 31484 6616
rect 31536 6604 31542 6656
rect 31941 6647 31999 6653
rect 31941 6613 31953 6647
rect 31987 6644 31999 6647
rect 33134 6644 33140 6656
rect 31987 6616 33140 6644
rect 31987 6613 31999 6616
rect 31941 6607 31999 6613
rect 33134 6604 33140 6616
rect 33192 6604 33198 6656
rect 33686 6644 33692 6656
rect 33647 6616 33692 6644
rect 33686 6604 33692 6616
rect 33744 6604 33750 6656
rect 36446 6644 36452 6656
rect 36407 6616 36452 6644
rect 36446 6604 36452 6616
rect 36504 6604 36510 6656
rect 1104 6554 38824 6576
rect 1104 6502 7648 6554
rect 7700 6502 7712 6554
rect 7764 6502 7776 6554
rect 7828 6502 7840 6554
rect 7892 6502 20982 6554
rect 21034 6502 21046 6554
rect 21098 6502 21110 6554
rect 21162 6502 21174 6554
rect 21226 6502 34315 6554
rect 34367 6502 34379 6554
rect 34431 6502 34443 6554
rect 34495 6502 34507 6554
rect 34559 6502 38824 6554
rect 1104 6480 38824 6502
rect 2866 6400 2872 6452
rect 2924 6440 2930 6452
rect 3145 6443 3203 6449
rect 3145 6440 3157 6443
rect 2924 6412 3157 6440
rect 2924 6400 2930 6412
rect 3145 6409 3157 6412
rect 3191 6409 3203 6443
rect 4154 6440 4160 6452
rect 4115 6412 4160 6440
rect 3145 6403 3203 6409
rect 4154 6400 4160 6412
rect 4212 6400 4218 6452
rect 6641 6443 6699 6449
rect 6641 6409 6653 6443
rect 6687 6440 6699 6443
rect 6822 6440 6828 6452
rect 6687 6412 6828 6440
rect 6687 6409 6699 6412
rect 6641 6403 6699 6409
rect 6822 6400 6828 6412
rect 6880 6400 6886 6452
rect 7285 6443 7343 6449
rect 7285 6409 7297 6443
rect 7331 6440 7343 6443
rect 8110 6440 8116 6452
rect 7331 6412 8116 6440
rect 7331 6409 7343 6412
rect 7285 6403 7343 6409
rect 5350 6264 5356 6316
rect 5408 6304 5414 6316
rect 7392 6313 7420 6412
rect 8110 6400 8116 6412
rect 8168 6400 8174 6452
rect 11330 6440 11336 6452
rect 11291 6412 11336 6440
rect 11330 6400 11336 6412
rect 11388 6400 11394 6452
rect 11790 6440 11796 6452
rect 11751 6412 11796 6440
rect 11790 6400 11796 6412
rect 11848 6400 11854 6452
rect 12158 6440 12164 6452
rect 12119 6412 12164 6440
rect 12158 6400 12164 6412
rect 12216 6400 12222 6452
rect 17770 6440 17776 6452
rect 17731 6412 17776 6440
rect 17770 6400 17776 6412
rect 17828 6400 17834 6452
rect 18690 6440 18696 6452
rect 18651 6412 18696 6440
rect 18690 6400 18696 6412
rect 18748 6400 18754 6452
rect 19334 6440 19340 6452
rect 19295 6412 19340 6440
rect 19334 6400 19340 6412
rect 19392 6400 19398 6452
rect 19610 6440 19616 6452
rect 19571 6412 19616 6440
rect 19610 6400 19616 6412
rect 19668 6400 19674 6452
rect 20806 6400 20812 6452
rect 20864 6440 20870 6452
rect 20993 6443 21051 6449
rect 20993 6440 21005 6443
rect 20864 6412 21005 6440
rect 20864 6400 20870 6412
rect 20993 6409 21005 6412
rect 21039 6440 21051 6443
rect 21266 6440 21272 6452
rect 21039 6412 21272 6440
rect 21039 6409 21051 6412
rect 20993 6403 21051 6409
rect 21266 6400 21272 6412
rect 21324 6400 21330 6452
rect 22462 6440 22468 6452
rect 22423 6412 22468 6440
rect 22462 6400 22468 6412
rect 22520 6400 22526 6452
rect 23106 6440 23112 6452
rect 23067 6412 23112 6440
rect 23106 6400 23112 6412
rect 23164 6400 23170 6452
rect 23474 6440 23480 6452
rect 23387 6412 23480 6440
rect 23474 6400 23480 6412
rect 23532 6440 23538 6452
rect 23934 6440 23940 6452
rect 23532 6412 23940 6440
rect 23532 6400 23538 6412
rect 23934 6400 23940 6412
rect 23992 6400 23998 6452
rect 24486 6440 24492 6452
rect 24447 6412 24492 6440
rect 24486 6400 24492 6412
rect 24544 6400 24550 6452
rect 25774 6440 25780 6452
rect 25735 6412 25780 6440
rect 25774 6400 25780 6412
rect 25832 6440 25838 6452
rect 26418 6440 26424 6452
rect 25832 6412 26424 6440
rect 25832 6400 25838 6412
rect 26418 6400 26424 6412
rect 26476 6400 26482 6452
rect 27062 6440 27068 6452
rect 27023 6412 27068 6440
rect 27062 6400 27068 6412
rect 27120 6400 27126 6452
rect 27338 6440 27344 6452
rect 27299 6412 27344 6440
rect 27338 6400 27344 6412
rect 27396 6400 27402 6452
rect 28994 6400 29000 6452
rect 29052 6440 29058 6452
rect 29457 6443 29515 6449
rect 29457 6440 29469 6443
rect 29052 6412 29469 6440
rect 29052 6400 29058 6412
rect 29457 6409 29469 6412
rect 29503 6440 29515 6443
rect 29914 6440 29920 6452
rect 29503 6412 29684 6440
rect 29875 6412 29920 6440
rect 29503 6409 29515 6412
rect 29457 6403 29515 6409
rect 9950 6372 9956 6384
rect 9911 6344 9956 6372
rect 9950 6332 9956 6344
rect 10008 6332 10014 6384
rect 12434 6332 12440 6384
rect 12492 6372 12498 6384
rect 12529 6375 12587 6381
rect 12529 6372 12541 6375
rect 12492 6344 12541 6372
rect 12492 6332 12498 6344
rect 12529 6341 12541 6344
rect 12575 6341 12587 6375
rect 12529 6335 12587 6341
rect 15562 6332 15568 6384
rect 15620 6372 15626 6384
rect 16758 6372 16764 6384
rect 15620 6344 16764 6372
rect 15620 6332 15626 6344
rect 16758 6332 16764 6344
rect 16816 6372 16822 6384
rect 16853 6375 16911 6381
rect 16853 6372 16865 6375
rect 16816 6344 16865 6372
rect 16816 6332 16822 6344
rect 16853 6341 16865 6344
rect 16899 6372 16911 6375
rect 17678 6372 17684 6384
rect 16899 6344 17684 6372
rect 16899 6341 16911 6344
rect 16853 6335 16911 6341
rect 17678 6332 17684 6344
rect 17736 6332 17742 6384
rect 7377 6307 7435 6313
rect 7377 6304 7389 6307
rect 5408 6276 7389 6304
rect 5408 6264 5414 6276
rect 7377 6273 7389 6276
rect 7423 6273 7435 6307
rect 19352 6304 19380 6400
rect 26053 6375 26111 6381
rect 26053 6341 26065 6375
rect 26099 6372 26111 6375
rect 26326 6372 26332 6384
rect 26099 6344 26332 6372
rect 26099 6341 26111 6344
rect 26053 6335 26111 6341
rect 26326 6332 26332 6344
rect 26384 6332 26390 6384
rect 19981 6307 20039 6313
rect 19981 6304 19993 6307
rect 19352 6276 19993 6304
rect 7377 6267 7435 6273
rect 19981 6273 19993 6276
rect 20027 6273 20039 6307
rect 20162 6304 20168 6316
rect 20123 6276 20168 6304
rect 19981 6267 20039 6273
rect 20162 6264 20168 6276
rect 20220 6264 20226 6316
rect 24949 6307 25007 6313
rect 24949 6273 24961 6307
rect 24995 6304 25007 6307
rect 25130 6304 25136 6316
rect 24995 6276 25136 6304
rect 24995 6273 25007 6276
rect 24949 6267 25007 6273
rect 25130 6264 25136 6276
rect 25188 6304 25194 6316
rect 26436 6313 26464 6400
rect 25409 6307 25467 6313
rect 25409 6304 25421 6307
rect 25188 6276 25421 6304
rect 25188 6264 25194 6276
rect 25409 6273 25421 6276
rect 25455 6273 25467 6307
rect 25409 6267 25467 6273
rect 26421 6307 26479 6313
rect 26421 6273 26433 6307
rect 26467 6273 26479 6307
rect 27080 6304 27108 6400
rect 27617 6375 27675 6381
rect 27617 6341 27629 6375
rect 27663 6372 27675 6375
rect 29546 6372 29552 6384
rect 27663 6344 29552 6372
rect 27663 6341 27675 6344
rect 27617 6335 27675 6341
rect 29546 6332 29552 6344
rect 29604 6332 29610 6384
rect 29656 6372 29684 6412
rect 29914 6400 29920 6412
rect 29972 6400 29978 6452
rect 32398 6440 32404 6452
rect 32359 6412 32404 6440
rect 32398 6400 32404 6412
rect 32456 6400 32462 6452
rect 33134 6400 33140 6452
rect 33192 6440 33198 6452
rect 33321 6443 33379 6449
rect 33321 6440 33333 6443
rect 33192 6412 33333 6440
rect 33192 6400 33198 6412
rect 33321 6409 33333 6412
rect 33367 6409 33379 6443
rect 36262 6440 36268 6452
rect 36223 6412 36268 6440
rect 33321 6403 33379 6409
rect 36262 6400 36268 6412
rect 36320 6400 36326 6452
rect 37553 6443 37611 6449
rect 37553 6409 37565 6443
rect 37599 6440 37611 6443
rect 37642 6440 37648 6452
rect 37599 6412 37648 6440
rect 37599 6409 37611 6412
rect 37553 6403 37611 6409
rect 37642 6400 37648 6412
rect 37700 6400 37706 6452
rect 30285 6375 30343 6381
rect 30285 6372 30297 6375
rect 29656 6344 30297 6372
rect 30285 6341 30297 6344
rect 30331 6372 30343 6375
rect 31849 6375 31907 6381
rect 30331 6344 30512 6372
rect 30331 6341 30343 6344
rect 30285 6335 30343 6341
rect 30484 6313 30512 6344
rect 31849 6341 31861 6375
rect 31895 6372 31907 6375
rect 33686 6372 33692 6384
rect 31895 6344 33692 6372
rect 31895 6341 31907 6344
rect 31849 6335 31907 6341
rect 33686 6332 33692 6344
rect 33744 6372 33750 6384
rect 33744 6344 33916 6372
rect 33744 6332 33750 6344
rect 27985 6307 28043 6313
rect 27985 6304 27997 6307
rect 27080 6276 27997 6304
rect 26421 6267 26479 6273
rect 27985 6273 27997 6276
rect 28031 6273 28043 6307
rect 27985 6267 28043 6273
rect 30469 6307 30527 6313
rect 30469 6273 30481 6307
rect 30515 6273 30527 6307
rect 33778 6304 33784 6316
rect 33739 6276 33784 6304
rect 30469 6267 30527 6273
rect 33778 6264 33784 6276
rect 33836 6264 33842 6316
rect 33888 6313 33916 6344
rect 33873 6307 33931 6313
rect 33873 6273 33885 6307
rect 33919 6273 33931 6307
rect 33873 6267 33931 6273
rect 1486 6196 1492 6248
rect 1544 6236 1550 6248
rect 1673 6239 1731 6245
rect 1673 6236 1685 6239
rect 1544 6208 1685 6236
rect 1544 6196 1550 6208
rect 1673 6205 1685 6208
rect 1719 6236 1731 6239
rect 1765 6239 1823 6245
rect 1765 6236 1777 6239
rect 1719 6208 1777 6236
rect 1719 6205 1731 6208
rect 1673 6199 1731 6205
rect 1765 6205 1777 6208
rect 1811 6236 1823 6239
rect 2958 6236 2964 6248
rect 1811 6208 2964 6236
rect 1811 6205 1823 6208
rect 1765 6199 1823 6205
rect 2958 6196 2964 6208
rect 3016 6236 3022 6248
rect 3789 6239 3847 6245
rect 3789 6236 3801 6239
rect 3016 6208 3801 6236
rect 3016 6196 3022 6208
rect 3789 6205 3801 6208
rect 3835 6236 3847 6239
rect 4249 6239 4307 6245
rect 4249 6236 4261 6239
rect 3835 6208 4261 6236
rect 3835 6205 3847 6208
rect 3789 6199 3847 6205
rect 4249 6205 4261 6208
rect 4295 6236 4307 6239
rect 5368 6236 5396 6264
rect 9674 6236 9680 6248
rect 4295 6208 5396 6236
rect 9635 6208 9680 6236
rect 4295 6205 4307 6208
rect 4249 6199 4307 6205
rect 9674 6196 9680 6208
rect 9732 6196 9738 6248
rect 10318 6196 10324 6248
rect 10376 6236 10382 6248
rect 10873 6239 10931 6245
rect 10873 6236 10885 6239
rect 10376 6208 10885 6236
rect 10376 6196 10382 6208
rect 10873 6205 10885 6208
rect 10919 6205 10931 6239
rect 10873 6199 10931 6205
rect 11790 6196 11796 6248
rect 11848 6236 11854 6248
rect 12805 6239 12863 6245
rect 12805 6236 12817 6239
rect 11848 6208 12817 6236
rect 11848 6196 11854 6208
rect 12805 6205 12817 6208
rect 12851 6205 12863 6239
rect 12805 6199 12863 6205
rect 12986 6196 12992 6248
rect 13044 6236 13050 6248
rect 13081 6239 13139 6245
rect 13081 6236 13093 6239
rect 13044 6208 13093 6236
rect 13044 6196 13050 6208
rect 13081 6205 13093 6208
rect 13127 6236 13139 6239
rect 13449 6239 13507 6245
rect 13449 6236 13461 6239
rect 13127 6208 13461 6236
rect 13127 6205 13139 6208
rect 13081 6199 13139 6205
rect 13449 6205 13461 6208
rect 13495 6205 13507 6239
rect 13449 6199 13507 6205
rect 13538 6196 13544 6248
rect 13596 6236 13602 6248
rect 14277 6239 14335 6245
rect 14277 6236 14289 6239
rect 13596 6208 14289 6236
rect 13596 6196 13602 6208
rect 14277 6205 14289 6208
rect 14323 6236 14335 6239
rect 14369 6239 14427 6245
rect 14369 6236 14381 6239
rect 14323 6208 14381 6236
rect 14323 6205 14335 6208
rect 14277 6199 14335 6205
rect 14369 6205 14381 6208
rect 14415 6236 14427 6239
rect 15562 6236 15568 6248
rect 14415 6208 15568 6236
rect 14415 6205 14427 6208
rect 14369 6199 14427 6205
rect 15562 6196 15568 6208
rect 15620 6196 15626 6248
rect 18966 6236 18972 6248
rect 18927 6208 18972 6236
rect 18966 6196 18972 6208
rect 19024 6236 19030 6248
rect 19794 6236 19800 6248
rect 19024 6208 19800 6236
rect 19024 6196 19030 6208
rect 19794 6196 19800 6208
rect 19852 6196 19858 6248
rect 21082 6236 21088 6248
rect 21043 6208 21088 6236
rect 21082 6196 21088 6208
rect 21140 6196 21146 6248
rect 21352 6239 21410 6245
rect 21352 6205 21364 6239
rect 21398 6236 21410 6239
rect 21634 6236 21640 6248
rect 21398 6208 21640 6236
rect 21398 6205 21410 6208
rect 21352 6199 21410 6205
rect 21634 6196 21640 6208
rect 21692 6196 21698 6248
rect 30742 6245 30748 6248
rect 30736 6236 30748 6245
rect 30703 6208 30748 6236
rect 30736 6199 30748 6208
rect 30742 6196 30748 6199
rect 30800 6196 30806 6248
rect 34609 6239 34667 6245
rect 34609 6205 34621 6239
rect 34655 6236 34667 6239
rect 34885 6239 34943 6245
rect 34885 6236 34897 6239
rect 34655 6208 34897 6236
rect 34655 6205 34667 6208
rect 34609 6199 34667 6205
rect 34885 6205 34897 6208
rect 34931 6236 34943 6239
rect 34974 6236 34980 6248
rect 34931 6208 34980 6236
rect 34931 6205 34943 6208
rect 34885 6199 34943 6205
rect 34974 6196 34980 6208
rect 35032 6196 35038 6248
rect 37366 6236 37372 6248
rect 37327 6208 37372 6236
rect 37366 6196 37372 6208
rect 37424 6236 37430 6248
rect 37921 6239 37979 6245
rect 37921 6236 37933 6239
rect 37424 6208 37933 6236
rect 37424 6196 37430 6208
rect 37921 6205 37933 6208
rect 37967 6205 37979 6239
rect 37921 6199 37979 6205
rect 2032 6171 2090 6177
rect 2032 6137 2044 6171
rect 2078 6168 2090 6171
rect 2222 6168 2228 6180
rect 2078 6140 2228 6168
rect 2078 6137 2090 6140
rect 2032 6131 2090 6137
rect 2222 6128 2228 6140
rect 2280 6128 2286 6180
rect 4516 6171 4574 6177
rect 4516 6137 4528 6171
rect 4562 6168 4574 6171
rect 4614 6168 4620 6180
rect 4562 6140 4620 6168
rect 4562 6137 4574 6140
rect 4516 6131 4574 6137
rect 4614 6128 4620 6140
rect 4672 6128 4678 6180
rect 7650 6177 7656 6180
rect 7644 6168 7656 6177
rect 7611 6140 7656 6168
rect 7644 6131 7656 6140
rect 7650 6128 7656 6131
rect 7708 6128 7714 6180
rect 9490 6128 9496 6180
rect 9548 6168 9554 6180
rect 10229 6171 10287 6177
rect 10229 6168 10241 6171
rect 9548 6140 10241 6168
rect 9548 6128 9554 6140
rect 10229 6137 10241 6140
rect 10275 6137 10287 6171
rect 10502 6168 10508 6180
rect 10463 6140 10508 6168
rect 10229 6131 10287 6137
rect 10502 6128 10508 6140
rect 10560 6128 10566 6180
rect 14636 6171 14694 6177
rect 14636 6137 14648 6171
rect 14682 6168 14694 6171
rect 14826 6168 14832 6180
rect 14682 6140 14832 6168
rect 14682 6137 14694 6140
rect 14636 6131 14694 6137
rect 14826 6128 14832 6140
rect 14884 6128 14890 6180
rect 20456 6140 24348 6168
rect 5534 6060 5540 6112
rect 5592 6100 5598 6112
rect 5629 6103 5687 6109
rect 5629 6100 5641 6103
rect 5592 6072 5641 6100
rect 5592 6060 5598 6072
rect 5629 6069 5641 6072
rect 5675 6069 5687 6103
rect 6178 6100 6184 6112
rect 6139 6072 6184 6100
rect 5629 6063 5687 6069
rect 6178 6060 6184 6072
rect 6236 6060 6242 6112
rect 8386 6060 8392 6112
rect 8444 6100 8450 6112
rect 8757 6103 8815 6109
rect 8757 6100 8769 6103
rect 8444 6072 8769 6100
rect 8444 6060 8450 6072
rect 8757 6069 8769 6072
rect 8803 6069 8815 6103
rect 9306 6100 9312 6112
rect 9267 6072 9312 6100
rect 8757 6063 8815 6069
rect 9306 6060 9312 6072
rect 9364 6060 9370 6112
rect 9766 6060 9772 6112
rect 9824 6100 9830 6112
rect 10413 6103 10471 6109
rect 10413 6100 10425 6103
rect 9824 6072 10425 6100
rect 9824 6060 9830 6072
rect 10413 6069 10425 6072
rect 10459 6069 10471 6103
rect 10413 6063 10471 6069
rect 12158 6060 12164 6112
rect 12216 6100 12222 6112
rect 12989 6103 13047 6109
rect 12989 6100 13001 6103
rect 12216 6072 13001 6100
rect 12216 6060 12222 6072
rect 12989 6069 13001 6072
rect 13035 6069 13047 6103
rect 15746 6100 15752 6112
rect 15707 6072 15752 6100
rect 12989 6063 13047 6069
rect 15746 6060 15752 6072
rect 15804 6060 15810 6112
rect 16850 6060 16856 6112
rect 16908 6100 16914 6112
rect 17129 6103 17187 6109
rect 17129 6100 17141 6103
rect 16908 6072 17141 6100
rect 16908 6060 16914 6072
rect 17129 6069 17141 6072
rect 17175 6069 17187 6103
rect 17129 6063 17187 6069
rect 18325 6103 18383 6109
rect 18325 6069 18337 6103
rect 18371 6100 18383 6103
rect 18506 6100 18512 6112
rect 18371 6072 18512 6100
rect 18371 6069 18383 6072
rect 18325 6063 18383 6069
rect 18506 6060 18512 6072
rect 18564 6060 18570 6112
rect 19518 6060 19524 6112
rect 19576 6100 19582 6112
rect 20073 6103 20131 6109
rect 20073 6100 20085 6103
rect 19576 6072 20085 6100
rect 19576 6060 19582 6072
rect 20073 6069 20085 6072
rect 20119 6100 20131 6103
rect 20456 6100 20484 6140
rect 20119 6072 20484 6100
rect 20119 6069 20131 6072
rect 20073 6063 20131 6069
rect 20530 6060 20536 6112
rect 20588 6100 20594 6112
rect 24118 6100 24124 6112
rect 20588 6072 20633 6100
rect 24079 6072 24124 6100
rect 20588 6060 20594 6072
rect 24118 6060 24124 6072
rect 24176 6060 24182 6112
rect 24320 6100 24348 6140
rect 24762 6128 24768 6180
rect 24820 6168 24826 6180
rect 25041 6171 25099 6177
rect 25041 6168 25053 6171
rect 24820 6140 25053 6168
rect 24820 6128 24826 6140
rect 25041 6137 25053 6140
rect 25087 6168 25099 6171
rect 26602 6168 26608 6180
rect 25087 6140 26608 6168
rect 25087 6137 25099 6140
rect 25041 6131 25099 6137
rect 26602 6128 26608 6140
rect 26660 6128 26666 6180
rect 27522 6168 27528 6180
rect 26712 6140 27528 6168
rect 24946 6100 24952 6112
rect 24320 6072 24952 6100
rect 24946 6060 24952 6072
rect 25004 6060 25010 6112
rect 25958 6060 25964 6112
rect 26016 6100 26022 6112
rect 26513 6103 26571 6109
rect 26513 6100 26525 6103
rect 26016 6072 26525 6100
rect 26016 6060 26022 6072
rect 26513 6069 26525 6072
rect 26559 6100 26571 6103
rect 26712 6100 26740 6140
rect 27522 6128 27528 6140
rect 27580 6128 27586 6180
rect 28169 6171 28227 6177
rect 28169 6137 28181 6171
rect 28215 6168 28227 6171
rect 28258 6168 28264 6180
rect 28215 6140 28264 6168
rect 28215 6137 28227 6140
rect 28169 6131 28227 6137
rect 28258 6128 28264 6140
rect 28316 6168 28322 6180
rect 28537 6171 28595 6177
rect 28537 6168 28549 6171
rect 28316 6140 28549 6168
rect 28316 6128 28322 6140
rect 28537 6137 28549 6140
rect 28583 6137 28595 6171
rect 28537 6131 28595 6137
rect 29822 6128 29828 6180
rect 29880 6168 29886 6180
rect 30282 6168 30288 6180
rect 29880 6140 30288 6168
rect 29880 6128 29886 6140
rect 30282 6128 30288 6140
rect 30340 6168 30346 6180
rect 35158 6177 35164 6180
rect 33137 6171 33195 6177
rect 33137 6168 33149 6171
rect 30340 6140 33149 6168
rect 30340 6128 30346 6140
rect 33137 6137 33149 6140
rect 33183 6168 33195 6171
rect 33781 6171 33839 6177
rect 33781 6168 33793 6171
rect 33183 6140 33793 6168
rect 33183 6137 33195 6140
rect 33137 6131 33195 6137
rect 33781 6137 33793 6140
rect 33827 6137 33839 6171
rect 35152 6168 35164 6177
rect 35119 6140 35164 6168
rect 33781 6131 33839 6137
rect 35152 6131 35164 6140
rect 35158 6128 35164 6131
rect 35216 6128 35222 6180
rect 26559 6072 26740 6100
rect 26559 6069 26571 6072
rect 26513 6063 26571 6069
rect 27338 6060 27344 6112
rect 27396 6100 27402 6112
rect 28077 6103 28135 6109
rect 28077 6100 28089 6103
rect 27396 6072 28089 6100
rect 27396 6060 27402 6072
rect 28077 6069 28089 6072
rect 28123 6069 28135 6103
rect 28077 6063 28135 6069
rect 1104 6010 38824 6032
rect 1104 5958 14315 6010
rect 14367 5958 14379 6010
rect 14431 5958 14443 6010
rect 14495 5958 14507 6010
rect 14559 5958 27648 6010
rect 27700 5958 27712 6010
rect 27764 5958 27776 6010
rect 27828 5958 27840 6010
rect 27892 5958 38824 6010
rect 1104 5936 38824 5958
rect 2866 5896 2872 5908
rect 2779 5868 2872 5896
rect 2866 5856 2872 5868
rect 2924 5896 2930 5908
rect 4614 5896 4620 5908
rect 2924 5868 4620 5896
rect 2924 5856 2930 5868
rect 4614 5856 4620 5868
rect 4672 5856 4678 5908
rect 5166 5896 5172 5908
rect 5127 5868 5172 5896
rect 5166 5856 5172 5868
rect 5224 5856 5230 5908
rect 6641 5899 6699 5905
rect 6641 5865 6653 5899
rect 6687 5896 6699 5899
rect 7285 5899 7343 5905
rect 7285 5896 7297 5899
rect 6687 5868 7297 5896
rect 6687 5865 6699 5868
rect 6641 5859 6699 5865
rect 7285 5865 7297 5868
rect 7331 5896 7343 5899
rect 7374 5896 7380 5908
rect 7331 5868 7380 5896
rect 7331 5865 7343 5868
rect 7285 5859 7343 5865
rect 7374 5856 7380 5868
rect 7432 5896 7438 5908
rect 7650 5896 7656 5908
rect 7432 5868 7656 5896
rect 7432 5856 7438 5868
rect 7650 5856 7656 5868
rect 7708 5856 7714 5908
rect 9493 5899 9551 5905
rect 9493 5865 9505 5899
rect 9539 5896 9551 5899
rect 9766 5896 9772 5908
rect 9539 5868 9772 5896
rect 9539 5865 9551 5868
rect 9493 5859 9551 5865
rect 9766 5856 9772 5868
rect 9824 5856 9830 5908
rect 10502 5856 10508 5908
rect 10560 5896 10566 5908
rect 10689 5899 10747 5905
rect 10689 5896 10701 5899
rect 10560 5868 10701 5896
rect 10560 5856 10566 5868
rect 10689 5865 10701 5868
rect 10735 5865 10747 5899
rect 11422 5896 11428 5908
rect 11383 5868 11428 5896
rect 10689 5859 10747 5865
rect 11422 5856 11428 5868
rect 11480 5856 11486 5908
rect 17954 5856 17960 5908
rect 18012 5896 18018 5908
rect 18509 5899 18567 5905
rect 18509 5896 18521 5899
rect 18012 5868 18521 5896
rect 18012 5856 18018 5868
rect 18509 5865 18521 5868
rect 18555 5896 18567 5899
rect 19058 5896 19064 5908
rect 18555 5868 19064 5896
rect 18555 5865 18567 5868
rect 18509 5859 18567 5865
rect 19058 5856 19064 5868
rect 19116 5856 19122 5908
rect 19518 5896 19524 5908
rect 19479 5868 19524 5896
rect 19518 5856 19524 5868
rect 19576 5856 19582 5908
rect 19981 5899 20039 5905
rect 19981 5865 19993 5899
rect 20027 5896 20039 5899
rect 20717 5899 20775 5905
rect 20717 5896 20729 5899
rect 20027 5868 20729 5896
rect 20027 5865 20039 5868
rect 19981 5859 20039 5865
rect 20717 5865 20729 5868
rect 20763 5896 20775 5899
rect 21634 5896 21640 5908
rect 20763 5868 21640 5896
rect 20763 5865 20775 5868
rect 20717 5859 20775 5865
rect 21634 5856 21640 5868
rect 21692 5856 21698 5908
rect 23382 5896 23388 5908
rect 23343 5868 23388 5896
rect 23382 5856 23388 5868
rect 23440 5856 23446 5908
rect 23842 5896 23848 5908
rect 23803 5868 23848 5896
rect 23842 5856 23848 5868
rect 23900 5856 23906 5908
rect 27699 5899 27757 5905
rect 27699 5865 27711 5899
rect 27745 5896 27757 5899
rect 29638 5896 29644 5908
rect 27745 5868 29644 5896
rect 27745 5865 27757 5868
rect 27699 5859 27757 5865
rect 29638 5856 29644 5868
rect 29696 5896 29702 5908
rect 29733 5899 29791 5905
rect 29733 5896 29745 5899
rect 29696 5868 29745 5896
rect 29696 5856 29702 5868
rect 29733 5865 29745 5868
rect 29779 5865 29791 5899
rect 29733 5859 29791 5865
rect 30561 5899 30619 5905
rect 30561 5865 30573 5899
rect 30607 5896 30619 5899
rect 30742 5896 30748 5908
rect 30607 5868 30748 5896
rect 30607 5865 30619 5868
rect 30561 5859 30619 5865
rect 30742 5856 30748 5868
rect 30800 5856 30806 5908
rect 31754 5856 31760 5908
rect 31812 5896 31818 5908
rect 31849 5899 31907 5905
rect 31849 5896 31861 5899
rect 31812 5868 31861 5896
rect 31812 5856 31818 5868
rect 31849 5865 31861 5868
rect 31895 5865 31907 5899
rect 31849 5859 31907 5865
rect 32401 5899 32459 5905
rect 32401 5865 32413 5899
rect 32447 5896 32459 5899
rect 32674 5896 32680 5908
rect 32447 5868 32680 5896
rect 32447 5865 32459 5868
rect 32401 5859 32459 5865
rect 32674 5856 32680 5868
rect 32732 5856 32738 5908
rect 33686 5856 33692 5908
rect 33744 5896 33750 5908
rect 34149 5899 34207 5905
rect 34149 5896 34161 5899
rect 33744 5868 34161 5896
rect 33744 5856 33750 5868
rect 34149 5865 34161 5868
rect 34195 5896 34207 5899
rect 35158 5896 35164 5908
rect 34195 5868 35164 5896
rect 34195 5865 34207 5868
rect 34149 5859 34207 5865
rect 1854 5788 1860 5840
rect 1912 5828 1918 5840
rect 3789 5831 3847 5837
rect 3789 5828 3801 5831
rect 1912 5800 3801 5828
rect 1912 5788 1918 5800
rect 3789 5797 3801 5800
rect 3835 5797 3847 5831
rect 3789 5791 3847 5797
rect 7098 5788 7104 5840
rect 7156 5828 7162 5840
rect 8297 5831 8355 5837
rect 8297 5828 8309 5831
rect 7156 5800 8309 5828
rect 7156 5788 7162 5800
rect 8297 5797 8309 5800
rect 8343 5797 8355 5831
rect 8297 5791 8355 5797
rect 8386 5788 8392 5840
rect 8444 5828 8450 5840
rect 8444 5800 8489 5828
rect 8444 5788 8450 5800
rect 8570 5788 8576 5840
rect 8628 5828 8634 5840
rect 9858 5828 9864 5840
rect 8628 5800 9864 5828
rect 8628 5788 8634 5800
rect 9858 5788 9864 5800
rect 9916 5828 9922 5840
rect 10045 5831 10103 5837
rect 10045 5828 10057 5831
rect 9916 5800 10057 5828
rect 9916 5788 9922 5800
rect 10045 5797 10057 5800
rect 10091 5797 10103 5831
rect 10045 5791 10103 5797
rect 10229 5831 10287 5837
rect 10229 5797 10241 5831
rect 10275 5828 10287 5831
rect 10594 5828 10600 5840
rect 10275 5800 10600 5828
rect 10275 5797 10287 5800
rect 10229 5791 10287 5797
rect 10594 5788 10600 5800
rect 10652 5788 10658 5840
rect 12526 5788 12532 5840
rect 12584 5828 12590 5840
rect 12621 5831 12679 5837
rect 12621 5828 12633 5831
rect 12584 5800 12633 5828
rect 12584 5788 12590 5800
rect 12621 5797 12633 5800
rect 12667 5828 12679 5831
rect 13081 5831 13139 5837
rect 13081 5828 13093 5831
rect 12667 5800 13093 5828
rect 12667 5797 12679 5800
rect 12621 5791 12679 5797
rect 13081 5797 13093 5800
rect 13127 5797 13139 5831
rect 13081 5791 13139 5797
rect 14185 5831 14243 5837
rect 14185 5797 14197 5831
rect 14231 5828 14243 5831
rect 14734 5828 14740 5840
rect 14231 5800 14740 5828
rect 14231 5797 14243 5800
rect 14185 5791 14243 5797
rect 14734 5788 14740 5800
rect 14792 5788 14798 5840
rect 18138 5788 18144 5840
rect 18196 5828 18202 5840
rect 18325 5831 18383 5837
rect 18325 5828 18337 5831
rect 18196 5800 18337 5828
rect 18196 5788 18202 5800
rect 18325 5797 18337 5800
rect 18371 5797 18383 5831
rect 18325 5791 18383 5797
rect 18601 5831 18659 5837
rect 18601 5797 18613 5831
rect 18647 5828 18659 5831
rect 20162 5828 20168 5840
rect 18647 5800 20168 5828
rect 18647 5797 18659 5800
rect 18601 5791 18659 5797
rect 1486 5760 1492 5772
rect 1447 5732 1492 5760
rect 1486 5720 1492 5732
rect 1544 5720 1550 5772
rect 1756 5763 1814 5769
rect 1756 5729 1768 5763
rect 1802 5760 1814 5763
rect 2774 5760 2780 5772
rect 1802 5732 2780 5760
rect 1802 5729 1814 5732
rect 1756 5723 1814 5729
rect 2774 5720 2780 5732
rect 2832 5720 2838 5772
rect 3510 5760 3516 5772
rect 3471 5732 3516 5760
rect 3510 5720 3516 5732
rect 3568 5720 3574 5772
rect 4065 5763 4123 5769
rect 4065 5760 4077 5763
rect 3988 5732 4077 5760
rect 3988 5704 4016 5732
rect 4065 5729 4077 5732
rect 4111 5729 4123 5763
rect 4065 5723 4123 5729
rect 5261 5763 5319 5769
rect 5261 5729 5273 5763
rect 5307 5760 5319 5763
rect 5350 5760 5356 5772
rect 5307 5732 5356 5760
rect 5307 5729 5319 5732
rect 5261 5723 5319 5729
rect 5350 5720 5356 5732
rect 5408 5720 5414 5772
rect 5534 5769 5540 5772
rect 5528 5760 5540 5769
rect 5495 5732 5540 5760
rect 5528 5723 5540 5732
rect 5534 5720 5540 5723
rect 5592 5720 5598 5772
rect 12342 5720 12348 5772
rect 12400 5760 12406 5772
rect 12437 5763 12495 5769
rect 12437 5760 12449 5763
rect 12400 5732 12449 5760
rect 12400 5720 12406 5732
rect 12437 5729 12449 5732
rect 12483 5760 12495 5763
rect 12802 5760 12808 5772
rect 12483 5732 12808 5760
rect 12483 5729 12495 5732
rect 12437 5723 12495 5729
rect 12802 5720 12808 5732
rect 12860 5720 12866 5772
rect 15746 5769 15752 5772
rect 15729 5763 15752 5769
rect 15729 5760 15741 5763
rect 14292 5732 15741 5760
rect 3970 5652 3976 5704
rect 4028 5652 4034 5704
rect 8202 5692 8208 5704
rect 8163 5664 8208 5692
rect 8202 5652 8208 5664
rect 8260 5652 8266 5704
rect 10318 5692 10324 5704
rect 10279 5664 10324 5692
rect 10318 5652 10324 5664
rect 10376 5652 10382 5704
rect 12710 5692 12716 5704
rect 12671 5664 12716 5692
rect 12710 5652 12716 5664
rect 12768 5652 12774 5704
rect 14093 5695 14151 5701
rect 14093 5692 14105 5695
rect 13464 5664 14105 5692
rect 4062 5584 4068 5636
rect 4120 5624 4126 5636
rect 4249 5627 4307 5633
rect 4249 5624 4261 5627
rect 4120 5596 4261 5624
rect 4120 5584 4126 5596
rect 4249 5593 4261 5596
rect 4295 5593 4307 5627
rect 4249 5587 4307 5593
rect 7190 5584 7196 5636
rect 7248 5624 7254 5636
rect 7837 5627 7895 5633
rect 7837 5624 7849 5627
rect 7248 5596 7849 5624
rect 7248 5584 7254 5596
rect 7837 5593 7849 5596
rect 7883 5593 7895 5627
rect 7837 5587 7895 5593
rect 9490 5584 9496 5636
rect 9548 5624 9554 5636
rect 13464 5633 13492 5664
rect 14093 5661 14105 5664
rect 14139 5661 14151 5695
rect 14093 5655 14151 5661
rect 14182 5652 14188 5704
rect 14240 5692 14246 5704
rect 14292 5701 14320 5732
rect 15729 5729 15741 5732
rect 15804 5760 15810 5772
rect 18340 5760 18368 5791
rect 20162 5788 20168 5800
rect 20220 5828 20226 5840
rect 20257 5831 20315 5837
rect 20257 5828 20269 5831
rect 20220 5800 20269 5828
rect 20220 5788 20226 5800
rect 20257 5797 20269 5800
rect 20303 5797 20315 5831
rect 20257 5791 20315 5797
rect 21720 5831 21778 5837
rect 21720 5797 21732 5831
rect 21766 5828 21778 5831
rect 21818 5828 21824 5840
rect 21766 5800 21824 5828
rect 21766 5797 21778 5800
rect 21720 5791 21778 5797
rect 21818 5788 21824 5800
rect 21876 5828 21882 5840
rect 22462 5828 22468 5840
rect 21876 5800 22468 5828
rect 21876 5788 21882 5800
rect 22462 5788 22468 5800
rect 22520 5788 22526 5840
rect 27798 5788 27804 5840
rect 27856 5828 27862 5840
rect 28169 5831 28227 5837
rect 28169 5828 28181 5831
rect 27856 5800 28181 5828
rect 27856 5788 27862 5800
rect 28169 5797 28181 5800
rect 28215 5828 28227 5831
rect 28534 5828 28540 5840
rect 28215 5800 28540 5828
rect 28215 5797 28227 5800
rect 28169 5791 28227 5797
rect 28534 5788 28540 5800
rect 28592 5788 28598 5840
rect 29546 5828 29552 5840
rect 29507 5800 29552 5828
rect 29546 5788 29552 5800
rect 29604 5828 29610 5840
rect 30374 5828 30380 5840
rect 29604 5800 30380 5828
rect 29604 5788 29610 5800
rect 30374 5788 30380 5800
rect 30432 5788 30438 5840
rect 33321 5831 33379 5837
rect 33321 5797 33333 5831
rect 33367 5828 33379 5831
rect 33410 5828 33416 5840
rect 33367 5800 33416 5828
rect 33367 5797 33379 5800
rect 33321 5791 33379 5797
rect 33410 5788 33416 5800
rect 33468 5788 33474 5840
rect 34238 5788 34244 5840
rect 34296 5828 34302 5840
rect 34992 5837 35020 5868
rect 35158 5856 35164 5868
rect 35216 5896 35222 5908
rect 35713 5899 35771 5905
rect 35713 5896 35725 5899
rect 35216 5868 35725 5896
rect 35216 5856 35222 5868
rect 35713 5865 35725 5868
rect 35759 5865 35771 5899
rect 36078 5896 36084 5908
rect 36039 5868 36084 5896
rect 35713 5859 35771 5865
rect 36078 5856 36084 5868
rect 36136 5856 36142 5908
rect 34885 5831 34943 5837
rect 34885 5828 34897 5831
rect 34296 5800 34897 5828
rect 34296 5788 34302 5800
rect 34885 5797 34897 5800
rect 34931 5797 34943 5831
rect 34885 5791 34943 5797
rect 34977 5831 35035 5837
rect 34977 5797 34989 5831
rect 35023 5797 35035 5831
rect 34977 5791 35035 5797
rect 19334 5760 19340 5772
rect 15804 5732 15877 5760
rect 18340 5732 19340 5760
rect 15729 5723 15752 5729
rect 15746 5720 15752 5723
rect 15804 5720 15810 5732
rect 19334 5720 19340 5732
rect 19392 5720 19398 5772
rect 24210 5769 24216 5772
rect 24204 5760 24216 5769
rect 24171 5732 24216 5760
rect 24204 5723 24216 5732
rect 24210 5720 24216 5723
rect 24268 5720 24274 5772
rect 27985 5763 28043 5769
rect 27985 5729 27997 5763
rect 28031 5760 28043 5763
rect 28350 5760 28356 5772
rect 28031 5732 28356 5760
rect 28031 5729 28043 5732
rect 27985 5723 28043 5729
rect 28350 5720 28356 5732
rect 28408 5720 28414 5772
rect 33226 5720 33232 5772
rect 33284 5760 33290 5772
rect 34422 5760 34428 5772
rect 33284 5732 34428 5760
rect 33284 5720 33290 5732
rect 14277 5695 14335 5701
rect 14277 5692 14289 5695
rect 14240 5664 14289 5692
rect 14240 5652 14246 5664
rect 14277 5661 14289 5664
rect 14323 5661 14335 5695
rect 15470 5692 15476 5704
rect 15431 5664 15476 5692
rect 14277 5655 14335 5661
rect 15470 5652 15476 5664
rect 15528 5652 15534 5704
rect 21082 5692 21088 5704
rect 20995 5664 21088 5692
rect 21082 5652 21088 5664
rect 21140 5692 21146 5704
rect 21450 5692 21456 5704
rect 21140 5664 21456 5692
rect 21140 5652 21146 5664
rect 21450 5652 21456 5664
rect 21508 5652 21514 5704
rect 23934 5692 23940 5704
rect 23895 5664 23940 5692
rect 23934 5652 23940 5664
rect 23992 5652 23998 5704
rect 26326 5652 26332 5704
rect 26384 5692 26390 5704
rect 28258 5692 28264 5704
rect 26384 5664 28120 5692
rect 28219 5664 28264 5692
rect 26384 5652 26390 5664
rect 9769 5627 9827 5633
rect 9769 5624 9781 5627
rect 9548 5596 9781 5624
rect 9548 5584 9554 5596
rect 9769 5593 9781 5596
rect 9815 5593 9827 5627
rect 9769 5587 9827 5593
rect 12161 5627 12219 5633
rect 12161 5593 12173 5627
rect 12207 5624 12219 5627
rect 13449 5627 13507 5633
rect 13449 5624 13461 5627
rect 12207 5596 13461 5624
rect 12207 5593 12219 5596
rect 12161 5587 12219 5593
rect 13449 5593 13461 5596
rect 13495 5593 13507 5627
rect 13449 5587 13507 5593
rect 17862 5584 17868 5636
rect 17920 5624 17926 5636
rect 18049 5627 18107 5633
rect 18049 5624 18061 5627
rect 17920 5596 18061 5624
rect 17920 5584 17926 5596
rect 18049 5593 18061 5596
rect 18095 5593 18107 5627
rect 18049 5587 18107 5593
rect 11054 5516 11060 5568
rect 11112 5556 11118 5568
rect 11698 5556 11704 5568
rect 11112 5528 11704 5556
rect 11112 5516 11118 5528
rect 11698 5516 11704 5528
rect 11756 5516 11762 5568
rect 13722 5556 13728 5568
rect 13683 5528 13728 5556
rect 13722 5516 13728 5528
rect 13780 5516 13786 5568
rect 16850 5556 16856 5568
rect 16811 5528 16856 5556
rect 16850 5516 16856 5528
rect 16908 5516 16914 5568
rect 18874 5516 18880 5568
rect 18932 5556 18938 5568
rect 19978 5556 19984 5568
rect 18932 5528 19984 5556
rect 18932 5516 18938 5528
rect 19978 5516 19984 5528
rect 20036 5556 20042 5568
rect 21100 5565 21128 5652
rect 26053 5627 26111 5633
rect 26053 5593 26065 5627
rect 26099 5624 26111 5627
rect 26602 5624 26608 5636
rect 26099 5596 26608 5624
rect 26099 5593 26111 5596
rect 26053 5587 26111 5593
rect 26602 5584 26608 5596
rect 26660 5624 26666 5636
rect 28092 5624 28120 5664
rect 28258 5652 28264 5664
rect 28316 5652 28322 5704
rect 29270 5652 29276 5704
rect 29328 5692 29334 5704
rect 29825 5695 29883 5701
rect 29825 5692 29837 5695
rect 29328 5664 29837 5692
rect 29328 5652 29334 5664
rect 29825 5661 29837 5664
rect 29871 5661 29883 5695
rect 33318 5692 33324 5704
rect 33279 5664 33324 5692
rect 29825 5655 29883 5661
rect 33318 5652 33324 5664
rect 33376 5652 33382 5704
rect 33428 5701 33456 5732
rect 34422 5720 34428 5732
rect 34480 5720 34486 5772
rect 34701 5763 34759 5769
rect 34701 5729 34713 5763
rect 34747 5760 34759 5763
rect 35710 5760 35716 5772
rect 34747 5732 35716 5760
rect 34747 5729 34759 5732
rect 34701 5723 34759 5729
rect 33413 5695 33471 5701
rect 33413 5661 33425 5695
rect 33459 5661 33471 5695
rect 33413 5655 33471 5661
rect 34606 5652 34612 5704
rect 34664 5692 34670 5704
rect 34716 5692 34744 5723
rect 35710 5720 35716 5732
rect 35768 5720 35774 5772
rect 35894 5760 35900 5772
rect 35855 5732 35900 5760
rect 35894 5720 35900 5732
rect 35952 5720 35958 5772
rect 34664 5664 34744 5692
rect 34664 5652 34670 5664
rect 34974 5652 34980 5704
rect 35032 5692 35038 5704
rect 35345 5695 35403 5701
rect 35345 5692 35357 5695
rect 35032 5664 35357 5692
rect 35032 5652 35038 5664
rect 35345 5661 35357 5664
rect 35391 5661 35403 5695
rect 35345 5655 35403 5661
rect 28810 5624 28816 5636
rect 26660 5596 27200 5624
rect 28092 5596 28816 5624
rect 26660 5584 26666 5596
rect 27172 5568 27200 5596
rect 28810 5584 28816 5596
rect 28868 5584 28874 5636
rect 32766 5584 32772 5636
rect 32824 5624 32830 5636
rect 32861 5627 32919 5633
rect 32861 5624 32873 5627
rect 32824 5596 32873 5624
rect 32824 5584 32830 5596
rect 32861 5593 32873 5596
rect 32907 5593 32919 5627
rect 32861 5587 32919 5593
rect 34054 5584 34060 5636
rect 34112 5624 34118 5636
rect 34425 5627 34483 5633
rect 34425 5624 34437 5627
rect 34112 5596 34437 5624
rect 34112 5584 34118 5596
rect 34425 5593 34437 5596
rect 34471 5593 34483 5627
rect 34425 5587 34483 5593
rect 21085 5559 21143 5565
rect 21085 5556 21097 5559
rect 20036 5528 21097 5556
rect 20036 5516 20042 5528
rect 21085 5525 21097 5528
rect 21131 5525 21143 5559
rect 22830 5556 22836 5568
rect 22791 5528 22836 5556
rect 21085 5519 21143 5525
rect 22830 5516 22836 5528
rect 22888 5516 22894 5568
rect 25317 5559 25375 5565
rect 25317 5525 25329 5559
rect 25363 5556 25375 5559
rect 25682 5556 25688 5568
rect 25363 5528 25688 5556
rect 25363 5525 25375 5528
rect 25317 5519 25375 5525
rect 25682 5516 25688 5528
rect 25740 5516 25746 5568
rect 26694 5556 26700 5568
rect 26655 5528 26700 5556
rect 26694 5516 26700 5528
rect 26752 5516 26758 5568
rect 27154 5556 27160 5568
rect 27115 5528 27160 5556
rect 27154 5516 27160 5528
rect 27212 5516 27218 5568
rect 29273 5559 29331 5565
rect 29273 5525 29285 5559
rect 29319 5556 29331 5559
rect 29822 5556 29828 5568
rect 29319 5528 29828 5556
rect 29319 5525 29331 5528
rect 29273 5519 29331 5525
rect 29822 5516 29828 5528
rect 29880 5516 29886 5568
rect 1104 5466 38824 5488
rect 1104 5414 7648 5466
rect 7700 5414 7712 5466
rect 7764 5414 7776 5466
rect 7828 5414 7840 5466
rect 7892 5414 20982 5466
rect 21034 5414 21046 5466
rect 21098 5414 21110 5466
rect 21162 5414 21174 5466
rect 21226 5414 34315 5466
rect 34367 5414 34379 5466
rect 34431 5414 34443 5466
rect 34495 5414 34507 5466
rect 34559 5414 38824 5466
rect 1104 5392 38824 5414
rect 1949 5355 2007 5361
rect 1949 5321 1961 5355
rect 1995 5352 2007 5355
rect 2590 5352 2596 5364
rect 1995 5324 2596 5352
rect 1995 5321 2007 5324
rect 1949 5315 2007 5321
rect 2590 5312 2596 5324
rect 2648 5312 2654 5364
rect 2958 5312 2964 5364
rect 3016 5352 3022 5364
rect 3053 5355 3111 5361
rect 3053 5352 3065 5355
rect 3016 5324 3065 5352
rect 3016 5312 3022 5324
rect 3053 5321 3065 5324
rect 3099 5321 3111 5355
rect 3053 5315 3111 5321
rect 3697 5355 3755 5361
rect 3697 5321 3709 5355
rect 3743 5352 3755 5355
rect 4062 5352 4068 5364
rect 3743 5324 4068 5352
rect 3743 5321 3755 5324
rect 3697 5315 3755 5321
rect 4062 5312 4068 5324
rect 4120 5312 4126 5364
rect 5350 5352 5356 5364
rect 5311 5324 5356 5352
rect 5350 5312 5356 5324
rect 5408 5312 5414 5364
rect 7006 5352 7012 5364
rect 6967 5324 7012 5352
rect 7006 5312 7012 5324
rect 7064 5312 7070 5364
rect 7098 5312 7104 5364
rect 7156 5352 7162 5364
rect 7377 5355 7435 5361
rect 7377 5352 7389 5355
rect 7156 5324 7389 5352
rect 7156 5312 7162 5324
rect 7377 5321 7389 5324
rect 7423 5321 7435 5355
rect 7377 5315 7435 5321
rect 8110 5312 8116 5364
rect 8168 5352 8174 5364
rect 8297 5355 8355 5361
rect 8297 5352 8309 5355
rect 8168 5324 8309 5352
rect 8168 5312 8174 5324
rect 8297 5321 8309 5324
rect 8343 5321 8355 5355
rect 8297 5315 8355 5321
rect 2133 5287 2191 5293
rect 2133 5253 2145 5287
rect 2179 5253 2191 5287
rect 3326 5284 3332 5296
rect 2133 5247 2191 5253
rect 2608 5256 3332 5284
rect 2148 5148 2176 5247
rect 2498 5176 2504 5228
rect 2556 5216 2562 5228
rect 2608 5225 2636 5256
rect 3326 5244 3332 5256
rect 3384 5244 3390 5296
rect 2593 5219 2651 5225
rect 2593 5216 2605 5219
rect 2556 5188 2605 5216
rect 2556 5176 2562 5188
rect 2593 5185 2605 5188
rect 2639 5185 2651 5219
rect 2593 5179 2651 5185
rect 2685 5219 2743 5225
rect 2685 5185 2697 5219
rect 2731 5216 2743 5219
rect 2866 5216 2872 5228
rect 2731 5188 2872 5216
rect 2731 5185 2743 5188
rect 2685 5179 2743 5185
rect 2866 5176 2872 5188
rect 2924 5176 2930 5228
rect 3878 5176 3884 5228
rect 3936 5216 3942 5228
rect 4249 5219 4307 5225
rect 4249 5216 4261 5219
rect 3936 5188 4261 5216
rect 3936 5176 3942 5188
rect 4249 5185 4261 5188
rect 4295 5216 4307 5219
rect 5534 5216 5540 5228
rect 4295 5188 5540 5216
rect 4295 5185 4307 5188
rect 4249 5179 4307 5185
rect 5534 5176 5540 5188
rect 5592 5216 5598 5228
rect 5629 5219 5687 5225
rect 5629 5216 5641 5219
rect 5592 5188 5641 5216
rect 5592 5176 5598 5188
rect 5629 5185 5641 5188
rect 5675 5185 5687 5219
rect 8312 5216 8340 5315
rect 10318 5312 10324 5364
rect 10376 5352 10382 5364
rect 10689 5355 10747 5361
rect 10689 5352 10701 5355
rect 10376 5324 10701 5352
rect 10376 5312 10382 5324
rect 10689 5321 10701 5324
rect 10735 5321 10747 5355
rect 10689 5315 10747 5321
rect 11425 5355 11483 5361
rect 11425 5321 11437 5355
rect 11471 5352 11483 5355
rect 12710 5352 12716 5364
rect 11471 5324 12716 5352
rect 11471 5321 11483 5324
rect 11425 5315 11483 5321
rect 12710 5312 12716 5324
rect 12768 5352 12774 5364
rect 13817 5355 13875 5361
rect 13817 5352 13829 5355
rect 12768 5324 13829 5352
rect 12768 5312 12774 5324
rect 13817 5321 13829 5324
rect 13863 5352 13875 5355
rect 14826 5352 14832 5364
rect 13863 5324 14832 5352
rect 13863 5321 13875 5324
rect 13817 5315 13875 5321
rect 14826 5312 14832 5324
rect 14884 5312 14890 5364
rect 15562 5352 15568 5364
rect 15523 5324 15568 5352
rect 15562 5312 15568 5324
rect 15620 5312 15626 5364
rect 17126 5352 17132 5364
rect 17087 5324 17132 5352
rect 17126 5312 17132 5324
rect 17184 5312 17190 5364
rect 17865 5355 17923 5361
rect 17865 5321 17877 5355
rect 17911 5352 17923 5355
rect 18322 5352 18328 5364
rect 17911 5324 18328 5352
rect 17911 5321 17923 5324
rect 17865 5315 17923 5321
rect 18322 5312 18328 5324
rect 18380 5312 18386 5364
rect 19058 5352 19064 5364
rect 19019 5324 19064 5352
rect 19058 5312 19064 5324
rect 19116 5312 19122 5364
rect 19334 5312 19340 5364
rect 19392 5352 19398 5364
rect 19429 5355 19487 5361
rect 19429 5352 19441 5355
rect 19392 5324 19441 5352
rect 19392 5312 19398 5324
rect 19429 5321 19441 5324
rect 19475 5321 19487 5355
rect 20254 5352 20260 5364
rect 20215 5324 20260 5352
rect 19429 5315 19487 5321
rect 20254 5312 20260 5324
rect 20312 5312 20318 5364
rect 21450 5312 21456 5364
rect 21508 5352 21514 5364
rect 22094 5352 22100 5364
rect 21508 5324 22100 5352
rect 21508 5312 21514 5324
rect 22094 5312 22100 5324
rect 22152 5352 22158 5364
rect 22189 5355 22247 5361
rect 22189 5352 22201 5355
rect 22152 5324 22201 5352
rect 22152 5312 22158 5324
rect 22189 5321 22201 5324
rect 22235 5352 22247 5355
rect 23934 5352 23940 5364
rect 22235 5324 23940 5352
rect 22235 5321 22247 5324
rect 22189 5315 22247 5321
rect 23934 5312 23940 5324
rect 23992 5312 23998 5364
rect 24762 5352 24768 5364
rect 24723 5324 24768 5352
rect 24762 5312 24768 5324
rect 24820 5312 24826 5364
rect 26694 5352 26700 5364
rect 25608 5324 26700 5352
rect 14642 5244 14648 5296
rect 14700 5284 14706 5296
rect 16025 5287 16083 5293
rect 16025 5284 16037 5287
rect 14700 5256 16037 5284
rect 14700 5244 14706 5256
rect 16025 5253 16037 5256
rect 16071 5253 16083 5287
rect 18141 5287 18199 5293
rect 18141 5284 18153 5287
rect 16025 5247 16083 5253
rect 16408 5256 18153 5284
rect 8389 5219 8447 5225
rect 8389 5216 8401 5219
rect 8312 5188 8401 5216
rect 5629 5179 5687 5185
rect 8389 5185 8401 5188
rect 8435 5185 8447 5219
rect 8389 5179 8447 5185
rect 16114 5176 16120 5228
rect 16172 5216 16178 5228
rect 16408 5225 16436 5256
rect 18141 5253 18153 5256
rect 18187 5253 18199 5287
rect 18141 5247 18199 5253
rect 21269 5287 21327 5293
rect 21269 5253 21281 5287
rect 21315 5284 21327 5287
rect 22370 5284 22376 5296
rect 21315 5256 22376 5284
rect 21315 5253 21327 5256
rect 21269 5247 21327 5253
rect 22370 5244 22376 5256
rect 22428 5244 22434 5296
rect 23952 5284 23980 5312
rect 25409 5287 25467 5293
rect 25409 5284 25421 5287
rect 23952 5256 25421 5284
rect 25409 5253 25421 5256
rect 25455 5284 25467 5287
rect 25608 5284 25636 5324
rect 26694 5312 26700 5324
rect 26752 5312 26758 5364
rect 26973 5355 27031 5361
rect 26973 5321 26985 5355
rect 27019 5352 27031 5355
rect 27154 5352 27160 5364
rect 27019 5324 27160 5352
rect 27019 5321 27031 5324
rect 26973 5315 27031 5321
rect 27154 5312 27160 5324
rect 27212 5312 27218 5364
rect 27709 5355 27767 5361
rect 27709 5321 27721 5355
rect 27755 5352 27767 5355
rect 27798 5352 27804 5364
rect 27755 5324 27804 5352
rect 27755 5321 27767 5324
rect 27709 5315 27767 5321
rect 27798 5312 27804 5324
rect 27856 5312 27862 5364
rect 28077 5355 28135 5361
rect 28077 5321 28089 5355
rect 28123 5352 28135 5355
rect 28350 5352 28356 5364
rect 28123 5324 28356 5352
rect 28123 5321 28135 5324
rect 28077 5315 28135 5321
rect 28350 5312 28356 5324
rect 28408 5312 28414 5364
rect 29362 5352 29368 5364
rect 29323 5324 29368 5352
rect 29362 5312 29368 5324
rect 29420 5312 29426 5364
rect 30374 5352 30380 5364
rect 30335 5324 30380 5352
rect 30374 5312 30380 5324
rect 30432 5312 30438 5364
rect 31757 5355 31815 5361
rect 31757 5321 31769 5355
rect 31803 5352 31815 5355
rect 33042 5352 33048 5364
rect 31803 5324 33048 5352
rect 31803 5321 31815 5324
rect 31757 5315 31815 5321
rect 33042 5312 33048 5324
rect 33100 5312 33106 5364
rect 34146 5312 34152 5364
rect 34204 5352 34210 5364
rect 34241 5355 34299 5361
rect 34241 5352 34253 5355
rect 34204 5324 34253 5352
rect 34204 5312 34210 5324
rect 34241 5321 34253 5324
rect 34287 5321 34299 5355
rect 34698 5352 34704 5364
rect 34659 5324 34704 5352
rect 34241 5315 34299 5321
rect 34698 5312 34704 5324
rect 34756 5312 34762 5364
rect 36630 5352 36636 5364
rect 36591 5324 36636 5352
rect 36630 5312 36636 5324
rect 36688 5312 36694 5364
rect 25455 5256 25636 5284
rect 25455 5253 25467 5256
rect 25409 5247 25467 5253
rect 16393 5219 16451 5225
rect 16393 5216 16405 5219
rect 16172 5188 16405 5216
rect 16172 5176 16178 5188
rect 16393 5185 16405 5188
rect 16439 5185 16451 5219
rect 16574 5216 16580 5228
rect 16535 5188 16580 5216
rect 16393 5179 16451 5185
rect 16574 5176 16580 5188
rect 16632 5176 16638 5228
rect 21085 5219 21143 5225
rect 21085 5185 21097 5219
rect 21131 5216 21143 5219
rect 21818 5216 21824 5228
rect 21131 5188 21824 5216
rect 21131 5185 21143 5188
rect 21085 5179 21143 5185
rect 21818 5176 21824 5188
rect 21876 5176 21882 5228
rect 25608 5225 25636 5256
rect 29089 5287 29147 5293
rect 29089 5253 29101 5287
rect 29135 5284 29147 5287
rect 29270 5284 29276 5296
rect 29135 5256 29276 5284
rect 29135 5253 29147 5256
rect 29089 5247 29147 5253
rect 29270 5244 29276 5256
rect 29328 5244 29334 5296
rect 32582 5244 32588 5296
rect 32640 5284 32646 5296
rect 32677 5287 32735 5293
rect 32677 5284 32689 5287
rect 32640 5256 32689 5284
rect 32640 5244 32646 5256
rect 32677 5253 32689 5256
rect 32723 5253 32735 5287
rect 33965 5287 34023 5293
rect 32677 5247 32735 5253
rect 32784 5256 33272 5284
rect 32784 5228 32812 5256
rect 33244 5228 33272 5256
rect 33965 5253 33977 5287
rect 34011 5284 34023 5287
rect 34606 5284 34612 5296
rect 34011 5256 34612 5284
rect 34011 5253 34023 5256
rect 33965 5247 34023 5253
rect 34606 5244 34612 5256
rect 34664 5244 34670 5296
rect 34974 5284 34980 5296
rect 34935 5256 34980 5284
rect 34974 5244 34980 5256
rect 35032 5244 35038 5296
rect 25593 5219 25651 5225
rect 25593 5185 25605 5219
rect 25639 5185 25651 5219
rect 29914 5216 29920 5228
rect 29875 5188 29920 5216
rect 25593 5179 25651 5185
rect 29914 5176 29920 5188
rect 29972 5176 29978 5228
rect 32493 5219 32551 5225
rect 32493 5185 32505 5219
rect 32539 5216 32551 5219
rect 32766 5216 32772 5228
rect 32539 5188 32772 5216
rect 32539 5185 32551 5188
rect 32493 5179 32551 5185
rect 32766 5176 32772 5188
rect 32824 5176 32830 5228
rect 32858 5176 32864 5228
rect 32916 5216 32922 5228
rect 33045 5219 33103 5225
rect 33045 5216 33057 5219
rect 32916 5188 33057 5216
rect 32916 5176 32922 5188
rect 33045 5185 33057 5188
rect 33091 5185 33103 5219
rect 33226 5216 33232 5228
rect 33187 5188 33232 5216
rect 33045 5179 33103 5185
rect 33226 5176 33232 5188
rect 33284 5176 33290 5228
rect 35158 5176 35164 5228
rect 35216 5216 35222 5228
rect 35529 5219 35587 5225
rect 35529 5216 35541 5219
rect 35216 5188 35541 5216
rect 35216 5176 35222 5188
rect 35529 5185 35541 5188
rect 35575 5185 35587 5219
rect 35529 5179 35587 5185
rect 11793 5151 11851 5157
rect 2148 5120 4200 5148
rect 4172 5092 4200 5120
rect 11793 5117 11805 5151
rect 11839 5148 11851 5151
rect 12437 5151 12495 5157
rect 12437 5148 12449 5151
rect 11839 5120 12449 5148
rect 11839 5117 11851 5120
rect 11793 5111 11851 5117
rect 12437 5117 12449 5120
rect 12483 5148 12495 5151
rect 13538 5148 13544 5160
rect 12483 5120 13544 5148
rect 12483 5117 12495 5120
rect 12437 5111 12495 5117
rect 13538 5108 13544 5120
rect 13596 5108 13602 5160
rect 20717 5151 20775 5157
rect 20717 5117 20729 5151
rect 20763 5148 20775 5151
rect 20763 5120 21772 5148
rect 20763 5117 20775 5120
rect 20717 5111 20775 5117
rect 21744 5092 21772 5120
rect 25682 5108 25688 5160
rect 25740 5148 25746 5160
rect 25849 5151 25907 5157
rect 25849 5148 25861 5151
rect 25740 5120 25861 5148
rect 25740 5108 25746 5120
rect 25849 5117 25861 5120
rect 25895 5117 25907 5151
rect 25849 5111 25907 5117
rect 28258 5108 28264 5160
rect 28316 5148 28322 5160
rect 28353 5151 28411 5157
rect 28353 5148 28365 5151
rect 28316 5120 28365 5148
rect 28316 5108 28322 5120
rect 28353 5117 28365 5120
rect 28399 5117 28411 5151
rect 28353 5111 28411 5117
rect 29546 5108 29552 5160
rect 29604 5148 29610 5160
rect 29641 5151 29699 5157
rect 29641 5148 29653 5151
rect 29604 5120 29653 5148
rect 29604 5108 29610 5120
rect 29641 5117 29653 5120
rect 29687 5148 29699 5151
rect 30653 5151 30711 5157
rect 30653 5148 30665 5151
rect 29687 5120 30665 5148
rect 29687 5117 29699 5120
rect 29641 5111 29699 5117
rect 30653 5117 30665 5120
rect 30699 5117 30711 5151
rect 30653 5111 30711 5117
rect 32125 5151 32183 5157
rect 32125 5117 32137 5151
rect 32171 5148 32183 5151
rect 33410 5148 33416 5160
rect 32171 5120 33416 5148
rect 32171 5117 32183 5120
rect 32125 5111 32183 5117
rect 33410 5108 33416 5120
rect 33468 5108 33474 5160
rect 34882 5108 34888 5160
rect 34940 5148 34946 5160
rect 35253 5151 35311 5157
rect 35253 5148 35265 5151
rect 34940 5120 35265 5148
rect 34940 5108 34946 5120
rect 35253 5117 35265 5120
rect 35299 5117 35311 5151
rect 35253 5111 35311 5117
rect 36449 5151 36507 5157
rect 36449 5117 36461 5151
rect 36495 5148 36507 5151
rect 37001 5151 37059 5157
rect 37001 5148 37013 5151
rect 36495 5120 37013 5148
rect 36495 5117 36507 5120
rect 36449 5111 36507 5117
rect 37001 5117 37013 5120
rect 37047 5117 37059 5151
rect 37001 5111 37059 5117
rect 2590 5040 2596 5092
rect 2648 5080 2654 5092
rect 2958 5080 2964 5092
rect 2648 5052 2964 5080
rect 2648 5040 2654 5052
rect 2958 5040 2964 5052
rect 3016 5080 3022 5092
rect 3142 5080 3148 5092
rect 3016 5052 3148 5080
rect 3016 5040 3022 5052
rect 3142 5040 3148 5052
rect 3200 5040 3206 5092
rect 3418 5040 3424 5092
rect 3476 5080 3482 5092
rect 3513 5083 3571 5089
rect 3513 5080 3525 5083
rect 3476 5052 3525 5080
rect 3476 5040 3482 5052
rect 3513 5049 3525 5052
rect 3559 5080 3571 5083
rect 3973 5083 4031 5089
rect 3973 5080 3985 5083
rect 3559 5052 3985 5080
rect 3559 5049 3571 5052
rect 3513 5043 3571 5049
rect 3973 5049 3985 5052
rect 4019 5049 4031 5083
rect 4154 5080 4160 5092
rect 4067 5052 4160 5080
rect 3973 5043 4031 5049
rect 3988 5012 4016 5043
rect 4154 5040 4160 5052
rect 4212 5040 4218 5092
rect 7837 5083 7895 5089
rect 7837 5049 7849 5083
rect 7883 5080 7895 5083
rect 8478 5080 8484 5092
rect 7883 5052 8484 5080
rect 7883 5049 7895 5052
rect 7837 5043 7895 5049
rect 8478 5040 8484 5052
rect 8536 5080 8542 5092
rect 8634 5083 8692 5089
rect 8634 5080 8646 5083
rect 8536 5052 8646 5080
rect 8536 5040 8542 5052
rect 8634 5049 8646 5052
rect 8680 5049 8692 5083
rect 8634 5043 8692 5049
rect 12250 5040 12256 5092
rect 12308 5080 12314 5092
rect 12682 5083 12740 5089
rect 12682 5080 12694 5083
rect 12308 5052 12694 5080
rect 12308 5040 12314 5052
rect 12682 5049 12694 5052
rect 12728 5080 12740 5083
rect 12986 5080 12992 5092
rect 12728 5052 12992 5080
rect 12728 5049 12740 5052
rect 12682 5043 12740 5049
rect 12986 5040 12992 5052
rect 13044 5040 13050 5092
rect 15105 5083 15163 5089
rect 15105 5080 15117 5083
rect 14384 5052 15117 5080
rect 4062 5012 4068 5024
rect 3988 4984 4068 5012
rect 4062 4972 4068 4984
rect 4120 4972 4126 5024
rect 4706 5012 4712 5024
rect 4667 4984 4712 5012
rect 4706 4972 4712 4984
rect 4764 4972 4770 5024
rect 9766 5012 9772 5024
rect 9727 4984 9772 5012
rect 9766 4972 9772 4984
rect 9824 4972 9830 5024
rect 10413 5015 10471 5021
rect 10413 4981 10425 5015
rect 10459 5012 10471 5015
rect 10594 5012 10600 5024
rect 10459 4984 10600 5012
rect 10459 4981 10471 4984
rect 10413 4975 10471 4981
rect 10594 4972 10600 4984
rect 10652 4972 10658 5024
rect 11974 4972 11980 5024
rect 12032 5012 12038 5024
rect 12069 5015 12127 5021
rect 12069 5012 12081 5015
rect 12032 4984 12081 5012
rect 12032 4972 12038 4984
rect 12069 4981 12081 4984
rect 12115 5012 12127 5015
rect 12342 5012 12348 5024
rect 12115 4984 12348 5012
rect 12115 4981 12127 4984
rect 12069 4975 12127 4981
rect 12342 4972 12348 4984
rect 12400 4972 12406 5024
rect 13538 4972 13544 5024
rect 13596 5012 13602 5024
rect 14182 5012 14188 5024
rect 13596 4984 14188 5012
rect 13596 4972 13602 4984
rect 14182 4972 14188 4984
rect 14240 5012 14246 5024
rect 14384 5021 14412 5052
rect 15105 5049 15117 5052
rect 15151 5049 15163 5083
rect 15105 5043 15163 5049
rect 18046 5040 18052 5092
rect 18104 5080 18110 5092
rect 18417 5083 18475 5089
rect 18417 5080 18429 5083
rect 18104 5052 18429 5080
rect 18104 5040 18110 5052
rect 18417 5049 18429 5052
rect 18463 5049 18475 5083
rect 18417 5043 18475 5049
rect 18506 5040 18512 5092
rect 18564 5080 18570 5092
rect 18693 5083 18751 5089
rect 18693 5080 18705 5083
rect 18564 5052 18705 5080
rect 18564 5040 18570 5052
rect 18693 5049 18705 5052
rect 18739 5080 18751 5083
rect 19150 5080 19156 5092
rect 18739 5052 19156 5080
rect 18739 5049 18751 5052
rect 18693 5043 18751 5049
rect 19150 5040 19156 5052
rect 19208 5040 19214 5092
rect 20254 5040 20260 5092
rect 20312 5080 20318 5092
rect 21545 5083 21603 5089
rect 21545 5080 21557 5083
rect 20312 5052 21557 5080
rect 20312 5040 20318 5052
rect 21545 5049 21557 5052
rect 21591 5049 21603 5083
rect 21726 5080 21732 5092
rect 21687 5052 21732 5080
rect 21545 5043 21603 5049
rect 21726 5040 21732 5052
rect 21784 5040 21790 5092
rect 22830 5040 22836 5092
rect 22888 5080 22894 5092
rect 24210 5080 24216 5092
rect 22888 5052 24216 5080
rect 22888 5040 22894 5052
rect 24210 5040 24216 5052
rect 24268 5080 24274 5092
rect 24305 5083 24363 5089
rect 24305 5080 24317 5083
rect 24268 5052 24317 5080
rect 24268 5040 24274 5052
rect 24305 5049 24317 5052
rect 24351 5049 24363 5083
rect 29822 5080 29828 5092
rect 29783 5052 29828 5080
rect 24305 5043 24363 5049
rect 29822 5040 29828 5052
rect 29880 5040 29886 5092
rect 33042 5040 33048 5092
rect 33100 5080 33106 5092
rect 33137 5083 33195 5089
rect 33137 5080 33149 5083
rect 33100 5052 33149 5080
rect 33100 5040 33106 5052
rect 33137 5049 33149 5052
rect 33183 5049 33195 5083
rect 36464 5080 36492 5111
rect 33137 5043 33195 5049
rect 34624 5052 36492 5080
rect 14369 5015 14427 5021
rect 14369 5012 14381 5015
rect 14240 4984 14381 5012
rect 14240 4972 14246 4984
rect 14369 4981 14381 4984
rect 14415 4981 14427 5015
rect 14734 5012 14740 5024
rect 14695 4984 14740 5012
rect 14369 4975 14427 4981
rect 14734 4972 14740 4984
rect 14792 4972 14798 5024
rect 16482 5012 16488 5024
rect 16443 4984 16488 5012
rect 16482 4972 16488 4984
rect 16540 4972 16546 5024
rect 17494 5012 17500 5024
rect 17455 4984 17500 5012
rect 17494 4972 17500 4984
rect 17552 4972 17558 5024
rect 18322 4972 18328 5024
rect 18380 5012 18386 5024
rect 18601 5015 18659 5021
rect 18601 5012 18613 5015
rect 18380 4984 18613 5012
rect 18380 4972 18386 4984
rect 18601 4981 18613 4984
rect 18647 4981 18659 5015
rect 18601 4975 18659 4981
rect 29178 4972 29184 5024
rect 29236 5012 29242 5024
rect 34624 5012 34652 5052
rect 29236 4984 34652 5012
rect 29236 4972 29242 4984
rect 34698 4972 34704 5024
rect 34756 5012 34762 5024
rect 35437 5015 35495 5021
rect 35437 5012 35449 5015
rect 34756 4984 35449 5012
rect 34756 4972 34762 4984
rect 35437 4981 35449 4984
rect 35483 5012 35495 5015
rect 35894 5012 35900 5024
rect 35483 4984 35900 5012
rect 35483 4981 35495 4984
rect 35437 4975 35495 4981
rect 35894 4972 35900 4984
rect 35952 4972 35958 5024
rect 1104 4922 38824 4944
rect 1104 4870 14315 4922
rect 14367 4870 14379 4922
rect 14431 4870 14443 4922
rect 14495 4870 14507 4922
rect 14559 4870 27648 4922
rect 27700 4870 27712 4922
rect 27764 4870 27776 4922
rect 27828 4870 27840 4922
rect 27892 4870 38824 4922
rect 1104 4848 38824 4870
rect 1394 4768 1400 4820
rect 1452 4808 1458 4820
rect 1581 4811 1639 4817
rect 1581 4808 1593 4811
rect 1452 4780 1593 4808
rect 1452 4768 1458 4780
rect 1581 4777 1593 4780
rect 1627 4777 1639 4811
rect 1581 4771 1639 4777
rect 2406 4768 2412 4820
rect 2464 4808 2470 4820
rect 2685 4811 2743 4817
rect 2685 4808 2697 4811
rect 2464 4780 2697 4808
rect 2464 4768 2470 4780
rect 2685 4777 2697 4780
rect 2731 4777 2743 4811
rect 2685 4771 2743 4777
rect 2866 4768 2872 4820
rect 2924 4808 2930 4820
rect 3421 4811 3479 4817
rect 3421 4808 3433 4811
rect 2924 4780 3433 4808
rect 2924 4768 2930 4780
rect 3421 4777 3433 4780
rect 3467 4777 3479 4811
rect 3878 4808 3884 4820
rect 3839 4780 3884 4808
rect 3421 4771 3479 4777
rect 3878 4768 3884 4780
rect 3936 4768 3942 4820
rect 4154 4768 4160 4820
rect 4212 4808 4218 4820
rect 4249 4811 4307 4817
rect 4249 4808 4261 4811
rect 4212 4780 4261 4808
rect 4212 4768 4218 4780
rect 4249 4777 4261 4780
rect 4295 4777 4307 4811
rect 4249 4771 4307 4777
rect 7469 4811 7527 4817
rect 7469 4777 7481 4811
rect 7515 4808 7527 4811
rect 8202 4808 8208 4820
rect 7515 4780 8208 4808
rect 7515 4777 7527 4780
rect 7469 4771 7527 4777
rect 8202 4768 8208 4780
rect 8260 4768 8266 4820
rect 8386 4768 8392 4820
rect 8444 4808 8450 4820
rect 8573 4811 8631 4817
rect 8573 4808 8585 4811
rect 8444 4780 8585 4808
rect 8444 4768 8450 4780
rect 8573 4777 8585 4780
rect 8619 4777 8631 4811
rect 9858 4808 9864 4820
rect 9819 4780 9864 4808
rect 8573 4771 8631 4777
rect 9858 4768 9864 4780
rect 9916 4768 9922 4820
rect 11885 4811 11943 4817
rect 11885 4777 11897 4811
rect 11931 4808 11943 4811
rect 12710 4808 12716 4820
rect 11931 4780 12716 4808
rect 11931 4777 11943 4780
rect 11885 4771 11943 4777
rect 12710 4768 12716 4780
rect 12768 4768 12774 4820
rect 12986 4808 12992 4820
rect 12947 4780 12992 4808
rect 12986 4768 12992 4780
rect 13044 4768 13050 4820
rect 13814 4768 13820 4820
rect 13872 4808 13878 4820
rect 14093 4811 14151 4817
rect 14093 4808 14105 4811
rect 13872 4780 14105 4808
rect 13872 4768 13878 4780
rect 14093 4777 14105 4780
rect 14139 4777 14151 4811
rect 14642 4808 14648 4820
rect 14603 4780 14648 4808
rect 14093 4771 14151 4777
rect 14642 4768 14648 4780
rect 14700 4768 14706 4820
rect 16117 4811 16175 4817
rect 16117 4777 16129 4811
rect 16163 4808 16175 4811
rect 16393 4811 16451 4817
rect 16393 4808 16405 4811
rect 16163 4780 16405 4808
rect 16163 4777 16175 4780
rect 16117 4771 16175 4777
rect 16393 4777 16405 4780
rect 16439 4808 16451 4811
rect 16574 4808 16580 4820
rect 16439 4780 16580 4808
rect 16439 4777 16451 4780
rect 16393 4771 16451 4777
rect 16574 4768 16580 4780
rect 16632 4768 16638 4820
rect 18046 4808 18052 4820
rect 18007 4780 18052 4808
rect 18046 4768 18052 4780
rect 18104 4768 18110 4820
rect 18966 4808 18972 4820
rect 18927 4780 18972 4808
rect 18966 4768 18972 4780
rect 19024 4768 19030 4820
rect 21545 4811 21603 4817
rect 21545 4777 21557 4811
rect 21591 4808 21603 4811
rect 21818 4808 21824 4820
rect 21591 4780 21824 4808
rect 21591 4777 21603 4780
rect 21545 4771 21603 4777
rect 21818 4768 21824 4780
rect 21876 4768 21882 4820
rect 22094 4768 22100 4820
rect 22152 4808 22158 4820
rect 22557 4811 22615 4817
rect 22557 4808 22569 4811
rect 22152 4780 22569 4808
rect 22152 4768 22158 4780
rect 22557 4777 22569 4780
rect 22603 4777 22615 4811
rect 25682 4808 25688 4820
rect 25643 4780 25688 4808
rect 22557 4771 22615 4777
rect 25682 4768 25688 4780
rect 25740 4808 25746 4820
rect 28258 4808 28264 4820
rect 25740 4780 28264 4808
rect 25740 4768 25746 4780
rect 2774 4700 2780 4752
rect 2832 4740 2838 4752
rect 3053 4743 3111 4749
rect 3053 4740 3065 4743
rect 2832 4712 3065 4740
rect 2832 4700 2838 4712
rect 3053 4709 3065 4712
rect 3099 4709 3111 4743
rect 8110 4740 8116 4752
rect 8071 4712 8116 4740
rect 3053 4703 3111 4709
rect 8110 4700 8116 4712
rect 8168 4700 8174 4752
rect 10962 4740 10968 4752
rect 10923 4712 10968 4740
rect 10962 4700 10968 4712
rect 11020 4700 11026 4752
rect 11517 4743 11575 4749
rect 11517 4709 11529 4743
rect 11563 4740 11575 4743
rect 12529 4743 12587 4749
rect 12529 4740 12541 4743
rect 11563 4712 12541 4740
rect 11563 4709 11575 4712
rect 11517 4703 11575 4709
rect 12529 4709 12541 4712
rect 12575 4740 12587 4743
rect 13615 4743 13673 4749
rect 13615 4740 13627 4743
rect 12575 4712 13627 4740
rect 12575 4709 12587 4712
rect 12529 4703 12587 4709
rect 13615 4709 13627 4712
rect 13661 4709 13673 4743
rect 13615 4703 13673 4709
rect 13909 4743 13967 4749
rect 13909 4709 13921 4743
rect 13955 4740 13967 4743
rect 13998 4740 14004 4752
rect 13955 4712 14004 4740
rect 13955 4709 13967 4712
rect 13909 4703 13967 4709
rect 13998 4700 14004 4712
rect 14056 4700 14062 4752
rect 15562 4700 15568 4752
rect 15620 4740 15626 4752
rect 15841 4743 15899 4749
rect 15841 4740 15853 4743
rect 15620 4712 15853 4740
rect 15620 4700 15626 4712
rect 15841 4709 15853 4712
rect 15887 4740 15899 4743
rect 16927 4743 16985 4749
rect 16927 4740 16939 4743
rect 15887 4712 16939 4740
rect 15887 4709 15899 4712
rect 15841 4703 15899 4709
rect 16927 4709 16939 4712
rect 16973 4709 16985 4743
rect 16927 4703 16985 4709
rect 17126 4700 17132 4752
rect 17184 4740 17190 4752
rect 17405 4743 17463 4749
rect 17405 4740 17417 4743
rect 17184 4712 17417 4740
rect 17184 4700 17190 4712
rect 17405 4709 17417 4712
rect 17451 4709 17463 4743
rect 18782 4740 18788 4752
rect 18743 4712 18788 4740
rect 17405 4703 17463 4709
rect 18782 4700 18788 4712
rect 18840 4700 18846 4752
rect 22370 4740 22376 4752
rect 22331 4712 22376 4740
rect 22370 4700 22376 4712
rect 22428 4700 22434 4752
rect 27706 4700 27712 4752
rect 27764 4740 27770 4752
rect 28074 4740 28080 4752
rect 27764 4712 28080 4740
rect 27764 4700 27770 4712
rect 28074 4700 28080 4712
rect 28132 4700 28138 4752
rect 28184 4749 28212 4780
rect 28258 4768 28264 4780
rect 28316 4768 28322 4820
rect 29638 4808 29644 4820
rect 29599 4780 29644 4808
rect 29638 4768 29644 4780
rect 29696 4768 29702 4820
rect 29822 4768 29828 4820
rect 29880 4808 29886 4820
rect 30009 4811 30067 4817
rect 30009 4808 30021 4811
rect 29880 4780 30021 4808
rect 29880 4768 29886 4780
rect 30009 4777 30021 4780
rect 30055 4777 30067 4811
rect 32766 4808 32772 4820
rect 32727 4780 32772 4808
rect 30009 4771 30067 4777
rect 32766 4768 32772 4780
rect 32824 4768 32830 4820
rect 32950 4808 32956 4820
rect 32911 4780 32956 4808
rect 32950 4768 32956 4780
rect 33008 4768 33014 4820
rect 33318 4768 33324 4820
rect 33376 4808 33382 4820
rect 33413 4811 33471 4817
rect 33413 4808 33425 4811
rect 33376 4780 33425 4808
rect 33376 4768 33382 4780
rect 33413 4777 33425 4780
rect 33459 4777 33471 4811
rect 33413 4771 33471 4777
rect 34517 4811 34575 4817
rect 34517 4777 34529 4811
rect 34563 4808 34575 4811
rect 34974 4808 34980 4820
rect 34563 4780 34980 4808
rect 34563 4777 34575 4780
rect 34517 4771 34575 4777
rect 34974 4768 34980 4780
rect 35032 4768 35038 4820
rect 35158 4768 35164 4820
rect 35216 4808 35222 4820
rect 35345 4811 35403 4817
rect 35345 4808 35357 4811
rect 35216 4780 35357 4808
rect 35216 4768 35222 4780
rect 35345 4777 35357 4780
rect 35391 4777 35403 4811
rect 35345 4771 35403 4777
rect 35526 4768 35532 4820
rect 35584 4808 35590 4820
rect 35713 4811 35771 4817
rect 35713 4808 35725 4811
rect 35584 4780 35725 4808
rect 35584 4768 35590 4780
rect 35713 4777 35725 4780
rect 35759 4777 35771 4811
rect 35713 4771 35771 4777
rect 28169 4743 28227 4749
rect 28169 4709 28181 4743
rect 28215 4709 28227 4743
rect 28169 4703 28227 4709
rect 29365 4743 29423 4749
rect 29365 4709 29377 4743
rect 29411 4740 29423 4743
rect 29914 4740 29920 4752
rect 29411 4712 29920 4740
rect 29411 4709 29423 4712
rect 29365 4703 29423 4709
rect 29914 4700 29920 4712
rect 29972 4700 29978 4752
rect 32493 4743 32551 4749
rect 32493 4709 32505 4743
rect 32539 4740 32551 4743
rect 32858 4740 32864 4752
rect 32539 4712 32864 4740
rect 32539 4709 32551 4712
rect 32493 4703 32551 4709
rect 32858 4700 32864 4712
rect 32916 4700 32922 4752
rect 34054 4700 34060 4752
rect 34112 4740 34118 4752
rect 34333 4743 34391 4749
rect 34333 4740 34345 4743
rect 34112 4712 34345 4740
rect 34112 4700 34118 4712
rect 34333 4709 34345 4712
rect 34379 4709 34391 4743
rect 34333 4703 34391 4709
rect 34609 4743 34667 4749
rect 34609 4709 34621 4743
rect 34655 4740 34667 4743
rect 34790 4740 34796 4752
rect 34655 4712 34796 4740
rect 34655 4709 34667 4712
rect 34609 4703 34667 4709
rect 34790 4700 34796 4712
rect 34848 4700 34854 4752
rect 1394 4672 1400 4684
rect 1355 4644 1400 4672
rect 1394 4632 1400 4644
rect 1452 4632 1458 4684
rect 2133 4675 2191 4681
rect 2133 4641 2145 4675
rect 2179 4672 2191 4675
rect 2498 4672 2504 4684
rect 2179 4644 2504 4672
rect 2179 4641 2191 4644
rect 2133 4635 2191 4641
rect 2498 4632 2504 4644
rect 2556 4632 2562 4684
rect 5534 4632 5540 4684
rect 5592 4672 5598 4684
rect 8205 4675 8263 4681
rect 8205 4672 8217 4675
rect 5592 4644 8217 4672
rect 5592 4632 5598 4644
rect 8205 4641 8217 4644
rect 8251 4672 8263 4675
rect 8294 4672 8300 4684
rect 8251 4644 8300 4672
rect 8251 4641 8263 4644
rect 8205 4635 8263 4641
rect 8294 4632 8300 4644
rect 8352 4632 8358 4684
rect 13357 4675 13415 4681
rect 13357 4672 13369 4675
rect 12452 4644 13369 4672
rect 12452 4616 12480 4644
rect 13357 4641 13369 4644
rect 13403 4641 13415 4675
rect 15654 4672 15660 4684
rect 15615 4644 15660 4672
rect 13357 4635 13415 4641
rect 15654 4632 15660 4644
rect 15712 4632 15718 4684
rect 15746 4632 15752 4684
rect 15804 4672 15810 4684
rect 15933 4675 15991 4681
rect 15933 4672 15945 4675
rect 15804 4644 15945 4672
rect 15804 4632 15810 4644
rect 15933 4641 15945 4644
rect 15979 4672 15991 4675
rect 16117 4675 16175 4681
rect 16117 4672 16129 4675
rect 15979 4644 16129 4672
rect 15979 4641 15991 4644
rect 15933 4635 15991 4641
rect 16117 4641 16129 4644
rect 16163 4641 16175 4675
rect 17218 4672 17224 4684
rect 17179 4644 17224 4672
rect 16117 4635 16175 4641
rect 17218 4632 17224 4644
rect 17276 4632 17282 4684
rect 27430 4632 27436 4684
rect 27488 4672 27494 4684
rect 27890 4672 27896 4684
rect 27488 4644 27896 4672
rect 27488 4632 27494 4644
rect 27890 4632 27896 4644
rect 27948 4632 27954 4684
rect 34882 4632 34888 4684
rect 34940 4672 34946 4684
rect 34977 4675 35035 4681
rect 34977 4672 34989 4675
rect 34940 4644 34989 4672
rect 34940 4632 34946 4644
rect 34977 4641 34989 4644
rect 35023 4641 35035 4675
rect 34977 4635 35035 4641
rect 35434 4632 35440 4684
rect 35492 4672 35498 4684
rect 35529 4675 35587 4681
rect 35529 4672 35541 4675
rect 35492 4644 35541 4672
rect 35492 4632 35498 4644
rect 35529 4641 35541 4644
rect 35575 4641 35587 4675
rect 35529 4635 35587 4641
rect 7374 4564 7380 4616
rect 7432 4604 7438 4616
rect 8018 4604 8024 4616
rect 7432 4576 8024 4604
rect 7432 4564 7438 4576
rect 8018 4564 8024 4576
rect 8076 4564 8082 4616
rect 10870 4604 10876 4616
rect 10831 4576 10876 4604
rect 10870 4564 10876 4576
rect 10928 4564 10934 4616
rect 11054 4604 11060 4616
rect 11015 4576 11060 4604
rect 11054 4564 11060 4576
rect 11112 4564 11118 4616
rect 12434 4564 12440 4616
rect 12492 4604 12498 4616
rect 12621 4607 12679 4613
rect 12492 4576 12537 4604
rect 12492 4564 12498 4576
rect 12621 4573 12633 4607
rect 12667 4604 12679 4607
rect 12710 4604 12716 4616
rect 12667 4576 12716 4604
rect 12667 4573 12679 4576
rect 12621 4567 12679 4573
rect 12710 4564 12716 4576
rect 12768 4564 12774 4616
rect 12986 4564 12992 4616
rect 13044 4604 13050 4616
rect 14090 4604 14096 4616
rect 13044 4576 14096 4604
rect 13044 4564 13050 4576
rect 14090 4564 14096 4576
rect 14148 4604 14154 4616
rect 14185 4607 14243 4613
rect 14185 4604 14197 4607
rect 14148 4576 14197 4604
rect 14148 4564 14154 4576
rect 14185 4573 14197 4576
rect 14231 4573 14243 4607
rect 17494 4604 17500 4616
rect 17455 4576 17500 4604
rect 14185 4567 14243 4573
rect 17494 4564 17500 4576
rect 17552 4564 17558 4616
rect 19061 4607 19119 4613
rect 19061 4573 19073 4607
rect 19107 4604 19119 4607
rect 19150 4604 19156 4616
rect 19107 4576 19156 4604
rect 19107 4573 19119 4576
rect 19061 4567 19119 4573
rect 19150 4564 19156 4576
rect 19208 4564 19214 4616
rect 22278 4564 22284 4616
rect 22336 4604 22342 4616
rect 22649 4607 22707 4613
rect 22649 4604 22661 4607
rect 22336 4576 22661 4604
rect 22336 4564 22342 4576
rect 22649 4573 22661 4576
rect 22695 4604 22707 4607
rect 22830 4604 22836 4616
rect 22695 4576 22836 4604
rect 22695 4573 22707 4576
rect 22649 4567 22707 4573
rect 22830 4564 22836 4576
rect 22888 4564 22894 4616
rect 7466 4496 7472 4548
rect 7524 4536 7530 4548
rect 7653 4539 7711 4545
rect 7653 4536 7665 4539
rect 7524 4508 7665 4536
rect 7524 4496 7530 4508
rect 7653 4505 7665 4508
rect 7699 4505 7711 4539
rect 7653 4499 7711 4505
rect 10505 4539 10563 4545
rect 10505 4505 10517 4539
rect 10551 4536 10563 4539
rect 10686 4536 10692 4548
rect 10551 4508 10692 4536
rect 10551 4505 10563 4508
rect 10505 4499 10563 4505
rect 10686 4496 10692 4508
rect 10744 4496 10750 4548
rect 16482 4496 16488 4548
rect 16540 4536 16546 4548
rect 16761 4539 16819 4545
rect 16761 4536 16773 4539
rect 16540 4508 16773 4536
rect 16540 4496 16546 4508
rect 16761 4505 16773 4508
rect 16807 4536 16819 4539
rect 18509 4539 18567 4545
rect 18509 4536 18521 4539
rect 16807 4508 18521 4536
rect 16807 4505 16819 4508
rect 16761 4499 16819 4505
rect 18509 4505 18521 4508
rect 18555 4505 18567 4539
rect 18509 4499 18567 4505
rect 27522 4496 27528 4548
rect 27580 4536 27586 4548
rect 27617 4539 27675 4545
rect 27617 4536 27629 4539
rect 27580 4508 27629 4536
rect 27580 4496 27586 4508
rect 27617 4505 27629 4508
rect 27663 4505 27675 4539
rect 27617 4499 27675 4505
rect 33410 4496 33416 4548
rect 33468 4536 33474 4548
rect 34057 4539 34115 4545
rect 34057 4536 34069 4539
rect 33468 4508 34069 4536
rect 33468 4496 33474 4508
rect 34057 4505 34069 4508
rect 34103 4505 34115 4539
rect 34057 4499 34115 4505
rect 12066 4468 12072 4480
rect 12027 4440 12072 4468
rect 12066 4428 12072 4440
rect 12124 4428 12130 4480
rect 15102 4428 15108 4480
rect 15160 4468 15166 4480
rect 15381 4471 15439 4477
rect 15381 4468 15393 4471
rect 15160 4440 15393 4468
rect 15160 4428 15166 4440
rect 15381 4437 15393 4440
rect 15427 4437 15439 4471
rect 15381 4431 15439 4437
rect 22097 4471 22155 4477
rect 22097 4437 22109 4471
rect 22143 4468 22155 4471
rect 22646 4468 22652 4480
rect 22143 4440 22652 4468
rect 22143 4437 22155 4440
rect 22097 4431 22155 4437
rect 22646 4428 22652 4440
rect 22704 4428 22710 4480
rect 1104 4378 38824 4400
rect 1104 4326 7648 4378
rect 7700 4326 7712 4378
rect 7764 4326 7776 4378
rect 7828 4326 7840 4378
rect 7892 4326 20982 4378
rect 21034 4326 21046 4378
rect 21098 4326 21110 4378
rect 21162 4326 21174 4378
rect 21226 4326 34315 4378
rect 34367 4326 34379 4378
rect 34431 4326 34443 4378
rect 34495 4326 34507 4378
rect 34559 4326 38824 4378
rect 1104 4304 38824 4326
rect 1394 4224 1400 4276
rect 1452 4264 1458 4276
rect 2314 4264 2320 4276
rect 1452 4236 2320 4264
rect 1452 4224 1458 4236
rect 2314 4224 2320 4236
rect 2372 4224 2378 4276
rect 2498 4224 2504 4276
rect 2556 4264 2562 4276
rect 2961 4267 3019 4273
rect 2961 4264 2973 4267
rect 2556 4236 2973 4264
rect 2556 4224 2562 4236
rect 2961 4233 2973 4236
rect 3007 4233 3019 4267
rect 2961 4227 3019 4233
rect 8021 4267 8079 4273
rect 8021 4233 8033 4267
rect 8067 4264 8079 4267
rect 8110 4264 8116 4276
rect 8067 4236 8116 4264
rect 8067 4233 8079 4236
rect 8021 4227 8079 4233
rect 8110 4224 8116 4236
rect 8168 4224 8174 4276
rect 9766 4224 9772 4276
rect 9824 4264 9830 4276
rect 11793 4267 11851 4273
rect 11793 4264 11805 4267
rect 9824 4236 11805 4264
rect 9824 4224 9830 4236
rect 11793 4233 11805 4236
rect 11839 4264 11851 4267
rect 12250 4264 12256 4276
rect 11839 4236 12256 4264
rect 11839 4233 11851 4236
rect 11793 4227 11851 4233
rect 12250 4224 12256 4236
rect 12308 4224 12314 4276
rect 12526 4264 12532 4276
rect 12487 4236 12532 4264
rect 12526 4224 12532 4236
rect 12584 4224 12590 4276
rect 13906 4224 13912 4276
rect 13964 4264 13970 4276
rect 14093 4267 14151 4273
rect 14093 4264 14105 4267
rect 13964 4236 14105 4264
rect 13964 4224 13970 4236
rect 14093 4233 14105 4236
rect 14139 4233 14151 4267
rect 16114 4264 16120 4276
rect 16075 4236 16120 4264
rect 14093 4227 14151 4233
rect 16114 4224 16120 4236
rect 16172 4224 16178 4276
rect 17310 4264 17316 4276
rect 17271 4236 17316 4264
rect 17310 4224 17316 4236
rect 17368 4224 17374 4276
rect 17494 4224 17500 4276
rect 17552 4264 17558 4276
rect 17681 4267 17739 4273
rect 17681 4264 17693 4267
rect 17552 4236 17693 4264
rect 17552 4224 17558 4236
rect 17681 4233 17693 4236
rect 17727 4264 17739 4267
rect 19150 4264 19156 4276
rect 17727 4236 19156 4264
rect 17727 4233 17739 4236
rect 17681 4227 17739 4233
rect 19150 4224 19156 4236
rect 19208 4224 19214 4276
rect 22094 4224 22100 4276
rect 22152 4264 22158 4276
rect 22373 4267 22431 4273
rect 22373 4264 22385 4267
rect 22152 4236 22385 4264
rect 22152 4224 22158 4236
rect 22373 4233 22385 4236
rect 22419 4233 22431 4267
rect 27706 4264 27712 4276
rect 27667 4236 27712 4264
rect 22373 4227 22431 4233
rect 27706 4224 27712 4236
rect 27764 4224 27770 4276
rect 27890 4224 27896 4276
rect 27948 4264 27954 4276
rect 27985 4267 28043 4273
rect 27985 4264 27997 4267
rect 27948 4236 27997 4264
rect 27948 4224 27954 4236
rect 27985 4233 27997 4236
rect 28031 4233 28043 4267
rect 27985 4227 28043 4233
rect 28258 4224 28264 4276
rect 28316 4264 28322 4276
rect 28353 4267 28411 4273
rect 28353 4264 28365 4267
rect 28316 4236 28365 4264
rect 28316 4224 28322 4236
rect 28353 4233 28365 4236
rect 28399 4233 28411 4267
rect 28353 4227 28411 4233
rect 33689 4267 33747 4273
rect 33689 4233 33701 4267
rect 33735 4264 33747 4267
rect 34054 4264 34060 4276
rect 33735 4236 34060 4264
rect 33735 4233 33747 4236
rect 33689 4227 33747 4233
rect 34054 4224 34060 4236
rect 34112 4224 34118 4276
rect 34425 4267 34483 4273
rect 34425 4233 34437 4267
rect 34471 4264 34483 4267
rect 34974 4264 34980 4276
rect 34471 4236 34980 4264
rect 34471 4233 34483 4236
rect 34425 4227 34483 4233
rect 34974 4224 34980 4236
rect 35032 4224 35038 4276
rect 10870 4196 10876 4208
rect 10783 4168 10876 4196
rect 10870 4156 10876 4168
rect 10928 4156 10934 4208
rect 13814 4156 13820 4208
rect 13872 4156 13878 4208
rect 15746 4196 15752 4208
rect 15707 4168 15752 4196
rect 15746 4156 15752 4168
rect 15804 4156 15810 4208
rect 18509 4199 18567 4205
rect 18509 4165 18521 4199
rect 18555 4196 18567 4199
rect 18966 4196 18972 4208
rect 18555 4168 18972 4196
rect 18555 4165 18567 4168
rect 18509 4159 18567 4165
rect 18966 4156 18972 4168
rect 19024 4156 19030 4208
rect 34790 4196 34796 4208
rect 34440 4168 34796 4196
rect 8294 4128 8300 4140
rect 8255 4100 8300 4128
rect 8294 4088 8300 4100
rect 8352 4088 8358 4140
rect 9585 4131 9643 4137
rect 9585 4097 9597 4131
rect 9631 4128 9643 4131
rect 10888 4128 10916 4156
rect 9631 4100 10916 4128
rect 9631 4097 9643 4100
rect 9585 4091 9643 4097
rect 12986 4088 12992 4140
rect 13044 4128 13050 4140
rect 13081 4131 13139 4137
rect 13081 4128 13093 4131
rect 13044 4100 13093 4128
rect 13044 4088 13050 4100
rect 13081 4097 13093 4100
rect 13127 4097 13139 4131
rect 13081 4091 13139 4097
rect 13633 4131 13691 4137
rect 13633 4097 13645 4131
rect 13679 4128 13691 4131
rect 13832 4128 13860 4156
rect 13679 4100 13860 4128
rect 13679 4097 13691 4100
rect 13633 4091 13691 4097
rect 14182 4088 14188 4140
rect 14240 4128 14246 4140
rect 14553 4131 14611 4137
rect 14553 4128 14565 4131
rect 14240 4100 14565 4128
rect 14240 4088 14246 4100
rect 14553 4097 14565 4100
rect 14599 4128 14611 4131
rect 15102 4128 15108 4140
rect 14599 4100 15108 4128
rect 14599 4097 14611 4100
rect 14553 4091 14611 4097
rect 15102 4088 15108 4100
rect 15160 4088 15166 4140
rect 18782 4128 18788 4140
rect 18743 4100 18788 4128
rect 18782 4088 18788 4100
rect 18840 4088 18846 4140
rect 22097 4131 22155 4137
rect 22097 4097 22109 4131
rect 22143 4128 22155 4131
rect 22278 4128 22284 4140
rect 22143 4100 22284 4128
rect 22143 4097 22155 4100
rect 22097 4091 22155 4097
rect 22278 4088 22284 4100
rect 22336 4088 22342 4140
rect 22370 4088 22376 4140
rect 22428 4128 22434 4140
rect 22741 4131 22799 4137
rect 22741 4128 22753 4131
rect 22428 4100 22753 4128
rect 22428 4088 22434 4100
rect 22741 4097 22753 4100
rect 22787 4097 22799 4131
rect 22741 4091 22799 4097
rect 26145 4131 26203 4137
rect 26145 4097 26157 4131
rect 26191 4128 26203 4131
rect 27157 4131 27215 4137
rect 27157 4128 27169 4131
rect 26191 4100 27169 4128
rect 26191 4097 26203 4100
rect 26145 4091 26203 4097
rect 27157 4097 27169 4100
rect 27203 4128 27215 4131
rect 27982 4128 27988 4140
rect 27203 4100 27988 4128
rect 27203 4097 27215 4100
rect 27157 4091 27215 4097
rect 27982 4088 27988 4100
rect 28040 4088 28046 4140
rect 34057 4131 34115 4137
rect 34057 4097 34069 4131
rect 34103 4128 34115 4131
rect 34440 4128 34468 4168
rect 34790 4156 34796 4168
rect 34848 4156 34854 4208
rect 35434 4156 35440 4208
rect 35492 4196 35498 4208
rect 35492 4168 35848 4196
rect 35492 4156 35498 4168
rect 34103 4100 34468 4128
rect 35820 4128 35848 4168
rect 36357 4131 36415 4137
rect 36357 4128 36369 4131
rect 35820 4100 36369 4128
rect 34103 4097 34115 4100
rect 34057 4091 34115 4097
rect 36357 4097 36369 4100
rect 36403 4097 36415 4131
rect 36357 4091 36415 4097
rect 1397 4063 1455 4069
rect 1397 4029 1409 4063
rect 1443 4060 1455 4063
rect 2501 4063 2559 4069
rect 1443 4032 2084 4060
rect 1443 4029 1455 4032
rect 1397 4023 1455 4029
rect 2056 4004 2084 4032
rect 2501 4029 2513 4063
rect 2547 4060 2559 4063
rect 2682 4060 2688 4072
rect 2547 4032 2688 4060
rect 2547 4029 2559 4032
rect 2501 4023 2559 4029
rect 2682 4020 2688 4032
rect 2740 4020 2746 4072
rect 10778 4020 10784 4072
rect 10836 4060 10842 4072
rect 11149 4063 11207 4069
rect 11149 4060 11161 4063
rect 10836 4032 11161 4060
rect 10836 4020 10842 4032
rect 11149 4029 11161 4032
rect 11195 4029 11207 4063
rect 11422 4060 11428 4072
rect 11383 4032 11428 4060
rect 11149 4023 11207 4029
rect 11422 4020 11428 4032
rect 11480 4020 11486 4072
rect 12342 4020 12348 4072
rect 12400 4060 12406 4072
rect 16853 4063 16911 4069
rect 16853 4060 16865 4063
rect 12400 4032 16865 4060
rect 12400 4020 12406 4032
rect 16853 4029 16865 4032
rect 16899 4060 16911 4063
rect 17126 4060 17132 4072
rect 16899 4032 17132 4060
rect 16899 4029 16911 4032
rect 16853 4023 16911 4029
rect 17126 4020 17132 4032
rect 17184 4020 17190 4072
rect 26679 4063 26737 4069
rect 26679 4029 26691 4063
rect 26725 4060 26737 4063
rect 27522 4060 27528 4072
rect 26725 4032 27528 4060
rect 26725 4029 26737 4032
rect 26679 4023 26737 4029
rect 27522 4020 27528 4032
rect 27580 4020 27586 4072
rect 35434 4060 35440 4072
rect 35395 4032 35440 4060
rect 35434 4020 35440 4032
rect 35492 4060 35498 4072
rect 35989 4063 36047 4069
rect 35989 4060 36001 4063
rect 35492 4032 36001 4060
rect 35492 4020 35498 4032
rect 35989 4029 36001 4032
rect 36035 4029 36047 4063
rect 35989 4023 36047 4029
rect 2038 3992 2044 4004
rect 1999 3964 2044 3992
rect 2038 3952 2044 3964
rect 2096 3952 2102 4004
rect 9953 3995 10011 4001
rect 9953 3961 9965 3995
rect 9999 3992 10011 3995
rect 10962 3992 10968 4004
rect 9999 3964 10968 3992
rect 9999 3961 10011 3964
rect 9953 3955 10011 3961
rect 10962 3952 10968 3964
rect 11020 3952 11026 4004
rect 12526 3952 12532 4004
rect 12584 3992 12590 4004
rect 12805 3995 12863 4001
rect 12805 3992 12817 3995
rect 12584 3964 12817 3992
rect 12584 3952 12590 3964
rect 12805 3961 12817 3964
rect 12851 3961 12863 3995
rect 14550 3992 14556 4004
rect 14511 3964 14556 3992
rect 12805 3955 12863 3961
rect 14550 3952 14556 3964
rect 14608 3952 14614 4004
rect 14642 3952 14648 4004
rect 14700 3992 14706 4004
rect 27246 3992 27252 4004
rect 14700 3964 14745 3992
rect 27207 3964 27252 3992
rect 14700 3952 14706 3964
rect 27246 3952 27252 3964
rect 27304 3952 27310 4004
rect 1578 3924 1584 3936
rect 1539 3896 1584 3924
rect 1578 3884 1584 3896
rect 1636 3884 1642 3936
rect 7466 3884 7472 3936
rect 7524 3924 7530 3936
rect 7561 3927 7619 3933
rect 7561 3924 7573 3927
rect 7524 3896 7573 3924
rect 7524 3884 7530 3896
rect 7561 3893 7573 3896
rect 7607 3893 7619 3927
rect 10318 3924 10324 3936
rect 10279 3896 10324 3924
rect 7561 3887 7619 3893
rect 10318 3884 10324 3896
rect 10376 3884 10382 3936
rect 10594 3924 10600 3936
rect 10555 3896 10600 3924
rect 10594 3884 10600 3896
rect 10652 3924 10658 3936
rect 11333 3927 11391 3933
rect 11333 3924 11345 3927
rect 10652 3896 11345 3924
rect 10652 3884 10658 3896
rect 11333 3893 11345 3896
rect 11379 3893 11391 3927
rect 12158 3924 12164 3936
rect 12119 3896 12164 3924
rect 11333 3887 11391 3893
rect 12158 3884 12164 3896
rect 12216 3924 12222 3936
rect 12986 3924 12992 3936
rect 12216 3896 12992 3924
rect 12216 3884 12222 3896
rect 12986 3884 12992 3896
rect 13044 3884 13050 3936
rect 13170 3884 13176 3936
rect 13228 3924 13234 3936
rect 15289 3927 15347 3933
rect 15289 3924 15301 3927
rect 13228 3896 15301 3924
rect 13228 3884 13234 3896
rect 15289 3893 15301 3896
rect 15335 3924 15347 3927
rect 15654 3924 15660 3936
rect 15335 3896 15660 3924
rect 15335 3893 15347 3896
rect 15289 3887 15347 3893
rect 15654 3884 15660 3896
rect 15712 3884 15718 3936
rect 26513 3927 26571 3933
rect 26513 3893 26525 3927
rect 26559 3924 26571 3927
rect 27157 3927 27215 3933
rect 27157 3924 27169 3927
rect 26559 3896 27169 3924
rect 26559 3893 26571 3896
rect 26513 3887 26571 3893
rect 27157 3893 27169 3896
rect 27203 3924 27215 3927
rect 27338 3924 27344 3936
rect 27203 3896 27344 3924
rect 27203 3893 27215 3896
rect 27157 3887 27215 3893
rect 27338 3884 27344 3896
rect 27396 3884 27402 3936
rect 35342 3884 35348 3936
rect 35400 3924 35406 3936
rect 35621 3927 35679 3933
rect 35621 3924 35633 3927
rect 35400 3896 35633 3924
rect 35400 3884 35406 3896
rect 35621 3893 35633 3896
rect 35667 3893 35679 3927
rect 35621 3887 35679 3893
rect 1104 3834 38824 3856
rect 1104 3782 14315 3834
rect 14367 3782 14379 3834
rect 14431 3782 14443 3834
rect 14495 3782 14507 3834
rect 14559 3782 27648 3834
rect 27700 3782 27712 3834
rect 27764 3782 27776 3834
rect 27828 3782 27840 3834
rect 27892 3782 38824 3834
rect 1104 3760 38824 3782
rect 1581 3723 1639 3729
rect 1581 3689 1593 3723
rect 1627 3720 1639 3723
rect 3050 3720 3056 3732
rect 1627 3692 3056 3720
rect 1627 3689 1639 3692
rect 1581 3683 1639 3689
rect 3050 3680 3056 3692
rect 3108 3680 3114 3732
rect 9582 3680 9588 3732
rect 9640 3680 9646 3732
rect 10778 3720 10784 3732
rect 10739 3692 10784 3720
rect 10778 3680 10784 3692
rect 10836 3680 10842 3732
rect 13357 3723 13415 3729
rect 13357 3689 13369 3723
rect 13403 3720 13415 3723
rect 13722 3720 13728 3732
rect 13403 3692 13728 3720
rect 13403 3689 13415 3692
rect 13357 3683 13415 3689
rect 13722 3680 13728 3692
rect 13780 3680 13786 3732
rect 13909 3723 13967 3729
rect 13909 3689 13921 3723
rect 13955 3720 13967 3723
rect 13998 3720 14004 3732
rect 13955 3692 14004 3720
rect 13955 3689 13967 3692
rect 13909 3683 13967 3689
rect 13998 3680 14004 3692
rect 14056 3680 14062 3732
rect 14090 3680 14096 3732
rect 14148 3720 14154 3732
rect 14185 3723 14243 3729
rect 14185 3720 14197 3723
rect 14148 3692 14197 3720
rect 14148 3680 14154 3692
rect 14185 3689 14197 3692
rect 14231 3689 14243 3723
rect 14642 3720 14648 3732
rect 14603 3692 14648 3720
rect 14185 3683 14243 3689
rect 14642 3680 14648 3692
rect 14700 3680 14706 3732
rect 15562 3720 15568 3732
rect 15523 3692 15568 3720
rect 15562 3680 15568 3692
rect 15620 3680 15626 3732
rect 26789 3723 26847 3729
rect 26789 3689 26801 3723
rect 26835 3720 26847 3723
rect 27246 3720 27252 3732
rect 26835 3692 27252 3720
rect 26835 3689 26847 3692
rect 26789 3683 26847 3689
rect 27246 3680 27252 3692
rect 27304 3680 27310 3732
rect 566 3612 572 3664
rect 624 3652 630 3664
rect 9600 3652 9628 3680
rect 624 3624 9628 3652
rect 10505 3655 10563 3661
rect 624 3612 630 3624
rect 10505 3621 10517 3655
rect 10551 3652 10563 3655
rect 11054 3652 11060 3664
rect 10551 3624 11060 3652
rect 10551 3621 10563 3624
rect 10505 3615 10563 3621
rect 11054 3612 11060 3624
rect 11112 3612 11118 3664
rect 11146 3612 11152 3664
rect 11204 3652 11210 3664
rect 11609 3655 11667 3661
rect 11609 3652 11621 3655
rect 11204 3624 11621 3652
rect 11204 3612 11210 3624
rect 11609 3621 11621 3624
rect 11655 3621 11667 3655
rect 11609 3615 11667 3621
rect 11698 3612 11704 3664
rect 11756 3652 11762 3664
rect 11793 3655 11851 3661
rect 11793 3652 11805 3655
rect 11756 3624 11805 3652
rect 11756 3612 11762 3624
rect 11793 3621 11805 3624
rect 11839 3621 11851 3655
rect 11793 3615 11851 3621
rect 1394 3584 1400 3596
rect 1355 3556 1400 3584
rect 1394 3544 1400 3556
rect 1452 3544 1458 3596
rect 11422 3544 11428 3596
rect 11480 3584 11486 3596
rect 11885 3587 11943 3593
rect 11885 3584 11897 3587
rect 11480 3556 11897 3584
rect 11480 3544 11486 3556
rect 11885 3553 11897 3556
rect 11931 3553 11943 3587
rect 11885 3547 11943 3553
rect 9674 3476 9680 3528
rect 9732 3516 9738 3528
rect 13170 3516 13176 3528
rect 9732 3488 13176 3516
rect 9732 3476 9738 3488
rect 13170 3476 13176 3488
rect 13228 3476 13234 3528
rect 13354 3516 13360 3528
rect 13315 3488 13360 3516
rect 13354 3476 13360 3488
rect 13412 3476 13418 3528
rect 13446 3476 13452 3528
rect 13504 3516 13510 3528
rect 13504 3488 13549 3516
rect 13504 3476 13510 3488
rect 10962 3408 10968 3460
rect 11020 3448 11026 3460
rect 11333 3451 11391 3457
rect 11333 3448 11345 3451
rect 11020 3420 11345 3448
rect 11020 3408 11026 3420
rect 11333 3417 11345 3420
rect 11379 3417 11391 3451
rect 12894 3448 12900 3460
rect 12855 3420 12900 3448
rect 11333 3411 11391 3417
rect 12894 3408 12900 3420
rect 12952 3408 12958 3460
rect 12526 3380 12532 3392
rect 12487 3352 12532 3380
rect 12526 3340 12532 3352
rect 12584 3340 12590 3392
rect 1104 3290 38824 3312
rect 1104 3238 7648 3290
rect 7700 3238 7712 3290
rect 7764 3238 7776 3290
rect 7828 3238 7840 3290
rect 7892 3238 20982 3290
rect 21034 3238 21046 3290
rect 21098 3238 21110 3290
rect 21162 3238 21174 3290
rect 21226 3238 34315 3290
rect 34367 3238 34379 3290
rect 34431 3238 34443 3290
rect 34495 3238 34507 3290
rect 34559 3238 38824 3290
rect 1104 3216 38824 3238
rect 1394 3136 1400 3188
rect 1452 3176 1458 3188
rect 1581 3179 1639 3185
rect 1581 3176 1593 3179
rect 1452 3148 1593 3176
rect 1452 3136 1458 3148
rect 1581 3145 1593 3148
rect 1627 3145 1639 3179
rect 1581 3139 1639 3145
rect 10318 3136 10324 3188
rect 10376 3176 10382 3188
rect 10965 3179 11023 3185
rect 10965 3176 10977 3179
rect 10376 3148 10977 3176
rect 10376 3136 10382 3148
rect 10965 3145 10977 3148
rect 11011 3176 11023 3179
rect 11422 3176 11428 3188
rect 11011 3148 11428 3176
rect 11011 3145 11023 3148
rect 10965 3139 11023 3145
rect 11422 3136 11428 3148
rect 11480 3136 11486 3188
rect 11606 3176 11612 3188
rect 11567 3148 11612 3176
rect 11606 3136 11612 3148
rect 11664 3136 11670 3188
rect 13446 3176 13452 3188
rect 13407 3148 13452 3176
rect 13446 3136 13452 3148
rect 13504 3136 13510 3188
rect 13722 3136 13728 3188
rect 13780 3176 13786 3188
rect 13817 3179 13875 3185
rect 13817 3176 13829 3179
rect 13780 3148 13829 3176
rect 13780 3136 13786 3148
rect 13817 3145 13829 3148
rect 13863 3145 13875 3179
rect 14182 3176 14188 3188
rect 14143 3148 14188 3176
rect 13817 3139 13875 3145
rect 14182 3136 14188 3148
rect 14240 3136 14246 3188
rect 11146 3068 11152 3120
rect 11204 3108 11210 3120
rect 11241 3111 11299 3117
rect 11241 3108 11253 3111
rect 11204 3080 11253 3108
rect 11204 3068 11210 3080
rect 11241 3077 11253 3080
rect 11287 3077 11299 3111
rect 11241 3071 11299 3077
rect 12529 3111 12587 3117
rect 12529 3077 12541 3111
rect 12575 3108 12587 3111
rect 13354 3108 13360 3120
rect 12575 3080 13360 3108
rect 12575 3077 12587 3080
rect 12529 3071 12587 3077
rect 13354 3068 13360 3080
rect 13412 3068 13418 3120
rect 12253 3043 12311 3049
rect 12253 3009 12265 3043
rect 12299 3040 12311 3043
rect 13081 3043 13139 3049
rect 13081 3040 13093 3043
rect 12299 3012 13093 3040
rect 12299 3009 12311 3012
rect 12253 3003 12311 3009
rect 13081 3009 13093 3012
rect 13127 3040 13139 3043
rect 13538 3040 13544 3052
rect 13127 3012 13544 3040
rect 13127 3009 13139 3012
rect 13081 3003 13139 3009
rect 13538 3000 13544 3012
rect 13596 3000 13602 3052
rect 12802 2972 12808 2984
rect 12763 2944 12808 2972
rect 12802 2932 12808 2944
rect 12860 2932 12866 2984
rect 13630 2972 13636 2984
rect 13004 2944 13636 2972
rect 12894 2864 12900 2916
rect 12952 2904 12958 2916
rect 13004 2913 13032 2944
rect 13630 2932 13636 2944
rect 13688 2932 13694 2984
rect 12989 2907 13047 2913
rect 12989 2904 13001 2907
rect 12952 2876 13001 2904
rect 12952 2864 12958 2876
rect 12989 2873 13001 2876
rect 13035 2873 13047 2907
rect 12989 2867 13047 2873
rect 1104 2746 38824 2768
rect 1104 2694 14315 2746
rect 14367 2694 14379 2746
rect 14431 2694 14443 2746
rect 14495 2694 14507 2746
rect 14559 2694 27648 2746
rect 27700 2694 27712 2746
rect 27764 2694 27776 2746
rect 27828 2694 27840 2746
rect 27892 2694 38824 2746
rect 1104 2672 38824 2694
rect 12894 2632 12900 2644
rect 12855 2604 12900 2632
rect 12894 2592 12900 2604
rect 12952 2592 12958 2644
rect 13354 2592 13360 2644
rect 13412 2632 13418 2644
rect 13541 2635 13599 2641
rect 13541 2632 13553 2635
rect 13412 2604 13553 2632
rect 13412 2592 13418 2604
rect 13541 2601 13553 2604
rect 13587 2601 13599 2635
rect 13541 2595 13599 2601
rect 12802 2524 12808 2576
rect 12860 2564 12866 2576
rect 13173 2567 13231 2573
rect 13173 2564 13185 2567
rect 12860 2536 13185 2564
rect 12860 2524 12866 2536
rect 13173 2533 13185 2536
rect 13219 2533 13231 2567
rect 13173 2527 13231 2533
rect 1104 2202 38824 2224
rect 1104 2150 7648 2202
rect 7700 2150 7712 2202
rect 7764 2150 7776 2202
rect 7828 2150 7840 2202
rect 7892 2150 20982 2202
rect 21034 2150 21046 2202
rect 21098 2150 21110 2202
rect 21162 2150 21174 2202
rect 21226 2150 34315 2202
rect 34367 2150 34379 2202
rect 34431 2150 34443 2202
rect 34495 2150 34507 2202
rect 34559 2150 38824 2202
rect 1104 2128 38824 2150
<< via1 >>
rect 3608 14084 3660 14136
rect 7472 14084 7524 14136
rect 3424 14016 3476 14068
rect 6920 14016 6972 14068
rect 3516 13948 3568 14000
rect 8392 13948 8444 14000
rect 3148 13880 3200 13932
rect 7104 13880 7156 13932
rect 33140 13880 33192 13932
rect 34796 13880 34848 13932
rect 3240 13812 3292 13864
rect 9864 13812 9916 13864
rect 9956 13812 10008 13864
rect 34520 13812 34572 13864
rect 31208 13676 31260 13728
rect 36176 13676 36228 13728
rect 14315 13574 14367 13626
rect 14379 13574 14431 13626
rect 14443 13574 14495 13626
rect 14507 13574 14559 13626
rect 27648 13574 27700 13626
rect 27712 13574 27764 13626
rect 27776 13574 27828 13626
rect 27840 13574 27892 13626
rect 2780 13472 2832 13524
rect 7104 13515 7156 13524
rect 7104 13481 7113 13515
rect 7113 13481 7147 13515
rect 7147 13481 7156 13515
rect 7104 13472 7156 13481
rect 34612 13472 34664 13524
rect 5816 13404 5868 13456
rect 17224 13404 17276 13456
rect 1584 13336 1636 13388
rect 2320 13336 2372 13388
rect 4160 13336 4212 13388
rect 5172 13379 5224 13388
rect 5172 13345 5181 13379
rect 5181 13345 5215 13379
rect 5215 13345 5224 13379
rect 5172 13336 5224 13345
rect 7104 13336 7156 13388
rect 23388 13336 23440 13388
rect 26976 13336 27028 13388
rect 33416 13336 33468 13388
rect 34152 13336 34204 13388
rect 35256 13336 35308 13388
rect 6092 13268 6144 13320
rect 32312 13268 32364 13320
rect 34796 13268 34848 13320
rect 37096 13268 37148 13320
rect 4528 13200 4580 13252
rect 11704 13200 11756 13252
rect 34704 13200 34756 13252
rect 2780 13132 2832 13184
rect 3516 13132 3568 13184
rect 24860 13175 24912 13184
rect 24860 13141 24869 13175
rect 24869 13141 24903 13175
rect 24903 13141 24912 13175
rect 24860 13132 24912 13141
rect 33968 13132 34020 13184
rect 34888 13175 34940 13184
rect 34888 13141 34897 13175
rect 34897 13141 34931 13175
rect 34931 13141 34940 13175
rect 34888 13132 34940 13141
rect 35440 13132 35492 13184
rect 35808 13132 35860 13184
rect 7648 13030 7700 13082
rect 7712 13030 7764 13082
rect 7776 13030 7828 13082
rect 7840 13030 7892 13082
rect 20982 13030 21034 13082
rect 21046 13030 21098 13082
rect 21110 13030 21162 13082
rect 21174 13030 21226 13082
rect 34315 13030 34367 13082
rect 34379 13030 34431 13082
rect 34443 13030 34495 13082
rect 34507 13030 34559 13082
rect 1584 12971 1636 12980
rect 1584 12937 1593 12971
rect 1593 12937 1627 12971
rect 1627 12937 1636 12971
rect 1584 12928 1636 12937
rect 4068 12928 4120 12980
rect 6644 12928 6696 12980
rect 7472 12928 7524 12980
rect 2964 12860 3016 12912
rect 3332 12792 3384 12844
rect 3424 12792 3476 12844
rect 7012 12792 7064 12844
rect 8116 12860 8168 12912
rect 25504 12928 25556 12980
rect 31116 12928 31168 12980
rect 34612 12928 34664 12980
rect 36452 12928 36504 12980
rect 37096 12971 37148 12980
rect 37096 12937 37105 12971
rect 37105 12937 37139 12971
rect 37139 12937 37148 12971
rect 37096 12928 37148 12937
rect 11704 12860 11756 12912
rect 19984 12860 20036 12912
rect 22928 12860 22980 12912
rect 25228 12860 25280 12912
rect 2044 12724 2096 12776
rect 4160 12724 4212 12776
rect 4620 12724 4672 12776
rect 7196 12724 7248 12776
rect 4068 12656 4120 12708
rect 4528 12699 4580 12708
rect 4528 12665 4537 12699
rect 4537 12665 4571 12699
rect 4571 12665 4580 12699
rect 4528 12656 4580 12665
rect 4804 12699 4856 12708
rect 4804 12665 4813 12699
rect 4813 12665 4847 12699
rect 4847 12665 4856 12699
rect 4804 12656 4856 12665
rect 5172 12656 5224 12708
rect 15200 12792 15252 12844
rect 17592 12792 17644 12844
rect 19892 12792 19944 12844
rect 22284 12792 22336 12844
rect 24860 12792 24912 12844
rect 26516 12792 26568 12844
rect 29368 12792 29420 12844
rect 31668 12792 31720 12844
rect 4712 12631 4764 12640
rect 4712 12597 4721 12631
rect 4721 12597 4755 12631
rect 4755 12597 4764 12631
rect 4712 12588 4764 12597
rect 5356 12588 5408 12640
rect 5724 12631 5776 12640
rect 5724 12597 5733 12631
rect 5733 12597 5767 12631
rect 5767 12597 5776 12631
rect 5724 12588 5776 12597
rect 7104 12588 7156 12640
rect 10508 12656 10560 12708
rect 12532 12724 12584 12776
rect 16856 12724 16908 12776
rect 19340 12724 19392 12776
rect 23480 12724 23532 12776
rect 33140 12860 33192 12912
rect 33508 12860 33560 12912
rect 34796 12860 34848 12912
rect 33784 12835 33836 12844
rect 33784 12801 33793 12835
rect 33793 12801 33827 12835
rect 33827 12801 33836 12835
rect 33784 12792 33836 12801
rect 36360 12792 36412 12844
rect 34888 12767 34940 12776
rect 12900 12656 12952 12708
rect 24768 12656 24820 12708
rect 34888 12733 34897 12767
rect 34897 12733 34931 12767
rect 34931 12733 34940 12767
rect 34888 12724 34940 12733
rect 36176 12767 36228 12776
rect 36176 12733 36185 12767
rect 36185 12733 36219 12767
rect 36219 12733 36228 12767
rect 36176 12724 36228 12733
rect 37280 12767 37332 12776
rect 37280 12733 37289 12767
rect 37289 12733 37323 12767
rect 37323 12733 37332 12767
rect 37280 12724 37332 12733
rect 32036 12656 32088 12708
rect 16212 12588 16264 12640
rect 22652 12588 22704 12640
rect 23388 12588 23440 12640
rect 25136 12588 25188 12640
rect 33508 12656 33560 12708
rect 36268 12656 36320 12708
rect 38752 12656 38804 12708
rect 33968 12588 34020 12640
rect 34336 12631 34388 12640
rect 34336 12597 34345 12631
rect 34345 12597 34379 12631
rect 34379 12597 34388 12631
rect 34336 12588 34388 12597
rect 35256 12588 35308 12640
rect 37464 12631 37516 12640
rect 37464 12597 37473 12631
rect 37473 12597 37507 12631
rect 37507 12597 37516 12631
rect 37464 12588 37516 12597
rect 14315 12486 14367 12538
rect 14379 12486 14431 12538
rect 14443 12486 14495 12538
rect 14507 12486 14559 12538
rect 27648 12486 27700 12538
rect 27712 12486 27764 12538
rect 27776 12486 27828 12538
rect 27840 12486 27892 12538
rect 4160 12384 4212 12436
rect 4712 12384 4764 12436
rect 6644 12427 6696 12436
rect 6644 12393 6653 12427
rect 6653 12393 6687 12427
rect 6687 12393 6696 12427
rect 6644 12384 6696 12393
rect 31116 12427 31168 12436
rect 31116 12393 31125 12427
rect 31125 12393 31159 12427
rect 31159 12393 31168 12427
rect 31116 12384 31168 12393
rect 32312 12427 32364 12436
rect 32312 12393 32321 12427
rect 32321 12393 32355 12427
rect 32355 12393 32364 12427
rect 32312 12384 32364 12393
rect 36268 12384 36320 12436
rect 1124 12316 1176 12368
rect 5264 12316 5316 12368
rect 2504 12291 2556 12300
rect 2504 12257 2513 12291
rect 2513 12257 2547 12291
rect 2547 12257 2556 12291
rect 2504 12248 2556 12257
rect 2688 12291 2740 12300
rect 2688 12257 2697 12291
rect 2697 12257 2731 12291
rect 2731 12257 2740 12291
rect 2688 12248 2740 12257
rect 6276 12248 6328 12300
rect 5356 12223 5408 12232
rect 5356 12189 5365 12223
rect 5365 12189 5399 12223
rect 5399 12189 5408 12223
rect 5356 12180 5408 12189
rect 5632 12180 5684 12232
rect 2596 12044 2648 12096
rect 2872 12087 2924 12096
rect 2872 12053 2881 12087
rect 2881 12053 2915 12087
rect 2915 12053 2924 12087
rect 2872 12044 2924 12053
rect 3608 12087 3660 12096
rect 3608 12053 3617 12087
rect 3617 12053 3651 12087
rect 3651 12053 3660 12087
rect 3608 12044 3660 12053
rect 4344 12087 4396 12096
rect 4344 12053 4353 12087
rect 4353 12053 4387 12087
rect 4387 12053 4396 12087
rect 4344 12044 4396 12053
rect 4804 12044 4856 12096
rect 4988 12087 5040 12096
rect 4988 12053 4997 12087
rect 4997 12053 5031 12087
rect 5031 12053 5040 12087
rect 4988 12044 5040 12053
rect 5908 12087 5960 12096
rect 5908 12053 5917 12087
rect 5917 12053 5951 12087
rect 5951 12053 5960 12087
rect 5908 12044 5960 12053
rect 7472 12044 7524 12096
rect 11704 12316 11756 12368
rect 17868 12316 17920 12368
rect 21364 12316 21416 12368
rect 25044 12316 25096 12368
rect 8300 12291 8352 12300
rect 8300 12257 8309 12291
rect 8309 12257 8343 12291
rect 8343 12257 8352 12291
rect 8300 12248 8352 12257
rect 31300 12248 31352 12300
rect 32956 12248 33008 12300
rect 33324 12248 33376 12300
rect 8576 12223 8628 12232
rect 8576 12189 8585 12223
rect 8585 12189 8619 12223
rect 8619 12189 8628 12223
rect 8576 12180 8628 12189
rect 11888 12223 11940 12232
rect 11888 12189 11897 12223
rect 11897 12189 11931 12223
rect 11931 12189 11940 12223
rect 11888 12180 11940 12189
rect 12256 12180 12308 12232
rect 17776 12223 17828 12232
rect 17776 12189 17785 12223
rect 17785 12189 17819 12223
rect 17819 12189 17828 12223
rect 17776 12180 17828 12189
rect 17500 12112 17552 12164
rect 21824 12180 21876 12232
rect 24952 12223 25004 12232
rect 24952 12189 24961 12223
rect 24961 12189 24995 12223
rect 24995 12189 25004 12223
rect 24952 12180 25004 12189
rect 25872 12180 25924 12232
rect 21732 12112 21784 12164
rect 24400 12112 24452 12164
rect 36268 12248 36320 12300
rect 33784 12112 33836 12164
rect 34612 12112 34664 12164
rect 8024 12087 8076 12096
rect 8024 12053 8033 12087
rect 8033 12053 8067 12087
rect 8067 12053 8076 12087
rect 8024 12044 8076 12053
rect 8944 12087 8996 12096
rect 8944 12053 8953 12087
rect 8953 12053 8987 12087
rect 8987 12053 8996 12087
rect 8944 12044 8996 12053
rect 11060 12044 11112 12096
rect 12992 12087 13044 12096
rect 12992 12053 13001 12087
rect 13001 12053 13035 12087
rect 13035 12053 13044 12087
rect 12992 12044 13044 12053
rect 15844 12044 15896 12096
rect 17408 12044 17460 12096
rect 18236 12044 18288 12096
rect 20628 12044 20680 12096
rect 24676 12044 24728 12096
rect 25504 12044 25556 12096
rect 25964 12044 26016 12096
rect 27436 12044 27488 12096
rect 30196 12087 30248 12096
rect 30196 12053 30205 12087
rect 30205 12053 30239 12087
rect 30239 12053 30248 12087
rect 30196 12044 30248 12053
rect 31024 12044 31076 12096
rect 32772 12087 32824 12096
rect 32772 12053 32781 12087
rect 32781 12053 32815 12087
rect 32815 12053 32824 12087
rect 32772 12044 32824 12053
rect 33692 12044 33744 12096
rect 35532 12044 35584 12096
rect 7648 11942 7700 11994
rect 7712 11942 7764 11994
rect 7776 11942 7828 11994
rect 7840 11942 7892 11994
rect 20982 11942 21034 11994
rect 21046 11942 21098 11994
rect 21110 11942 21162 11994
rect 21174 11942 21226 11994
rect 34315 11942 34367 11994
rect 34379 11942 34431 11994
rect 34443 11942 34495 11994
rect 34507 11942 34559 11994
rect 2504 11840 2556 11892
rect 4712 11840 4764 11892
rect 7012 11883 7064 11892
rect 7012 11849 7021 11883
rect 7021 11849 7055 11883
rect 7055 11849 7064 11883
rect 7012 11840 7064 11849
rect 1676 11772 1728 11824
rect 2688 11772 2740 11824
rect 2504 11747 2556 11756
rect 2504 11713 2513 11747
rect 2513 11713 2547 11747
rect 2547 11713 2556 11747
rect 2504 11704 2556 11713
rect 2596 11747 2648 11756
rect 2596 11713 2605 11747
rect 2605 11713 2639 11747
rect 2639 11713 2648 11747
rect 2596 11704 2648 11713
rect 3608 11704 3660 11756
rect 4988 11704 5040 11756
rect 5908 11704 5960 11756
rect 7380 11704 7432 11756
rect 8300 11840 8352 11892
rect 10692 11883 10744 11892
rect 10692 11849 10701 11883
rect 10701 11849 10735 11883
rect 10735 11849 10744 11883
rect 10692 11840 10744 11849
rect 10968 11840 11020 11892
rect 17500 11883 17552 11892
rect 17500 11849 17509 11883
rect 17509 11849 17543 11883
rect 17543 11849 17552 11883
rect 17500 11840 17552 11849
rect 25044 11883 25096 11892
rect 25044 11849 25053 11883
rect 25053 11849 25087 11883
rect 25087 11849 25096 11883
rect 25044 11840 25096 11849
rect 26516 11883 26568 11892
rect 26516 11849 26525 11883
rect 26525 11849 26559 11883
rect 26559 11849 26568 11883
rect 29552 11883 29604 11892
rect 26516 11840 26568 11849
rect 8024 11772 8076 11824
rect 13176 11772 13228 11824
rect 16488 11815 16540 11824
rect 16488 11781 16497 11815
rect 16497 11781 16531 11815
rect 16531 11781 16540 11815
rect 16488 11772 16540 11781
rect 23756 11772 23808 11824
rect 8116 11704 8168 11756
rect 12808 11704 12860 11756
rect 16948 11747 17000 11756
rect 16948 11713 16957 11747
rect 16957 11713 16991 11747
rect 16991 11713 17000 11747
rect 16948 11704 17000 11713
rect 24400 11747 24452 11756
rect 24400 11713 24409 11747
rect 24409 11713 24443 11747
rect 24443 11713 24452 11747
rect 24400 11704 24452 11713
rect 5632 11636 5684 11688
rect 6828 11679 6880 11688
rect 6828 11645 6837 11679
rect 6837 11645 6871 11679
rect 6871 11645 6880 11679
rect 11060 11679 11112 11688
rect 6828 11636 6880 11645
rect 2412 11568 2464 11620
rect 4160 11611 4212 11620
rect 4160 11577 4169 11611
rect 4169 11577 4203 11611
rect 4203 11577 4212 11611
rect 4160 11568 4212 11577
rect 6000 11568 6052 11620
rect 3608 11500 3660 11552
rect 4896 11543 4948 11552
rect 4896 11509 4905 11543
rect 4905 11509 4939 11543
rect 4939 11509 4948 11543
rect 4896 11500 4948 11509
rect 6276 11500 6328 11552
rect 11060 11645 11069 11679
rect 11069 11645 11103 11679
rect 11103 11645 11112 11679
rect 11060 11636 11112 11645
rect 13452 11636 13504 11688
rect 20904 11636 20956 11688
rect 8576 11568 8628 11620
rect 12992 11568 13044 11620
rect 15844 11568 15896 11620
rect 17684 11568 17736 11620
rect 17776 11568 17828 11620
rect 19524 11568 19576 11620
rect 19616 11568 19668 11620
rect 27160 11815 27212 11824
rect 27160 11781 27169 11815
rect 27169 11781 27203 11815
rect 27203 11781 27212 11815
rect 27160 11772 27212 11781
rect 24676 11704 24728 11756
rect 7564 11500 7616 11552
rect 8300 11500 8352 11552
rect 8944 11500 8996 11552
rect 9128 11543 9180 11552
rect 9128 11509 9137 11543
rect 9137 11509 9171 11543
rect 9171 11509 9180 11543
rect 9128 11500 9180 11509
rect 12256 11500 12308 11552
rect 12624 11500 12676 11552
rect 15936 11543 15988 11552
rect 15936 11509 15945 11543
rect 15945 11509 15979 11543
rect 15979 11509 15988 11543
rect 15936 11500 15988 11509
rect 16212 11500 16264 11552
rect 17132 11500 17184 11552
rect 17868 11543 17920 11552
rect 17868 11509 17877 11543
rect 17877 11509 17911 11543
rect 17911 11509 17920 11543
rect 17868 11500 17920 11509
rect 20812 11543 20864 11552
rect 20812 11509 20821 11543
rect 20821 11509 20855 11543
rect 20855 11509 20864 11543
rect 20812 11500 20864 11509
rect 21364 11543 21416 11552
rect 21364 11509 21373 11543
rect 21373 11509 21407 11543
rect 21407 11509 21416 11543
rect 21364 11500 21416 11509
rect 21732 11543 21784 11552
rect 21732 11509 21741 11543
rect 21741 11509 21775 11543
rect 21775 11509 21784 11543
rect 21732 11500 21784 11509
rect 21824 11500 21876 11552
rect 23296 11500 23348 11552
rect 23572 11500 23624 11552
rect 24400 11500 24452 11552
rect 27252 11704 27304 11756
rect 29552 11849 29561 11883
rect 29561 11849 29595 11883
rect 29595 11849 29604 11883
rect 29552 11840 29604 11849
rect 31944 11883 31996 11892
rect 31944 11849 31953 11883
rect 31953 11849 31987 11883
rect 31987 11849 31996 11883
rect 31944 11840 31996 11849
rect 33324 11883 33376 11892
rect 33324 11849 33333 11883
rect 33333 11849 33367 11883
rect 33367 11849 33376 11883
rect 33324 11840 33376 11849
rect 30380 11772 30432 11824
rect 32864 11772 32916 11824
rect 34612 11840 34664 11892
rect 36268 11883 36320 11892
rect 36268 11849 36277 11883
rect 36277 11849 36311 11883
rect 36311 11849 36320 11883
rect 36268 11840 36320 11849
rect 34152 11772 34204 11824
rect 33784 11747 33836 11756
rect 33784 11713 33793 11747
rect 33793 11713 33827 11747
rect 33827 11713 33836 11747
rect 33784 11704 33836 11713
rect 37556 11747 37608 11756
rect 37556 11713 37565 11747
rect 37565 11713 37599 11747
rect 37599 11713 37608 11747
rect 37556 11704 37608 11713
rect 29368 11679 29420 11688
rect 29368 11645 29377 11679
rect 29377 11645 29411 11679
rect 29411 11645 29420 11679
rect 29920 11679 29972 11688
rect 29368 11636 29420 11645
rect 29920 11645 29929 11679
rect 29929 11645 29963 11679
rect 29963 11645 29972 11679
rect 29920 11636 29972 11645
rect 30196 11636 30248 11688
rect 31668 11636 31720 11688
rect 31944 11636 31996 11688
rect 33876 11679 33928 11688
rect 33876 11645 33885 11679
rect 33885 11645 33919 11679
rect 33919 11645 33928 11679
rect 33876 11636 33928 11645
rect 25872 11568 25924 11620
rect 27436 11611 27488 11620
rect 27436 11577 27445 11611
rect 27445 11577 27479 11611
rect 27479 11577 27488 11611
rect 27436 11568 27488 11577
rect 31024 11611 31076 11620
rect 31024 11577 31033 11611
rect 31033 11577 31067 11611
rect 31067 11577 31076 11611
rect 31024 11568 31076 11577
rect 34612 11611 34664 11620
rect 25964 11500 26016 11552
rect 28264 11500 28316 11552
rect 34612 11577 34621 11611
rect 34621 11577 34655 11611
rect 34655 11577 34664 11611
rect 35992 11636 36044 11688
rect 34612 11568 34664 11577
rect 31208 11500 31260 11552
rect 31300 11500 31352 11552
rect 32312 11543 32364 11552
rect 32312 11509 32321 11543
rect 32321 11509 32355 11543
rect 32355 11509 32364 11543
rect 32312 11500 32364 11509
rect 32956 11500 33008 11552
rect 33140 11543 33192 11552
rect 33140 11509 33149 11543
rect 33149 11509 33183 11543
rect 33183 11509 33192 11543
rect 33784 11543 33836 11552
rect 33140 11500 33192 11509
rect 33784 11509 33793 11543
rect 33793 11509 33827 11543
rect 33827 11509 33836 11543
rect 33784 11500 33836 11509
rect 34888 11500 34940 11552
rect 36084 11500 36136 11552
rect 36820 11500 36872 11552
rect 14315 11398 14367 11450
rect 14379 11398 14431 11450
rect 14443 11398 14495 11450
rect 14507 11398 14559 11450
rect 27648 11398 27700 11450
rect 27712 11398 27764 11450
rect 27776 11398 27828 11450
rect 27840 11398 27892 11450
rect 2412 11296 2464 11348
rect 4160 11296 4212 11348
rect 5540 11296 5592 11348
rect 8392 11296 8444 11348
rect 15108 11296 15160 11348
rect 16028 11296 16080 11348
rect 16948 11296 17000 11348
rect 17408 11339 17460 11348
rect 17408 11305 17417 11339
rect 17417 11305 17451 11339
rect 17451 11305 17460 11339
rect 17408 11296 17460 11305
rect 17500 11296 17552 11348
rect 22928 11339 22980 11348
rect 22928 11305 22937 11339
rect 22937 11305 22971 11339
rect 22971 11305 22980 11339
rect 22928 11296 22980 11305
rect 23296 11296 23348 11348
rect 23848 11296 23900 11348
rect 3424 11228 3476 11280
rect 7104 11271 7156 11280
rect 7104 11237 7113 11271
rect 7113 11237 7147 11271
rect 7147 11237 7156 11271
rect 7104 11228 7156 11237
rect 9956 11271 10008 11280
rect 9956 11237 9990 11271
rect 9990 11237 10008 11271
rect 9956 11228 10008 11237
rect 12440 11228 12492 11280
rect 15936 11228 15988 11280
rect 3700 11160 3752 11212
rect 4160 11160 4212 11212
rect 5632 11160 5684 11212
rect 5816 11160 5868 11212
rect 1400 11135 1452 11144
rect 1400 11101 1409 11135
rect 1409 11101 1443 11135
rect 1443 11101 1452 11135
rect 1400 11092 1452 11101
rect 2964 11135 3016 11144
rect 2964 11101 2973 11135
rect 2973 11101 3007 11135
rect 3007 11101 3016 11135
rect 2964 11092 3016 11101
rect 3976 11092 4028 11144
rect 8392 11160 8444 11212
rect 10692 11160 10744 11212
rect 11888 11160 11940 11212
rect 12808 11203 12860 11212
rect 12808 11169 12817 11203
rect 12817 11169 12851 11203
rect 12851 11169 12860 11203
rect 12808 11160 12860 11169
rect 2504 11067 2556 11076
rect 2504 11033 2513 11067
rect 2513 11033 2547 11067
rect 2547 11033 2556 11067
rect 2504 11024 2556 11033
rect 2688 11024 2740 11076
rect 3608 11067 3660 11076
rect 3608 11033 3617 11067
rect 3617 11033 3651 11067
rect 3651 11033 3660 11067
rect 3608 11024 3660 11033
rect 5356 11024 5408 11076
rect 3148 10956 3200 11008
rect 4344 10956 4396 11008
rect 6828 10956 6880 11008
rect 8300 11092 8352 11144
rect 8668 11092 8720 11144
rect 9680 11135 9732 11144
rect 9680 11101 9689 11135
rect 9689 11101 9723 11135
rect 9723 11101 9732 11135
rect 9680 11092 9732 11101
rect 11704 11135 11756 11144
rect 11704 11101 11713 11135
rect 11713 11101 11747 11135
rect 11747 11101 11756 11135
rect 11704 11092 11756 11101
rect 13084 11135 13136 11144
rect 13084 11101 13093 11135
rect 13093 11101 13127 11135
rect 13127 11101 13136 11135
rect 13084 11092 13136 11101
rect 11152 11024 11204 11076
rect 12532 11067 12584 11076
rect 12532 11033 12541 11067
rect 12541 11033 12575 11067
rect 12575 11033 12584 11067
rect 12532 11024 12584 11033
rect 18788 11160 18840 11212
rect 19064 11271 19116 11280
rect 19064 11237 19073 11271
rect 19073 11237 19107 11271
rect 19107 11237 19116 11271
rect 19064 11228 19116 11237
rect 20812 11228 20864 11280
rect 21640 11228 21692 11280
rect 24400 11228 24452 11280
rect 24584 11228 24636 11280
rect 26332 11228 26384 11280
rect 27160 11228 27212 11280
rect 30932 11271 30984 11280
rect 30932 11237 30941 11271
rect 30941 11237 30975 11271
rect 30975 11237 30984 11271
rect 30932 11228 30984 11237
rect 32680 11228 32732 11280
rect 33876 11228 33928 11280
rect 35716 11228 35768 11280
rect 36360 11228 36412 11280
rect 20720 11160 20772 11212
rect 20904 11203 20956 11212
rect 20904 11169 20913 11203
rect 20913 11169 20947 11203
rect 20947 11169 20956 11203
rect 20904 11160 20956 11169
rect 23756 11203 23808 11212
rect 23756 11169 23765 11203
rect 23765 11169 23799 11203
rect 23799 11169 23808 11203
rect 23756 11160 23808 11169
rect 24860 11160 24912 11212
rect 26240 11203 26292 11212
rect 26240 11169 26249 11203
rect 26249 11169 26283 11203
rect 26283 11169 26292 11203
rect 26240 11160 26292 11169
rect 28448 11203 28500 11212
rect 28448 11169 28482 11203
rect 28482 11169 28500 11203
rect 28448 11160 28500 11169
rect 30380 11160 30432 11212
rect 33048 11160 33100 11212
rect 15752 11135 15804 11144
rect 9128 10999 9180 11008
rect 9128 10965 9137 10999
rect 9137 10965 9171 10999
rect 9171 10965 9180 10999
rect 9128 10956 9180 10965
rect 9588 10956 9640 11008
rect 15016 10956 15068 11008
rect 15752 11101 15761 11135
rect 15761 11101 15795 11135
rect 15795 11101 15804 11135
rect 15752 11092 15804 11101
rect 15844 11092 15896 11144
rect 17132 11092 17184 11144
rect 17684 11092 17736 11144
rect 18236 11092 18288 11144
rect 18880 11135 18932 11144
rect 18880 11101 18889 11135
rect 18889 11101 18923 11135
rect 18923 11101 18932 11135
rect 18880 11092 18932 11101
rect 24032 11135 24084 11144
rect 24032 11101 24041 11135
rect 24041 11101 24075 11135
rect 24075 11101 24084 11135
rect 24032 11092 24084 11101
rect 26700 11092 26752 11144
rect 28172 11135 28224 11144
rect 28172 11101 28181 11135
rect 28181 11101 28215 11135
rect 28215 11101 28224 11135
rect 28172 11092 28224 11101
rect 32864 11092 32916 11144
rect 36084 11135 36136 11144
rect 36084 11101 36093 11135
rect 36093 11101 36127 11135
rect 36127 11101 36136 11135
rect 36084 11092 36136 11101
rect 16856 11024 16908 11076
rect 19616 11067 19668 11076
rect 19616 11033 19625 11067
rect 19625 11033 19659 11067
rect 19659 11033 19668 11067
rect 19616 11024 19668 11033
rect 22284 11067 22336 11076
rect 22284 11033 22293 11067
rect 22293 11033 22327 11067
rect 22327 11033 22336 11067
rect 22284 11024 22336 11033
rect 23480 11067 23532 11076
rect 23480 11033 23489 11067
rect 23489 11033 23523 11067
rect 23523 11033 23532 11067
rect 23480 11024 23532 11033
rect 24952 11024 25004 11076
rect 25320 11024 25372 11076
rect 26608 11067 26660 11076
rect 26608 11033 26617 11067
rect 26617 11033 26651 11067
rect 26651 11033 26660 11067
rect 26608 11024 26660 11033
rect 29552 11067 29604 11076
rect 29552 11033 29561 11067
rect 29561 11033 29595 11067
rect 29595 11033 29604 11067
rect 29552 11024 29604 11033
rect 24308 10956 24360 11008
rect 25044 10956 25096 11008
rect 25872 10956 25924 11008
rect 30840 10956 30892 11008
rect 34520 11024 34572 11076
rect 34888 11067 34940 11076
rect 34888 11033 34897 11067
rect 34897 11033 34931 11067
rect 34931 11033 34940 11067
rect 34888 11024 34940 11033
rect 35532 11067 35584 11076
rect 35532 11033 35541 11067
rect 35541 11033 35575 11067
rect 35575 11033 35584 11067
rect 35532 11024 35584 11033
rect 33692 10956 33744 11008
rect 33876 10956 33928 11008
rect 35624 10956 35676 11008
rect 7648 10854 7700 10906
rect 7712 10854 7764 10906
rect 7776 10854 7828 10906
rect 7840 10854 7892 10906
rect 20982 10854 21034 10906
rect 21046 10854 21098 10906
rect 21110 10854 21162 10906
rect 21174 10854 21226 10906
rect 34315 10854 34367 10906
rect 34379 10854 34431 10906
rect 34443 10854 34495 10906
rect 34507 10854 34559 10906
rect 1400 10752 1452 10804
rect 3884 10795 3936 10804
rect 3884 10761 3893 10795
rect 3893 10761 3927 10795
rect 3927 10761 3936 10795
rect 3884 10752 3936 10761
rect 5264 10795 5316 10804
rect 5264 10761 5273 10795
rect 5273 10761 5307 10795
rect 5307 10761 5316 10795
rect 5264 10752 5316 10761
rect 5724 10752 5776 10804
rect 6828 10752 6880 10804
rect 6920 10752 6972 10804
rect 2228 10727 2280 10736
rect 2228 10693 2237 10727
rect 2237 10693 2271 10727
rect 2271 10693 2280 10727
rect 2228 10684 2280 10693
rect 4160 10684 4212 10736
rect 7932 10684 7984 10736
rect 8392 10752 8444 10804
rect 9956 10752 10008 10804
rect 10784 10795 10836 10804
rect 10784 10761 10793 10795
rect 10793 10761 10827 10795
rect 10827 10761 10836 10795
rect 10784 10752 10836 10761
rect 15108 10752 15160 10804
rect 17868 10752 17920 10804
rect 19064 10795 19116 10804
rect 19064 10761 19073 10795
rect 19073 10761 19107 10795
rect 19107 10761 19116 10795
rect 19064 10752 19116 10761
rect 19524 10752 19576 10804
rect 20812 10752 20864 10804
rect 23848 10795 23900 10804
rect 23848 10761 23857 10795
rect 23857 10761 23891 10795
rect 23891 10761 23900 10795
rect 23848 10752 23900 10761
rect 25872 10795 25924 10804
rect 25872 10761 25881 10795
rect 25881 10761 25915 10795
rect 25915 10761 25924 10795
rect 25872 10752 25924 10761
rect 27804 10795 27856 10804
rect 27804 10761 27813 10795
rect 27813 10761 27847 10795
rect 27847 10761 27856 10795
rect 27804 10752 27856 10761
rect 28448 10752 28500 10804
rect 30288 10752 30340 10804
rect 31208 10752 31260 10804
rect 31668 10795 31720 10804
rect 31668 10761 31677 10795
rect 31677 10761 31711 10795
rect 31711 10761 31720 10795
rect 31668 10752 31720 10761
rect 32680 10795 32732 10804
rect 32680 10761 32689 10795
rect 32689 10761 32723 10795
rect 32723 10761 32732 10795
rect 32680 10752 32732 10761
rect 32864 10752 32916 10804
rect 33968 10752 34020 10804
rect 35716 10752 35768 10804
rect 9496 10684 9548 10736
rect 14096 10684 14148 10736
rect 15016 10727 15068 10736
rect 15016 10693 15025 10727
rect 15025 10693 15059 10727
rect 15059 10693 15068 10727
rect 15016 10684 15068 10693
rect 20720 10684 20772 10736
rect 23572 10684 23624 10736
rect 4988 10616 5040 10668
rect 5632 10659 5684 10668
rect 5632 10625 5641 10659
rect 5641 10625 5675 10659
rect 5675 10625 5684 10659
rect 5632 10616 5684 10625
rect 5816 10659 5868 10668
rect 5816 10625 5825 10659
rect 5825 10625 5859 10659
rect 5859 10625 5868 10659
rect 5816 10616 5868 10625
rect 9680 10616 9732 10668
rect 4804 10548 4856 10600
rect 6552 10548 6604 10600
rect 8300 10548 8352 10600
rect 9588 10548 9640 10600
rect 11060 10591 11112 10600
rect 11060 10557 11069 10591
rect 11069 10557 11103 10591
rect 11103 10557 11112 10591
rect 11060 10548 11112 10557
rect 18236 10616 18288 10668
rect 19616 10616 19668 10668
rect 23020 10659 23072 10668
rect 23020 10625 23029 10659
rect 23029 10625 23063 10659
rect 23063 10625 23072 10659
rect 23020 10616 23072 10625
rect 24032 10616 24084 10668
rect 24400 10659 24452 10668
rect 24400 10625 24409 10659
rect 24409 10625 24443 10659
rect 24443 10625 24452 10659
rect 24400 10616 24452 10625
rect 24768 10616 24820 10668
rect 25320 10659 25372 10668
rect 25320 10625 25329 10659
rect 25329 10625 25363 10659
rect 25363 10625 25372 10659
rect 25320 10616 25372 10625
rect 33692 10684 33744 10736
rect 35164 10684 35216 10736
rect 35992 10684 36044 10736
rect 12716 10548 12768 10600
rect 15108 10591 15160 10600
rect 15108 10557 15117 10591
rect 15117 10557 15151 10591
rect 15151 10557 15160 10591
rect 15108 10548 15160 10557
rect 16948 10548 17000 10600
rect 18328 10548 18380 10600
rect 19984 10591 20036 10600
rect 19984 10557 19993 10591
rect 19993 10557 20027 10591
rect 20027 10557 20036 10591
rect 19984 10548 20036 10557
rect 26700 10591 26752 10600
rect 26700 10557 26723 10591
rect 26723 10557 26752 10591
rect 3148 10480 3200 10532
rect 4620 10480 4672 10532
rect 3700 10412 3752 10464
rect 5356 10412 5408 10464
rect 10324 10480 10376 10532
rect 11336 10523 11388 10532
rect 11336 10489 11345 10523
rect 11345 10489 11379 10523
rect 11379 10489 11388 10523
rect 11336 10480 11388 10489
rect 13544 10480 13596 10532
rect 5816 10412 5868 10464
rect 6828 10412 6880 10464
rect 11796 10455 11848 10464
rect 11796 10421 11805 10455
rect 11805 10421 11839 10455
rect 11839 10421 11848 10455
rect 11796 10412 11848 10421
rect 13084 10412 13136 10464
rect 16488 10455 16540 10464
rect 16488 10421 16497 10455
rect 16497 10421 16531 10455
rect 16531 10421 16540 10455
rect 16488 10412 16540 10421
rect 17132 10455 17184 10464
rect 17132 10421 17141 10455
rect 17141 10421 17175 10455
rect 17175 10421 17184 10455
rect 17132 10412 17184 10421
rect 17408 10455 17460 10464
rect 17408 10421 17417 10455
rect 17417 10421 17451 10455
rect 17451 10421 17460 10455
rect 17408 10412 17460 10421
rect 24308 10523 24360 10532
rect 20168 10455 20220 10464
rect 20168 10421 20177 10455
rect 20177 10421 20211 10455
rect 20211 10421 20220 10455
rect 20168 10412 20220 10421
rect 22008 10412 22060 10464
rect 24308 10489 24317 10523
rect 24317 10489 24351 10523
rect 24351 10489 24360 10523
rect 24308 10480 24360 10489
rect 24492 10480 24544 10532
rect 26700 10548 26752 10557
rect 27068 10480 27120 10532
rect 28172 10480 28224 10532
rect 29092 10480 29144 10532
rect 33140 10616 33192 10668
rect 34152 10616 34204 10668
rect 32772 10548 32824 10600
rect 33876 10591 33928 10600
rect 33876 10557 33885 10591
rect 33885 10557 33919 10591
rect 33919 10557 33928 10591
rect 33876 10548 33928 10557
rect 30840 10480 30892 10532
rect 33692 10480 33744 10532
rect 22928 10412 22980 10464
rect 24860 10412 24912 10464
rect 30012 10412 30064 10464
rect 36268 10616 36320 10668
rect 37280 10616 37332 10668
rect 35992 10548 36044 10600
rect 35532 10523 35584 10532
rect 34612 10455 34664 10464
rect 34612 10421 34621 10455
rect 34621 10421 34655 10455
rect 34655 10421 34664 10455
rect 34612 10412 34664 10421
rect 35164 10412 35216 10464
rect 35532 10489 35541 10523
rect 35541 10489 35575 10523
rect 35575 10489 35584 10523
rect 35532 10480 35584 10489
rect 35624 10412 35676 10464
rect 36360 10455 36412 10464
rect 36360 10421 36369 10455
rect 36369 10421 36403 10455
rect 36403 10421 36412 10455
rect 36360 10412 36412 10421
rect 36912 10412 36964 10464
rect 14315 10310 14367 10362
rect 14379 10310 14431 10362
rect 14443 10310 14495 10362
rect 14507 10310 14559 10362
rect 27648 10310 27700 10362
rect 27712 10310 27764 10362
rect 27776 10310 27828 10362
rect 27840 10310 27892 10362
rect 1676 10208 1728 10260
rect 4068 10208 4120 10260
rect 5908 10208 5960 10260
rect 6644 10251 6696 10260
rect 6644 10217 6653 10251
rect 6653 10217 6687 10251
rect 6687 10217 6696 10251
rect 6644 10208 6696 10217
rect 9128 10251 9180 10260
rect 2228 10140 2280 10192
rect 5540 10183 5592 10192
rect 5540 10149 5574 10183
rect 5574 10149 5592 10183
rect 5540 10140 5592 10149
rect 8300 10140 8352 10192
rect 9128 10217 9137 10251
rect 9137 10217 9171 10251
rect 9171 10217 9180 10251
rect 9128 10208 9180 10217
rect 9864 10251 9916 10260
rect 9864 10217 9873 10251
rect 9873 10217 9907 10251
rect 9907 10217 9916 10251
rect 9864 10208 9916 10217
rect 10324 10251 10376 10260
rect 10324 10217 10333 10251
rect 10333 10217 10367 10251
rect 10367 10217 10376 10251
rect 10324 10208 10376 10217
rect 13084 10208 13136 10260
rect 16488 10251 16540 10260
rect 16488 10217 16497 10251
rect 16497 10217 16531 10251
rect 16531 10217 16540 10251
rect 16488 10208 16540 10217
rect 18236 10251 18288 10260
rect 18236 10217 18245 10251
rect 18245 10217 18279 10251
rect 18279 10217 18288 10251
rect 18236 10208 18288 10217
rect 18788 10251 18840 10260
rect 18788 10217 18797 10251
rect 18797 10217 18831 10251
rect 18831 10217 18840 10251
rect 18788 10208 18840 10217
rect 18880 10208 18932 10260
rect 21824 10251 21876 10260
rect 21824 10217 21833 10251
rect 21833 10217 21867 10251
rect 21867 10217 21876 10251
rect 21824 10208 21876 10217
rect 24400 10208 24452 10260
rect 9496 10140 9548 10192
rect 11336 10140 11388 10192
rect 11704 10183 11756 10192
rect 11704 10149 11713 10183
rect 11713 10149 11747 10183
rect 11747 10149 11756 10183
rect 11704 10140 11756 10149
rect 15292 10140 15344 10192
rect 17040 10140 17092 10192
rect 22376 10140 22428 10192
rect 4344 10072 4396 10124
rect 5356 10072 5408 10124
rect 10508 10072 10560 10124
rect 11520 10115 11572 10124
rect 11520 10081 11529 10115
rect 11529 10081 11563 10115
rect 11563 10081 11572 10115
rect 11520 10072 11572 10081
rect 12164 10072 12216 10124
rect 15660 10115 15712 10124
rect 15660 10081 15669 10115
rect 15669 10081 15703 10115
rect 15703 10081 15712 10115
rect 15660 10072 15712 10081
rect 1952 10004 2004 10056
rect 2596 10047 2648 10056
rect 2596 10013 2605 10047
rect 2605 10013 2639 10047
rect 2639 10013 2648 10047
rect 2596 10004 2648 10013
rect 4620 10047 4672 10056
rect 4620 10013 4629 10047
rect 4629 10013 4663 10047
rect 4663 10013 4672 10047
rect 4620 10004 4672 10013
rect 8484 10047 8536 10056
rect 8484 10013 8493 10047
rect 8493 10013 8527 10047
rect 8527 10013 8536 10047
rect 8484 10004 8536 10013
rect 11796 10047 11848 10056
rect 11796 10013 11805 10047
rect 11805 10013 11839 10047
rect 11839 10013 11848 10047
rect 11796 10004 11848 10013
rect 12716 10047 12768 10056
rect 12716 10013 12725 10047
rect 12725 10013 12759 10047
rect 12759 10013 12768 10047
rect 12716 10004 12768 10013
rect 13728 10004 13780 10056
rect 15108 10047 15160 10056
rect 15108 10013 15117 10047
rect 15117 10013 15151 10047
rect 15151 10013 15160 10047
rect 17684 10072 17736 10124
rect 24400 10072 24452 10124
rect 26148 10208 26200 10260
rect 26332 10251 26384 10260
rect 26332 10217 26341 10251
rect 26341 10217 26375 10251
rect 26375 10217 26384 10251
rect 26332 10208 26384 10217
rect 26700 10251 26752 10260
rect 26700 10217 26709 10251
rect 26709 10217 26743 10251
rect 26743 10217 26752 10251
rect 26700 10208 26752 10217
rect 35532 10208 35584 10260
rect 36084 10208 36136 10260
rect 25412 10140 25464 10192
rect 26516 10140 26568 10192
rect 27344 10183 27396 10192
rect 27344 10149 27378 10183
rect 27378 10149 27396 10183
rect 27344 10140 27396 10149
rect 28908 10140 28960 10192
rect 29000 10140 29052 10192
rect 30012 10140 30064 10192
rect 30932 10140 30984 10192
rect 31668 10140 31720 10192
rect 31852 10140 31904 10192
rect 27068 10115 27120 10124
rect 27068 10081 27077 10115
rect 27077 10081 27111 10115
rect 27111 10081 27120 10115
rect 27068 10072 27120 10081
rect 15936 10047 15988 10056
rect 15108 10004 15160 10013
rect 15936 10013 15945 10047
rect 15945 10013 15979 10047
rect 15979 10013 15988 10047
rect 15936 10004 15988 10013
rect 20720 10004 20772 10056
rect 25228 10047 25280 10056
rect 25228 10013 25237 10047
rect 25237 10013 25271 10047
rect 25271 10013 25280 10047
rect 25228 10004 25280 10013
rect 25320 10004 25372 10056
rect 30564 10115 30616 10124
rect 30564 10081 30573 10115
rect 30573 10081 30607 10115
rect 30607 10081 30616 10115
rect 30564 10072 30616 10081
rect 32864 10072 32916 10124
rect 30840 10047 30892 10056
rect 30840 10013 30849 10047
rect 30849 10013 30883 10047
rect 30883 10013 30892 10047
rect 30840 10004 30892 10013
rect 31668 10004 31720 10056
rect 3148 9936 3200 9988
rect 3700 9936 3752 9988
rect 8116 9979 8168 9988
rect 8116 9945 8125 9979
rect 8125 9945 8159 9979
rect 8159 9945 8168 9979
rect 8116 9936 8168 9945
rect 12348 9936 12400 9988
rect 24676 9936 24728 9988
rect 30196 9936 30248 9988
rect 35532 10072 35584 10124
rect 2412 9868 2464 9920
rect 3424 9911 3476 9920
rect 3424 9877 3433 9911
rect 3433 9877 3467 9911
rect 3467 9877 3476 9911
rect 3424 9868 3476 9877
rect 4068 9868 4120 9920
rect 5080 9911 5132 9920
rect 5080 9877 5089 9911
rect 5089 9877 5123 9911
rect 5123 9877 5132 9911
rect 5080 9868 5132 9877
rect 13636 9868 13688 9920
rect 15384 9911 15436 9920
rect 15384 9877 15393 9911
rect 15393 9877 15427 9911
rect 15427 9877 15436 9911
rect 15384 9868 15436 9877
rect 20168 9868 20220 9920
rect 20536 9868 20588 9920
rect 23480 9868 23532 9920
rect 24492 9911 24544 9920
rect 24492 9877 24501 9911
rect 24501 9877 24535 9911
rect 24535 9877 24544 9911
rect 24492 9868 24544 9877
rect 28448 9911 28500 9920
rect 28448 9877 28457 9911
rect 28457 9877 28491 9911
rect 28491 9877 28500 9911
rect 28448 9868 28500 9877
rect 31024 9868 31076 9920
rect 32588 9868 32640 9920
rect 33876 9868 33928 9920
rect 34704 9868 34756 9920
rect 7648 9766 7700 9818
rect 7712 9766 7764 9818
rect 7776 9766 7828 9818
rect 7840 9766 7892 9818
rect 20982 9766 21034 9818
rect 21046 9766 21098 9818
rect 21110 9766 21162 9818
rect 21174 9766 21226 9818
rect 34315 9766 34367 9818
rect 34379 9766 34431 9818
rect 34443 9766 34495 9818
rect 34507 9766 34559 9818
rect 3792 9664 3844 9716
rect 4528 9664 4580 9716
rect 5540 9664 5592 9716
rect 10508 9707 10560 9716
rect 10508 9673 10517 9707
rect 10517 9673 10551 9707
rect 10551 9673 10560 9707
rect 10508 9664 10560 9673
rect 11796 9664 11848 9716
rect 15292 9707 15344 9716
rect 15292 9673 15301 9707
rect 15301 9673 15335 9707
rect 15335 9673 15344 9707
rect 15292 9664 15344 9673
rect 17408 9664 17460 9716
rect 20720 9664 20772 9716
rect 2044 9639 2096 9648
rect 2044 9605 2053 9639
rect 2053 9605 2087 9639
rect 2087 9605 2096 9639
rect 2044 9596 2096 9605
rect 2964 9639 3016 9648
rect 2964 9605 2973 9639
rect 2973 9605 3007 9639
rect 3007 9605 3016 9639
rect 2964 9596 3016 9605
rect 7472 9596 7524 9648
rect 9588 9596 9640 9648
rect 11520 9596 11572 9648
rect 2412 9571 2464 9580
rect 2412 9537 2421 9571
rect 2421 9537 2455 9571
rect 2455 9537 2464 9571
rect 2412 9528 2464 9537
rect 2688 9528 2740 9580
rect 4528 9528 4580 9580
rect 7380 9528 7432 9580
rect 17040 9571 17092 9580
rect 3424 9460 3476 9512
rect 2504 9435 2556 9444
rect 2504 9401 2513 9435
rect 2513 9401 2547 9435
rect 2547 9401 2556 9435
rect 2504 9392 2556 9401
rect 3608 9460 3660 9512
rect 5356 9460 5408 9512
rect 17040 9537 17049 9571
rect 17049 9537 17083 9571
rect 17083 9537 17092 9571
rect 17040 9528 17092 9537
rect 17132 9528 17184 9580
rect 2596 9324 2648 9376
rect 3700 9392 3752 9444
rect 6092 9392 6144 9444
rect 7288 9435 7340 9444
rect 7288 9401 7297 9435
rect 7297 9401 7331 9435
rect 7331 9401 7340 9435
rect 7288 9392 7340 9401
rect 9128 9460 9180 9512
rect 12716 9460 12768 9512
rect 8668 9392 8720 9444
rect 13452 9392 13504 9444
rect 13728 9392 13780 9444
rect 16580 9392 16632 9444
rect 4252 9324 4304 9376
rect 5908 9324 5960 9376
rect 7932 9324 7984 9376
rect 8300 9324 8352 9376
rect 10784 9324 10836 9376
rect 11704 9324 11756 9376
rect 11980 9324 12032 9376
rect 12164 9367 12216 9376
rect 12164 9333 12173 9367
rect 12173 9333 12207 9367
rect 12207 9333 12216 9367
rect 12164 9324 12216 9333
rect 13360 9324 13412 9376
rect 14924 9324 14976 9376
rect 15660 9367 15712 9376
rect 15660 9333 15669 9367
rect 15669 9333 15703 9367
rect 15703 9333 15712 9367
rect 15660 9324 15712 9333
rect 17316 9324 17368 9376
rect 17684 9324 17736 9376
rect 19064 9460 19116 9512
rect 24032 9639 24084 9648
rect 24032 9605 24041 9639
rect 24041 9605 24075 9639
rect 24075 9605 24084 9639
rect 25228 9664 25280 9716
rect 25872 9707 25924 9716
rect 25872 9673 25881 9707
rect 25881 9673 25915 9707
rect 25915 9673 25924 9707
rect 25872 9664 25924 9673
rect 27344 9664 27396 9716
rect 29092 9664 29144 9716
rect 30288 9664 30340 9716
rect 24032 9596 24084 9605
rect 26056 9596 26108 9648
rect 29828 9639 29880 9648
rect 29828 9605 29837 9639
rect 29837 9605 29871 9639
rect 29871 9605 29880 9639
rect 29828 9596 29880 9605
rect 30748 9664 30800 9716
rect 35624 9664 35676 9716
rect 22376 9528 22428 9580
rect 28908 9528 28960 9580
rect 35808 9596 35860 9648
rect 36268 9639 36320 9648
rect 36268 9605 36277 9639
rect 36277 9605 36311 9639
rect 36311 9605 36320 9639
rect 36268 9596 36320 9605
rect 36544 9639 36596 9648
rect 36544 9605 36553 9639
rect 36553 9605 36587 9639
rect 36587 9605 36596 9639
rect 36544 9596 36596 9605
rect 30380 9528 30432 9580
rect 35532 9571 35584 9580
rect 21640 9460 21692 9512
rect 23388 9460 23440 9512
rect 24492 9503 24544 9512
rect 24492 9469 24501 9503
rect 24501 9469 24535 9503
rect 24535 9469 24544 9503
rect 27068 9503 27120 9512
rect 24492 9460 24544 9469
rect 27068 9469 27077 9503
rect 27077 9469 27111 9503
rect 27111 9469 27120 9503
rect 27068 9460 27120 9469
rect 35532 9537 35541 9571
rect 35541 9537 35575 9571
rect 35575 9537 35584 9571
rect 35532 9528 35584 9537
rect 19984 9324 20036 9376
rect 20168 9324 20220 9376
rect 23020 9392 23072 9444
rect 25412 9392 25464 9444
rect 28172 9392 28224 9444
rect 31024 9435 31076 9444
rect 31024 9401 31058 9435
rect 31058 9401 31076 9435
rect 31024 9392 31076 9401
rect 22376 9367 22428 9376
rect 22376 9333 22385 9367
rect 22385 9333 22419 9367
rect 22419 9333 22428 9367
rect 22376 9324 22428 9333
rect 24124 9324 24176 9376
rect 24400 9324 24452 9376
rect 28540 9367 28592 9376
rect 28540 9333 28549 9367
rect 28549 9333 28583 9367
rect 28583 9333 28592 9367
rect 28540 9324 28592 9333
rect 28908 9367 28960 9376
rect 28908 9333 28917 9367
rect 28917 9333 28951 9367
rect 28951 9333 28960 9367
rect 28908 9324 28960 9333
rect 30288 9367 30340 9376
rect 30288 9333 30297 9367
rect 30297 9333 30331 9367
rect 30331 9333 30340 9367
rect 30288 9324 30340 9333
rect 31668 9324 31720 9376
rect 31944 9324 31996 9376
rect 33692 9392 33744 9444
rect 33876 9435 33928 9444
rect 33876 9401 33885 9435
rect 33885 9401 33919 9435
rect 33919 9401 33928 9435
rect 33876 9392 33928 9401
rect 34704 9392 34756 9444
rect 34888 9392 34940 9444
rect 36268 9392 36320 9444
rect 32956 9324 33008 9376
rect 33140 9367 33192 9376
rect 33140 9333 33149 9367
rect 33149 9333 33183 9367
rect 33183 9333 33192 9367
rect 33140 9324 33192 9333
rect 34612 9367 34664 9376
rect 34612 9333 34621 9367
rect 34621 9333 34655 9367
rect 34655 9333 34664 9367
rect 34612 9324 34664 9333
rect 35900 9367 35952 9376
rect 35900 9333 35909 9367
rect 35909 9333 35943 9367
rect 35943 9333 35952 9367
rect 35900 9324 35952 9333
rect 37004 9367 37056 9376
rect 37004 9333 37013 9367
rect 37013 9333 37047 9367
rect 37047 9333 37056 9367
rect 37004 9324 37056 9333
rect 14315 9222 14367 9274
rect 14379 9222 14431 9274
rect 14443 9222 14495 9274
rect 14507 9222 14559 9274
rect 27648 9222 27700 9274
rect 27712 9222 27764 9274
rect 27776 9222 27828 9274
rect 27840 9222 27892 9274
rect 1676 9163 1728 9172
rect 1676 9129 1685 9163
rect 1685 9129 1719 9163
rect 1719 9129 1728 9163
rect 1676 9120 1728 9129
rect 1952 9163 2004 9172
rect 1952 9129 1961 9163
rect 1961 9129 1995 9163
rect 1995 9129 2004 9163
rect 1952 9120 2004 9129
rect 5080 9120 5132 9172
rect 7288 9120 7340 9172
rect 7932 9120 7984 9172
rect 8760 9120 8812 9172
rect 13452 9120 13504 9172
rect 14004 9120 14056 9172
rect 14924 9120 14976 9172
rect 5448 9052 5500 9104
rect 6644 9052 6696 9104
rect 7380 9095 7432 9104
rect 1676 8984 1728 9036
rect 2688 8984 2740 9036
rect 3700 8984 3752 9036
rect 5264 8984 5316 9036
rect 2872 8959 2924 8968
rect 2872 8925 2881 8959
rect 2881 8925 2915 8959
rect 2915 8925 2924 8959
rect 2872 8916 2924 8925
rect 5356 8959 5408 8968
rect 5356 8925 5365 8959
rect 5365 8925 5399 8959
rect 5399 8925 5408 8959
rect 5356 8916 5408 8925
rect 6368 8984 6420 9036
rect 7380 9061 7389 9095
rect 7389 9061 7423 9095
rect 7423 9061 7432 9095
rect 7380 9052 7432 9061
rect 8116 9052 8168 9104
rect 8668 9095 8720 9104
rect 8668 9061 8677 9095
rect 8677 9061 8711 9095
rect 8711 9061 8720 9095
rect 8668 9052 8720 9061
rect 9128 9052 9180 9104
rect 10232 9052 10284 9104
rect 11704 9095 11756 9104
rect 11704 9061 11713 9095
rect 11713 9061 11747 9095
rect 11747 9061 11756 9095
rect 11704 9052 11756 9061
rect 8484 8984 8536 9036
rect 12164 8984 12216 9036
rect 17040 9120 17092 9172
rect 18052 9163 18104 9172
rect 18052 9129 18061 9163
rect 18061 9129 18095 9163
rect 18095 9129 18104 9163
rect 18052 9120 18104 9129
rect 19524 9120 19576 9172
rect 23020 9163 23072 9172
rect 23020 9129 23029 9163
rect 23029 9129 23063 9163
rect 23063 9129 23072 9163
rect 23020 9120 23072 9129
rect 23480 9120 23532 9172
rect 25412 9163 25464 9172
rect 25412 9129 25421 9163
rect 25421 9129 25455 9163
rect 25455 9129 25464 9163
rect 25412 9120 25464 9129
rect 35808 9163 35860 9172
rect 35808 9129 35817 9163
rect 35817 9129 35851 9163
rect 35851 9129 35860 9163
rect 35808 9120 35860 9129
rect 15752 9052 15804 9104
rect 19892 9095 19944 9104
rect 19892 9061 19901 9095
rect 19901 9061 19935 9095
rect 19935 9061 19944 9095
rect 19892 9052 19944 9061
rect 21916 9095 21968 9104
rect 21916 9061 21950 9095
rect 21950 9061 21968 9095
rect 21916 9052 21968 9061
rect 24952 9052 25004 9104
rect 26976 9095 27028 9104
rect 26976 9061 26985 9095
rect 26985 9061 27019 9095
rect 27019 9061 27028 9095
rect 26976 9052 27028 9061
rect 27712 9052 27764 9104
rect 28448 9052 28500 9104
rect 30748 9052 30800 9104
rect 31852 9095 31904 9104
rect 31852 9061 31861 9095
rect 31861 9061 31895 9095
rect 31895 9061 31904 9095
rect 31852 9052 31904 9061
rect 34152 9052 34204 9104
rect 34888 9095 34940 9104
rect 34888 9061 34897 9095
rect 34897 9061 34931 9095
rect 34931 9061 34940 9095
rect 34888 9052 34940 9061
rect 15936 9027 15988 9036
rect 15936 8993 15945 9027
rect 15945 8993 15979 9027
rect 15979 8993 15988 9027
rect 15936 8984 15988 8993
rect 26056 8984 26108 9036
rect 27068 8984 27120 9036
rect 28080 8984 28132 9036
rect 30840 9027 30892 9036
rect 30840 8993 30849 9027
rect 30849 8993 30883 9027
rect 30883 8993 30892 9027
rect 30840 8984 30892 8993
rect 31944 8984 31996 9036
rect 33140 8984 33192 9036
rect 35624 9027 35676 9036
rect 35624 8993 35633 9027
rect 35633 8993 35667 9027
rect 35667 8993 35676 9027
rect 35624 8984 35676 8993
rect 35992 8984 36044 9036
rect 8576 8959 8628 8968
rect 2320 8891 2372 8900
rect 2320 8857 2329 8891
rect 2329 8857 2363 8891
rect 2363 8857 2372 8891
rect 2320 8848 2372 8857
rect 4160 8848 4212 8900
rect 6736 8848 6788 8900
rect 8576 8925 8585 8959
rect 8585 8925 8619 8959
rect 8619 8925 8628 8959
rect 8576 8916 8628 8925
rect 11612 8959 11664 8968
rect 11612 8925 11621 8959
rect 11621 8925 11655 8959
rect 11655 8925 11664 8959
rect 11612 8916 11664 8925
rect 13268 8959 13320 8968
rect 13268 8925 13277 8959
rect 13277 8925 13311 8959
rect 13311 8925 13320 8959
rect 13268 8916 13320 8925
rect 13544 8916 13596 8968
rect 15292 8916 15344 8968
rect 8208 8848 8260 8900
rect 11520 8848 11572 8900
rect 12808 8891 12860 8900
rect 12808 8857 12817 8891
rect 12817 8857 12851 8891
rect 12851 8857 12860 8891
rect 12808 8848 12860 8857
rect 18052 8916 18104 8968
rect 19800 8959 19852 8968
rect 18236 8848 18288 8900
rect 4344 8823 4396 8832
rect 4344 8789 4353 8823
rect 4353 8789 4387 8823
rect 4387 8789 4396 8823
rect 4344 8780 4396 8789
rect 5724 8780 5776 8832
rect 6460 8823 6512 8832
rect 6460 8789 6469 8823
rect 6469 8789 6503 8823
rect 6503 8789 6512 8823
rect 6460 8780 6512 8789
rect 10324 8780 10376 8832
rect 12164 8780 12216 8832
rect 13268 8780 13320 8832
rect 16580 8780 16632 8832
rect 16948 8780 17000 8832
rect 17868 8780 17920 8832
rect 18604 8823 18656 8832
rect 18604 8789 18613 8823
rect 18613 8789 18647 8823
rect 18647 8789 18656 8823
rect 18604 8780 18656 8789
rect 19800 8925 19809 8959
rect 19809 8925 19843 8959
rect 19843 8925 19852 8959
rect 19800 8916 19852 8925
rect 21640 8959 21692 8968
rect 21640 8925 21649 8959
rect 21649 8925 21683 8959
rect 21683 8925 21692 8959
rect 21640 8916 21692 8925
rect 25044 8916 25096 8968
rect 31024 8916 31076 8968
rect 31484 8916 31536 8968
rect 32680 8959 32732 8968
rect 32680 8925 32689 8959
rect 32689 8925 32723 8959
rect 32723 8925 32732 8959
rect 32680 8916 32732 8925
rect 33600 8916 33652 8968
rect 35900 8959 35952 8968
rect 35900 8925 35909 8959
rect 35909 8925 35943 8959
rect 35943 8925 35952 8959
rect 35900 8916 35952 8925
rect 36268 8916 36320 8968
rect 19340 8891 19392 8900
rect 19340 8857 19349 8891
rect 19349 8857 19383 8891
rect 19383 8857 19392 8891
rect 19340 8848 19392 8857
rect 30564 8891 30616 8900
rect 30564 8857 30573 8891
rect 30573 8857 30607 8891
rect 30607 8857 30616 8891
rect 30564 8848 30616 8857
rect 31760 8848 31812 8900
rect 33692 8848 33744 8900
rect 33968 8848 34020 8900
rect 34520 8848 34572 8900
rect 19984 8780 20036 8832
rect 20260 8823 20312 8832
rect 20260 8789 20269 8823
rect 20269 8789 20303 8823
rect 20303 8789 20312 8823
rect 20260 8780 20312 8789
rect 23756 8823 23808 8832
rect 23756 8789 23765 8823
rect 23765 8789 23799 8823
rect 23799 8789 23808 8823
rect 23756 8780 23808 8789
rect 24768 8780 24820 8832
rect 28172 8780 28224 8832
rect 29184 8780 29236 8832
rect 33784 8823 33836 8832
rect 33784 8789 33793 8823
rect 33793 8789 33827 8823
rect 33827 8789 33836 8823
rect 33784 8780 33836 8789
rect 35900 8780 35952 8832
rect 37004 8780 37056 8832
rect 7648 8678 7700 8730
rect 7712 8678 7764 8730
rect 7776 8678 7828 8730
rect 7840 8678 7892 8730
rect 20982 8678 21034 8730
rect 21046 8678 21098 8730
rect 21110 8678 21162 8730
rect 21174 8678 21226 8730
rect 34315 8678 34367 8730
rect 34379 8678 34431 8730
rect 34443 8678 34495 8730
rect 34507 8678 34559 8730
rect 1952 8576 2004 8628
rect 2504 8576 2556 8628
rect 3424 8576 3476 8628
rect 4160 8576 4212 8628
rect 5080 8576 5132 8628
rect 8576 8576 8628 8628
rect 9680 8619 9732 8628
rect 9680 8585 9689 8619
rect 9689 8585 9723 8619
rect 9723 8585 9732 8619
rect 9680 8576 9732 8585
rect 10232 8619 10284 8628
rect 10232 8585 10241 8619
rect 10241 8585 10275 8619
rect 10275 8585 10284 8619
rect 10232 8576 10284 8585
rect 10876 8619 10928 8628
rect 10876 8585 10885 8619
rect 10885 8585 10919 8619
rect 10919 8585 10928 8619
rect 10876 8576 10928 8585
rect 11612 8576 11664 8628
rect 14004 8619 14056 8628
rect 14004 8585 14013 8619
rect 14013 8585 14047 8619
rect 14047 8585 14056 8619
rect 14004 8576 14056 8585
rect 14924 8619 14976 8628
rect 14924 8585 14933 8619
rect 14933 8585 14967 8619
rect 14967 8585 14976 8619
rect 14924 8576 14976 8585
rect 17960 8576 18012 8628
rect 19800 8576 19852 8628
rect 23388 8619 23440 8628
rect 23388 8585 23397 8619
rect 23397 8585 23431 8619
rect 23431 8585 23440 8619
rect 23388 8576 23440 8585
rect 25044 8619 25096 8628
rect 25044 8585 25053 8619
rect 25053 8585 25087 8619
rect 25087 8585 25096 8619
rect 25044 8576 25096 8585
rect 26056 8619 26108 8628
rect 26056 8585 26065 8619
rect 26065 8585 26099 8619
rect 26099 8585 26108 8619
rect 26056 8576 26108 8585
rect 26516 8619 26568 8628
rect 26516 8585 26525 8619
rect 26525 8585 26559 8619
rect 26559 8585 26568 8619
rect 28080 8619 28132 8628
rect 26516 8576 26568 8585
rect 3976 8508 4028 8560
rect 7840 8508 7892 8560
rect 15752 8551 15804 8560
rect 15752 8517 15761 8551
rect 15761 8517 15795 8551
rect 15795 8517 15804 8551
rect 15752 8508 15804 8517
rect 16396 8508 16448 8560
rect 18144 8551 18196 8560
rect 18144 8517 18153 8551
rect 18153 8517 18187 8551
rect 18187 8517 18196 8551
rect 18144 8508 18196 8517
rect 19892 8508 19944 8560
rect 22008 8508 22060 8560
rect 5264 8440 5316 8492
rect 5540 8440 5592 8492
rect 6460 8440 6512 8492
rect 10324 8440 10376 8492
rect 16948 8483 17000 8492
rect 16948 8449 16957 8483
rect 16957 8449 16991 8483
rect 16991 8449 17000 8483
rect 16948 8440 17000 8449
rect 19064 8483 19116 8492
rect 19064 8449 19073 8483
rect 19073 8449 19107 8483
rect 19107 8449 19116 8483
rect 19064 8440 19116 8449
rect 20628 8483 20680 8492
rect 20628 8449 20637 8483
rect 20637 8449 20671 8483
rect 20671 8449 20680 8483
rect 20628 8440 20680 8449
rect 26884 8551 26936 8560
rect 26884 8517 26893 8551
rect 26893 8517 26927 8551
rect 26927 8517 26936 8551
rect 26884 8508 26936 8517
rect 27160 8551 27212 8560
rect 27160 8517 27169 8551
rect 27169 8517 27203 8551
rect 27203 8517 27212 8551
rect 27160 8508 27212 8517
rect 28080 8585 28089 8619
rect 28089 8585 28123 8619
rect 28123 8585 28132 8619
rect 28080 8576 28132 8585
rect 28540 8576 28592 8628
rect 30932 8619 30984 8628
rect 30932 8585 30941 8619
rect 30941 8585 30975 8619
rect 30975 8585 30984 8619
rect 30932 8576 30984 8585
rect 37280 8619 37332 8628
rect 37280 8585 37289 8619
rect 37289 8585 37323 8619
rect 37323 8585 37332 8619
rect 37280 8576 37332 8585
rect 23664 8483 23716 8492
rect 23664 8449 23673 8483
rect 23673 8449 23707 8483
rect 23707 8449 23716 8483
rect 23664 8440 23716 8449
rect 28356 8508 28408 8560
rect 30840 8508 30892 8560
rect 32772 8551 32824 8560
rect 32772 8517 32781 8551
rect 32781 8517 32815 8551
rect 32815 8517 32824 8551
rect 32772 8508 32824 8517
rect 33048 8551 33100 8560
rect 33048 8517 33057 8551
rect 33057 8517 33091 8551
rect 33091 8517 33100 8551
rect 33048 8508 33100 8517
rect 36268 8551 36320 8560
rect 36268 8517 36277 8551
rect 36277 8517 36311 8551
rect 36311 8517 36320 8551
rect 36268 8508 36320 8517
rect 37556 8551 37608 8560
rect 37556 8517 37565 8551
rect 37565 8517 37599 8551
rect 37599 8517 37608 8551
rect 37556 8508 37608 8517
rect 27712 8483 27764 8492
rect 27712 8449 27721 8483
rect 27721 8449 27755 8483
rect 27755 8449 27764 8483
rect 27712 8440 27764 8449
rect 30012 8440 30064 8492
rect 31484 8483 31536 8492
rect 31484 8449 31493 8483
rect 31493 8449 31527 8483
rect 31527 8449 31536 8483
rect 31484 8440 31536 8449
rect 33416 8483 33468 8492
rect 33416 8449 33425 8483
rect 33425 8449 33459 8483
rect 33459 8449 33468 8483
rect 33416 8440 33468 8449
rect 1952 8372 2004 8424
rect 5356 8372 5408 8424
rect 6828 8415 6880 8424
rect 6828 8381 6837 8415
rect 6837 8381 6871 8415
rect 6871 8381 6880 8415
rect 6828 8372 6880 8381
rect 5448 8304 5500 8356
rect 5724 8347 5776 8356
rect 5724 8313 5733 8347
rect 5733 8313 5767 8347
rect 5767 8313 5776 8347
rect 5724 8304 5776 8313
rect 6368 8347 6420 8356
rect 6368 8313 6377 8347
rect 6377 8313 6411 8347
rect 6411 8313 6420 8347
rect 6368 8304 6420 8313
rect 8392 8372 8444 8424
rect 10416 8372 10468 8424
rect 11888 8372 11940 8424
rect 18420 8415 18472 8424
rect 18420 8381 18429 8415
rect 18429 8381 18463 8415
rect 18463 8381 18472 8415
rect 18420 8372 18472 8381
rect 19984 8372 20036 8424
rect 20168 8372 20220 8424
rect 20904 8372 20956 8424
rect 21916 8372 21968 8424
rect 22100 8372 22152 8424
rect 8760 8304 8812 8356
rect 10968 8304 11020 8356
rect 11336 8347 11388 8356
rect 11336 8313 11345 8347
rect 11345 8313 11379 8347
rect 11379 8313 11388 8347
rect 11336 8304 11388 8313
rect 12532 8304 12584 8356
rect 15292 8347 15344 8356
rect 15292 8313 15301 8347
rect 15301 8313 15335 8347
rect 15335 8313 15344 8347
rect 15292 8304 15344 8313
rect 16304 8347 16356 8356
rect 16304 8313 16313 8347
rect 16313 8313 16347 8347
rect 16347 8313 16356 8347
rect 17040 8347 17092 8356
rect 16304 8304 16356 8313
rect 6460 8236 6512 8288
rect 6644 8236 6696 8288
rect 7012 8236 7064 8288
rect 7196 8236 7248 8288
rect 7472 8236 7524 8288
rect 8116 8236 8168 8288
rect 17040 8313 17049 8347
rect 17049 8313 17083 8347
rect 17083 8313 17092 8347
rect 17040 8304 17092 8313
rect 17224 8304 17276 8356
rect 18604 8347 18656 8356
rect 18604 8313 18613 8347
rect 18613 8313 18647 8347
rect 18647 8313 18656 8347
rect 18604 8304 18656 8313
rect 19616 8304 19668 8356
rect 20260 8304 20312 8356
rect 22468 8347 22520 8356
rect 21640 8279 21692 8288
rect 21640 8245 21649 8279
rect 21649 8245 21683 8279
rect 21683 8245 21692 8279
rect 21640 8236 21692 8245
rect 21916 8236 21968 8288
rect 22468 8313 22477 8347
rect 22477 8313 22511 8347
rect 22511 8313 22520 8347
rect 22468 8304 22520 8313
rect 23756 8304 23808 8356
rect 22376 8279 22428 8288
rect 22376 8245 22385 8279
rect 22385 8245 22419 8279
rect 22419 8245 22428 8279
rect 22376 8236 22428 8245
rect 24952 8304 25004 8356
rect 26884 8304 26936 8356
rect 28540 8372 28592 8424
rect 29184 8372 29236 8424
rect 30656 8415 30708 8424
rect 30656 8381 30665 8415
rect 30665 8381 30699 8415
rect 30699 8381 30708 8415
rect 30656 8372 30708 8381
rect 31116 8372 31168 8424
rect 32956 8372 33008 8424
rect 34060 8415 34112 8424
rect 34060 8381 34069 8415
rect 34069 8381 34103 8415
rect 34103 8381 34112 8415
rect 34060 8372 34112 8381
rect 34704 8372 34756 8424
rect 27712 8304 27764 8356
rect 32496 8347 32548 8356
rect 32496 8313 32505 8347
rect 32505 8313 32539 8347
rect 32539 8313 32548 8347
rect 33600 8347 33652 8356
rect 32496 8304 32548 8313
rect 25504 8236 25556 8288
rect 30380 8279 30432 8288
rect 30380 8245 30389 8279
rect 30389 8245 30423 8279
rect 30423 8245 30432 8279
rect 30380 8236 30432 8245
rect 32220 8236 32272 8288
rect 33600 8313 33609 8347
rect 33609 8313 33643 8347
rect 33643 8313 33652 8347
rect 33600 8304 33652 8313
rect 33876 8304 33928 8356
rect 34336 8304 34388 8356
rect 37372 8415 37424 8424
rect 37372 8381 37381 8415
rect 37381 8381 37415 8415
rect 37415 8381 37424 8415
rect 37372 8372 37424 8381
rect 33508 8279 33560 8288
rect 33508 8245 33517 8279
rect 33517 8245 33551 8279
rect 33551 8245 33560 8279
rect 33508 8236 33560 8245
rect 34704 8279 34756 8288
rect 34704 8245 34713 8279
rect 34713 8245 34747 8279
rect 34747 8245 34756 8279
rect 34704 8236 34756 8245
rect 35164 8236 35216 8288
rect 14315 8134 14367 8186
rect 14379 8134 14431 8186
rect 14443 8134 14495 8186
rect 14507 8134 14559 8186
rect 27648 8134 27700 8186
rect 27712 8134 27764 8186
rect 27776 8134 27828 8186
rect 27840 8134 27892 8186
rect 2780 8032 2832 8084
rect 3884 8075 3936 8084
rect 3884 8041 3893 8075
rect 3893 8041 3927 8075
rect 3927 8041 3936 8075
rect 3884 8032 3936 8041
rect 7472 8032 7524 8084
rect 8668 8075 8720 8084
rect 8668 8041 8677 8075
rect 8677 8041 8711 8075
rect 8711 8041 8720 8075
rect 8668 8032 8720 8041
rect 10968 8032 11020 8084
rect 12532 8032 12584 8084
rect 13544 8075 13596 8084
rect 13544 8041 13553 8075
rect 13553 8041 13587 8075
rect 13587 8041 13596 8075
rect 13544 8032 13596 8041
rect 17592 8075 17644 8084
rect 17592 8041 17601 8075
rect 17601 8041 17635 8075
rect 17635 8041 17644 8075
rect 17592 8032 17644 8041
rect 19524 8032 19576 8084
rect 20628 8075 20680 8084
rect 20628 8041 20637 8075
rect 20637 8041 20671 8075
rect 20671 8041 20680 8075
rect 20628 8032 20680 8041
rect 21732 8032 21784 8084
rect 21916 8075 21968 8084
rect 21916 8041 21925 8075
rect 21925 8041 21959 8075
rect 21959 8041 21968 8075
rect 21916 8032 21968 8041
rect 2320 8007 2372 8016
rect 2320 7973 2329 8007
rect 2329 7973 2363 8007
rect 2363 7973 2372 8007
rect 2320 7964 2372 7973
rect 2872 8007 2924 8016
rect 2872 7973 2881 8007
rect 2881 7973 2915 8007
rect 2915 7973 2924 8007
rect 2872 7964 2924 7973
rect 4160 7964 4212 8016
rect 5080 7964 5132 8016
rect 6644 7964 6696 8016
rect 7840 7964 7892 8016
rect 8392 7964 8444 8016
rect 9312 7964 9364 8016
rect 9680 7964 9732 8016
rect 2504 7896 2556 7948
rect 10324 7939 10376 7948
rect 10324 7905 10333 7939
rect 10333 7905 10367 7939
rect 10367 7905 10376 7939
rect 10324 7896 10376 7905
rect 11888 7964 11940 8016
rect 16672 8007 16724 8016
rect 16672 7973 16681 8007
rect 16681 7973 16715 8007
rect 16715 7973 16724 8007
rect 16672 7964 16724 7973
rect 17040 7964 17092 8016
rect 17776 7964 17828 8016
rect 18052 7964 18104 8016
rect 21364 7964 21416 8016
rect 22100 7964 22152 8016
rect 11520 7939 11572 7948
rect 11520 7905 11554 7939
rect 11554 7905 11572 7939
rect 11520 7896 11572 7905
rect 13728 7939 13780 7948
rect 13728 7905 13737 7939
rect 13737 7905 13771 7939
rect 13771 7905 13780 7939
rect 13728 7896 13780 7905
rect 16488 7939 16540 7948
rect 16488 7905 16497 7939
rect 16497 7905 16531 7939
rect 16531 7905 16540 7939
rect 16488 7896 16540 7905
rect 20168 7939 20220 7948
rect 2688 7828 2740 7880
rect 4712 7871 4764 7880
rect 4712 7837 4721 7871
rect 4721 7837 4755 7871
rect 4755 7837 4764 7871
rect 4712 7828 4764 7837
rect 8024 7828 8076 7880
rect 8116 7828 8168 7880
rect 8760 7828 8812 7880
rect 10048 7828 10100 7880
rect 15936 7828 15988 7880
rect 20168 7905 20177 7939
rect 20177 7905 20211 7939
rect 20211 7905 20220 7939
rect 20168 7896 20220 7905
rect 21548 7896 21600 7948
rect 25044 8032 25096 8084
rect 27160 8032 27212 8084
rect 28448 8032 28500 8084
rect 30472 8075 30524 8084
rect 30472 8041 30481 8075
rect 30481 8041 30515 8075
rect 30515 8041 30524 8075
rect 30472 8032 30524 8041
rect 30748 8032 30800 8084
rect 31484 8075 31536 8084
rect 31484 8041 31493 8075
rect 31493 8041 31527 8075
rect 31527 8041 31536 8075
rect 31484 8032 31536 8041
rect 31944 8075 31996 8084
rect 31944 8041 31953 8075
rect 31953 8041 31987 8075
rect 31987 8041 31996 8075
rect 31944 8032 31996 8041
rect 33600 8032 33652 8084
rect 34336 8075 34388 8084
rect 34336 8041 34345 8075
rect 34345 8041 34379 8075
rect 34379 8041 34388 8075
rect 34336 8032 34388 8041
rect 36268 8032 36320 8084
rect 35992 8007 36044 8016
rect 35992 7973 36001 8007
rect 36001 7973 36035 8007
rect 36035 7973 36044 8007
rect 35992 7964 36044 7973
rect 25504 7939 25556 7948
rect 25504 7905 25513 7939
rect 25513 7905 25547 7939
rect 25547 7905 25556 7939
rect 25504 7896 25556 7905
rect 26332 7896 26384 7948
rect 27344 7896 27396 7948
rect 28908 7896 28960 7948
rect 29092 7939 29144 7948
rect 29092 7905 29101 7939
rect 29101 7905 29135 7939
rect 29135 7905 29144 7939
rect 29092 7896 29144 7905
rect 29184 7896 29236 7948
rect 32404 7896 32456 7948
rect 34980 7896 35032 7948
rect 35532 7896 35584 7948
rect 17684 7871 17736 7880
rect 17684 7837 17693 7871
rect 17693 7837 17727 7871
rect 17727 7837 17736 7871
rect 17684 7828 17736 7837
rect 21640 7828 21692 7880
rect 21916 7828 21968 7880
rect 25412 7871 25464 7880
rect 25412 7837 25421 7871
rect 25421 7837 25455 7871
rect 25455 7837 25464 7871
rect 25412 7828 25464 7837
rect 27160 7871 27212 7880
rect 27160 7837 27169 7871
rect 27169 7837 27203 7871
rect 27203 7837 27212 7871
rect 27160 7828 27212 7837
rect 28080 7871 28132 7880
rect 28080 7837 28089 7871
rect 28089 7837 28123 7871
rect 28123 7837 28132 7871
rect 28080 7828 28132 7837
rect 32956 7871 33008 7880
rect 32956 7837 32965 7871
rect 32965 7837 32999 7871
rect 32999 7837 33008 7871
rect 32956 7828 33008 7837
rect 36452 7896 36504 7948
rect 35992 7828 36044 7880
rect 6828 7760 6880 7812
rect 8208 7760 8260 7812
rect 16212 7803 16264 7812
rect 16212 7769 16221 7803
rect 16221 7769 16255 7803
rect 16255 7769 16264 7803
rect 16212 7760 16264 7769
rect 24952 7803 25004 7812
rect 24952 7769 24961 7803
rect 24961 7769 24995 7803
rect 24995 7769 25004 7803
rect 24952 7760 25004 7769
rect 34796 7760 34848 7812
rect 1860 7735 1912 7744
rect 1860 7701 1869 7735
rect 1869 7701 1903 7735
rect 1903 7701 1912 7735
rect 1860 7692 1912 7701
rect 4344 7735 4396 7744
rect 4344 7701 4353 7735
rect 4353 7701 4387 7735
rect 4387 7701 4396 7735
rect 4344 7692 4396 7701
rect 6092 7735 6144 7744
rect 6092 7701 6101 7735
rect 6101 7701 6135 7735
rect 6135 7701 6144 7735
rect 6092 7692 6144 7701
rect 6460 7692 6512 7744
rect 7012 7692 7064 7744
rect 9772 7735 9824 7744
rect 9772 7701 9781 7735
rect 9781 7701 9815 7735
rect 9815 7701 9824 7735
rect 9772 7692 9824 7701
rect 14096 7692 14148 7744
rect 14648 7692 14700 7744
rect 17592 7692 17644 7744
rect 19248 7692 19300 7744
rect 21364 7692 21416 7744
rect 23388 7735 23440 7744
rect 23388 7701 23397 7735
rect 23397 7701 23431 7735
rect 23431 7701 23440 7735
rect 23388 7692 23440 7701
rect 32956 7692 33008 7744
rect 33140 7692 33192 7744
rect 34980 7735 35032 7744
rect 34980 7701 34989 7735
rect 34989 7701 35023 7735
rect 35023 7701 35032 7735
rect 34980 7692 35032 7701
rect 35256 7735 35308 7744
rect 35256 7701 35265 7735
rect 35265 7701 35299 7735
rect 35299 7701 35308 7735
rect 35256 7692 35308 7701
rect 35624 7692 35676 7744
rect 7648 7590 7700 7642
rect 7712 7590 7764 7642
rect 7776 7590 7828 7642
rect 7840 7590 7892 7642
rect 20982 7590 21034 7642
rect 21046 7590 21098 7642
rect 21110 7590 21162 7642
rect 21174 7590 21226 7642
rect 34315 7590 34367 7642
rect 34379 7590 34431 7642
rect 34443 7590 34495 7642
rect 34507 7590 34559 7642
rect 2688 7488 2740 7540
rect 5356 7488 5408 7540
rect 5540 7488 5592 7540
rect 6644 7531 6696 7540
rect 6644 7497 6653 7531
rect 6653 7497 6687 7531
rect 6687 7497 6696 7531
rect 6644 7488 6696 7497
rect 7380 7488 7432 7540
rect 8116 7488 8168 7540
rect 9312 7531 9364 7540
rect 9312 7497 9321 7531
rect 9321 7497 9355 7531
rect 9355 7497 9364 7531
rect 9312 7488 9364 7497
rect 11888 7531 11940 7540
rect 11888 7497 11897 7531
rect 11897 7497 11931 7531
rect 11931 7497 11940 7531
rect 11888 7488 11940 7497
rect 11980 7488 12032 7540
rect 15936 7531 15988 7540
rect 15936 7497 15945 7531
rect 15945 7497 15979 7531
rect 15979 7497 15988 7531
rect 15936 7488 15988 7497
rect 16488 7531 16540 7540
rect 16488 7497 16497 7531
rect 16497 7497 16531 7531
rect 16531 7497 16540 7531
rect 16488 7488 16540 7497
rect 19800 7488 19852 7540
rect 21548 7531 21600 7540
rect 21548 7497 21557 7531
rect 21557 7497 21591 7531
rect 21591 7497 21600 7531
rect 21548 7488 21600 7497
rect 22376 7488 22428 7540
rect 23664 7488 23716 7540
rect 2136 7420 2188 7472
rect 2320 7420 2372 7472
rect 3148 7420 3200 7472
rect 10968 7420 11020 7472
rect 13636 7420 13688 7472
rect 2780 7352 2832 7404
rect 6092 7352 6144 7404
rect 12164 7395 12216 7404
rect 12164 7361 12173 7395
rect 12173 7361 12207 7395
rect 12207 7361 12216 7395
rect 12164 7352 12216 7361
rect 13360 7352 13412 7404
rect 14096 7395 14148 7404
rect 14096 7361 14105 7395
rect 14105 7361 14139 7395
rect 14139 7361 14148 7395
rect 14740 7395 14792 7404
rect 14096 7352 14148 7361
rect 14740 7361 14749 7395
rect 14749 7361 14783 7395
rect 14783 7361 14792 7395
rect 14740 7352 14792 7361
rect 16212 7352 16264 7404
rect 17132 7352 17184 7404
rect 17592 7352 17644 7404
rect 20812 7352 20864 7404
rect 25412 7488 25464 7540
rect 27988 7488 28040 7540
rect 29000 7488 29052 7540
rect 32404 7531 32456 7540
rect 32404 7497 32413 7531
rect 32413 7497 32447 7531
rect 32447 7497 32456 7531
rect 32404 7488 32456 7497
rect 35992 7488 36044 7540
rect 26332 7463 26384 7472
rect 26332 7429 26341 7463
rect 26341 7429 26375 7463
rect 26375 7429 26384 7463
rect 26332 7420 26384 7429
rect 29092 7463 29144 7472
rect 29092 7429 29101 7463
rect 29101 7429 29135 7463
rect 29135 7429 29144 7463
rect 29092 7420 29144 7429
rect 31760 7420 31812 7472
rect 32864 7420 32916 7472
rect 33324 7463 33376 7472
rect 33324 7429 33333 7463
rect 33333 7429 33367 7463
rect 33367 7429 33376 7463
rect 33324 7420 33376 7429
rect 33600 7420 33652 7472
rect 26056 7395 26108 7404
rect 4344 7327 4396 7336
rect 4344 7293 4378 7327
rect 4378 7293 4396 7327
rect 2504 7259 2556 7268
rect 2504 7225 2513 7259
rect 2513 7225 2547 7259
rect 2547 7225 2556 7259
rect 2504 7216 2556 7225
rect 2964 7216 3016 7268
rect 4344 7284 4396 7293
rect 7380 7327 7432 7336
rect 7380 7293 7389 7327
rect 7389 7293 7423 7327
rect 7423 7293 7432 7327
rect 7380 7284 7432 7293
rect 7472 7284 7524 7336
rect 8024 7284 8076 7336
rect 11244 7284 11296 7336
rect 4712 7216 4764 7268
rect 6828 7216 6880 7268
rect 2596 7148 2648 7200
rect 3148 7148 3200 7200
rect 6644 7148 6696 7200
rect 7012 7148 7064 7200
rect 7564 7148 7616 7200
rect 11060 7216 11112 7268
rect 11336 7259 11388 7268
rect 11336 7225 11345 7259
rect 11345 7225 11379 7259
rect 11379 7225 11388 7259
rect 11336 7216 11388 7225
rect 12256 7216 12308 7268
rect 13176 7259 13228 7268
rect 13176 7225 13185 7259
rect 13185 7225 13219 7259
rect 13219 7225 13228 7259
rect 13176 7216 13228 7225
rect 13268 7259 13320 7268
rect 13268 7225 13277 7259
rect 13277 7225 13311 7259
rect 13311 7225 13320 7259
rect 16396 7284 16448 7336
rect 13268 7216 13320 7225
rect 14832 7259 14884 7268
rect 14832 7225 14841 7259
rect 14841 7225 14875 7259
rect 14875 7225 14884 7259
rect 14832 7216 14884 7225
rect 17684 7284 17736 7336
rect 18880 7284 18932 7336
rect 26056 7361 26065 7395
rect 26065 7361 26099 7395
rect 26099 7361 26108 7395
rect 27068 7395 27120 7404
rect 26056 7352 26108 7361
rect 27068 7361 27077 7395
rect 27077 7361 27111 7395
rect 27111 7361 27120 7395
rect 27068 7352 27120 7361
rect 29184 7352 29236 7404
rect 31576 7352 31628 7404
rect 33968 7352 34020 7404
rect 24124 7284 24176 7336
rect 28080 7284 28132 7336
rect 33232 7284 33284 7336
rect 35072 7284 35124 7336
rect 36084 7284 36136 7336
rect 18512 7216 18564 7268
rect 22744 7216 22796 7268
rect 9680 7191 9732 7200
rect 9680 7157 9689 7191
rect 9689 7157 9723 7191
rect 9723 7157 9732 7191
rect 9680 7148 9732 7157
rect 10048 7191 10100 7200
rect 10048 7157 10057 7191
rect 10057 7157 10091 7191
rect 10091 7157 10100 7191
rect 10048 7148 10100 7157
rect 10140 7148 10192 7200
rect 27160 7259 27212 7268
rect 27160 7225 27169 7259
rect 27169 7225 27203 7259
rect 27203 7225 27212 7259
rect 27160 7216 27212 7225
rect 29092 7216 29144 7268
rect 29828 7259 29880 7268
rect 29828 7225 29837 7259
rect 29837 7225 29871 7259
rect 29871 7225 29880 7259
rect 29828 7216 29880 7225
rect 31484 7259 31536 7268
rect 31484 7225 31493 7259
rect 31493 7225 31527 7259
rect 31527 7225 31536 7259
rect 31484 7216 31536 7225
rect 34612 7216 34664 7268
rect 34980 7216 35032 7268
rect 35716 7216 35768 7268
rect 14740 7191 14792 7200
rect 14740 7157 14749 7191
rect 14749 7157 14783 7191
rect 14783 7157 14792 7191
rect 14740 7148 14792 7157
rect 16212 7191 16264 7200
rect 16212 7157 16221 7191
rect 16221 7157 16255 7191
rect 16255 7157 16264 7191
rect 16212 7148 16264 7157
rect 19432 7191 19484 7200
rect 19432 7157 19441 7191
rect 19441 7157 19475 7191
rect 19475 7157 19484 7191
rect 19432 7148 19484 7157
rect 20904 7191 20956 7200
rect 20904 7157 20913 7191
rect 20913 7157 20947 7191
rect 20947 7157 20956 7191
rect 20904 7148 20956 7157
rect 22560 7191 22612 7200
rect 22560 7157 22569 7191
rect 22569 7157 22603 7191
rect 22603 7157 22612 7191
rect 22560 7148 22612 7157
rect 23388 7191 23440 7200
rect 23388 7157 23397 7191
rect 23397 7157 23431 7191
rect 23431 7157 23440 7191
rect 23388 7148 23440 7157
rect 25412 7191 25464 7200
rect 25412 7157 25421 7191
rect 25421 7157 25455 7191
rect 25455 7157 25464 7191
rect 25412 7148 25464 7157
rect 27068 7191 27120 7200
rect 27068 7157 27077 7191
rect 27077 7157 27111 7191
rect 27111 7157 27120 7191
rect 27528 7191 27580 7200
rect 27068 7148 27120 7157
rect 27528 7157 27537 7191
rect 27537 7157 27571 7191
rect 27571 7157 27580 7191
rect 27528 7148 27580 7157
rect 27988 7148 28040 7200
rect 31392 7191 31444 7200
rect 31392 7157 31401 7191
rect 31401 7157 31435 7191
rect 31435 7157 31444 7191
rect 31392 7148 31444 7157
rect 33140 7148 33192 7200
rect 35072 7191 35124 7200
rect 35072 7157 35081 7191
rect 35081 7157 35115 7191
rect 35115 7157 35124 7191
rect 35072 7148 35124 7157
rect 14315 7046 14367 7098
rect 14379 7046 14431 7098
rect 14443 7046 14495 7098
rect 14507 7046 14559 7098
rect 27648 7046 27700 7098
rect 27712 7046 27764 7098
rect 27776 7046 27828 7098
rect 27840 7046 27892 7098
rect 2596 6987 2648 6996
rect 2596 6953 2605 6987
rect 2605 6953 2639 6987
rect 2639 6953 2648 6987
rect 2596 6944 2648 6953
rect 4252 6987 4304 6996
rect 4252 6953 4261 6987
rect 4261 6953 4295 6987
rect 4295 6953 4304 6987
rect 4252 6944 4304 6953
rect 5080 6987 5132 6996
rect 5080 6953 5089 6987
rect 5089 6953 5123 6987
rect 5123 6953 5132 6987
rect 5080 6944 5132 6953
rect 7472 6944 7524 6996
rect 8116 6987 8168 6996
rect 8116 6953 8125 6987
rect 8125 6953 8159 6987
rect 8159 6953 8168 6987
rect 8116 6944 8168 6953
rect 11244 6987 11296 6996
rect 11244 6953 11253 6987
rect 11253 6953 11287 6987
rect 11287 6953 11296 6987
rect 11244 6944 11296 6953
rect 13176 6944 13228 6996
rect 14832 6944 14884 6996
rect 17132 6944 17184 6996
rect 19800 6987 19852 6996
rect 19800 6953 19809 6987
rect 19809 6953 19843 6987
rect 19843 6953 19852 6987
rect 19800 6944 19852 6953
rect 2136 6919 2188 6928
rect 2136 6885 2145 6919
rect 2145 6885 2179 6919
rect 2179 6885 2188 6919
rect 2136 6876 2188 6885
rect 1860 6808 1912 6860
rect 2228 6783 2280 6792
rect 2228 6749 2237 6783
rect 2237 6749 2271 6783
rect 2271 6749 2280 6783
rect 2228 6740 2280 6749
rect 3516 6740 3568 6792
rect 5356 6876 5408 6928
rect 5172 6808 5224 6860
rect 6644 6808 6696 6860
rect 7012 6808 7064 6860
rect 7380 6808 7432 6860
rect 9312 6808 9364 6860
rect 10508 6876 10560 6928
rect 11060 6876 11112 6928
rect 11888 6876 11940 6928
rect 12532 6876 12584 6928
rect 13268 6919 13320 6928
rect 13268 6885 13277 6919
rect 13277 6885 13311 6919
rect 13311 6885 13320 6919
rect 13268 6876 13320 6885
rect 11336 6851 11388 6860
rect 11336 6817 11345 6851
rect 11345 6817 11379 6851
rect 11379 6817 11388 6851
rect 11336 6808 11388 6817
rect 11428 6808 11480 6860
rect 13820 6851 13872 6860
rect 13820 6817 13829 6851
rect 13829 6817 13863 6851
rect 13863 6817 13872 6851
rect 13820 6808 13872 6817
rect 16672 6876 16724 6928
rect 17868 6876 17920 6928
rect 16856 6808 16908 6860
rect 18696 6808 18748 6860
rect 20904 6876 20956 6928
rect 21272 6876 21324 6928
rect 25504 6987 25556 6996
rect 25504 6953 25513 6987
rect 25513 6953 25547 6987
rect 25547 6953 25556 6987
rect 25504 6944 25556 6953
rect 27160 6944 27212 6996
rect 29184 6944 29236 6996
rect 21548 6919 21600 6928
rect 21548 6885 21557 6919
rect 21557 6885 21591 6919
rect 21591 6885 21600 6919
rect 21548 6876 21600 6885
rect 23112 6919 23164 6928
rect 23112 6885 23121 6919
rect 23121 6885 23155 6919
rect 23155 6885 23164 6919
rect 23112 6876 23164 6885
rect 24676 6919 24728 6928
rect 24676 6885 24685 6919
rect 24685 6885 24719 6919
rect 24719 6885 24728 6919
rect 24676 6876 24728 6885
rect 4160 6740 4212 6792
rect 5448 6740 5500 6792
rect 7472 6783 7524 6792
rect 1676 6715 1728 6724
rect 1676 6681 1685 6715
rect 1685 6681 1719 6715
rect 1719 6681 1728 6715
rect 1676 6672 1728 6681
rect 2964 6672 3016 6724
rect 4344 6672 4396 6724
rect 5724 6672 5776 6724
rect 4712 6604 4764 6656
rect 5356 6604 5408 6656
rect 7472 6749 7481 6783
rect 7481 6749 7515 6783
rect 7515 6749 7524 6783
rect 7472 6740 7524 6749
rect 8576 6783 8628 6792
rect 8576 6749 8585 6783
rect 8585 6749 8619 6783
rect 8619 6749 8628 6783
rect 8576 6740 8628 6749
rect 9680 6740 9732 6792
rect 10324 6783 10376 6792
rect 6828 6672 6880 6724
rect 10324 6749 10333 6783
rect 10333 6749 10367 6783
rect 10367 6749 10376 6783
rect 10324 6740 10376 6749
rect 16764 6783 16816 6792
rect 16764 6749 16773 6783
rect 16773 6749 16807 6783
rect 16807 6749 16816 6783
rect 16764 6740 16816 6749
rect 21640 6783 21692 6792
rect 21640 6749 21649 6783
rect 21649 6749 21683 6783
rect 21683 6749 21692 6783
rect 22744 6808 22796 6860
rect 23848 6808 23900 6860
rect 25412 6876 25464 6928
rect 25688 6876 25740 6928
rect 28908 6876 28960 6928
rect 26608 6808 26660 6860
rect 21640 6740 21692 6749
rect 11152 6672 11204 6724
rect 21364 6672 21416 6724
rect 22560 6672 22612 6724
rect 23388 6740 23440 6792
rect 24124 6740 24176 6792
rect 26700 6783 26752 6792
rect 26700 6749 26709 6783
rect 26709 6749 26743 6783
rect 26743 6749 26752 6783
rect 26700 6740 26752 6749
rect 23480 6672 23532 6724
rect 24032 6715 24084 6724
rect 24032 6681 24041 6715
rect 24041 6681 24075 6715
rect 24075 6681 24084 6715
rect 24032 6672 24084 6681
rect 24676 6672 24728 6724
rect 29920 6808 29972 6860
rect 31484 6944 31536 6996
rect 33968 6987 34020 6996
rect 33968 6953 33977 6987
rect 33977 6953 34011 6987
rect 34011 6953 34020 6987
rect 33968 6944 34020 6953
rect 31760 6808 31812 6860
rect 32680 6919 32732 6928
rect 32680 6885 32689 6919
rect 32689 6885 32723 6919
rect 32723 6885 32732 6919
rect 32680 6876 32732 6885
rect 35716 6944 35768 6996
rect 34520 6876 34572 6928
rect 34980 6876 35032 6928
rect 34796 6851 34848 6860
rect 34796 6817 34819 6851
rect 34819 6817 34848 6851
rect 34796 6808 34848 6817
rect 36268 6808 36320 6860
rect 29000 6740 29052 6792
rect 30748 6740 30800 6792
rect 32404 6740 32456 6792
rect 34520 6783 34572 6792
rect 34520 6749 34529 6783
rect 34529 6749 34563 6783
rect 34563 6749 34572 6783
rect 34520 6740 34572 6749
rect 6184 6604 6236 6656
rect 7104 6647 7156 6656
rect 7104 6613 7113 6647
rect 7113 6613 7147 6647
rect 7147 6613 7156 6647
rect 7104 6604 7156 6613
rect 9496 6647 9548 6656
rect 9496 6613 9505 6647
rect 9505 6613 9539 6647
rect 9539 6613 9548 6647
rect 9496 6604 9548 6613
rect 9772 6647 9824 6656
rect 9772 6613 9781 6647
rect 9781 6613 9815 6647
rect 9815 6613 9824 6647
rect 9772 6604 9824 6613
rect 11704 6604 11756 6656
rect 18512 6604 18564 6656
rect 18880 6604 18932 6656
rect 20260 6604 20312 6656
rect 20536 6604 20588 6656
rect 21548 6604 21600 6656
rect 21916 6604 21968 6656
rect 22100 6647 22152 6656
rect 22100 6613 22109 6647
rect 22109 6613 22143 6647
rect 22143 6613 22152 6647
rect 22100 6604 22152 6613
rect 24216 6647 24268 6656
rect 24216 6613 24225 6647
rect 24225 6613 24259 6647
rect 24259 6613 24268 6647
rect 24216 6604 24268 6613
rect 24952 6604 25004 6656
rect 25964 6647 26016 6656
rect 25964 6613 25973 6647
rect 25973 6613 26007 6647
rect 26007 6613 26016 6647
rect 25964 6604 26016 6613
rect 32036 6672 32088 6724
rect 33784 6672 33836 6724
rect 28816 6604 28868 6656
rect 31484 6647 31536 6656
rect 31484 6613 31493 6647
rect 31493 6613 31527 6647
rect 31527 6613 31536 6647
rect 31484 6604 31536 6613
rect 33140 6604 33192 6656
rect 33692 6647 33744 6656
rect 33692 6613 33701 6647
rect 33701 6613 33735 6647
rect 33735 6613 33744 6647
rect 33692 6604 33744 6613
rect 36452 6647 36504 6656
rect 36452 6613 36461 6647
rect 36461 6613 36495 6647
rect 36495 6613 36504 6647
rect 36452 6604 36504 6613
rect 7648 6502 7700 6554
rect 7712 6502 7764 6554
rect 7776 6502 7828 6554
rect 7840 6502 7892 6554
rect 20982 6502 21034 6554
rect 21046 6502 21098 6554
rect 21110 6502 21162 6554
rect 21174 6502 21226 6554
rect 34315 6502 34367 6554
rect 34379 6502 34431 6554
rect 34443 6502 34495 6554
rect 34507 6502 34559 6554
rect 2872 6400 2924 6452
rect 4160 6443 4212 6452
rect 4160 6409 4169 6443
rect 4169 6409 4203 6443
rect 4203 6409 4212 6443
rect 4160 6400 4212 6409
rect 6828 6400 6880 6452
rect 5356 6264 5408 6316
rect 8116 6400 8168 6452
rect 11336 6443 11388 6452
rect 11336 6409 11345 6443
rect 11345 6409 11379 6443
rect 11379 6409 11388 6443
rect 11336 6400 11388 6409
rect 11796 6443 11848 6452
rect 11796 6409 11805 6443
rect 11805 6409 11839 6443
rect 11839 6409 11848 6443
rect 11796 6400 11848 6409
rect 12164 6443 12216 6452
rect 12164 6409 12173 6443
rect 12173 6409 12207 6443
rect 12207 6409 12216 6443
rect 12164 6400 12216 6409
rect 17776 6443 17828 6452
rect 17776 6409 17785 6443
rect 17785 6409 17819 6443
rect 17819 6409 17828 6443
rect 17776 6400 17828 6409
rect 18696 6443 18748 6452
rect 18696 6409 18705 6443
rect 18705 6409 18739 6443
rect 18739 6409 18748 6443
rect 18696 6400 18748 6409
rect 19340 6443 19392 6452
rect 19340 6409 19349 6443
rect 19349 6409 19383 6443
rect 19383 6409 19392 6443
rect 19340 6400 19392 6409
rect 19616 6443 19668 6452
rect 19616 6409 19625 6443
rect 19625 6409 19659 6443
rect 19659 6409 19668 6443
rect 19616 6400 19668 6409
rect 20812 6400 20864 6452
rect 21272 6400 21324 6452
rect 22468 6443 22520 6452
rect 22468 6409 22477 6443
rect 22477 6409 22511 6443
rect 22511 6409 22520 6443
rect 22468 6400 22520 6409
rect 23112 6443 23164 6452
rect 23112 6409 23121 6443
rect 23121 6409 23155 6443
rect 23155 6409 23164 6443
rect 23112 6400 23164 6409
rect 23480 6443 23532 6452
rect 23480 6409 23489 6443
rect 23489 6409 23523 6443
rect 23523 6409 23532 6443
rect 23480 6400 23532 6409
rect 23940 6400 23992 6452
rect 24492 6443 24544 6452
rect 24492 6409 24501 6443
rect 24501 6409 24535 6443
rect 24535 6409 24544 6443
rect 24492 6400 24544 6409
rect 25780 6443 25832 6452
rect 25780 6409 25789 6443
rect 25789 6409 25823 6443
rect 25823 6409 25832 6443
rect 25780 6400 25832 6409
rect 26424 6400 26476 6452
rect 27068 6443 27120 6452
rect 27068 6409 27077 6443
rect 27077 6409 27111 6443
rect 27111 6409 27120 6443
rect 27068 6400 27120 6409
rect 27344 6443 27396 6452
rect 27344 6409 27353 6443
rect 27353 6409 27387 6443
rect 27387 6409 27396 6443
rect 27344 6400 27396 6409
rect 29000 6400 29052 6452
rect 29920 6443 29972 6452
rect 9956 6375 10008 6384
rect 9956 6341 9965 6375
rect 9965 6341 9999 6375
rect 9999 6341 10008 6375
rect 9956 6332 10008 6341
rect 12440 6332 12492 6384
rect 15568 6332 15620 6384
rect 16764 6332 16816 6384
rect 17684 6332 17736 6384
rect 26332 6332 26384 6384
rect 20168 6307 20220 6316
rect 20168 6273 20177 6307
rect 20177 6273 20211 6307
rect 20211 6273 20220 6307
rect 20168 6264 20220 6273
rect 25136 6264 25188 6316
rect 29552 6332 29604 6384
rect 29920 6409 29929 6443
rect 29929 6409 29963 6443
rect 29963 6409 29972 6443
rect 29920 6400 29972 6409
rect 32404 6443 32456 6452
rect 32404 6409 32413 6443
rect 32413 6409 32447 6443
rect 32447 6409 32456 6443
rect 32404 6400 32456 6409
rect 33140 6400 33192 6452
rect 36268 6443 36320 6452
rect 36268 6409 36277 6443
rect 36277 6409 36311 6443
rect 36311 6409 36320 6443
rect 36268 6400 36320 6409
rect 37648 6400 37700 6452
rect 33692 6332 33744 6384
rect 33784 6307 33836 6316
rect 33784 6273 33793 6307
rect 33793 6273 33827 6307
rect 33827 6273 33836 6307
rect 33784 6264 33836 6273
rect 1492 6196 1544 6248
rect 2964 6196 3016 6248
rect 9680 6239 9732 6248
rect 9680 6205 9689 6239
rect 9689 6205 9723 6239
rect 9723 6205 9732 6239
rect 9680 6196 9732 6205
rect 10324 6196 10376 6248
rect 11796 6196 11848 6248
rect 12992 6196 13044 6248
rect 13544 6196 13596 6248
rect 15568 6196 15620 6248
rect 18972 6239 19024 6248
rect 18972 6205 18981 6239
rect 18981 6205 19015 6239
rect 19015 6205 19024 6239
rect 18972 6196 19024 6205
rect 19800 6196 19852 6248
rect 21088 6239 21140 6248
rect 21088 6205 21097 6239
rect 21097 6205 21131 6239
rect 21131 6205 21140 6239
rect 21088 6196 21140 6205
rect 21640 6196 21692 6248
rect 30748 6239 30800 6248
rect 30748 6205 30782 6239
rect 30782 6205 30800 6239
rect 30748 6196 30800 6205
rect 34980 6196 35032 6248
rect 37372 6239 37424 6248
rect 37372 6205 37381 6239
rect 37381 6205 37415 6239
rect 37415 6205 37424 6239
rect 37372 6196 37424 6205
rect 2228 6128 2280 6180
rect 4620 6128 4672 6180
rect 7656 6171 7708 6180
rect 7656 6137 7690 6171
rect 7690 6137 7708 6171
rect 7656 6128 7708 6137
rect 9496 6128 9548 6180
rect 10508 6171 10560 6180
rect 10508 6137 10517 6171
rect 10517 6137 10551 6171
rect 10551 6137 10560 6171
rect 10508 6128 10560 6137
rect 14832 6128 14884 6180
rect 5540 6060 5592 6112
rect 6184 6103 6236 6112
rect 6184 6069 6193 6103
rect 6193 6069 6227 6103
rect 6227 6069 6236 6103
rect 6184 6060 6236 6069
rect 8392 6060 8444 6112
rect 9312 6103 9364 6112
rect 9312 6069 9321 6103
rect 9321 6069 9355 6103
rect 9355 6069 9364 6103
rect 9312 6060 9364 6069
rect 9772 6060 9824 6112
rect 12164 6060 12216 6112
rect 15752 6103 15804 6112
rect 15752 6069 15761 6103
rect 15761 6069 15795 6103
rect 15795 6069 15804 6103
rect 15752 6060 15804 6069
rect 16856 6060 16908 6112
rect 18512 6060 18564 6112
rect 19524 6060 19576 6112
rect 20536 6103 20588 6112
rect 20536 6069 20545 6103
rect 20545 6069 20579 6103
rect 20579 6069 20588 6103
rect 24124 6103 24176 6112
rect 20536 6060 20588 6069
rect 24124 6069 24133 6103
rect 24133 6069 24167 6103
rect 24167 6069 24176 6103
rect 24124 6060 24176 6069
rect 24768 6128 24820 6180
rect 26608 6171 26660 6180
rect 26608 6137 26617 6171
rect 26617 6137 26651 6171
rect 26651 6137 26660 6171
rect 26608 6128 26660 6137
rect 24952 6103 25004 6112
rect 24952 6069 24961 6103
rect 24961 6069 24995 6103
rect 24995 6069 25004 6103
rect 24952 6060 25004 6069
rect 25964 6060 26016 6112
rect 27528 6128 27580 6180
rect 28264 6128 28316 6180
rect 29828 6128 29880 6180
rect 30288 6128 30340 6180
rect 35164 6171 35216 6180
rect 35164 6137 35198 6171
rect 35198 6137 35216 6171
rect 35164 6128 35216 6137
rect 27344 6060 27396 6112
rect 14315 5958 14367 6010
rect 14379 5958 14431 6010
rect 14443 5958 14495 6010
rect 14507 5958 14559 6010
rect 27648 5958 27700 6010
rect 27712 5958 27764 6010
rect 27776 5958 27828 6010
rect 27840 5958 27892 6010
rect 2872 5899 2924 5908
rect 2872 5865 2881 5899
rect 2881 5865 2915 5899
rect 2915 5865 2924 5899
rect 4620 5899 4672 5908
rect 2872 5856 2924 5865
rect 4620 5865 4629 5899
rect 4629 5865 4663 5899
rect 4663 5865 4672 5899
rect 4620 5856 4672 5865
rect 5172 5899 5224 5908
rect 5172 5865 5181 5899
rect 5181 5865 5215 5899
rect 5215 5865 5224 5899
rect 5172 5856 5224 5865
rect 7380 5856 7432 5908
rect 7656 5899 7708 5908
rect 7656 5865 7665 5899
rect 7665 5865 7699 5899
rect 7699 5865 7708 5899
rect 7656 5856 7708 5865
rect 9772 5856 9824 5908
rect 10508 5856 10560 5908
rect 11428 5899 11480 5908
rect 11428 5865 11437 5899
rect 11437 5865 11471 5899
rect 11471 5865 11480 5899
rect 11428 5856 11480 5865
rect 17960 5856 18012 5908
rect 19064 5856 19116 5908
rect 19524 5899 19576 5908
rect 19524 5865 19533 5899
rect 19533 5865 19567 5899
rect 19567 5865 19576 5899
rect 19524 5856 19576 5865
rect 21640 5856 21692 5908
rect 23388 5899 23440 5908
rect 23388 5865 23397 5899
rect 23397 5865 23431 5899
rect 23431 5865 23440 5899
rect 23388 5856 23440 5865
rect 23848 5899 23900 5908
rect 23848 5865 23857 5899
rect 23857 5865 23891 5899
rect 23891 5865 23900 5899
rect 23848 5856 23900 5865
rect 29644 5856 29696 5908
rect 30748 5856 30800 5908
rect 31760 5856 31812 5908
rect 32680 5856 32732 5908
rect 33692 5856 33744 5908
rect 1860 5788 1912 5840
rect 7104 5788 7156 5840
rect 8392 5831 8444 5840
rect 8392 5797 8401 5831
rect 8401 5797 8435 5831
rect 8435 5797 8444 5831
rect 8392 5788 8444 5797
rect 8576 5788 8628 5840
rect 9864 5788 9916 5840
rect 10600 5788 10652 5840
rect 12532 5788 12584 5840
rect 14740 5788 14792 5840
rect 18144 5788 18196 5840
rect 1492 5763 1544 5772
rect 1492 5729 1501 5763
rect 1501 5729 1535 5763
rect 1535 5729 1544 5763
rect 1492 5720 1544 5729
rect 2780 5720 2832 5772
rect 3516 5763 3568 5772
rect 3516 5729 3525 5763
rect 3525 5729 3559 5763
rect 3559 5729 3568 5763
rect 3516 5720 3568 5729
rect 5356 5720 5408 5772
rect 5540 5763 5592 5772
rect 5540 5729 5574 5763
rect 5574 5729 5592 5763
rect 5540 5720 5592 5729
rect 12348 5720 12400 5772
rect 12808 5720 12860 5772
rect 15752 5763 15804 5772
rect 3976 5652 4028 5704
rect 8208 5695 8260 5704
rect 8208 5661 8217 5695
rect 8217 5661 8251 5695
rect 8251 5661 8260 5695
rect 8208 5652 8260 5661
rect 10324 5695 10376 5704
rect 10324 5661 10333 5695
rect 10333 5661 10367 5695
rect 10367 5661 10376 5695
rect 10324 5652 10376 5661
rect 12716 5695 12768 5704
rect 12716 5661 12725 5695
rect 12725 5661 12759 5695
rect 12759 5661 12768 5695
rect 12716 5652 12768 5661
rect 4068 5584 4120 5636
rect 7196 5584 7248 5636
rect 9496 5584 9548 5636
rect 14188 5652 14240 5704
rect 15752 5729 15775 5763
rect 15775 5729 15804 5763
rect 20168 5788 20220 5840
rect 21824 5788 21876 5840
rect 22468 5788 22520 5840
rect 27804 5788 27856 5840
rect 28540 5788 28592 5840
rect 29552 5831 29604 5840
rect 29552 5797 29561 5831
rect 29561 5797 29595 5831
rect 29595 5797 29604 5831
rect 29552 5788 29604 5797
rect 30380 5788 30432 5840
rect 33416 5788 33468 5840
rect 34244 5788 34296 5840
rect 35164 5856 35216 5908
rect 36084 5899 36136 5908
rect 36084 5865 36093 5899
rect 36093 5865 36127 5899
rect 36127 5865 36136 5899
rect 36084 5856 36136 5865
rect 15752 5720 15804 5729
rect 19340 5720 19392 5772
rect 24216 5763 24268 5772
rect 24216 5729 24250 5763
rect 24250 5729 24268 5763
rect 24216 5720 24268 5729
rect 28356 5720 28408 5772
rect 33232 5720 33284 5772
rect 15476 5695 15528 5704
rect 15476 5661 15485 5695
rect 15485 5661 15519 5695
rect 15519 5661 15528 5695
rect 15476 5652 15528 5661
rect 21088 5652 21140 5704
rect 21456 5695 21508 5704
rect 21456 5661 21465 5695
rect 21465 5661 21499 5695
rect 21499 5661 21508 5695
rect 21456 5652 21508 5661
rect 23940 5695 23992 5704
rect 23940 5661 23949 5695
rect 23949 5661 23983 5695
rect 23983 5661 23992 5695
rect 23940 5652 23992 5661
rect 26332 5652 26384 5704
rect 28264 5695 28316 5704
rect 17868 5584 17920 5636
rect 11060 5516 11112 5568
rect 11704 5559 11756 5568
rect 11704 5525 11713 5559
rect 11713 5525 11747 5559
rect 11747 5525 11756 5559
rect 11704 5516 11756 5525
rect 13728 5559 13780 5568
rect 13728 5525 13737 5559
rect 13737 5525 13771 5559
rect 13771 5525 13780 5559
rect 13728 5516 13780 5525
rect 16856 5559 16908 5568
rect 16856 5525 16865 5559
rect 16865 5525 16899 5559
rect 16899 5525 16908 5559
rect 16856 5516 16908 5525
rect 18880 5516 18932 5568
rect 19984 5516 20036 5568
rect 26608 5584 26660 5636
rect 28264 5661 28273 5695
rect 28273 5661 28307 5695
rect 28307 5661 28316 5695
rect 28264 5652 28316 5661
rect 29276 5652 29328 5704
rect 33324 5695 33376 5704
rect 33324 5661 33333 5695
rect 33333 5661 33367 5695
rect 33367 5661 33376 5695
rect 33324 5652 33376 5661
rect 34428 5720 34480 5772
rect 34612 5652 34664 5704
rect 35716 5720 35768 5772
rect 35900 5763 35952 5772
rect 35900 5729 35909 5763
rect 35909 5729 35943 5763
rect 35943 5729 35952 5763
rect 35900 5720 35952 5729
rect 34980 5652 35032 5704
rect 28816 5584 28868 5636
rect 32772 5584 32824 5636
rect 34060 5584 34112 5636
rect 22836 5559 22888 5568
rect 22836 5525 22845 5559
rect 22845 5525 22879 5559
rect 22879 5525 22888 5559
rect 22836 5516 22888 5525
rect 25688 5516 25740 5568
rect 26700 5559 26752 5568
rect 26700 5525 26709 5559
rect 26709 5525 26743 5559
rect 26743 5525 26752 5559
rect 26700 5516 26752 5525
rect 27160 5559 27212 5568
rect 27160 5525 27169 5559
rect 27169 5525 27203 5559
rect 27203 5525 27212 5559
rect 27160 5516 27212 5525
rect 29828 5516 29880 5568
rect 7648 5414 7700 5466
rect 7712 5414 7764 5466
rect 7776 5414 7828 5466
rect 7840 5414 7892 5466
rect 20982 5414 21034 5466
rect 21046 5414 21098 5466
rect 21110 5414 21162 5466
rect 21174 5414 21226 5466
rect 34315 5414 34367 5466
rect 34379 5414 34431 5466
rect 34443 5414 34495 5466
rect 34507 5414 34559 5466
rect 2596 5312 2648 5364
rect 2964 5312 3016 5364
rect 4068 5312 4120 5364
rect 5356 5355 5408 5364
rect 5356 5321 5365 5355
rect 5365 5321 5399 5355
rect 5399 5321 5408 5355
rect 5356 5312 5408 5321
rect 7012 5355 7064 5364
rect 7012 5321 7021 5355
rect 7021 5321 7055 5355
rect 7055 5321 7064 5355
rect 7012 5312 7064 5321
rect 7104 5312 7156 5364
rect 8116 5312 8168 5364
rect 2504 5176 2556 5228
rect 3332 5244 3384 5296
rect 2872 5176 2924 5228
rect 3884 5176 3936 5228
rect 5540 5176 5592 5228
rect 10324 5312 10376 5364
rect 12716 5312 12768 5364
rect 14832 5312 14884 5364
rect 15568 5355 15620 5364
rect 15568 5321 15577 5355
rect 15577 5321 15611 5355
rect 15611 5321 15620 5355
rect 15568 5312 15620 5321
rect 17132 5355 17184 5364
rect 17132 5321 17141 5355
rect 17141 5321 17175 5355
rect 17175 5321 17184 5355
rect 17132 5312 17184 5321
rect 18328 5312 18380 5364
rect 19064 5355 19116 5364
rect 19064 5321 19073 5355
rect 19073 5321 19107 5355
rect 19107 5321 19116 5355
rect 19064 5312 19116 5321
rect 19340 5312 19392 5364
rect 20260 5355 20312 5364
rect 20260 5321 20269 5355
rect 20269 5321 20303 5355
rect 20303 5321 20312 5355
rect 20260 5312 20312 5321
rect 21456 5312 21508 5364
rect 22100 5312 22152 5364
rect 23940 5355 23992 5364
rect 23940 5321 23949 5355
rect 23949 5321 23983 5355
rect 23983 5321 23992 5355
rect 23940 5312 23992 5321
rect 24768 5355 24820 5364
rect 24768 5321 24777 5355
rect 24777 5321 24811 5355
rect 24811 5321 24820 5355
rect 24768 5312 24820 5321
rect 14648 5244 14700 5296
rect 16120 5176 16172 5228
rect 22376 5244 22428 5296
rect 26700 5312 26752 5364
rect 27160 5312 27212 5364
rect 27804 5312 27856 5364
rect 28356 5312 28408 5364
rect 29368 5355 29420 5364
rect 29368 5321 29377 5355
rect 29377 5321 29411 5355
rect 29411 5321 29420 5355
rect 29368 5312 29420 5321
rect 30380 5355 30432 5364
rect 30380 5321 30389 5355
rect 30389 5321 30423 5355
rect 30423 5321 30432 5355
rect 30380 5312 30432 5321
rect 33048 5312 33100 5364
rect 34152 5312 34204 5364
rect 34704 5355 34756 5364
rect 34704 5321 34713 5355
rect 34713 5321 34747 5355
rect 34747 5321 34756 5355
rect 34704 5312 34756 5321
rect 36636 5355 36688 5364
rect 36636 5321 36645 5355
rect 36645 5321 36679 5355
rect 36679 5321 36688 5355
rect 36636 5312 36688 5321
rect 16580 5219 16632 5228
rect 16580 5185 16589 5219
rect 16589 5185 16623 5219
rect 16623 5185 16632 5219
rect 16580 5176 16632 5185
rect 21824 5219 21876 5228
rect 21824 5185 21833 5219
rect 21833 5185 21867 5219
rect 21867 5185 21876 5219
rect 21824 5176 21876 5185
rect 29276 5244 29328 5296
rect 32588 5244 32640 5296
rect 34612 5244 34664 5296
rect 34980 5287 35032 5296
rect 34980 5253 34989 5287
rect 34989 5253 35023 5287
rect 35023 5253 35032 5287
rect 34980 5244 35032 5253
rect 29920 5219 29972 5228
rect 29920 5185 29929 5219
rect 29929 5185 29963 5219
rect 29963 5185 29972 5219
rect 29920 5176 29972 5185
rect 32772 5176 32824 5228
rect 32864 5176 32916 5228
rect 33232 5219 33284 5228
rect 33232 5185 33241 5219
rect 33241 5185 33275 5219
rect 33275 5185 33284 5219
rect 33232 5176 33284 5185
rect 35164 5176 35216 5228
rect 13544 5108 13596 5160
rect 25688 5108 25740 5160
rect 28264 5108 28316 5160
rect 29552 5108 29604 5160
rect 33416 5108 33468 5160
rect 34888 5108 34940 5160
rect 2596 5083 2648 5092
rect 2596 5049 2605 5083
rect 2605 5049 2639 5083
rect 2639 5049 2648 5083
rect 2596 5040 2648 5049
rect 2964 5040 3016 5092
rect 3148 5040 3200 5092
rect 3424 5040 3476 5092
rect 4160 5083 4212 5092
rect 4160 5049 4169 5083
rect 4169 5049 4203 5083
rect 4203 5049 4212 5083
rect 4160 5040 4212 5049
rect 8484 5040 8536 5092
rect 12256 5040 12308 5092
rect 12992 5040 13044 5092
rect 4068 4972 4120 5024
rect 4712 5015 4764 5024
rect 4712 4981 4721 5015
rect 4721 4981 4755 5015
rect 4755 4981 4764 5015
rect 4712 4972 4764 4981
rect 9772 5015 9824 5024
rect 9772 4981 9781 5015
rect 9781 4981 9815 5015
rect 9815 4981 9824 5015
rect 9772 4972 9824 4981
rect 10600 4972 10652 5024
rect 11980 4972 12032 5024
rect 12348 4972 12400 5024
rect 13544 4972 13596 5024
rect 14188 4972 14240 5024
rect 18052 5040 18104 5092
rect 18512 5040 18564 5092
rect 19156 5040 19208 5092
rect 20260 5040 20312 5092
rect 21732 5083 21784 5092
rect 21732 5049 21741 5083
rect 21741 5049 21775 5083
rect 21775 5049 21784 5083
rect 21732 5040 21784 5049
rect 22836 5040 22888 5092
rect 24216 5040 24268 5092
rect 29828 5083 29880 5092
rect 29828 5049 29837 5083
rect 29837 5049 29871 5083
rect 29871 5049 29880 5083
rect 29828 5040 29880 5049
rect 33048 5040 33100 5092
rect 14740 5015 14792 5024
rect 14740 4981 14749 5015
rect 14749 4981 14783 5015
rect 14783 4981 14792 5015
rect 14740 4972 14792 4981
rect 16488 5015 16540 5024
rect 16488 4981 16497 5015
rect 16497 4981 16531 5015
rect 16531 4981 16540 5015
rect 16488 4972 16540 4981
rect 17500 5015 17552 5024
rect 17500 4981 17509 5015
rect 17509 4981 17543 5015
rect 17543 4981 17552 5015
rect 17500 4972 17552 4981
rect 18328 4972 18380 5024
rect 29184 4972 29236 5024
rect 34704 4972 34756 5024
rect 35900 5015 35952 5024
rect 35900 4981 35909 5015
rect 35909 4981 35943 5015
rect 35943 4981 35952 5015
rect 35900 4972 35952 4981
rect 14315 4870 14367 4922
rect 14379 4870 14431 4922
rect 14443 4870 14495 4922
rect 14507 4870 14559 4922
rect 27648 4870 27700 4922
rect 27712 4870 27764 4922
rect 27776 4870 27828 4922
rect 27840 4870 27892 4922
rect 1400 4768 1452 4820
rect 2412 4768 2464 4820
rect 2872 4768 2924 4820
rect 3884 4811 3936 4820
rect 3884 4777 3893 4811
rect 3893 4777 3927 4811
rect 3927 4777 3936 4811
rect 3884 4768 3936 4777
rect 4160 4768 4212 4820
rect 8208 4768 8260 4820
rect 8392 4768 8444 4820
rect 9864 4811 9916 4820
rect 9864 4777 9873 4811
rect 9873 4777 9907 4811
rect 9907 4777 9916 4811
rect 9864 4768 9916 4777
rect 12716 4768 12768 4820
rect 12992 4811 13044 4820
rect 12992 4777 13001 4811
rect 13001 4777 13035 4811
rect 13035 4777 13044 4811
rect 12992 4768 13044 4777
rect 13820 4768 13872 4820
rect 14648 4811 14700 4820
rect 14648 4777 14657 4811
rect 14657 4777 14691 4811
rect 14691 4777 14700 4811
rect 14648 4768 14700 4777
rect 16580 4768 16632 4820
rect 18052 4811 18104 4820
rect 18052 4777 18061 4811
rect 18061 4777 18095 4811
rect 18095 4777 18104 4811
rect 18052 4768 18104 4777
rect 18972 4811 19024 4820
rect 18972 4777 18981 4811
rect 18981 4777 19015 4811
rect 19015 4777 19024 4811
rect 18972 4768 19024 4777
rect 21824 4768 21876 4820
rect 22100 4768 22152 4820
rect 25688 4811 25740 4820
rect 25688 4777 25697 4811
rect 25697 4777 25731 4811
rect 25731 4777 25740 4811
rect 25688 4768 25740 4777
rect 2780 4700 2832 4752
rect 8116 4743 8168 4752
rect 8116 4709 8125 4743
rect 8125 4709 8159 4743
rect 8159 4709 8168 4743
rect 8116 4700 8168 4709
rect 10968 4743 11020 4752
rect 10968 4709 10977 4743
rect 10977 4709 11011 4743
rect 11011 4709 11020 4743
rect 10968 4700 11020 4709
rect 14004 4700 14056 4752
rect 15568 4700 15620 4752
rect 17132 4700 17184 4752
rect 18788 4743 18840 4752
rect 18788 4709 18797 4743
rect 18797 4709 18831 4743
rect 18831 4709 18840 4743
rect 18788 4700 18840 4709
rect 22376 4743 22428 4752
rect 22376 4709 22385 4743
rect 22385 4709 22419 4743
rect 22419 4709 22428 4743
rect 22376 4700 22428 4709
rect 27712 4700 27764 4752
rect 28080 4743 28132 4752
rect 28080 4709 28089 4743
rect 28089 4709 28123 4743
rect 28123 4709 28132 4743
rect 28080 4700 28132 4709
rect 28264 4768 28316 4820
rect 29644 4811 29696 4820
rect 29644 4777 29653 4811
rect 29653 4777 29687 4811
rect 29687 4777 29696 4811
rect 29644 4768 29696 4777
rect 29828 4768 29880 4820
rect 32772 4811 32824 4820
rect 32772 4777 32781 4811
rect 32781 4777 32815 4811
rect 32815 4777 32824 4811
rect 32772 4768 32824 4777
rect 32956 4811 33008 4820
rect 32956 4777 32965 4811
rect 32965 4777 32999 4811
rect 32999 4777 33008 4811
rect 32956 4768 33008 4777
rect 33324 4768 33376 4820
rect 34980 4768 35032 4820
rect 35164 4768 35216 4820
rect 35532 4768 35584 4820
rect 29920 4700 29972 4752
rect 32864 4700 32916 4752
rect 34060 4700 34112 4752
rect 34796 4700 34848 4752
rect 1400 4675 1452 4684
rect 1400 4641 1409 4675
rect 1409 4641 1443 4675
rect 1443 4641 1452 4675
rect 1400 4632 1452 4641
rect 2504 4675 2556 4684
rect 2504 4641 2513 4675
rect 2513 4641 2547 4675
rect 2547 4641 2556 4675
rect 2504 4632 2556 4641
rect 5540 4632 5592 4684
rect 8300 4632 8352 4684
rect 15660 4675 15712 4684
rect 15660 4641 15669 4675
rect 15669 4641 15703 4675
rect 15703 4641 15712 4675
rect 15660 4632 15712 4641
rect 15752 4632 15804 4684
rect 17224 4675 17276 4684
rect 17224 4641 17233 4675
rect 17233 4641 17267 4675
rect 17267 4641 17276 4675
rect 17224 4632 17276 4641
rect 27436 4632 27488 4684
rect 27896 4675 27948 4684
rect 27896 4641 27905 4675
rect 27905 4641 27939 4675
rect 27939 4641 27948 4675
rect 27896 4632 27948 4641
rect 34888 4632 34940 4684
rect 35440 4632 35492 4684
rect 7380 4564 7432 4616
rect 8024 4607 8076 4616
rect 8024 4573 8033 4607
rect 8033 4573 8067 4607
rect 8067 4573 8076 4607
rect 8024 4564 8076 4573
rect 10876 4607 10928 4616
rect 10876 4573 10885 4607
rect 10885 4573 10919 4607
rect 10919 4573 10928 4607
rect 10876 4564 10928 4573
rect 11060 4607 11112 4616
rect 11060 4573 11069 4607
rect 11069 4573 11103 4607
rect 11103 4573 11112 4607
rect 11060 4564 11112 4573
rect 12440 4607 12492 4616
rect 12440 4573 12449 4607
rect 12449 4573 12483 4607
rect 12483 4573 12492 4607
rect 12440 4564 12492 4573
rect 12716 4564 12768 4616
rect 12992 4564 13044 4616
rect 14096 4564 14148 4616
rect 17500 4607 17552 4616
rect 17500 4573 17509 4607
rect 17509 4573 17543 4607
rect 17543 4573 17552 4607
rect 17500 4564 17552 4573
rect 19156 4564 19208 4616
rect 22284 4564 22336 4616
rect 22836 4564 22888 4616
rect 7472 4496 7524 4548
rect 10692 4496 10744 4548
rect 16488 4496 16540 4548
rect 27528 4496 27580 4548
rect 33416 4496 33468 4548
rect 12072 4471 12124 4480
rect 12072 4437 12081 4471
rect 12081 4437 12115 4471
rect 12115 4437 12124 4471
rect 12072 4428 12124 4437
rect 15108 4428 15160 4480
rect 22652 4428 22704 4480
rect 7648 4326 7700 4378
rect 7712 4326 7764 4378
rect 7776 4326 7828 4378
rect 7840 4326 7892 4378
rect 20982 4326 21034 4378
rect 21046 4326 21098 4378
rect 21110 4326 21162 4378
rect 21174 4326 21226 4378
rect 34315 4326 34367 4378
rect 34379 4326 34431 4378
rect 34443 4326 34495 4378
rect 34507 4326 34559 4378
rect 1400 4224 1452 4276
rect 2320 4267 2372 4276
rect 2320 4233 2329 4267
rect 2329 4233 2363 4267
rect 2363 4233 2372 4267
rect 2320 4224 2372 4233
rect 2504 4224 2556 4276
rect 8116 4224 8168 4276
rect 9772 4224 9824 4276
rect 12256 4224 12308 4276
rect 12532 4267 12584 4276
rect 12532 4233 12541 4267
rect 12541 4233 12575 4267
rect 12575 4233 12584 4267
rect 12532 4224 12584 4233
rect 13912 4224 13964 4276
rect 16120 4267 16172 4276
rect 16120 4233 16129 4267
rect 16129 4233 16163 4267
rect 16163 4233 16172 4267
rect 16120 4224 16172 4233
rect 17316 4267 17368 4276
rect 17316 4233 17325 4267
rect 17325 4233 17359 4267
rect 17359 4233 17368 4267
rect 17316 4224 17368 4233
rect 17500 4224 17552 4276
rect 19156 4267 19208 4276
rect 19156 4233 19165 4267
rect 19165 4233 19199 4267
rect 19199 4233 19208 4267
rect 19156 4224 19208 4233
rect 22100 4224 22152 4276
rect 27712 4267 27764 4276
rect 27712 4233 27721 4267
rect 27721 4233 27755 4267
rect 27755 4233 27764 4267
rect 27712 4224 27764 4233
rect 27896 4224 27948 4276
rect 28264 4224 28316 4276
rect 34060 4224 34112 4276
rect 34980 4224 35032 4276
rect 10876 4199 10928 4208
rect 10876 4165 10885 4199
rect 10885 4165 10919 4199
rect 10919 4165 10928 4199
rect 10876 4156 10928 4165
rect 13820 4156 13872 4208
rect 15752 4199 15804 4208
rect 15752 4165 15761 4199
rect 15761 4165 15795 4199
rect 15795 4165 15804 4199
rect 15752 4156 15804 4165
rect 18972 4156 19024 4208
rect 8300 4131 8352 4140
rect 8300 4097 8309 4131
rect 8309 4097 8343 4131
rect 8343 4097 8352 4131
rect 8300 4088 8352 4097
rect 12992 4088 13044 4140
rect 14188 4088 14240 4140
rect 15108 4088 15160 4140
rect 18788 4131 18840 4140
rect 18788 4097 18797 4131
rect 18797 4097 18831 4131
rect 18831 4097 18840 4131
rect 18788 4088 18840 4097
rect 22284 4088 22336 4140
rect 22376 4088 22428 4140
rect 27988 4088 28040 4140
rect 34796 4156 34848 4208
rect 35440 4156 35492 4208
rect 2688 4020 2740 4072
rect 10784 4020 10836 4072
rect 11428 4063 11480 4072
rect 11428 4029 11437 4063
rect 11437 4029 11471 4063
rect 11471 4029 11480 4063
rect 11428 4020 11480 4029
rect 12348 4020 12400 4072
rect 17132 4020 17184 4072
rect 27528 4020 27580 4072
rect 35440 4063 35492 4072
rect 35440 4029 35449 4063
rect 35449 4029 35483 4063
rect 35483 4029 35492 4063
rect 35440 4020 35492 4029
rect 2044 3995 2096 4004
rect 2044 3961 2053 3995
rect 2053 3961 2087 3995
rect 2087 3961 2096 3995
rect 2044 3952 2096 3961
rect 10968 3952 11020 4004
rect 12532 3952 12584 4004
rect 14556 3995 14608 4004
rect 14556 3961 14565 3995
rect 14565 3961 14599 3995
rect 14599 3961 14608 3995
rect 14556 3952 14608 3961
rect 14648 3995 14700 4004
rect 14648 3961 14657 3995
rect 14657 3961 14691 3995
rect 14691 3961 14700 3995
rect 27252 3995 27304 4004
rect 14648 3952 14700 3961
rect 27252 3961 27261 3995
rect 27261 3961 27295 3995
rect 27295 3961 27304 3995
rect 27252 3952 27304 3961
rect 1584 3927 1636 3936
rect 1584 3893 1593 3927
rect 1593 3893 1627 3927
rect 1627 3893 1636 3927
rect 1584 3884 1636 3893
rect 7472 3884 7524 3936
rect 10324 3927 10376 3936
rect 10324 3893 10333 3927
rect 10333 3893 10367 3927
rect 10367 3893 10376 3927
rect 10324 3884 10376 3893
rect 10600 3927 10652 3936
rect 10600 3893 10609 3927
rect 10609 3893 10643 3927
rect 10643 3893 10652 3927
rect 10600 3884 10652 3893
rect 12164 3927 12216 3936
rect 12164 3893 12173 3927
rect 12173 3893 12207 3927
rect 12207 3893 12216 3927
rect 12992 3927 13044 3936
rect 12164 3884 12216 3893
rect 12992 3893 13001 3927
rect 13001 3893 13035 3927
rect 13035 3893 13044 3927
rect 12992 3884 13044 3893
rect 13176 3884 13228 3936
rect 15660 3884 15712 3936
rect 27344 3884 27396 3936
rect 35348 3884 35400 3936
rect 14315 3782 14367 3834
rect 14379 3782 14431 3834
rect 14443 3782 14495 3834
rect 14507 3782 14559 3834
rect 27648 3782 27700 3834
rect 27712 3782 27764 3834
rect 27776 3782 27828 3834
rect 27840 3782 27892 3834
rect 3056 3680 3108 3732
rect 9588 3680 9640 3732
rect 10784 3723 10836 3732
rect 10784 3689 10793 3723
rect 10793 3689 10827 3723
rect 10827 3689 10836 3723
rect 10784 3680 10836 3689
rect 13728 3680 13780 3732
rect 14004 3680 14056 3732
rect 14096 3680 14148 3732
rect 14648 3723 14700 3732
rect 14648 3689 14657 3723
rect 14657 3689 14691 3723
rect 14691 3689 14700 3723
rect 14648 3680 14700 3689
rect 15568 3723 15620 3732
rect 15568 3689 15577 3723
rect 15577 3689 15611 3723
rect 15611 3689 15620 3723
rect 15568 3680 15620 3689
rect 27252 3680 27304 3732
rect 572 3612 624 3664
rect 11060 3612 11112 3664
rect 11152 3612 11204 3664
rect 11704 3612 11756 3664
rect 1400 3587 1452 3596
rect 1400 3553 1409 3587
rect 1409 3553 1443 3587
rect 1443 3553 1452 3587
rect 1400 3544 1452 3553
rect 11428 3544 11480 3596
rect 9680 3476 9732 3528
rect 13176 3476 13228 3528
rect 13360 3519 13412 3528
rect 13360 3485 13369 3519
rect 13369 3485 13403 3519
rect 13403 3485 13412 3519
rect 13360 3476 13412 3485
rect 13452 3519 13504 3528
rect 13452 3485 13461 3519
rect 13461 3485 13495 3519
rect 13495 3485 13504 3519
rect 13452 3476 13504 3485
rect 10968 3408 11020 3460
rect 12900 3451 12952 3460
rect 12900 3417 12909 3451
rect 12909 3417 12943 3451
rect 12943 3417 12952 3451
rect 12900 3408 12952 3417
rect 12532 3383 12584 3392
rect 12532 3349 12541 3383
rect 12541 3349 12575 3383
rect 12575 3349 12584 3383
rect 12532 3340 12584 3349
rect 7648 3238 7700 3290
rect 7712 3238 7764 3290
rect 7776 3238 7828 3290
rect 7840 3238 7892 3290
rect 20982 3238 21034 3290
rect 21046 3238 21098 3290
rect 21110 3238 21162 3290
rect 21174 3238 21226 3290
rect 34315 3238 34367 3290
rect 34379 3238 34431 3290
rect 34443 3238 34495 3290
rect 34507 3238 34559 3290
rect 1400 3136 1452 3188
rect 10324 3136 10376 3188
rect 11428 3136 11480 3188
rect 11612 3179 11664 3188
rect 11612 3145 11621 3179
rect 11621 3145 11655 3179
rect 11655 3145 11664 3179
rect 11612 3136 11664 3145
rect 13452 3179 13504 3188
rect 13452 3145 13461 3179
rect 13461 3145 13495 3179
rect 13495 3145 13504 3179
rect 13452 3136 13504 3145
rect 13728 3136 13780 3188
rect 14188 3179 14240 3188
rect 14188 3145 14197 3179
rect 14197 3145 14231 3179
rect 14231 3145 14240 3179
rect 14188 3136 14240 3145
rect 11152 3068 11204 3120
rect 13360 3068 13412 3120
rect 13544 3000 13596 3052
rect 12808 2975 12860 2984
rect 12808 2941 12817 2975
rect 12817 2941 12851 2975
rect 12851 2941 12860 2975
rect 12808 2932 12860 2941
rect 12900 2864 12952 2916
rect 13636 2932 13688 2984
rect 14315 2694 14367 2746
rect 14379 2694 14431 2746
rect 14443 2694 14495 2746
rect 14507 2694 14559 2746
rect 27648 2694 27700 2746
rect 27712 2694 27764 2746
rect 27776 2694 27828 2746
rect 27840 2694 27892 2746
rect 12900 2635 12952 2644
rect 12900 2601 12909 2635
rect 12909 2601 12943 2635
rect 12943 2601 12952 2635
rect 12900 2592 12952 2601
rect 13360 2592 13412 2644
rect 12808 2524 12860 2576
rect 7648 2150 7700 2202
rect 7712 2150 7764 2202
rect 7776 2150 7828 2202
rect 7840 2150 7892 2202
rect 20982 2150 21034 2202
rect 21046 2150 21098 2202
rect 21110 2150 21162 2202
rect 21174 2150 21226 2202
rect 34315 2150 34367 2202
rect 34379 2150 34431 2202
rect 34443 2150 34495 2202
rect 34507 2150 34559 2202
<< metal2 >>
rect 1122 15520 1178 16000
rect 3422 15520 3478 16000
rect 3606 15872 3662 15881
rect 3606 15807 3662 15816
rect 1136 12374 1164 15520
rect 3238 15464 3294 15473
rect 3238 15399 3294 15408
rect 3146 14648 3202 14657
rect 3146 14583 3202 14592
rect 3054 14240 3110 14249
rect 3054 14175 3110 14184
rect 2780 13524 2832 13530
rect 2780 13466 2832 13472
rect 2792 13433 2820 13466
rect 2778 13424 2834 13433
rect 1584 13388 1636 13394
rect 1584 13330 1636 13336
rect 2320 13388 2372 13394
rect 2778 13359 2834 13368
rect 2320 13330 2372 13336
rect 1596 12986 1624 13330
rect 1584 12980 1636 12986
rect 1584 12922 1636 12928
rect 2044 12776 2096 12782
rect 2044 12718 2096 12724
rect 1124 12368 1176 12374
rect 1124 12310 1176 12316
rect 1676 11824 1728 11830
rect 1676 11766 1728 11772
rect 1400 11144 1452 11150
rect 1400 11086 1452 11092
rect 1306 10976 1362 10985
rect 1306 10911 1362 10920
rect 1320 9636 1348 10911
rect 1412 10810 1440 11086
rect 1400 10804 1452 10810
rect 1400 10746 1452 10752
rect 1688 10266 1716 11766
rect 1676 10260 1728 10266
rect 1676 10202 1728 10208
rect 1320 9608 1440 9636
rect 1412 4826 1440 9608
rect 1688 9178 1716 10202
rect 1952 10056 2004 10062
rect 1952 9998 2004 10004
rect 1964 9178 1992 9998
rect 2056 9654 2084 12718
rect 2228 10736 2280 10742
rect 2228 10678 2280 10684
rect 2240 10198 2268 10678
rect 2228 10192 2280 10198
rect 2228 10134 2280 10140
rect 2044 9648 2096 9654
rect 2044 9590 2096 9596
rect 1676 9172 1728 9178
rect 1676 9114 1728 9120
rect 1952 9172 2004 9178
rect 1952 9114 2004 9120
rect 1676 9036 1728 9042
rect 1676 8978 1728 8984
rect 1582 8936 1638 8945
rect 1582 8871 1638 8880
rect 1492 6248 1544 6254
rect 1492 6190 1544 6196
rect 1504 5778 1532 6190
rect 1492 5772 1544 5778
rect 1492 5714 1544 5720
rect 1400 4820 1452 4826
rect 1400 4762 1452 4768
rect 1400 4684 1452 4690
rect 1400 4626 1452 4632
rect 1412 4282 1440 4626
rect 1400 4276 1452 4282
rect 1400 4218 1452 4224
rect 1596 3942 1624 8871
rect 1688 6730 1716 8978
rect 1964 8634 1992 9114
rect 2332 8906 2360 13330
rect 2780 13184 2832 13190
rect 2780 13126 2832 13132
rect 2504 12300 2556 12306
rect 2504 12242 2556 12248
rect 2688 12300 2740 12306
rect 2688 12242 2740 12248
rect 2516 11898 2544 12242
rect 2596 12096 2648 12102
rect 2596 12038 2648 12044
rect 2504 11892 2556 11898
rect 2504 11834 2556 11840
rect 2608 11762 2636 12038
rect 2700 11830 2728 12242
rect 2688 11824 2740 11830
rect 2688 11766 2740 11772
rect 2504 11756 2556 11762
rect 2504 11698 2556 11704
rect 2596 11756 2648 11762
rect 2596 11698 2648 11704
rect 2410 11656 2466 11665
rect 2410 11591 2412 11600
rect 2464 11591 2466 11600
rect 2412 11562 2464 11568
rect 2424 11354 2452 11562
rect 2516 11529 2544 11698
rect 2502 11520 2558 11529
rect 2502 11455 2558 11464
rect 2412 11348 2464 11354
rect 2412 11290 2464 11296
rect 2608 11098 2636 11698
rect 2608 11082 2728 11098
rect 2504 11076 2556 11082
rect 2608 11076 2740 11082
rect 2608 11070 2688 11076
rect 2504 11018 2556 11024
rect 2688 11018 2740 11024
rect 2516 10033 2544 11018
rect 2596 10056 2648 10062
rect 2502 10024 2558 10033
rect 2596 9998 2648 10004
rect 2502 9959 2558 9968
rect 2412 9920 2464 9926
rect 2412 9862 2464 9868
rect 2424 9586 2452 9862
rect 2412 9580 2464 9586
rect 2412 9522 2464 9528
rect 2516 9450 2544 9959
rect 2608 9897 2636 9998
rect 2594 9888 2650 9897
rect 2594 9823 2650 9832
rect 2792 9761 2820 13126
rect 2964 12912 3016 12918
rect 2964 12854 3016 12860
rect 2872 12096 2924 12102
rect 2872 12038 2924 12044
rect 2884 10169 2912 12038
rect 2976 11150 3004 12854
rect 2964 11144 3016 11150
rect 2964 11086 3016 11092
rect 2870 10160 2926 10169
rect 2870 10095 2926 10104
rect 2778 9752 2834 9761
rect 2778 9687 2834 9696
rect 2976 9654 3004 11086
rect 2964 9648 3016 9654
rect 2964 9590 3016 9596
rect 2688 9580 2740 9586
rect 2688 9522 2740 9528
rect 2700 9466 2728 9522
rect 2504 9444 2556 9450
rect 2700 9438 2820 9466
rect 2504 9386 2556 9392
rect 2596 9376 2648 9382
rect 2596 9318 2648 9324
rect 2320 8900 2372 8906
rect 2320 8842 2372 8848
rect 2608 8650 2636 9318
rect 2686 9072 2742 9081
rect 2686 9007 2688 9016
rect 2740 9007 2742 9016
rect 2688 8978 2740 8984
rect 2516 8634 2636 8650
rect 1952 8628 2004 8634
rect 1952 8570 2004 8576
rect 2504 8628 2636 8634
rect 2556 8622 2636 8628
rect 2504 8570 2556 8576
rect 1964 8430 1992 8570
rect 2410 8528 2466 8537
rect 2410 8463 2466 8472
rect 1952 8424 2004 8430
rect 1952 8366 2004 8372
rect 2320 8016 2372 8022
rect 2320 7958 2372 7964
rect 1860 7744 1912 7750
rect 1860 7686 1912 7692
rect 1872 6866 1900 7686
rect 2332 7478 2360 7958
rect 2136 7472 2188 7478
rect 2136 7414 2188 7420
rect 2320 7472 2372 7478
rect 2320 7414 2372 7420
rect 2148 6934 2176 7414
rect 2136 6928 2188 6934
rect 2136 6870 2188 6876
rect 1860 6860 1912 6866
rect 1860 6802 1912 6808
rect 1676 6724 1728 6730
rect 1676 6666 1728 6672
rect 1872 5846 1900 6802
rect 2228 6792 2280 6798
rect 2228 6734 2280 6740
rect 2240 6186 2268 6734
rect 2228 6180 2280 6186
rect 2228 6122 2280 6128
rect 1860 5840 1912 5846
rect 1860 5782 1912 5788
rect 2424 4826 2452 8463
rect 2792 8090 2820 9438
rect 2872 8968 2924 8974
rect 2872 8910 2924 8916
rect 2780 8084 2832 8090
rect 2780 8026 2832 8032
rect 2884 8022 2912 8910
rect 2872 8016 2924 8022
rect 2872 7958 2924 7964
rect 2504 7948 2556 7954
rect 2504 7890 2556 7896
rect 2516 7274 2544 7890
rect 2688 7880 2740 7886
rect 2688 7822 2740 7828
rect 2594 7576 2650 7585
rect 2700 7546 2728 7822
rect 2594 7511 2650 7520
rect 2688 7540 2740 7546
rect 2504 7268 2556 7274
rect 2504 7210 2556 7216
rect 2608 7206 2636 7511
rect 2688 7482 2740 7488
rect 2596 7200 2648 7206
rect 2596 7142 2648 7148
rect 2608 7002 2636 7142
rect 2596 6996 2648 7002
rect 2596 6938 2648 6944
rect 2596 5364 2648 5370
rect 2596 5306 2648 5312
rect 2504 5228 2556 5234
rect 2504 5170 2556 5176
rect 2412 4820 2464 4826
rect 2412 4762 2464 4768
rect 2516 4690 2544 5170
rect 2608 5098 2636 5306
rect 2596 5092 2648 5098
rect 2596 5034 2648 5040
rect 2504 4684 2556 4690
rect 2504 4626 2556 4632
rect 2516 4282 2544 4626
rect 2320 4276 2372 4282
rect 2320 4218 2372 4224
rect 2504 4276 2556 4282
rect 2504 4218 2556 4224
rect 2332 4185 2360 4218
rect 2318 4176 2374 4185
rect 2318 4111 2374 4120
rect 2700 4078 2728 7482
rect 2780 7404 2832 7410
rect 2780 7346 2832 7352
rect 2792 7041 2820 7346
rect 2778 7032 2834 7041
rect 2778 6967 2834 6976
rect 2884 6458 2912 7958
rect 2964 7268 3016 7274
rect 2964 7210 3016 7216
rect 2976 6730 3004 7210
rect 2964 6724 3016 6730
rect 2964 6666 3016 6672
rect 2872 6452 2924 6458
rect 2872 6394 2924 6400
rect 2884 6066 2912 6394
rect 2964 6248 3016 6254
rect 2964 6190 3016 6196
rect 2792 6038 2912 6066
rect 2792 5778 2820 6038
rect 2872 5908 2924 5914
rect 2872 5850 2924 5856
rect 2780 5772 2832 5778
rect 2780 5714 2832 5720
rect 2792 4758 2820 5714
rect 2884 5234 2912 5850
rect 2976 5370 3004 6190
rect 2964 5364 3016 5370
rect 2964 5306 3016 5312
rect 2872 5228 2924 5234
rect 2872 5170 2924 5176
rect 2884 4826 2912 5170
rect 2964 5092 3016 5098
rect 2964 5034 3016 5040
rect 2872 4820 2924 4826
rect 2872 4762 2924 4768
rect 2780 4752 2832 4758
rect 2780 4694 2832 4700
rect 2688 4072 2740 4078
rect 2042 4040 2098 4049
rect 2688 4014 2740 4020
rect 2042 3975 2044 3984
rect 2096 3975 2098 3984
rect 2044 3946 2096 3952
rect 1584 3936 1636 3942
rect 1584 3878 1636 3884
rect 570 3768 626 3777
rect 570 3703 626 3712
rect 584 3670 612 3703
rect 572 3664 624 3670
rect 572 3606 624 3612
rect 1398 3632 1454 3641
rect 1398 3567 1400 3576
rect 1452 3567 1454 3576
rect 1400 3538 1452 3544
rect 1412 3194 1440 3538
rect 1400 3188 1452 3194
rect 1400 3130 1452 3136
rect 2976 513 3004 5034
rect 3068 3738 3096 14175
rect 3160 13938 3188 14583
rect 3148 13932 3200 13938
rect 3148 13874 3200 13880
rect 3252 13870 3280 15399
rect 3436 14226 3464 15520
rect 3514 15056 3570 15065
rect 3514 14991 3570 15000
rect 3344 14198 3464 14226
rect 3240 13864 3292 13870
rect 3240 13806 3292 13812
rect 3344 12850 3372 14198
rect 3424 14068 3476 14074
rect 3424 14010 3476 14016
rect 3436 13841 3464 14010
rect 3528 14006 3556 14991
rect 3620 14142 3648 15807
rect 5814 15520 5870 16000
rect 8114 15520 8170 16000
rect 10506 15520 10562 16000
rect 12806 15520 12862 16000
rect 15198 15520 15254 16000
rect 17590 15520 17646 16000
rect 19890 15520 19946 16000
rect 22282 15520 22338 16000
rect 24582 15520 24638 16000
rect 26974 15520 27030 16000
rect 29366 15520 29422 16000
rect 31666 15520 31722 16000
rect 34058 15520 34114 16000
rect 34518 15872 34574 15881
rect 34518 15807 34574 15816
rect 3608 14136 3660 14142
rect 3608 14078 3660 14084
rect 3516 14000 3568 14006
rect 3516 13942 3568 13948
rect 3422 13832 3478 13841
rect 3422 13767 3478 13776
rect 5828 13462 5856 15520
rect 7472 14136 7524 14142
rect 7472 14078 7524 14084
rect 6920 14068 6972 14074
rect 6920 14010 6972 14016
rect 5816 13456 5868 13462
rect 5816 13398 5868 13404
rect 4160 13388 4212 13394
rect 4160 13330 4212 13336
rect 5172 13388 5224 13394
rect 5172 13330 5224 13336
rect 3516 13184 3568 13190
rect 3516 13126 3568 13132
rect 3332 12844 3384 12850
rect 3332 12786 3384 12792
rect 3424 12844 3476 12850
rect 3424 12786 3476 12792
rect 3436 12617 3464 12786
rect 3422 12608 3478 12617
rect 3422 12543 3478 12552
rect 3528 12209 3556 13126
rect 4066 13016 4122 13025
rect 4066 12951 4068 12960
rect 4120 12951 4122 12960
rect 4068 12922 4120 12928
rect 4172 12782 4200 13330
rect 4528 13252 4580 13258
rect 4528 13194 4580 13200
rect 4160 12776 4212 12782
rect 4160 12718 4212 12724
rect 4540 12714 4568 13194
rect 4620 12776 4672 12782
rect 4620 12718 4672 12724
rect 4068 12708 4120 12714
rect 4068 12650 4120 12656
rect 4528 12708 4580 12714
rect 4528 12650 4580 12656
rect 4080 12594 4108 12650
rect 4080 12566 4200 12594
rect 4172 12442 4200 12566
rect 4160 12436 4212 12442
rect 4160 12378 4212 12384
rect 3514 12200 3570 12209
rect 3514 12135 3570 12144
rect 3608 12096 3660 12102
rect 3608 12038 3660 12044
rect 4344 12096 4396 12102
rect 4344 12038 4396 12044
rect 3620 11762 3648 12038
rect 3882 11792 3938 11801
rect 3608 11756 3660 11762
rect 3882 11727 3938 11736
rect 3608 11698 3660 11704
rect 3608 11552 3660 11558
rect 3608 11494 3660 11500
rect 3424 11280 3476 11286
rect 3424 11222 3476 11228
rect 3148 11008 3200 11014
rect 3148 10950 3200 10956
rect 3160 10538 3188 10950
rect 3148 10532 3200 10538
rect 3148 10474 3200 10480
rect 3160 9994 3188 10474
rect 3148 9988 3200 9994
rect 3148 9930 3200 9936
rect 3436 9926 3464 11222
rect 3620 11121 3648 11494
rect 3700 11212 3752 11218
rect 3700 11154 3752 11160
rect 3606 11112 3662 11121
rect 3606 11047 3608 11056
rect 3660 11047 3662 11056
rect 3608 11018 3660 11024
rect 3712 10470 3740 11154
rect 3896 10810 3924 11727
rect 4160 11620 4212 11626
rect 4160 11562 4212 11568
rect 4066 11384 4122 11393
rect 4172 11354 4200 11562
rect 4066 11319 4122 11328
rect 4160 11348 4212 11354
rect 3976 11144 4028 11150
rect 3976 11086 4028 11092
rect 3884 10804 3936 10810
rect 3884 10746 3936 10752
rect 3882 10568 3938 10577
rect 3882 10503 3938 10512
rect 3700 10464 3752 10470
rect 3620 10424 3700 10452
rect 3424 9920 3476 9926
rect 3424 9862 3476 9868
rect 3620 9518 3648 10424
rect 3700 10406 3752 10412
rect 3700 9988 3752 9994
rect 3700 9930 3752 9936
rect 3424 9512 3476 9518
rect 3424 9454 3476 9460
rect 3608 9512 3660 9518
rect 3608 9454 3660 9460
rect 3436 8634 3464 9454
rect 3712 9450 3740 9930
rect 3792 9716 3844 9722
rect 3792 9658 3844 9664
rect 3700 9444 3752 9450
rect 3700 9386 3752 9392
rect 3712 9042 3740 9386
rect 3700 9036 3752 9042
rect 3700 8978 3752 8984
rect 3424 8628 3476 8634
rect 3424 8570 3476 8576
rect 3148 7472 3200 7478
rect 3148 7414 3200 7420
rect 3160 7206 3188 7414
rect 3148 7200 3200 7206
rect 3146 7168 3148 7177
rect 3200 7168 3202 7177
rect 3146 7103 3202 7112
rect 3146 6896 3202 6905
rect 3146 6831 3202 6840
rect 3160 5098 3188 6831
rect 3516 6792 3568 6798
rect 3516 6734 3568 6740
rect 3606 6760 3662 6769
rect 3238 6080 3294 6089
rect 3238 6015 3294 6024
rect 3148 5092 3200 5098
rect 3148 5034 3200 5040
rect 3056 3732 3108 3738
rect 3056 3674 3108 3680
rect 3252 921 3280 6015
rect 3528 5778 3556 6734
rect 3606 6695 3662 6704
rect 3516 5772 3568 5778
rect 3516 5714 3568 5720
rect 3332 5296 3384 5302
rect 3332 5238 3384 5244
rect 3344 5137 3372 5238
rect 3330 5128 3386 5137
rect 3330 5063 3386 5072
rect 3424 5092 3476 5098
rect 3424 5034 3476 5040
rect 3436 1329 3464 5034
rect 3422 1320 3478 1329
rect 3422 1255 3478 1264
rect 3238 912 3294 921
rect 3238 847 3294 856
rect 2962 504 3018 513
rect 2962 439 3018 448
rect 3620 241 3648 6695
rect 3804 4593 3832 9658
rect 3896 9602 3924 10503
rect 3988 10146 4016 11086
rect 4080 10266 4108 11319
rect 4160 11290 4212 11296
rect 4160 11212 4212 11218
rect 4160 11154 4212 11160
rect 4172 10742 4200 11154
rect 4356 11014 4384 12038
rect 4344 11008 4396 11014
rect 4344 10950 4396 10956
rect 4160 10736 4212 10742
rect 4160 10678 4212 10684
rect 4068 10260 4120 10266
rect 4068 10202 4120 10208
rect 3988 10118 4292 10146
rect 3988 9897 4016 10118
rect 4068 9920 4120 9926
rect 3974 9888 4030 9897
rect 4120 9880 4200 9908
rect 4068 9862 4120 9868
rect 3974 9823 4030 9832
rect 3896 9574 4016 9602
rect 3988 8566 4016 9574
rect 4066 9344 4122 9353
rect 4066 9279 4122 9288
rect 3976 8560 4028 8566
rect 3976 8502 4028 8508
rect 3882 8392 3938 8401
rect 3882 8327 3938 8336
rect 3896 8090 3924 8327
rect 3884 8084 3936 8090
rect 3884 8026 3936 8032
rect 3974 7032 4030 7041
rect 3974 6967 4030 6976
rect 3988 5817 4016 6967
rect 3974 5808 4030 5817
rect 3974 5743 4030 5752
rect 3976 5704 4028 5710
rect 3976 5646 4028 5652
rect 3884 5228 3936 5234
rect 3884 5170 3936 5176
rect 3896 4826 3924 5170
rect 3988 5001 4016 5646
rect 4080 5642 4108 9279
rect 4172 8906 4200 9880
rect 4264 9382 4292 10118
rect 4344 10124 4396 10130
rect 4344 10066 4396 10072
rect 4252 9376 4304 9382
rect 4252 9318 4304 9324
rect 4160 8900 4212 8906
rect 4160 8842 4212 8848
rect 4356 8838 4384 10066
rect 4540 9722 4568 12650
rect 4632 10538 4660 12718
rect 5184 12714 5212 13330
rect 6092 13320 6144 13326
rect 6092 13262 6144 13268
rect 4804 12708 4856 12714
rect 4804 12650 4856 12656
rect 5172 12708 5224 12714
rect 5172 12650 5224 12656
rect 4712 12640 4764 12646
rect 4712 12582 4764 12588
rect 4724 12442 4752 12582
rect 4712 12436 4764 12442
rect 4712 12378 4764 12384
rect 4724 11898 4752 12378
rect 4816 12102 4844 12650
rect 5356 12640 5408 12646
rect 5356 12582 5408 12588
rect 5724 12640 5776 12646
rect 5724 12582 5776 12588
rect 5264 12368 5316 12374
rect 5264 12310 5316 12316
rect 4804 12096 4856 12102
rect 4804 12038 4856 12044
rect 4988 12096 5040 12102
rect 4988 12038 5040 12044
rect 4712 11892 4764 11898
rect 4712 11834 4764 11840
rect 5000 11762 5028 12038
rect 4988 11756 5040 11762
rect 4988 11698 5040 11704
rect 4896 11552 4948 11558
rect 4896 11494 4948 11500
rect 4804 10600 4856 10606
rect 4804 10542 4856 10548
rect 4620 10532 4672 10538
rect 4620 10474 4672 10480
rect 4620 10056 4672 10062
rect 4618 10024 4620 10033
rect 4672 10024 4674 10033
rect 4618 9959 4674 9968
rect 4528 9716 4580 9722
rect 4528 9658 4580 9664
rect 4528 9580 4580 9586
rect 4528 9522 4580 9528
rect 4344 8832 4396 8838
rect 4344 8774 4396 8780
rect 4160 8628 4212 8634
rect 4160 8570 4212 8576
rect 4172 8022 4200 8570
rect 4250 8256 4306 8265
rect 4250 8191 4306 8200
rect 4160 8016 4212 8022
rect 4160 7958 4212 7964
rect 4264 7002 4292 8191
rect 4356 8129 4384 8774
rect 4342 8120 4398 8129
rect 4342 8055 4398 8064
rect 4344 7744 4396 7750
rect 4342 7712 4344 7721
rect 4396 7712 4398 7721
rect 4342 7647 4398 7656
rect 4356 7342 4384 7647
rect 4344 7336 4396 7342
rect 4344 7278 4396 7284
rect 4252 6996 4304 7002
rect 4252 6938 4304 6944
rect 4160 6792 4212 6798
rect 4160 6734 4212 6740
rect 4172 6458 4200 6734
rect 4356 6730 4384 7278
rect 4344 6724 4396 6730
rect 4344 6666 4396 6672
rect 4160 6452 4212 6458
rect 4160 6394 4212 6400
rect 4068 5636 4120 5642
rect 4068 5578 4120 5584
rect 4066 5400 4122 5409
rect 4066 5335 4068 5344
rect 4120 5335 4122 5344
rect 4068 5306 4120 5312
rect 4160 5092 4212 5098
rect 4160 5034 4212 5040
rect 4068 5024 4120 5030
rect 3974 4992 4030 5001
rect 4068 4966 4120 4972
rect 3974 4927 4030 4936
rect 4080 4865 4108 4966
rect 4066 4856 4122 4865
rect 3884 4820 3936 4826
rect 4172 4826 4200 5034
rect 4066 4791 4122 4800
rect 4160 4820 4212 4826
rect 3884 4762 3936 4768
rect 4160 4762 4212 4768
rect 3790 4584 3846 4593
rect 3790 4519 3846 4528
rect 4540 4321 4568 9522
rect 4712 7880 4764 7886
rect 4712 7822 4764 7828
rect 4724 7274 4752 7822
rect 4712 7268 4764 7274
rect 4712 7210 4764 7216
rect 4724 6662 4752 7210
rect 4712 6656 4764 6662
rect 4712 6598 4764 6604
rect 4620 6180 4672 6186
rect 4620 6122 4672 6128
rect 4632 5914 4660 6122
rect 4620 5908 4672 5914
rect 4620 5850 4672 5856
rect 4712 5024 4764 5030
rect 4710 4992 4712 5001
rect 4764 4992 4766 5001
rect 4710 4927 4766 4936
rect 4526 4312 4582 4321
rect 4526 4247 4582 4256
rect 4816 2825 4844 10542
rect 4908 3097 4936 11494
rect 5276 10810 5304 12310
rect 5368 12238 5396 12582
rect 5356 12232 5408 12238
rect 5356 12174 5408 12180
rect 5632 12232 5684 12238
rect 5632 12174 5684 12180
rect 5368 11082 5396 12174
rect 5644 11694 5672 12174
rect 5632 11688 5684 11694
rect 5632 11630 5684 11636
rect 5540 11348 5592 11354
rect 5540 11290 5592 11296
rect 5356 11076 5408 11082
rect 5356 11018 5408 11024
rect 5264 10804 5316 10810
rect 5264 10746 5316 10752
rect 4988 10668 5040 10674
rect 4988 10610 5040 10616
rect 5000 6633 5028 10610
rect 5356 10464 5408 10470
rect 5356 10406 5408 10412
rect 5368 10130 5396 10406
rect 5552 10198 5580 11290
rect 5644 11218 5672 11630
rect 5632 11212 5684 11218
rect 5632 11154 5684 11160
rect 5644 10849 5672 11154
rect 5630 10840 5686 10849
rect 5736 10810 5764 12582
rect 5908 12096 5960 12102
rect 5908 12038 5960 12044
rect 5920 11762 5948 12038
rect 5908 11756 5960 11762
rect 5908 11698 5960 11704
rect 5816 11212 5868 11218
rect 5816 11154 5868 11160
rect 5630 10775 5686 10784
rect 5724 10804 5776 10810
rect 5724 10746 5776 10752
rect 5828 10674 5856 11154
rect 5632 10668 5684 10674
rect 5632 10610 5684 10616
rect 5816 10668 5868 10674
rect 5816 10610 5868 10616
rect 5644 10577 5672 10610
rect 5630 10568 5686 10577
rect 5630 10503 5686 10512
rect 5816 10464 5868 10470
rect 5816 10406 5868 10412
rect 5540 10192 5592 10198
rect 5540 10134 5592 10140
rect 5356 10124 5408 10130
rect 5356 10066 5408 10072
rect 5080 9920 5132 9926
rect 5080 9862 5132 9868
rect 5092 9178 5120 9862
rect 5368 9518 5396 10066
rect 5552 9722 5580 10134
rect 5540 9716 5592 9722
rect 5540 9658 5592 9664
rect 5356 9512 5408 9518
rect 5356 9454 5408 9460
rect 5262 9208 5318 9217
rect 5080 9172 5132 9178
rect 5262 9143 5318 9152
rect 5080 9114 5132 9120
rect 5092 8634 5120 9114
rect 5276 9042 5304 9143
rect 5448 9104 5500 9110
rect 5448 9046 5500 9052
rect 5264 9036 5316 9042
rect 5264 8978 5316 8984
rect 5080 8628 5132 8634
rect 5080 8570 5132 8576
rect 5276 8498 5304 8978
rect 5356 8968 5408 8974
rect 5354 8936 5356 8945
rect 5408 8936 5410 8945
rect 5354 8871 5410 8880
rect 5264 8492 5316 8498
rect 5264 8434 5316 8440
rect 5356 8424 5408 8430
rect 5356 8366 5408 8372
rect 5080 8016 5132 8022
rect 5080 7958 5132 7964
rect 5092 7002 5120 7958
rect 5368 7546 5396 8366
rect 5460 8362 5488 9046
rect 5724 8832 5776 8838
rect 5724 8774 5776 8780
rect 5540 8492 5592 8498
rect 5540 8434 5592 8440
rect 5552 8401 5580 8434
rect 5538 8392 5594 8401
rect 5448 8356 5500 8362
rect 5736 8362 5764 8774
rect 5828 8537 5856 10406
rect 5920 10266 5948 11698
rect 6000 11620 6052 11626
rect 6000 11562 6052 11568
rect 5908 10260 5960 10266
rect 5908 10202 5960 10208
rect 5908 9376 5960 9382
rect 5908 9318 5960 9324
rect 5814 8528 5870 8537
rect 5814 8463 5870 8472
rect 5538 8327 5594 8336
rect 5724 8356 5776 8362
rect 5448 8298 5500 8304
rect 5724 8298 5776 8304
rect 5356 7540 5408 7546
rect 5356 7482 5408 7488
rect 5080 6996 5132 7002
rect 5080 6938 5132 6944
rect 5368 6934 5396 7482
rect 5460 7449 5488 8298
rect 5540 7540 5592 7546
rect 5540 7482 5592 7488
rect 5446 7440 5502 7449
rect 5446 7375 5502 7384
rect 5356 6928 5408 6934
rect 5552 6882 5580 7482
rect 5356 6870 5408 6876
rect 5172 6860 5224 6866
rect 5172 6802 5224 6808
rect 5460 6854 5580 6882
rect 4986 6624 5042 6633
rect 4986 6559 5042 6568
rect 5184 5914 5212 6802
rect 5460 6798 5488 6854
rect 5448 6792 5500 6798
rect 5448 6734 5500 6740
rect 5736 6730 5764 8298
rect 5724 6724 5776 6730
rect 5724 6666 5776 6672
rect 5356 6656 5408 6662
rect 5356 6598 5408 6604
rect 5368 6322 5396 6598
rect 5356 6316 5408 6322
rect 5356 6258 5408 6264
rect 5172 5908 5224 5914
rect 5172 5850 5224 5856
rect 5368 5778 5396 6258
rect 5540 6112 5592 6118
rect 5540 6054 5592 6060
rect 5552 5778 5580 6054
rect 5356 5772 5408 5778
rect 5356 5714 5408 5720
rect 5540 5772 5592 5778
rect 5540 5714 5592 5720
rect 5368 5370 5396 5714
rect 5356 5364 5408 5370
rect 5356 5306 5408 5312
rect 5552 5234 5580 5714
rect 5540 5228 5592 5234
rect 5540 5170 5592 5176
rect 5552 4690 5580 5170
rect 5540 4684 5592 4690
rect 5540 4626 5592 4632
rect 5920 3913 5948 9318
rect 6012 4593 6040 11562
rect 6104 9450 6132 13262
rect 6644 12980 6696 12986
rect 6644 12922 6696 12928
rect 6656 12442 6684 12922
rect 6644 12436 6696 12442
rect 6644 12378 6696 12384
rect 6276 12300 6328 12306
rect 6276 12242 6328 12248
rect 6288 11558 6316 12242
rect 6828 11688 6880 11694
rect 6826 11656 6828 11665
rect 6880 11656 6882 11665
rect 6826 11591 6882 11600
rect 6276 11552 6328 11558
rect 6276 11494 6328 11500
rect 6092 9444 6144 9450
rect 6092 9386 6144 9392
rect 6182 8256 6238 8265
rect 6182 8191 6238 8200
rect 6092 7744 6144 7750
rect 6092 7686 6144 7692
rect 6104 7410 6132 7686
rect 6092 7404 6144 7410
rect 6092 7346 6144 7352
rect 6196 6662 6224 8191
rect 6184 6656 6236 6662
rect 6184 6598 6236 6604
rect 6196 6118 6224 6598
rect 6184 6112 6236 6118
rect 6182 6080 6184 6089
rect 6236 6080 6238 6089
rect 6182 6015 6238 6024
rect 6288 5817 6316 11494
rect 6828 11008 6880 11014
rect 6828 10950 6880 10956
rect 6840 10810 6868 10950
rect 6932 10810 6960 14010
rect 7104 13932 7156 13938
rect 7104 13874 7156 13880
rect 7116 13530 7144 13874
rect 7104 13524 7156 13530
rect 7104 13466 7156 13472
rect 7104 13388 7156 13394
rect 7104 13330 7156 13336
rect 7012 12844 7064 12850
rect 7012 12786 7064 12792
rect 7024 11898 7052 12786
rect 7116 12646 7144 13330
rect 7484 12986 7512 14078
rect 7622 13084 7918 13104
rect 7678 13082 7702 13084
rect 7758 13082 7782 13084
rect 7838 13082 7862 13084
rect 7700 13030 7702 13082
rect 7764 13030 7776 13082
rect 7838 13030 7840 13082
rect 7678 13028 7702 13030
rect 7758 13028 7782 13030
rect 7838 13028 7862 13030
rect 7622 13008 7918 13028
rect 7472 12980 7524 12986
rect 7472 12922 7524 12928
rect 8128 12918 8156 15520
rect 8392 14000 8444 14006
rect 8392 13942 8444 13948
rect 8116 12912 8168 12918
rect 8116 12854 8168 12860
rect 7196 12776 7248 12782
rect 7196 12718 7248 12724
rect 7104 12640 7156 12646
rect 7104 12582 7156 12588
rect 7012 11892 7064 11898
rect 7012 11834 7064 11840
rect 7116 11286 7144 12582
rect 7104 11280 7156 11286
rect 7104 11222 7156 11228
rect 6828 10804 6880 10810
rect 6828 10746 6880 10752
rect 6920 10804 6972 10810
rect 6920 10746 6972 10752
rect 6552 10600 6604 10606
rect 6552 10542 6604 10548
rect 6368 9036 6420 9042
rect 6368 8978 6420 8984
rect 6380 8362 6408 8978
rect 6460 8832 6512 8838
rect 6460 8774 6512 8780
rect 6472 8498 6500 8774
rect 6460 8492 6512 8498
rect 6460 8434 6512 8440
rect 6368 8356 6420 8362
rect 6368 8298 6420 8304
rect 6380 7313 6408 8298
rect 6460 8288 6512 8294
rect 6460 8230 6512 8236
rect 6472 7750 6500 8230
rect 6460 7744 6512 7750
rect 6460 7686 6512 7692
rect 6366 7304 6422 7313
rect 6366 7239 6422 7248
rect 6274 5808 6330 5817
rect 6274 5743 6330 5752
rect 5998 4584 6054 4593
rect 5998 4519 6054 4528
rect 5906 3904 5962 3913
rect 5906 3839 5962 3848
rect 4894 3088 4950 3097
rect 4894 3023 4950 3032
rect 4802 2816 4858 2825
rect 4802 2751 4858 2760
rect 4908 2145 4936 3023
rect 4894 2136 4950 2145
rect 4894 2071 4950 2080
rect 5920 1737 5948 3839
rect 6380 2553 6408 7239
rect 6472 4049 6500 7686
rect 6564 7177 6592 10542
rect 6828 10464 6880 10470
rect 7116 10418 7144 11222
rect 6880 10412 7144 10418
rect 6828 10406 7144 10412
rect 6840 10390 7144 10406
rect 6644 10260 6696 10266
rect 6644 10202 6696 10208
rect 6656 10033 6684 10202
rect 6642 10024 6698 10033
rect 6642 9959 6698 9968
rect 6644 9104 6696 9110
rect 6644 9046 6696 9052
rect 6656 8294 6684 9046
rect 6736 8900 6788 8906
rect 6736 8842 6788 8848
rect 6644 8288 6696 8294
rect 6644 8230 6696 8236
rect 6644 8016 6696 8022
rect 6644 7958 6696 7964
rect 6656 7546 6684 7958
rect 6748 7721 6776 8842
rect 6828 8424 6880 8430
rect 6828 8366 6880 8372
rect 6840 7818 6868 8366
rect 7012 8288 7064 8294
rect 7012 8230 7064 8236
rect 7024 7834 7052 8230
rect 7116 7936 7144 10390
rect 7208 8294 7236 12718
rect 8300 12300 8352 12306
rect 8300 12242 8352 12248
rect 7472 12096 7524 12102
rect 7472 12038 7524 12044
rect 8024 12096 8076 12102
rect 8024 12038 8076 12044
rect 7380 11756 7432 11762
rect 7380 11698 7432 11704
rect 7392 9586 7420 11698
rect 7484 9654 7512 12038
rect 7622 11996 7918 12016
rect 7678 11994 7702 11996
rect 7758 11994 7782 11996
rect 7838 11994 7862 11996
rect 7700 11942 7702 11994
rect 7764 11942 7776 11994
rect 7838 11942 7840 11994
rect 7678 11940 7702 11942
rect 7758 11940 7782 11942
rect 7838 11940 7862 11942
rect 7622 11920 7918 11940
rect 8036 11937 8064 12038
rect 8022 11928 8078 11937
rect 8312 11898 8340 12242
rect 8022 11863 8078 11872
rect 8300 11892 8352 11898
rect 8300 11834 8352 11840
rect 8024 11824 8076 11830
rect 8024 11766 8076 11772
rect 7564 11552 7616 11558
rect 7564 11494 7616 11500
rect 7576 11257 7604 11494
rect 7562 11248 7618 11257
rect 7562 11183 7618 11192
rect 7622 10908 7918 10928
rect 7678 10906 7702 10908
rect 7758 10906 7782 10908
rect 7838 10906 7862 10908
rect 7700 10854 7702 10906
rect 7764 10854 7776 10906
rect 7838 10854 7840 10906
rect 7678 10852 7702 10854
rect 7758 10852 7782 10854
rect 7838 10852 7862 10854
rect 7622 10832 7918 10852
rect 7932 10736 7984 10742
rect 7932 10678 7984 10684
rect 7944 10180 7972 10678
rect 8036 10305 8064 11766
rect 8116 11756 8168 11762
rect 8116 11698 8168 11704
rect 8022 10296 8078 10305
rect 8022 10231 8078 10240
rect 7944 10152 8064 10180
rect 7622 9820 7918 9840
rect 7678 9818 7702 9820
rect 7758 9818 7782 9820
rect 7838 9818 7862 9820
rect 7700 9766 7702 9818
rect 7764 9766 7776 9818
rect 7838 9766 7840 9818
rect 7678 9764 7702 9766
rect 7758 9764 7782 9766
rect 7838 9764 7862 9766
rect 7622 9744 7918 9764
rect 7472 9648 7524 9654
rect 7472 9590 7524 9596
rect 7380 9580 7432 9586
rect 7380 9522 7432 9528
rect 7288 9444 7340 9450
rect 7288 9386 7340 9392
rect 7300 9353 7328 9386
rect 7932 9376 7984 9382
rect 7286 9344 7342 9353
rect 7932 9318 7984 9324
rect 7286 9279 7342 9288
rect 7944 9178 7972 9318
rect 7288 9172 7340 9178
rect 7288 9114 7340 9120
rect 7932 9172 7984 9178
rect 7932 9114 7984 9120
rect 7196 8288 7248 8294
rect 7300 8265 7328 9114
rect 7380 9104 7432 9110
rect 7378 9072 7380 9081
rect 7432 9072 7434 9081
rect 7378 9007 7434 9016
rect 8036 8809 8064 10152
rect 8128 9994 8156 11698
rect 8312 11665 8340 11834
rect 8298 11656 8354 11665
rect 8298 11591 8354 11600
rect 8300 11552 8352 11558
rect 8220 11512 8300 11540
rect 8116 9988 8168 9994
rect 8116 9930 8168 9936
rect 8114 9480 8170 9489
rect 8114 9415 8170 9424
rect 8128 9110 8156 9415
rect 8116 9104 8168 9110
rect 8116 9046 8168 9052
rect 8022 8800 8078 8809
rect 7622 8732 7918 8752
rect 8022 8735 8078 8744
rect 7678 8730 7702 8732
rect 7758 8730 7782 8732
rect 7838 8730 7862 8732
rect 7700 8678 7702 8730
rect 7764 8678 7776 8730
rect 7838 8678 7840 8730
rect 7678 8676 7702 8678
rect 7758 8676 7782 8678
rect 7838 8676 7862 8678
rect 7622 8656 7918 8676
rect 7840 8560 7892 8566
rect 7840 8502 7892 8508
rect 7472 8288 7524 8294
rect 7196 8230 7248 8236
rect 7286 8256 7342 8265
rect 7472 8230 7524 8236
rect 7562 8256 7618 8265
rect 7286 8191 7342 8200
rect 7484 8090 7512 8230
rect 7562 8191 7618 8200
rect 7472 8084 7524 8090
rect 7472 8026 7524 8032
rect 7116 7908 7328 7936
rect 6828 7812 6880 7818
rect 7024 7806 7236 7834
rect 6828 7754 6880 7760
rect 6734 7712 6790 7721
rect 6734 7647 6790 7656
rect 6644 7540 6696 7546
rect 6644 7482 6696 7488
rect 6748 7256 6776 7647
rect 6840 7585 6868 7754
rect 7012 7744 7064 7750
rect 7012 7686 7064 7692
rect 6826 7576 6882 7585
rect 6826 7511 6882 7520
rect 6828 7268 6880 7274
rect 6748 7228 6828 7256
rect 6828 7210 6880 7216
rect 6644 7200 6696 7206
rect 6550 7168 6606 7177
rect 6644 7142 6696 7148
rect 6550 7103 6606 7112
rect 6656 6866 6684 7142
rect 6644 6860 6696 6866
rect 6644 6802 6696 6808
rect 6840 6730 6868 7210
rect 7024 7206 7052 7686
rect 7012 7200 7064 7206
rect 7012 7142 7064 7148
rect 7012 6860 7064 6866
rect 7012 6802 7064 6808
rect 6828 6724 6880 6730
rect 6828 6666 6880 6672
rect 6840 6458 6868 6666
rect 6828 6452 6880 6458
rect 6828 6394 6880 6400
rect 7024 5409 7052 6802
rect 7104 6656 7156 6662
rect 7104 6598 7156 6604
rect 7116 5846 7144 6598
rect 7104 5840 7156 5846
rect 7104 5782 7156 5788
rect 7010 5400 7066 5409
rect 7116 5370 7144 5782
rect 7208 5642 7236 7806
rect 7300 6089 7328 7908
rect 7380 7540 7432 7546
rect 7484 7528 7512 8026
rect 7576 7857 7604 8191
rect 7852 8022 7880 8502
rect 8128 8294 8156 9046
rect 8220 8906 8248 11512
rect 8300 11494 8352 11500
rect 8404 11354 8432 13942
rect 9864 13864 9916 13870
rect 9864 13806 9916 13812
rect 9956 13864 10008 13870
rect 9956 13806 10008 13812
rect 8576 12232 8628 12238
rect 8576 12174 8628 12180
rect 8588 11626 8616 12174
rect 8944 12096 8996 12102
rect 8944 12038 8996 12044
rect 8576 11620 8628 11626
rect 8576 11562 8628 11568
rect 8956 11558 8984 12038
rect 8944 11552 8996 11558
rect 8944 11494 8996 11500
rect 9128 11552 9180 11558
rect 9128 11494 9180 11500
rect 8392 11348 8444 11354
rect 8392 11290 8444 11296
rect 8392 11212 8444 11218
rect 8392 11154 8444 11160
rect 8300 11144 8352 11150
rect 8300 11086 8352 11092
rect 8312 10606 8340 11086
rect 8404 10810 8432 11154
rect 8668 11144 8720 11150
rect 8668 11086 8720 11092
rect 8392 10804 8444 10810
rect 8392 10746 8444 10752
rect 8300 10600 8352 10606
rect 8300 10542 8352 10548
rect 8300 10192 8352 10198
rect 8300 10134 8352 10140
rect 8312 9382 8340 10134
rect 8484 10056 8536 10062
rect 8390 10024 8446 10033
rect 8484 9998 8536 10004
rect 8390 9959 8446 9968
rect 8300 9376 8352 9382
rect 8300 9318 8352 9324
rect 8208 8900 8260 8906
rect 8208 8842 8260 8848
rect 8116 8288 8168 8294
rect 8116 8230 8168 8236
rect 7840 8016 7892 8022
rect 7840 7958 7892 7964
rect 8024 7880 8076 7886
rect 7562 7848 7618 7857
rect 8024 7822 8076 7828
rect 8116 7880 8168 7886
rect 8116 7822 8168 7828
rect 8206 7848 8262 7857
rect 7562 7783 7618 7792
rect 7622 7644 7918 7664
rect 7678 7642 7702 7644
rect 7758 7642 7782 7644
rect 7838 7642 7862 7644
rect 7700 7590 7702 7642
rect 7764 7590 7776 7642
rect 7838 7590 7840 7642
rect 7678 7588 7702 7590
rect 7758 7588 7782 7590
rect 7838 7588 7862 7590
rect 7622 7568 7918 7588
rect 7484 7500 7604 7528
rect 7380 7482 7432 7488
rect 7392 7342 7420 7482
rect 7380 7336 7432 7342
rect 7380 7278 7432 7284
rect 7472 7336 7524 7342
rect 7472 7278 7524 7284
rect 7484 7002 7512 7278
rect 7576 7206 7604 7500
rect 8036 7342 8064 7822
rect 8128 7546 8156 7822
rect 8206 7783 8208 7792
rect 8260 7783 8262 7792
rect 8208 7754 8260 7760
rect 8312 7585 8340 9318
rect 8404 8430 8432 9959
rect 8496 9042 8524 9998
rect 8574 9616 8630 9625
rect 8574 9551 8630 9560
rect 8484 9036 8536 9042
rect 8484 8978 8536 8984
rect 8496 8673 8524 8978
rect 8588 8974 8616 9551
rect 8680 9450 8708 11086
rect 9140 11014 9168 11494
rect 9680 11144 9732 11150
rect 9680 11086 9732 11092
rect 9128 11008 9180 11014
rect 9128 10950 9180 10956
rect 9588 11008 9640 11014
rect 9588 10950 9640 10956
rect 9496 10736 9548 10742
rect 9494 10704 9496 10713
rect 9548 10704 9550 10713
rect 9494 10639 9550 10648
rect 9126 10432 9182 10441
rect 9126 10367 9182 10376
rect 9140 10266 9168 10367
rect 9128 10260 9180 10266
rect 9128 10202 9180 10208
rect 9140 9518 9168 10202
rect 9508 10198 9536 10639
rect 9600 10606 9628 10950
rect 9692 10674 9720 11086
rect 9680 10668 9732 10674
rect 9680 10610 9732 10616
rect 9588 10600 9640 10606
rect 9588 10542 9640 10548
rect 9496 10192 9548 10198
rect 9496 10134 9548 10140
rect 9600 9654 9628 10542
rect 9876 10266 9904 13806
rect 9968 11286 9996 13806
rect 10520 12714 10548 15520
rect 11704 13252 11756 13258
rect 11704 13194 11756 13200
rect 11716 12918 11744 13194
rect 11704 12912 11756 12918
rect 11704 12854 11756 12860
rect 12532 12776 12584 12782
rect 12532 12718 12584 12724
rect 10508 12708 10560 12714
rect 10508 12650 10560 12656
rect 11704 12368 11756 12374
rect 11704 12310 11756 12316
rect 11060 12096 11112 12102
rect 11060 12038 11112 12044
rect 10690 11928 10746 11937
rect 10690 11863 10692 11872
rect 10744 11863 10746 11872
rect 10968 11892 11020 11898
rect 10692 11834 10744 11840
rect 10968 11834 11020 11840
rect 10980 11370 11008 11834
rect 11072 11694 11100 12038
rect 11060 11688 11112 11694
rect 11060 11630 11112 11636
rect 11610 11656 11666 11665
rect 11610 11591 11666 11600
rect 10980 11342 11100 11370
rect 9956 11280 10008 11286
rect 9956 11222 10008 11228
rect 9968 10810 9996 11222
rect 10692 11212 10744 11218
rect 10692 11154 10744 11160
rect 9956 10804 10008 10810
rect 9956 10746 10008 10752
rect 10324 10532 10376 10538
rect 10324 10474 10376 10480
rect 10336 10305 10364 10474
rect 10322 10296 10378 10305
rect 9864 10260 9916 10266
rect 10322 10231 10324 10240
rect 9864 10202 9916 10208
rect 10376 10231 10378 10240
rect 10324 10202 10376 10208
rect 10508 10124 10560 10130
rect 10508 10066 10560 10072
rect 10520 9761 10548 10066
rect 10506 9752 10562 9761
rect 10506 9687 10508 9696
rect 10560 9687 10562 9696
rect 10508 9658 10560 9664
rect 9588 9648 9640 9654
rect 9588 9590 9640 9596
rect 9128 9512 9180 9518
rect 9128 9454 9180 9460
rect 8668 9444 8720 9450
rect 8720 9404 8800 9432
rect 8668 9386 8720 9392
rect 8772 9178 8800 9404
rect 8760 9172 8812 9178
rect 8760 9114 8812 9120
rect 8668 9104 8720 9110
rect 8668 9046 8720 9052
rect 8576 8968 8628 8974
rect 8576 8910 8628 8916
rect 8482 8664 8538 8673
rect 8588 8634 8616 8910
rect 8482 8599 8538 8608
rect 8576 8628 8628 8634
rect 8576 8570 8628 8576
rect 8392 8424 8444 8430
rect 8392 8366 8444 8372
rect 8404 8022 8432 8366
rect 8680 8090 8708 9046
rect 8772 8362 8800 9114
rect 9140 9110 9168 9454
rect 9678 9208 9734 9217
rect 9678 9143 9734 9152
rect 9128 9104 9180 9110
rect 9128 9046 9180 9052
rect 9692 8634 9720 9143
rect 10232 9104 10284 9110
rect 10232 9046 10284 9052
rect 10244 8673 10272 9046
rect 10324 8832 10376 8838
rect 10324 8774 10376 8780
rect 10230 8664 10286 8673
rect 9680 8628 9732 8634
rect 10230 8599 10232 8608
rect 9680 8570 9732 8576
rect 10284 8599 10286 8608
rect 10232 8570 10284 8576
rect 10336 8498 10364 8774
rect 10324 8492 10376 8498
rect 10324 8434 10376 8440
rect 8760 8356 8812 8362
rect 8760 8298 8812 8304
rect 8668 8084 8720 8090
rect 8668 8026 8720 8032
rect 8392 8016 8444 8022
rect 8392 7958 8444 7964
rect 8772 7886 8800 8298
rect 9312 8016 9364 8022
rect 9312 7958 9364 7964
rect 9680 8016 9732 8022
rect 9680 7958 9732 7964
rect 8760 7880 8812 7886
rect 8760 7822 8812 7828
rect 8298 7576 8354 7585
rect 8116 7540 8168 7546
rect 9324 7546 9352 7958
rect 8298 7511 8354 7520
rect 9312 7540 9364 7546
rect 8116 7482 8168 7488
rect 9312 7482 9364 7488
rect 8024 7336 8076 7342
rect 8024 7278 8076 7284
rect 7564 7200 7616 7206
rect 7564 7142 7616 7148
rect 7472 6996 7524 7002
rect 7472 6938 7524 6944
rect 7380 6860 7432 6866
rect 7380 6802 7432 6808
rect 7286 6080 7342 6089
rect 7286 6015 7342 6024
rect 7392 5914 7420 6802
rect 7472 6792 7524 6798
rect 7576 6769 7604 7142
rect 8128 7002 8156 7482
rect 9692 7206 9720 7958
rect 10336 7954 10364 8434
rect 10416 8424 10468 8430
rect 10416 8366 10468 8372
rect 10324 7948 10376 7954
rect 10324 7890 10376 7896
rect 10048 7880 10100 7886
rect 10048 7822 10100 7828
rect 9772 7744 9824 7750
rect 9772 7686 9824 7692
rect 9784 7449 9812 7686
rect 9770 7440 9826 7449
rect 9770 7375 9826 7384
rect 10060 7206 10088 7822
rect 9680 7200 9732 7206
rect 9680 7142 9732 7148
rect 10048 7200 10100 7206
rect 10140 7200 10192 7206
rect 10048 7142 10100 7148
rect 10138 7168 10140 7177
rect 10192 7168 10194 7177
rect 8116 6996 8168 7002
rect 8116 6938 8168 6944
rect 7472 6734 7524 6740
rect 7562 6760 7618 6769
rect 7380 5908 7432 5914
rect 7380 5850 7432 5856
rect 7196 5636 7248 5642
rect 7196 5578 7248 5584
rect 7010 5335 7012 5344
rect 7064 5335 7066 5344
rect 7104 5364 7156 5370
rect 7012 5306 7064 5312
rect 7104 5306 7156 5312
rect 7380 4616 7432 4622
rect 7380 4558 7432 4564
rect 7392 4434 7420 4558
rect 7484 4554 7512 6734
rect 7562 6695 7618 6704
rect 7622 6556 7918 6576
rect 7678 6554 7702 6556
rect 7758 6554 7782 6556
rect 7838 6554 7862 6556
rect 7700 6502 7702 6554
rect 7764 6502 7776 6554
rect 7838 6502 7840 6554
rect 7678 6500 7702 6502
rect 7758 6500 7782 6502
rect 7838 6500 7862 6502
rect 7622 6480 7918 6500
rect 8128 6458 8156 6938
rect 9692 6905 9720 7142
rect 9678 6896 9734 6905
rect 9312 6860 9364 6866
rect 9678 6831 9734 6840
rect 9312 6802 9364 6808
rect 8576 6792 8628 6798
rect 8576 6734 8628 6740
rect 8116 6452 8168 6458
rect 8116 6394 8168 6400
rect 7656 6180 7708 6186
rect 7656 6122 7708 6128
rect 7668 5953 7696 6122
rect 7654 5944 7710 5953
rect 7654 5879 7656 5888
rect 7708 5879 7710 5888
rect 7656 5850 7708 5856
rect 7622 5468 7918 5488
rect 7678 5466 7702 5468
rect 7758 5466 7782 5468
rect 7838 5466 7862 5468
rect 7700 5414 7702 5466
rect 7764 5414 7776 5466
rect 7838 5414 7840 5466
rect 7678 5412 7702 5414
rect 7758 5412 7782 5414
rect 7838 5412 7862 5414
rect 7622 5392 7918 5412
rect 8022 5400 8078 5409
rect 8128 5370 8156 6394
rect 8392 6112 8444 6118
rect 8392 6054 8444 6060
rect 8404 5846 8432 6054
rect 8588 5846 8616 6734
rect 9324 6118 9352 6802
rect 9680 6792 9732 6798
rect 9680 6734 9732 6740
rect 9496 6656 9548 6662
rect 9496 6598 9548 6604
rect 9508 6186 9536 6598
rect 9692 6254 9720 6734
rect 9772 6656 9824 6662
rect 9772 6598 9824 6604
rect 9680 6248 9732 6254
rect 9678 6216 9680 6225
rect 9732 6216 9734 6225
rect 9496 6180 9548 6186
rect 9678 6151 9734 6160
rect 9496 6122 9548 6128
rect 9312 6112 9364 6118
rect 9312 6054 9364 6060
rect 8392 5840 8444 5846
rect 8206 5808 8262 5817
rect 8392 5782 8444 5788
rect 8576 5840 8628 5846
rect 8576 5782 8628 5788
rect 8206 5743 8262 5752
rect 8220 5710 8248 5743
rect 8208 5704 8260 5710
rect 8208 5646 8260 5652
rect 8022 5335 8078 5344
rect 8116 5364 8168 5370
rect 8036 4622 8064 5335
rect 8116 5306 8168 5312
rect 8114 4992 8170 5001
rect 8114 4927 8170 4936
rect 8128 4758 8156 4927
rect 8220 4826 8248 5646
rect 8298 5536 8354 5545
rect 8298 5471 8354 5480
rect 8208 4820 8260 4826
rect 8208 4762 8260 4768
rect 8116 4752 8168 4758
rect 8116 4694 8168 4700
rect 8024 4616 8076 4622
rect 8024 4558 8076 4564
rect 7472 4548 7524 4554
rect 7472 4490 7524 4496
rect 7392 4406 7512 4434
rect 6458 4040 6514 4049
rect 6458 3975 6514 3984
rect 7484 3942 7512 4406
rect 7622 4380 7918 4400
rect 7678 4378 7702 4380
rect 7758 4378 7782 4380
rect 7838 4378 7862 4380
rect 7700 4326 7702 4378
rect 7764 4326 7776 4378
rect 7838 4326 7840 4378
rect 7678 4324 7702 4326
rect 7758 4324 7782 4326
rect 7838 4324 7862 4326
rect 7622 4304 7918 4324
rect 8128 4282 8156 4694
rect 8312 4690 8340 5471
rect 8404 5080 8432 5782
rect 8484 5092 8536 5098
rect 8404 5052 8484 5080
rect 8404 4826 8432 5052
rect 8484 5034 8536 5040
rect 8392 4820 8444 4826
rect 8392 4762 8444 4768
rect 8300 4684 8352 4690
rect 8300 4626 8352 4632
rect 8116 4276 8168 4282
rect 8116 4218 8168 4224
rect 8312 4146 8340 4626
rect 9324 4185 9352 6054
rect 9508 5642 9536 6122
rect 9784 6118 9812 6598
rect 9956 6384 10008 6390
rect 9956 6326 10008 6332
rect 9772 6112 9824 6118
rect 9772 6054 9824 6060
rect 9784 5914 9812 6054
rect 9772 5908 9824 5914
rect 9772 5850 9824 5856
rect 9864 5840 9916 5846
rect 9968 5817 9996 6326
rect 9864 5782 9916 5788
rect 9954 5808 10010 5817
rect 9496 5636 9548 5642
rect 9496 5578 9548 5584
rect 9772 5024 9824 5030
rect 9772 4966 9824 4972
rect 9784 4282 9812 4966
rect 9876 4826 9904 5782
rect 9954 5743 10010 5752
rect 10060 5681 10088 7142
rect 10138 7103 10194 7112
rect 10324 6792 10376 6798
rect 10324 6734 10376 6740
rect 10336 6254 10364 6734
rect 10324 6248 10376 6254
rect 10324 6190 10376 6196
rect 10336 5710 10364 6190
rect 10324 5704 10376 5710
rect 10046 5672 10102 5681
rect 10324 5646 10376 5652
rect 10046 5607 10102 5616
rect 10060 5137 10088 5607
rect 10336 5545 10364 5646
rect 10322 5536 10378 5545
rect 10322 5471 10378 5480
rect 10336 5370 10364 5471
rect 10324 5364 10376 5370
rect 10324 5306 10376 5312
rect 10046 5128 10102 5137
rect 10046 5063 10102 5072
rect 10428 4865 10456 8366
rect 10508 6928 10560 6934
rect 10508 6870 10560 6876
rect 10520 6769 10548 6870
rect 10506 6760 10562 6769
rect 10506 6695 10562 6704
rect 10598 6216 10654 6225
rect 10508 6180 10560 6186
rect 10598 6151 10654 6160
rect 10508 6122 10560 6128
rect 10520 5953 10548 6122
rect 10506 5944 10562 5953
rect 10506 5879 10508 5888
rect 10560 5879 10562 5888
rect 10508 5850 10560 5856
rect 10520 5819 10548 5850
rect 10612 5846 10640 6151
rect 10600 5840 10652 5846
rect 10600 5782 10652 5788
rect 10612 5030 10640 5782
rect 10600 5024 10652 5030
rect 10600 4966 10652 4972
rect 10414 4856 10470 4865
rect 9864 4820 9916 4826
rect 10414 4791 10470 4800
rect 9864 4762 9916 4768
rect 9772 4276 9824 4282
rect 9772 4218 9824 4224
rect 9310 4176 9366 4185
rect 8300 4140 8352 4146
rect 9310 4111 9366 4120
rect 8300 4082 8352 4088
rect 10612 3942 10640 4966
rect 10704 4554 10732 11154
rect 10782 11112 10838 11121
rect 10782 11047 10838 11056
rect 10796 10810 10824 11047
rect 10784 10804 10836 10810
rect 10784 10746 10836 10752
rect 11072 10606 11100 11342
rect 11152 11076 11204 11082
rect 11152 11018 11204 11024
rect 11060 10600 11112 10606
rect 11060 10542 11112 10548
rect 11164 10441 11192 11018
rect 11336 10532 11388 10538
rect 11336 10474 11388 10480
rect 11150 10432 11206 10441
rect 11150 10367 11206 10376
rect 11348 10198 11376 10474
rect 11336 10192 11388 10198
rect 11336 10134 11388 10140
rect 11520 10124 11572 10130
rect 11520 10066 11572 10072
rect 11532 9654 11560 10066
rect 11624 10033 11652 11591
rect 11716 11150 11744 12310
rect 11888 12232 11940 12238
rect 11888 12174 11940 12180
rect 12256 12232 12308 12238
rect 12256 12174 12308 12180
rect 11900 11218 11928 12174
rect 12268 11558 12296 12174
rect 12256 11552 12308 11558
rect 12256 11494 12308 11500
rect 11888 11212 11940 11218
rect 11888 11154 11940 11160
rect 11704 11144 11756 11150
rect 11702 11112 11704 11121
rect 11756 11112 11758 11121
rect 11702 11047 11758 11056
rect 11796 10464 11848 10470
rect 11796 10406 11848 10412
rect 11704 10192 11756 10198
rect 11704 10134 11756 10140
rect 11610 10024 11666 10033
rect 11610 9959 11666 9968
rect 11520 9648 11572 9654
rect 11520 9590 11572 9596
rect 10784 9376 10836 9382
rect 10784 9318 10836 9324
rect 10692 4548 10744 4554
rect 10692 4490 10744 4496
rect 10796 4078 10824 9318
rect 10874 8936 10930 8945
rect 10874 8871 10930 8880
rect 11334 8936 11390 8945
rect 11532 8906 11560 9590
rect 11624 8974 11652 9959
rect 11716 9382 11744 10134
rect 11808 10062 11836 10406
rect 12164 10124 12216 10130
rect 12164 10066 12216 10072
rect 11796 10056 11848 10062
rect 11796 9998 11848 10004
rect 11808 9722 11836 9998
rect 11796 9716 11848 9722
rect 11796 9658 11848 9664
rect 12176 9382 12204 10066
rect 12268 9738 12296 11494
rect 12440 11280 12492 11286
rect 12360 11228 12440 11234
rect 12360 11222 12492 11228
rect 12360 11206 12480 11222
rect 12360 9994 12388 11206
rect 12544 11082 12572 12718
rect 12820 11762 12848 15520
rect 14289 13628 14585 13648
rect 14345 13626 14369 13628
rect 14425 13626 14449 13628
rect 14505 13626 14529 13628
rect 14367 13574 14369 13626
rect 14431 13574 14443 13626
rect 14505 13574 14507 13626
rect 14345 13572 14369 13574
rect 14425 13572 14449 13574
rect 14505 13572 14529 13574
rect 14289 13552 14585 13572
rect 15212 12850 15240 15520
rect 17224 13456 17276 13462
rect 17224 13398 17276 13404
rect 15200 12844 15252 12850
rect 15200 12786 15252 12792
rect 16856 12776 16908 12782
rect 16856 12718 16908 12724
rect 12900 12708 12952 12714
rect 12900 12650 12952 12656
rect 12808 11756 12860 11762
rect 12808 11698 12860 11704
rect 12624 11552 12676 11558
rect 12624 11494 12676 11500
rect 12532 11076 12584 11082
rect 12532 11018 12584 11024
rect 12348 9988 12400 9994
rect 12348 9930 12400 9936
rect 12268 9710 12572 9738
rect 11704 9376 11756 9382
rect 11704 9318 11756 9324
rect 11980 9376 12032 9382
rect 11980 9318 12032 9324
rect 12164 9376 12216 9382
rect 12164 9318 12216 9324
rect 11704 9104 11756 9110
rect 11704 9046 11756 9052
rect 11612 8968 11664 8974
rect 11612 8910 11664 8916
rect 11334 8871 11390 8880
rect 11520 8900 11572 8906
rect 10888 8634 10916 8871
rect 10876 8628 10928 8634
rect 10876 8570 10928 8576
rect 11348 8362 11376 8871
rect 11520 8842 11572 8848
rect 11624 8634 11652 8910
rect 11716 8673 11744 9046
rect 11702 8664 11758 8673
rect 11612 8628 11664 8634
rect 11702 8599 11758 8608
rect 11612 8570 11664 8576
rect 10968 8356 11020 8362
rect 10968 8298 11020 8304
rect 11336 8356 11388 8362
rect 11336 8298 11388 8304
rect 10980 8090 11008 8298
rect 10968 8084 11020 8090
rect 10888 8044 10968 8072
rect 10888 5409 10916 8044
rect 10968 8026 11020 8032
rect 11716 8004 11744 8599
rect 11888 8424 11940 8430
rect 11888 8366 11940 8372
rect 11900 8022 11928 8366
rect 11888 8016 11940 8022
rect 11716 7976 11836 8004
rect 11520 7948 11572 7954
rect 11572 7908 11744 7936
rect 11520 7890 11572 7896
rect 11334 7712 11390 7721
rect 11334 7647 11390 7656
rect 10968 7472 11020 7478
rect 10968 7414 11020 7420
rect 10874 5400 10930 5409
rect 10874 5335 10930 5344
rect 10888 5001 10916 5335
rect 10874 4992 10930 5001
rect 10874 4927 10930 4936
rect 10980 4865 11008 7414
rect 11244 7336 11296 7342
rect 11244 7278 11296 7284
rect 11060 7268 11112 7274
rect 11060 7210 11112 7216
rect 11072 6934 11100 7210
rect 11256 7002 11284 7278
rect 11348 7274 11376 7647
rect 11336 7268 11388 7274
rect 11336 7210 11388 7216
rect 11244 6996 11296 7002
rect 11244 6938 11296 6944
rect 11060 6928 11112 6934
rect 11058 6896 11060 6905
rect 11112 6896 11114 6905
rect 11058 6831 11114 6840
rect 11336 6860 11388 6866
rect 11336 6802 11388 6808
rect 11428 6860 11480 6866
rect 11428 6802 11480 6808
rect 11152 6724 11204 6730
rect 11152 6666 11204 6672
rect 11060 5568 11112 5574
rect 11060 5510 11112 5516
rect 10966 4856 11022 4865
rect 10966 4791 11022 4800
rect 10968 4752 11020 4758
rect 10968 4694 11020 4700
rect 10876 4616 10928 4622
rect 10876 4558 10928 4564
rect 10888 4214 10916 4558
rect 10876 4208 10928 4214
rect 10876 4150 10928 4156
rect 10784 4072 10836 4078
rect 10784 4014 10836 4020
rect 7472 3936 7524 3942
rect 7472 3878 7524 3884
rect 10324 3936 10376 3942
rect 10324 3878 10376 3884
rect 10600 3936 10652 3942
rect 10600 3878 10652 3884
rect 7484 2961 7512 3878
rect 9588 3732 9640 3738
rect 9640 3692 9720 3720
rect 9588 3674 9640 3680
rect 9692 3534 9720 3692
rect 9680 3528 9732 3534
rect 9680 3470 9732 3476
rect 7622 3292 7918 3312
rect 7678 3290 7702 3292
rect 7758 3290 7782 3292
rect 7838 3290 7862 3292
rect 7700 3238 7702 3290
rect 7764 3238 7776 3290
rect 7838 3238 7840 3290
rect 7678 3236 7702 3238
rect 7758 3236 7782 3238
rect 7838 3236 7862 3238
rect 7622 3216 7918 3236
rect 10336 3194 10364 3878
rect 10612 3641 10640 3878
rect 10796 3738 10824 4014
rect 10980 4010 11008 4694
rect 11072 4622 11100 5510
rect 11060 4616 11112 4622
rect 11060 4558 11112 4564
rect 11072 4049 11100 4558
rect 11164 4457 11192 6666
rect 11348 6458 11376 6802
rect 11336 6452 11388 6458
rect 11336 6394 11388 6400
rect 11440 5914 11468 6802
rect 11716 6662 11744 7908
rect 11704 6656 11756 6662
rect 11704 6598 11756 6604
rect 11428 5908 11480 5914
rect 11428 5850 11480 5856
rect 11150 4448 11206 4457
rect 11150 4383 11206 4392
rect 11058 4040 11114 4049
rect 10968 4004 11020 4010
rect 11058 3975 11114 3984
rect 10968 3946 11020 3952
rect 10784 3732 10836 3738
rect 10784 3674 10836 3680
rect 10598 3632 10654 3641
rect 10598 3567 10654 3576
rect 10980 3466 11008 3946
rect 11072 3670 11100 3975
rect 11164 3670 11192 4383
rect 11440 4321 11468 5850
rect 11716 5574 11744 6598
rect 11808 6458 11836 7976
rect 11888 7958 11940 7964
rect 11900 7546 11928 7958
rect 11992 7546 12020 9318
rect 12176 9042 12204 9318
rect 12164 9036 12216 9042
rect 12164 8978 12216 8984
rect 12176 8838 12204 8978
rect 12164 8832 12216 8838
rect 12164 8774 12216 8780
rect 12544 8362 12572 9710
rect 12636 9489 12664 11494
rect 12808 11212 12860 11218
rect 12808 11154 12860 11160
rect 12716 10600 12768 10606
rect 12716 10542 12768 10548
rect 12728 10062 12756 10542
rect 12716 10056 12768 10062
rect 12716 9998 12768 10004
rect 12728 9518 12756 9998
rect 12716 9512 12768 9518
rect 12622 9480 12678 9489
rect 12716 9454 12768 9460
rect 12622 9415 12678 9424
rect 12820 8906 12848 11154
rect 12808 8900 12860 8906
rect 12808 8842 12860 8848
rect 12532 8356 12584 8362
rect 12532 8298 12584 8304
rect 12544 8090 12572 8298
rect 12532 8084 12584 8090
rect 12532 8026 12584 8032
rect 12162 7576 12218 7585
rect 11888 7540 11940 7546
rect 11888 7482 11940 7488
rect 11980 7540 12032 7546
rect 12162 7511 12218 7520
rect 11980 7482 12032 7488
rect 11900 6934 11928 7482
rect 12176 7410 12204 7511
rect 12164 7404 12216 7410
rect 12164 7346 12216 7352
rect 12176 7256 12204 7346
rect 12256 7268 12308 7274
rect 12176 7228 12256 7256
rect 11888 6928 11940 6934
rect 11888 6870 11940 6876
rect 12176 6458 12204 7228
rect 12256 7210 12308 7216
rect 12532 6928 12584 6934
rect 12532 6870 12584 6876
rect 11796 6452 11848 6458
rect 11796 6394 11848 6400
rect 12164 6452 12216 6458
rect 12164 6394 12216 6400
rect 11808 6254 11836 6394
rect 11796 6248 11848 6254
rect 11796 6190 11848 6196
rect 12176 6118 12204 6394
rect 12440 6384 12492 6390
rect 12544 6361 12572 6870
rect 12806 6624 12862 6633
rect 12806 6559 12862 6568
rect 12440 6326 12492 6332
rect 12530 6352 12586 6361
rect 12164 6112 12216 6118
rect 12164 6054 12216 6060
rect 12348 5772 12400 5778
rect 12348 5714 12400 5720
rect 11704 5568 11756 5574
rect 11704 5510 11756 5516
rect 12256 5092 12308 5098
rect 12256 5034 12308 5040
rect 11980 5024 12032 5030
rect 11980 4966 12032 4972
rect 11426 4312 11482 4321
rect 11426 4247 11482 4256
rect 11440 4078 11468 4247
rect 11428 4072 11480 4078
rect 11428 4014 11480 4020
rect 11060 3664 11112 3670
rect 11060 3606 11112 3612
rect 11152 3664 11204 3670
rect 11152 3606 11204 3612
rect 10968 3460 11020 3466
rect 10968 3402 11020 3408
rect 10324 3188 10376 3194
rect 10324 3130 10376 3136
rect 11164 3126 11192 3606
rect 11440 3602 11468 4014
rect 11704 3664 11756 3670
rect 11702 3632 11704 3641
rect 11756 3632 11758 3641
rect 11428 3596 11480 3602
rect 11428 3538 11480 3544
rect 11624 3590 11702 3618
rect 11440 3194 11468 3538
rect 11624 3194 11652 3590
rect 11702 3567 11758 3576
rect 11716 3507 11744 3567
rect 11992 3505 12020 4966
rect 12070 4720 12126 4729
rect 12070 4655 12126 4664
rect 12084 4486 12112 4655
rect 12072 4480 12124 4486
rect 12072 4422 12124 4428
rect 12268 4282 12296 5034
rect 12360 5030 12388 5714
rect 12348 5024 12400 5030
rect 12348 4966 12400 4972
rect 12452 4622 12480 6326
rect 12530 6287 12586 6296
rect 12532 5840 12584 5846
rect 12532 5782 12584 5788
rect 12440 4616 12492 4622
rect 12440 4558 12492 4564
rect 12544 4282 12572 5782
rect 12820 5778 12848 6559
rect 12808 5772 12860 5778
rect 12808 5714 12860 5720
rect 12716 5704 12768 5710
rect 12716 5646 12768 5652
rect 12728 5370 12756 5646
rect 12716 5364 12768 5370
rect 12716 5306 12768 5312
rect 12728 4826 12756 5306
rect 12806 4856 12862 4865
rect 12716 4820 12768 4826
rect 12806 4791 12862 4800
rect 12716 4762 12768 4768
rect 12728 4622 12756 4762
rect 12716 4616 12768 4622
rect 12716 4558 12768 4564
rect 12256 4276 12308 4282
rect 12256 4218 12308 4224
rect 12532 4276 12584 4282
rect 12532 4218 12584 4224
rect 12530 4176 12586 4185
rect 12530 4111 12586 4120
rect 12348 4072 12400 4078
rect 12348 4014 12400 4020
rect 12164 3936 12216 3942
rect 12162 3904 12164 3913
rect 12216 3904 12218 3913
rect 12162 3839 12218 3848
rect 11978 3496 12034 3505
rect 11978 3431 12034 3440
rect 11428 3188 11480 3194
rect 11428 3130 11480 3136
rect 11612 3188 11664 3194
rect 11612 3130 11664 3136
rect 11152 3120 11204 3126
rect 11152 3062 11204 3068
rect 7470 2952 7526 2961
rect 7470 2887 7526 2896
rect 11624 2825 11652 3130
rect 12360 3097 12388 4014
rect 12544 4010 12572 4111
rect 12532 4004 12584 4010
rect 12532 3946 12584 3952
rect 12544 3398 12572 3946
rect 12532 3392 12584 3398
rect 12532 3334 12584 3340
rect 12346 3088 12402 3097
rect 12346 3023 12402 3032
rect 11610 2816 11666 2825
rect 11610 2751 11666 2760
rect 6366 2544 6422 2553
rect 6366 2479 6422 2488
rect 7622 2204 7918 2224
rect 7678 2202 7702 2204
rect 7758 2202 7782 2204
rect 7838 2202 7862 2204
rect 7700 2150 7702 2202
rect 7764 2150 7776 2202
rect 7838 2150 7840 2202
rect 7678 2148 7702 2150
rect 7758 2148 7782 2150
rect 7838 2148 7862 2150
rect 7622 2128 7918 2148
rect 12544 1873 12572 3334
rect 12820 2990 12848 4791
rect 12912 3466 12940 12650
rect 16212 12640 16264 12646
rect 16212 12582 16264 12588
rect 14289 12540 14585 12560
rect 14345 12538 14369 12540
rect 14425 12538 14449 12540
rect 14505 12538 14529 12540
rect 14367 12486 14369 12538
rect 14431 12486 14443 12538
rect 14505 12486 14507 12538
rect 14345 12484 14369 12486
rect 14425 12484 14449 12486
rect 14505 12484 14529 12486
rect 14289 12464 14585 12484
rect 12992 12096 13044 12102
rect 12992 12038 13044 12044
rect 15844 12096 15896 12102
rect 15844 12038 15896 12044
rect 13004 11626 13032 12038
rect 13176 11824 13228 11830
rect 13176 11766 13228 11772
rect 12992 11620 13044 11626
rect 12992 11562 13044 11568
rect 13004 9625 13032 11562
rect 13084 11144 13136 11150
rect 13084 11086 13136 11092
rect 13096 10470 13124 11086
rect 13084 10464 13136 10470
rect 13084 10406 13136 10412
rect 13096 10266 13124 10406
rect 13084 10260 13136 10266
rect 13084 10202 13136 10208
rect 12990 9616 13046 9625
rect 12990 9551 13046 9560
rect 13188 7274 13216 11766
rect 13452 11688 13504 11694
rect 13452 11630 13504 11636
rect 13464 9450 13492 11630
rect 15856 11626 15884 12038
rect 15844 11620 15896 11626
rect 15844 11562 15896 11568
rect 14289 11452 14585 11472
rect 14345 11450 14369 11452
rect 14425 11450 14449 11452
rect 14505 11450 14529 11452
rect 14367 11398 14369 11450
rect 14431 11398 14443 11450
rect 14505 11398 14507 11450
rect 14345 11396 14369 11398
rect 14425 11396 14449 11398
rect 14505 11396 14529 11398
rect 14289 11376 14585 11396
rect 15108 11348 15160 11354
rect 15108 11290 15160 11296
rect 15120 11257 15148 11290
rect 15106 11248 15162 11257
rect 15106 11183 15162 11192
rect 15750 11248 15806 11257
rect 15750 11183 15806 11192
rect 13910 11112 13966 11121
rect 13910 11047 13966 11056
rect 13544 10532 13596 10538
rect 13544 10474 13596 10480
rect 13556 9874 13584 10474
rect 13728 10056 13780 10062
rect 13728 9998 13780 10004
rect 13636 9920 13688 9926
rect 13556 9868 13636 9874
rect 13556 9862 13688 9868
rect 13556 9846 13676 9862
rect 13452 9444 13504 9450
rect 13452 9386 13504 9392
rect 13360 9376 13412 9382
rect 13360 9318 13412 9324
rect 13266 9072 13322 9081
rect 13266 9007 13322 9016
rect 13280 8974 13308 9007
rect 13268 8968 13320 8974
rect 13268 8910 13320 8916
rect 13268 8832 13320 8838
rect 13372 8820 13400 9318
rect 13464 9178 13492 9386
rect 13452 9172 13504 9178
rect 13452 9114 13504 9120
rect 13556 8974 13584 9846
rect 13634 9480 13690 9489
rect 13740 9450 13768 9998
rect 13634 9415 13690 9424
rect 13728 9444 13780 9450
rect 13544 8968 13596 8974
rect 13544 8910 13596 8916
rect 13320 8792 13400 8820
rect 13268 8774 13320 8780
rect 13280 7274 13308 8774
rect 13556 8090 13584 8910
rect 13544 8084 13596 8090
rect 13544 8026 13596 8032
rect 13358 7576 13414 7585
rect 13648 7562 13676 9415
rect 13728 9386 13780 9392
rect 13726 7984 13782 7993
rect 13726 7919 13728 7928
rect 13780 7919 13782 7928
rect 13728 7890 13780 7896
rect 13648 7534 13768 7562
rect 13358 7511 13414 7520
rect 13372 7410 13400 7511
rect 13636 7472 13688 7478
rect 13636 7414 13688 7420
rect 13360 7404 13412 7410
rect 13360 7346 13412 7352
rect 13176 7268 13228 7274
rect 13176 7210 13228 7216
rect 13268 7268 13320 7274
rect 13268 7210 13320 7216
rect 13188 7002 13216 7210
rect 13176 6996 13228 7002
rect 13176 6938 13228 6944
rect 13280 6934 13308 7210
rect 13268 6928 13320 6934
rect 13268 6870 13320 6876
rect 13542 6352 13598 6361
rect 13542 6287 13598 6296
rect 13556 6254 13584 6287
rect 12992 6248 13044 6254
rect 12992 6190 13044 6196
rect 13544 6248 13596 6254
rect 13544 6190 13596 6196
rect 13004 5098 13032 6190
rect 13450 5536 13506 5545
rect 13450 5471 13506 5480
rect 13174 5400 13230 5409
rect 13174 5335 13230 5344
rect 13188 5137 13216 5335
rect 13174 5128 13230 5137
rect 12992 5092 13044 5098
rect 13174 5063 13230 5072
rect 12992 5034 13044 5040
rect 13004 4826 13032 5034
rect 12992 4820 13044 4826
rect 12992 4762 13044 4768
rect 13004 4622 13032 4762
rect 12992 4616 13044 4622
rect 12992 4558 13044 4564
rect 13004 4146 13032 4558
rect 12992 4140 13044 4146
rect 12992 4082 13044 4088
rect 12992 3936 13044 3942
rect 12992 3878 13044 3884
rect 13176 3936 13228 3942
rect 13176 3878 13228 3884
rect 13004 3641 13032 3878
rect 12990 3632 13046 3641
rect 12990 3567 13046 3576
rect 13188 3534 13216 3878
rect 13464 3534 13492 5471
rect 13556 5166 13584 6190
rect 13544 5160 13596 5166
rect 13544 5102 13596 5108
rect 13544 5024 13596 5030
rect 13544 4966 13596 4972
rect 13176 3528 13228 3534
rect 13176 3470 13228 3476
rect 13360 3528 13412 3534
rect 13360 3470 13412 3476
rect 13452 3528 13504 3534
rect 13452 3470 13504 3476
rect 12900 3460 12952 3466
rect 12900 3402 12952 3408
rect 13372 3126 13400 3470
rect 13464 3194 13492 3470
rect 13452 3188 13504 3194
rect 13452 3130 13504 3136
rect 13360 3120 13412 3126
rect 13360 3062 13412 3068
rect 12808 2984 12860 2990
rect 12808 2926 12860 2932
rect 12820 2582 12848 2926
rect 12900 2916 12952 2922
rect 12900 2858 12952 2864
rect 12912 2650 12940 2858
rect 13372 2650 13400 3062
rect 13556 3058 13584 4966
rect 13544 3052 13596 3058
rect 13544 2994 13596 3000
rect 13648 2990 13676 7414
rect 13740 5658 13768 7534
rect 13818 6896 13874 6905
rect 13818 6831 13820 6840
rect 13872 6831 13874 6840
rect 13820 6802 13872 6808
rect 13740 5630 13860 5658
rect 13728 5568 13780 5574
rect 13728 5510 13780 5516
rect 13740 3738 13768 5510
rect 13832 4826 13860 5630
rect 13820 4820 13872 4826
rect 13820 4762 13872 4768
rect 13832 4214 13860 4762
rect 13924 4282 13952 11047
rect 15016 11008 15068 11014
rect 15016 10950 15068 10956
rect 15028 10742 15056 10950
rect 15120 10810 15148 11183
rect 15764 11150 15792 11183
rect 15856 11150 15884 11562
rect 16224 11558 16252 12582
rect 16488 11824 16540 11830
rect 16488 11766 16540 11772
rect 15936 11552 15988 11558
rect 15936 11494 15988 11500
rect 16212 11552 16264 11558
rect 16212 11494 16264 11500
rect 15948 11286 15976 11494
rect 16500 11393 16528 11766
rect 16486 11384 16542 11393
rect 16028 11348 16080 11354
rect 16486 11319 16542 11328
rect 16028 11290 16080 11296
rect 15936 11280 15988 11286
rect 15936 11222 15988 11228
rect 15752 11144 15804 11150
rect 15752 11086 15804 11092
rect 15844 11144 15896 11150
rect 15844 11086 15896 11092
rect 15108 10804 15160 10810
rect 15108 10746 15160 10752
rect 14096 10736 14148 10742
rect 14096 10678 14148 10684
rect 15016 10736 15068 10742
rect 15016 10678 15068 10684
rect 14004 9172 14056 9178
rect 14004 9114 14056 9120
rect 14016 8634 14044 9114
rect 14004 8628 14056 8634
rect 14004 8570 14056 8576
rect 14108 8265 14136 10678
rect 15108 10600 15160 10606
rect 15108 10542 15160 10548
rect 14289 10364 14585 10384
rect 14345 10362 14369 10364
rect 14425 10362 14449 10364
rect 14505 10362 14529 10364
rect 14367 10310 14369 10362
rect 14431 10310 14443 10362
rect 14505 10310 14507 10362
rect 14345 10308 14369 10310
rect 14425 10308 14449 10310
rect 14505 10308 14529 10310
rect 14289 10288 14585 10308
rect 15120 10062 15148 10542
rect 15292 10192 15344 10198
rect 15292 10134 15344 10140
rect 15108 10056 15160 10062
rect 15108 9998 15160 10004
rect 15304 9761 15332 10134
rect 15660 10124 15712 10130
rect 15660 10066 15712 10072
rect 15384 9920 15436 9926
rect 15384 9862 15436 9868
rect 15290 9752 15346 9761
rect 15290 9687 15292 9696
rect 15344 9687 15346 9696
rect 15292 9658 15344 9664
rect 14186 9616 14242 9625
rect 14186 9551 14242 9560
rect 14094 8256 14150 8265
rect 14094 8191 14150 8200
rect 14094 8120 14150 8129
rect 14094 8055 14150 8064
rect 14108 7750 14136 8055
rect 14096 7744 14148 7750
rect 14096 7686 14148 7692
rect 14200 7562 14228 9551
rect 14924 9376 14976 9382
rect 14924 9318 14976 9324
rect 14289 9276 14585 9296
rect 14345 9274 14369 9276
rect 14425 9274 14449 9276
rect 14505 9274 14529 9276
rect 14367 9222 14369 9274
rect 14431 9222 14443 9274
rect 14505 9222 14507 9274
rect 14345 9220 14369 9222
rect 14425 9220 14449 9222
rect 14505 9220 14529 9222
rect 14289 9200 14585 9220
rect 14936 9178 14964 9318
rect 14924 9172 14976 9178
rect 14924 9114 14976 9120
rect 14936 8634 14964 9114
rect 15396 9081 15424 9862
rect 15672 9382 15700 10066
rect 15936 10056 15988 10062
rect 15936 9998 15988 10004
rect 15660 9376 15712 9382
rect 15660 9318 15712 9324
rect 15382 9072 15438 9081
rect 15382 9007 15438 9016
rect 15292 8968 15344 8974
rect 15292 8910 15344 8916
rect 14924 8628 14976 8634
rect 14924 8570 14976 8576
rect 15304 8401 15332 8910
rect 15290 8392 15346 8401
rect 15290 8327 15292 8336
rect 15344 8327 15346 8336
rect 15292 8298 15344 8304
rect 14289 8188 14585 8208
rect 14345 8186 14369 8188
rect 14425 8186 14449 8188
rect 14505 8186 14529 8188
rect 14367 8134 14369 8186
rect 14431 8134 14443 8186
rect 14505 8134 14507 8186
rect 14345 8132 14369 8134
rect 14425 8132 14449 8134
rect 14505 8132 14529 8134
rect 14289 8112 14585 8132
rect 15672 7993 15700 9318
rect 15752 9104 15804 9110
rect 15752 9046 15804 9052
rect 15764 8566 15792 9046
rect 15948 9042 15976 9998
rect 16040 9761 16068 11290
rect 16868 11082 16896 12718
rect 16948 11756 17000 11762
rect 16948 11698 17000 11704
rect 16960 11354 16988 11698
rect 17130 11656 17186 11665
rect 17130 11591 17186 11600
rect 17144 11558 17172 11591
rect 17132 11552 17184 11558
rect 17132 11494 17184 11500
rect 16948 11348 17000 11354
rect 16948 11290 17000 11296
rect 17132 11144 17184 11150
rect 17132 11086 17184 11092
rect 16856 11076 16908 11082
rect 16856 11018 16908 11024
rect 16948 10600 17000 10606
rect 16948 10542 17000 10548
rect 16488 10464 16540 10470
rect 16488 10406 16540 10412
rect 16500 10266 16528 10406
rect 16488 10260 16540 10266
rect 16488 10202 16540 10208
rect 16026 9752 16082 9761
rect 16026 9687 16082 9696
rect 16580 9444 16632 9450
rect 16580 9386 16632 9392
rect 15936 9036 15988 9042
rect 15936 8978 15988 8984
rect 16592 8838 16620 9386
rect 16960 8945 16988 10542
rect 17144 10470 17172 11086
rect 17132 10464 17184 10470
rect 17132 10406 17184 10412
rect 17040 10192 17092 10198
rect 17040 10134 17092 10140
rect 17052 9586 17080 10134
rect 17144 9586 17172 10406
rect 17040 9580 17092 9586
rect 17040 9522 17092 9528
rect 17132 9580 17184 9586
rect 17132 9522 17184 9528
rect 17052 9178 17080 9522
rect 17040 9172 17092 9178
rect 17040 9114 17092 9120
rect 16946 8936 17002 8945
rect 16946 8871 17002 8880
rect 16580 8832 16632 8838
rect 16580 8774 16632 8780
rect 16948 8832 17000 8838
rect 16948 8774 17000 8780
rect 15752 8560 15804 8566
rect 15750 8528 15752 8537
rect 16396 8560 16448 8566
rect 15804 8528 15806 8537
rect 16396 8502 16448 8508
rect 15750 8463 15806 8472
rect 16304 8356 16356 8362
rect 16304 8298 16356 8304
rect 16210 8120 16266 8129
rect 16210 8055 16266 8064
rect 15658 7984 15714 7993
rect 15658 7919 15714 7928
rect 15936 7880 15988 7886
rect 15936 7822 15988 7828
rect 14648 7744 14700 7750
rect 14648 7686 14700 7692
rect 14016 7534 14228 7562
rect 14016 4758 14044 7534
rect 14096 7404 14148 7410
rect 14096 7346 14148 7352
rect 14108 7041 14136 7346
rect 14660 7290 14688 7686
rect 15948 7546 15976 7822
rect 16224 7818 16252 8055
rect 16212 7812 16264 7818
rect 16212 7754 16264 7760
rect 15936 7540 15988 7546
rect 15936 7482 15988 7488
rect 14738 7440 14794 7449
rect 14738 7375 14740 7384
rect 14792 7375 14794 7384
rect 16212 7404 16264 7410
rect 14740 7346 14792 7352
rect 16212 7346 16264 7352
rect 14660 7262 14780 7290
rect 14752 7206 14780 7262
rect 14832 7268 14884 7274
rect 14832 7210 14884 7216
rect 14740 7200 14792 7206
rect 14738 7168 14740 7177
rect 14792 7168 14794 7177
rect 14289 7100 14585 7120
rect 14738 7103 14794 7112
rect 14345 7098 14369 7100
rect 14425 7098 14449 7100
rect 14505 7098 14529 7100
rect 14367 7046 14369 7098
rect 14431 7046 14443 7098
rect 14505 7046 14507 7098
rect 14345 7044 14369 7046
rect 14425 7044 14449 7046
rect 14505 7044 14529 7046
rect 14094 7032 14150 7041
rect 14289 7024 14585 7044
rect 14844 7002 14872 7210
rect 16224 7206 16252 7346
rect 16212 7200 16264 7206
rect 16212 7142 16264 7148
rect 14094 6967 14150 6976
rect 14832 6996 14884 7002
rect 14832 6938 14884 6944
rect 14844 6186 14872 6938
rect 16224 6905 16252 7142
rect 16210 6896 16266 6905
rect 16210 6831 16266 6840
rect 15568 6384 15620 6390
rect 15568 6326 15620 6332
rect 15580 6254 15608 6326
rect 15568 6248 15620 6254
rect 15568 6190 15620 6196
rect 14832 6180 14884 6186
rect 14832 6122 14884 6128
rect 14289 6012 14585 6032
rect 14345 6010 14369 6012
rect 14425 6010 14449 6012
rect 14505 6010 14529 6012
rect 14367 5958 14369 6010
rect 14431 5958 14443 6010
rect 14505 5958 14507 6010
rect 14345 5956 14369 5958
rect 14425 5956 14449 5958
rect 14505 5956 14529 5958
rect 14289 5936 14585 5956
rect 14740 5840 14792 5846
rect 14740 5782 14792 5788
rect 14188 5704 14240 5710
rect 14188 5646 14240 5652
rect 14200 5030 14228 5646
rect 14648 5296 14700 5302
rect 14648 5238 14700 5244
rect 14188 5024 14240 5030
rect 14188 4966 14240 4972
rect 14289 4924 14585 4944
rect 14345 4922 14369 4924
rect 14425 4922 14449 4924
rect 14505 4922 14529 4924
rect 14367 4870 14369 4922
rect 14431 4870 14443 4922
rect 14505 4870 14507 4922
rect 14345 4868 14369 4870
rect 14425 4868 14449 4870
rect 14505 4868 14529 4870
rect 14289 4848 14585 4868
rect 14660 4826 14688 5238
rect 14752 5030 14780 5782
rect 14844 5370 14872 6122
rect 15476 5704 15528 5710
rect 15580 5692 15608 6190
rect 15752 6112 15804 6118
rect 15752 6054 15804 6060
rect 15764 5778 15792 6054
rect 15752 5772 15804 5778
rect 15752 5714 15804 5720
rect 15528 5664 15608 5692
rect 15476 5646 15528 5652
rect 15580 5370 15608 5664
rect 14832 5364 14884 5370
rect 14832 5306 14884 5312
rect 15568 5364 15620 5370
rect 15568 5306 15620 5312
rect 16224 5273 16252 6831
rect 16316 6633 16344 8298
rect 16408 7342 16436 8502
rect 16488 7948 16540 7954
rect 16488 7890 16540 7896
rect 16500 7546 16528 7890
rect 16488 7540 16540 7546
rect 16488 7482 16540 7488
rect 16396 7336 16448 7342
rect 16396 7278 16448 7284
rect 16302 6624 16358 6633
rect 16302 6559 16358 6568
rect 16592 5953 16620 8774
rect 16960 8498 16988 8774
rect 16948 8492 17000 8498
rect 16948 8434 17000 8440
rect 16672 8016 16724 8022
rect 16672 7958 16724 7964
rect 16684 6934 16712 7958
rect 16960 7177 16988 8434
rect 17236 8362 17264 13398
rect 17604 12850 17632 15520
rect 19904 12850 19932 15520
rect 20956 13084 21252 13104
rect 21012 13082 21036 13084
rect 21092 13082 21116 13084
rect 21172 13082 21196 13084
rect 21034 13030 21036 13082
rect 21098 13030 21110 13082
rect 21172 13030 21174 13082
rect 21012 13028 21036 13030
rect 21092 13028 21116 13030
rect 21172 13028 21196 13030
rect 20956 13008 21252 13028
rect 19984 12912 20036 12918
rect 19984 12854 20036 12860
rect 17592 12844 17644 12850
rect 17592 12786 17644 12792
rect 19892 12844 19944 12850
rect 19892 12786 19944 12792
rect 19340 12776 19392 12782
rect 19340 12718 19392 12724
rect 17868 12368 17920 12374
rect 17868 12310 17920 12316
rect 17776 12232 17828 12238
rect 17776 12174 17828 12180
rect 17500 12164 17552 12170
rect 17500 12106 17552 12112
rect 17408 12096 17460 12102
rect 17408 12038 17460 12044
rect 17420 11354 17448 12038
rect 17512 11898 17540 12106
rect 17500 11892 17552 11898
rect 17500 11834 17552 11840
rect 17512 11354 17540 11834
rect 17788 11626 17816 12174
rect 17684 11620 17736 11626
rect 17684 11562 17736 11568
rect 17776 11620 17828 11626
rect 17776 11562 17828 11568
rect 17408 11348 17460 11354
rect 17408 11290 17460 11296
rect 17500 11348 17552 11354
rect 17500 11290 17552 11296
rect 17696 11150 17724 11562
rect 17880 11558 17908 12310
rect 18236 12096 18288 12102
rect 18236 12038 18288 12044
rect 17868 11552 17920 11558
rect 17868 11494 17920 11500
rect 17684 11144 17736 11150
rect 17684 11086 17736 11092
rect 17880 10810 17908 11494
rect 18248 11150 18276 12038
rect 19062 11520 19118 11529
rect 19062 11455 19118 11464
rect 18878 11384 18934 11393
rect 18878 11319 18934 11328
rect 18788 11212 18840 11218
rect 18788 11154 18840 11160
rect 18236 11144 18288 11150
rect 18236 11086 18288 11092
rect 17868 10804 17920 10810
rect 17868 10746 17920 10752
rect 18248 10674 18276 11086
rect 18236 10668 18288 10674
rect 18236 10610 18288 10616
rect 17408 10464 17460 10470
rect 17408 10406 17460 10412
rect 17420 9722 17448 10406
rect 18248 10266 18276 10610
rect 18328 10600 18380 10606
rect 18328 10542 18380 10548
rect 18236 10260 18288 10266
rect 18236 10202 18288 10208
rect 17684 10124 17736 10130
rect 17684 10066 17736 10072
rect 17408 9716 17460 9722
rect 17408 9658 17460 9664
rect 17590 9616 17646 9625
rect 17590 9551 17646 9560
rect 17316 9376 17368 9382
rect 17316 9318 17368 9324
rect 17040 8356 17092 8362
rect 17040 8298 17092 8304
rect 17224 8356 17276 8362
rect 17224 8298 17276 8304
rect 17052 8022 17080 8298
rect 17040 8016 17092 8022
rect 17040 7958 17092 7964
rect 17132 7404 17184 7410
rect 17132 7346 17184 7352
rect 16946 7168 17002 7177
rect 16946 7103 17002 7112
rect 16672 6928 16724 6934
rect 16672 6870 16724 6876
rect 16856 6860 16908 6866
rect 16856 6802 16908 6808
rect 16764 6792 16816 6798
rect 16764 6734 16816 6740
rect 16776 6390 16804 6734
rect 16764 6384 16816 6390
rect 16764 6326 16816 6332
rect 16868 6118 16896 6802
rect 16856 6112 16908 6118
rect 16856 6054 16908 6060
rect 16578 5944 16634 5953
rect 16578 5879 16634 5888
rect 16592 5681 16620 5879
rect 16578 5672 16634 5681
rect 16578 5607 16634 5616
rect 16868 5574 16896 6054
rect 16856 5568 16908 5574
rect 16854 5536 16856 5545
rect 16908 5536 16910 5545
rect 16854 5471 16910 5480
rect 16210 5264 16266 5273
rect 16120 5228 16172 5234
rect 16210 5199 16266 5208
rect 16578 5264 16634 5273
rect 16578 5199 16580 5208
rect 16120 5170 16172 5176
rect 16632 5199 16634 5208
rect 16580 5170 16632 5176
rect 14740 5024 14792 5030
rect 14740 4966 14792 4972
rect 15658 4992 15714 5001
rect 14648 4820 14700 4826
rect 14568 4780 14648 4808
rect 14004 4752 14056 4758
rect 14004 4694 14056 4700
rect 13912 4276 13964 4282
rect 13912 4218 13964 4224
rect 13820 4208 13872 4214
rect 13820 4150 13872 4156
rect 14016 3738 14044 4694
rect 14096 4616 14148 4622
rect 14096 4558 14148 4564
rect 14108 3738 14136 4558
rect 14188 4140 14240 4146
rect 14188 4082 14240 4088
rect 13728 3732 13780 3738
rect 13728 3674 13780 3680
rect 14004 3732 14056 3738
rect 14004 3674 14056 3680
rect 14096 3732 14148 3738
rect 14096 3674 14148 3680
rect 13740 3194 13768 3674
rect 14200 3194 14228 4082
rect 14568 4010 14596 4780
rect 14648 4762 14700 4768
rect 14752 4729 14780 4966
rect 15658 4927 15714 4936
rect 15568 4752 15620 4758
rect 14738 4720 14794 4729
rect 15568 4694 15620 4700
rect 14738 4655 14794 4664
rect 15108 4480 15160 4486
rect 15108 4422 15160 4428
rect 15120 4146 15148 4422
rect 15108 4140 15160 4146
rect 15108 4082 15160 4088
rect 14646 4040 14702 4049
rect 14556 4004 14608 4010
rect 14646 3975 14648 3984
rect 14556 3946 14608 3952
rect 14700 3975 14702 3984
rect 14648 3946 14700 3952
rect 14289 3836 14585 3856
rect 14345 3834 14369 3836
rect 14425 3834 14449 3836
rect 14505 3834 14529 3836
rect 14367 3782 14369 3834
rect 14431 3782 14443 3834
rect 14505 3782 14507 3834
rect 14345 3780 14369 3782
rect 14425 3780 14449 3782
rect 14505 3780 14529 3782
rect 14289 3760 14585 3780
rect 14660 3738 14688 3946
rect 15580 3738 15608 4694
rect 15672 4690 15700 4927
rect 15660 4684 15712 4690
rect 15660 4626 15712 4632
rect 15752 4684 15804 4690
rect 15752 4626 15804 4632
rect 15672 3942 15700 4626
rect 15764 4321 15792 4626
rect 15750 4312 15806 4321
rect 16132 4282 16160 5170
rect 16488 5024 16540 5030
rect 16488 4966 16540 4972
rect 16500 4554 16528 4966
rect 16592 4826 16620 5170
rect 16580 4820 16632 4826
rect 16580 4762 16632 4768
rect 16488 4548 16540 4554
rect 16488 4490 16540 4496
rect 15750 4247 15806 4256
rect 16120 4276 16172 4282
rect 15764 4214 15792 4247
rect 16120 4218 16172 4224
rect 15752 4208 15804 4214
rect 15752 4150 15804 4156
rect 15660 3936 15712 3942
rect 15660 3878 15712 3884
rect 14648 3732 14700 3738
rect 14648 3674 14700 3680
rect 15568 3732 15620 3738
rect 15568 3674 15620 3680
rect 13728 3188 13780 3194
rect 13728 3130 13780 3136
rect 14188 3188 14240 3194
rect 14188 3130 14240 3136
rect 13636 2984 13688 2990
rect 16960 2961 16988 7103
rect 17144 7002 17172 7346
rect 17132 6996 17184 7002
rect 17132 6938 17184 6944
rect 17144 5370 17172 6938
rect 17328 6497 17356 9318
rect 17604 8401 17632 9551
rect 17696 9382 17724 10066
rect 18050 9480 18106 9489
rect 18050 9415 18106 9424
rect 17684 9376 17736 9382
rect 17684 9318 17736 9324
rect 17590 8392 17646 8401
rect 17590 8327 17646 8336
rect 17604 8090 17632 8327
rect 17592 8084 17644 8090
rect 17592 8026 17644 8032
rect 17696 7886 17724 9318
rect 18064 9178 18092 9415
rect 18052 9172 18104 9178
rect 17972 9132 18052 9160
rect 17868 8832 17920 8838
rect 17868 8774 17920 8780
rect 17776 8016 17828 8022
rect 17776 7958 17828 7964
rect 17684 7880 17736 7886
rect 17684 7822 17736 7828
rect 17592 7744 17644 7750
rect 17592 7686 17644 7692
rect 17604 7410 17632 7686
rect 17592 7404 17644 7410
rect 17592 7346 17644 7352
rect 17696 7342 17724 7822
rect 17684 7336 17736 7342
rect 17684 7278 17736 7284
rect 17314 6488 17370 6497
rect 17314 6423 17370 6432
rect 17328 5681 17356 6423
rect 17696 6390 17724 7278
rect 17788 6458 17816 7958
rect 17880 7018 17908 8774
rect 17972 8634 18000 9132
rect 18052 9114 18104 9120
rect 18052 8968 18104 8974
rect 18052 8910 18104 8916
rect 17960 8628 18012 8634
rect 17960 8570 18012 8576
rect 18064 8022 18092 8910
rect 18236 8900 18288 8906
rect 18236 8842 18288 8848
rect 18144 8560 18196 8566
rect 18144 8502 18196 8508
rect 18052 8016 18104 8022
rect 18052 7958 18104 7964
rect 17880 6990 18000 7018
rect 17868 6928 17920 6934
rect 17868 6870 17920 6876
rect 17776 6452 17828 6458
rect 17776 6394 17828 6400
rect 17684 6384 17736 6390
rect 17684 6326 17736 6332
rect 17314 5672 17370 5681
rect 17880 5642 17908 6870
rect 17972 5914 18000 6990
rect 17960 5908 18012 5914
rect 17960 5850 18012 5856
rect 18156 5846 18184 8502
rect 18248 8401 18276 8842
rect 18234 8392 18290 8401
rect 18234 8327 18290 8336
rect 18340 7721 18368 10542
rect 18800 10266 18828 11154
rect 18892 11150 18920 11319
rect 19076 11286 19104 11455
rect 19064 11280 19116 11286
rect 19064 11222 19116 11228
rect 18880 11144 18932 11150
rect 18880 11086 18932 11092
rect 18892 10266 18920 11086
rect 19076 10810 19104 11222
rect 19064 10804 19116 10810
rect 19064 10746 19116 10752
rect 19062 10704 19118 10713
rect 19062 10639 19118 10648
rect 18788 10260 18840 10266
rect 18788 10202 18840 10208
rect 18880 10260 18932 10266
rect 18880 10202 18932 10208
rect 19076 9518 19104 10639
rect 19064 9512 19116 9518
rect 19064 9454 19116 9460
rect 19352 8906 19380 12718
rect 19996 11801 20024 12854
rect 22296 12850 22324 15520
rect 23388 13388 23440 13394
rect 23388 13330 23440 13336
rect 22928 12912 22980 12918
rect 22928 12854 22980 12860
rect 22284 12844 22336 12850
rect 22284 12786 22336 12792
rect 22652 12640 22704 12646
rect 22652 12582 22704 12588
rect 21364 12368 21416 12374
rect 21364 12310 21416 12316
rect 20628 12096 20680 12102
rect 20628 12038 20680 12044
rect 19982 11792 20038 11801
rect 19982 11727 20038 11736
rect 19524 11620 19576 11626
rect 19524 11562 19576 11568
rect 19616 11620 19668 11626
rect 19616 11562 19668 11568
rect 19536 10810 19564 11562
rect 19628 11082 19656 11562
rect 19616 11076 19668 11082
rect 19616 11018 19668 11024
rect 19524 10804 19576 10810
rect 19524 10746 19576 10752
rect 19628 10674 19656 11018
rect 19616 10668 19668 10674
rect 19616 10610 19668 10616
rect 19996 10606 20024 11727
rect 19984 10600 20036 10606
rect 19984 10542 20036 10548
rect 20168 10464 20220 10470
rect 20168 10406 20220 10412
rect 20180 9926 20208 10406
rect 20168 9920 20220 9926
rect 20168 9862 20220 9868
rect 20536 9920 20588 9926
rect 20536 9862 20588 9868
rect 19984 9376 20036 9382
rect 19890 9344 19946 9353
rect 19984 9318 20036 9324
rect 20168 9376 20220 9382
rect 20168 9318 20220 9324
rect 19890 9279 19946 9288
rect 19524 9172 19576 9178
rect 19524 9114 19576 9120
rect 19340 8900 19392 8906
rect 19340 8842 19392 8848
rect 18604 8832 18656 8838
rect 18604 8774 18656 8780
rect 18418 8664 18474 8673
rect 18418 8599 18474 8608
rect 18432 8430 18460 8599
rect 18420 8424 18472 8430
rect 18420 8366 18472 8372
rect 18616 8362 18644 8774
rect 19064 8492 19116 8498
rect 19064 8434 19116 8440
rect 18604 8356 18656 8362
rect 18604 8298 18656 8304
rect 18616 8265 18644 8298
rect 18602 8256 18658 8265
rect 18602 8191 18658 8200
rect 18326 7712 18382 7721
rect 18326 7647 18382 7656
rect 18144 5840 18196 5846
rect 18144 5782 18196 5788
rect 17314 5607 17370 5616
rect 17868 5636 17920 5642
rect 17868 5578 17920 5584
rect 18340 5370 18368 7647
rect 18616 7585 18644 8191
rect 18602 7576 18658 7585
rect 18602 7511 18658 7520
rect 18880 7336 18932 7342
rect 18880 7278 18932 7284
rect 18512 7268 18564 7274
rect 18512 7210 18564 7216
rect 18524 6662 18552 7210
rect 18696 6860 18748 6866
rect 18696 6802 18748 6808
rect 18512 6656 18564 6662
rect 18512 6598 18564 6604
rect 18524 6118 18552 6598
rect 18708 6458 18736 6802
rect 18892 6662 18920 7278
rect 19076 7041 19104 8434
rect 19536 8129 19564 9114
rect 19904 9110 19932 9279
rect 19892 9104 19944 9110
rect 19892 9046 19944 9052
rect 19800 8968 19852 8974
rect 19800 8910 19852 8916
rect 19812 8634 19840 8910
rect 19800 8628 19852 8634
rect 19800 8570 19852 8576
rect 19616 8356 19668 8362
rect 19616 8298 19668 8304
rect 19522 8120 19578 8129
rect 19522 8055 19524 8064
rect 19576 8055 19578 8064
rect 19524 8026 19576 8032
rect 19248 7744 19300 7750
rect 19246 7712 19248 7721
rect 19300 7712 19302 7721
rect 19246 7647 19302 7656
rect 19432 7200 19484 7206
rect 19338 7168 19394 7177
rect 19432 7142 19484 7148
rect 19338 7103 19394 7112
rect 19062 7032 19118 7041
rect 19062 6967 19118 6976
rect 18880 6656 18932 6662
rect 18880 6598 18932 6604
rect 18696 6452 18748 6458
rect 18696 6394 18748 6400
rect 18512 6112 18564 6118
rect 18512 6054 18564 6060
rect 17132 5364 17184 5370
rect 17132 5306 17184 5312
rect 18328 5364 18380 5370
rect 18328 5306 18380 5312
rect 18050 5128 18106 5137
rect 18050 5063 18052 5072
rect 18104 5063 18106 5072
rect 18052 5034 18104 5040
rect 17500 5024 17552 5030
rect 17500 4966 17552 4972
rect 17132 4752 17184 4758
rect 17130 4720 17132 4729
rect 17184 4720 17186 4729
rect 17130 4655 17186 4664
rect 17224 4684 17276 4690
rect 17144 4078 17172 4655
rect 17224 4626 17276 4632
rect 17236 4593 17264 4626
rect 17512 4622 17540 4966
rect 18064 4826 18092 5034
rect 18340 5030 18368 5306
rect 18524 5098 18552 6054
rect 18786 5944 18842 5953
rect 18786 5879 18842 5888
rect 18512 5092 18564 5098
rect 18512 5034 18564 5040
rect 18328 5024 18380 5030
rect 18328 4966 18380 4972
rect 18052 4820 18104 4826
rect 18052 4762 18104 4768
rect 18800 4758 18828 5879
rect 18892 5574 18920 6598
rect 19352 6458 19380 7103
rect 19340 6452 19392 6458
rect 19340 6394 19392 6400
rect 18972 6248 19024 6254
rect 18970 6216 18972 6225
rect 19024 6216 19026 6225
rect 18970 6151 19026 6160
rect 19064 5908 19116 5914
rect 19064 5850 19116 5856
rect 18970 5672 19026 5681
rect 18970 5607 19026 5616
rect 18880 5568 18932 5574
rect 18880 5510 18932 5516
rect 18984 4826 19012 5607
rect 19076 5370 19104 5850
rect 19340 5772 19392 5778
rect 19340 5714 19392 5720
rect 19352 5370 19380 5714
rect 19064 5364 19116 5370
rect 19064 5306 19116 5312
rect 19340 5364 19392 5370
rect 19340 5306 19392 5312
rect 19444 5273 19472 7142
rect 19628 6458 19656 8298
rect 19812 7546 19840 8570
rect 19904 8566 19932 9046
rect 19996 8838 20024 9318
rect 19984 8832 20036 8838
rect 19984 8774 20036 8780
rect 19892 8560 19944 8566
rect 19892 8502 19944 8508
rect 19996 8430 20024 8774
rect 20180 8430 20208 9318
rect 20548 9217 20576 9862
rect 20534 9208 20590 9217
rect 20534 9143 20590 9152
rect 20260 8832 20312 8838
rect 20260 8774 20312 8780
rect 19984 8424 20036 8430
rect 19984 8366 20036 8372
rect 20168 8424 20220 8430
rect 20168 8366 20220 8372
rect 20180 7954 20208 8366
rect 20272 8362 20300 8774
rect 20260 8356 20312 8362
rect 20260 8298 20312 8304
rect 20168 7948 20220 7954
rect 20168 7890 20220 7896
rect 20166 7712 20222 7721
rect 20166 7647 20222 7656
rect 19800 7540 19852 7546
rect 19800 7482 19852 7488
rect 19798 7168 19854 7177
rect 19798 7103 19854 7112
rect 19812 7002 19840 7103
rect 19800 6996 19852 7002
rect 19800 6938 19852 6944
rect 19616 6452 19668 6458
rect 19616 6394 19668 6400
rect 19812 6254 19840 6938
rect 20180 6322 20208 7647
rect 20548 6662 20576 9143
rect 20640 8498 20668 12038
rect 20956 11996 21252 12016
rect 21012 11994 21036 11996
rect 21092 11994 21116 11996
rect 21172 11994 21196 11996
rect 21034 11942 21036 11994
rect 21098 11942 21110 11994
rect 21172 11942 21174 11994
rect 21012 11940 21036 11942
rect 21092 11940 21116 11942
rect 21172 11940 21196 11942
rect 20956 11920 21252 11940
rect 20904 11688 20956 11694
rect 20904 11630 20956 11636
rect 20812 11552 20864 11558
rect 20810 11520 20812 11529
rect 20864 11520 20866 11529
rect 20810 11455 20866 11464
rect 20824 11286 20852 11455
rect 20812 11280 20864 11286
rect 20812 11222 20864 11228
rect 20720 11212 20772 11218
rect 20720 11154 20772 11160
rect 20732 10742 20760 11154
rect 20824 10810 20852 11222
rect 20916 11218 20944 11630
rect 21376 11558 21404 12310
rect 21824 12232 21876 12238
rect 21824 12174 21876 12180
rect 21732 12164 21784 12170
rect 21732 12106 21784 12112
rect 21744 11558 21772 12106
rect 21836 11558 21864 12174
rect 21364 11552 21416 11558
rect 21364 11494 21416 11500
rect 21732 11552 21784 11558
rect 21732 11494 21784 11500
rect 21824 11552 21876 11558
rect 21824 11494 21876 11500
rect 20904 11212 20956 11218
rect 20904 11154 20956 11160
rect 20956 10908 21252 10928
rect 21012 10906 21036 10908
rect 21092 10906 21116 10908
rect 21172 10906 21196 10908
rect 21034 10854 21036 10906
rect 21098 10854 21110 10906
rect 21172 10854 21174 10906
rect 21012 10852 21036 10854
rect 21092 10852 21116 10854
rect 21172 10852 21196 10854
rect 20956 10832 21252 10852
rect 20812 10804 20864 10810
rect 20812 10746 20864 10752
rect 20720 10736 20772 10742
rect 20720 10678 20772 10684
rect 20732 10062 20760 10678
rect 20720 10056 20772 10062
rect 20720 9998 20772 10004
rect 20732 9722 20760 9998
rect 20810 9888 20866 9897
rect 20810 9823 20866 9832
rect 20720 9716 20772 9722
rect 20720 9658 20772 9664
rect 20824 9081 20852 9823
rect 20956 9820 21252 9840
rect 21012 9818 21036 9820
rect 21092 9818 21116 9820
rect 21172 9818 21196 9820
rect 21034 9766 21036 9818
rect 21098 9766 21110 9818
rect 21172 9766 21174 9818
rect 21012 9764 21036 9766
rect 21092 9764 21116 9766
rect 21172 9764 21196 9766
rect 20956 9744 21252 9764
rect 21376 9081 21404 11494
rect 21640 11280 21692 11286
rect 21638 11248 21640 11257
rect 21692 11248 21694 11257
rect 21638 11183 21694 11192
rect 21640 9512 21692 9518
rect 21640 9454 21692 9460
rect 20810 9072 20866 9081
rect 20810 9007 20866 9016
rect 21362 9072 21418 9081
rect 21362 9007 21418 9016
rect 21652 8974 21680 9454
rect 21640 8968 21692 8974
rect 21640 8910 21692 8916
rect 20956 8732 21252 8752
rect 21012 8730 21036 8732
rect 21092 8730 21116 8732
rect 21172 8730 21196 8732
rect 21034 8678 21036 8730
rect 21098 8678 21110 8730
rect 21172 8678 21174 8730
rect 21012 8676 21036 8678
rect 21092 8676 21116 8678
rect 21172 8676 21196 8678
rect 20956 8656 21252 8676
rect 20628 8492 20680 8498
rect 20628 8434 20680 8440
rect 20640 8090 20668 8434
rect 20904 8424 20956 8430
rect 20824 8384 20904 8412
rect 20628 8084 20680 8090
rect 20628 8026 20680 8032
rect 20824 7721 20852 8384
rect 20904 8366 20956 8372
rect 21652 8294 21680 8910
rect 21640 8288 21692 8294
rect 21640 8230 21692 8236
rect 21364 8016 21416 8022
rect 21364 7958 21416 7964
rect 21376 7750 21404 7958
rect 21548 7948 21600 7954
rect 21548 7890 21600 7896
rect 21364 7744 21416 7750
rect 20810 7712 20866 7721
rect 21364 7686 21416 7692
rect 20810 7647 20866 7656
rect 20956 7644 21252 7664
rect 21012 7642 21036 7644
rect 21092 7642 21116 7644
rect 21172 7642 21196 7644
rect 21034 7590 21036 7642
rect 21098 7590 21110 7642
rect 21172 7590 21174 7642
rect 21012 7588 21036 7590
rect 21092 7588 21116 7590
rect 21172 7588 21196 7590
rect 20810 7576 20866 7585
rect 20956 7568 21252 7588
rect 20810 7511 20866 7520
rect 20824 7410 20852 7511
rect 20812 7404 20864 7410
rect 20812 7346 20864 7352
rect 20904 7200 20956 7206
rect 20904 7142 20956 7148
rect 20916 6934 20944 7142
rect 20904 6928 20956 6934
rect 20904 6870 20956 6876
rect 21272 6928 21324 6934
rect 21272 6870 21324 6876
rect 20260 6656 20312 6662
rect 20260 6598 20312 6604
rect 20536 6656 20588 6662
rect 20536 6598 20588 6604
rect 20168 6316 20220 6322
rect 20168 6258 20220 6264
rect 19800 6248 19852 6254
rect 19800 6190 19852 6196
rect 19524 6112 19576 6118
rect 19524 6054 19576 6060
rect 19536 5953 19564 6054
rect 19522 5944 19578 5953
rect 19522 5879 19524 5888
rect 19576 5879 19578 5888
rect 19524 5850 19576 5856
rect 20180 5846 20208 6258
rect 20168 5840 20220 5846
rect 20168 5782 20220 5788
rect 19984 5568 20036 5574
rect 19984 5510 20036 5516
rect 19430 5264 19486 5273
rect 19430 5199 19486 5208
rect 19156 5092 19208 5098
rect 19156 5034 19208 5040
rect 18972 4820 19024 4826
rect 18972 4762 19024 4768
rect 18788 4752 18840 4758
rect 18788 4694 18840 4700
rect 17500 4616 17552 4622
rect 17222 4584 17278 4593
rect 17278 4542 17356 4570
rect 17500 4558 17552 4564
rect 17222 4519 17278 4528
rect 17328 4282 17356 4542
rect 17512 4282 17540 4558
rect 17316 4276 17368 4282
rect 17500 4276 17552 4282
rect 17368 4236 17448 4264
rect 17316 4218 17368 4224
rect 17132 4072 17184 4078
rect 17132 4014 17184 4020
rect 13636 2926 13688 2932
rect 16946 2952 17002 2961
rect 16946 2887 17002 2896
rect 14289 2748 14585 2768
rect 14345 2746 14369 2748
rect 14425 2746 14449 2748
rect 14505 2746 14529 2748
rect 14367 2694 14369 2746
rect 14431 2694 14443 2746
rect 14505 2694 14507 2746
rect 14345 2692 14369 2694
rect 14425 2692 14449 2694
rect 14505 2692 14529 2694
rect 14289 2672 14585 2692
rect 12900 2644 12952 2650
rect 12900 2586 12952 2592
rect 13360 2644 13412 2650
rect 13360 2586 13412 2592
rect 12808 2576 12860 2582
rect 12808 2518 12860 2524
rect 12530 1864 12586 1873
rect 12530 1799 12586 1808
rect 17420 1737 17448 4236
rect 17500 4218 17552 4224
rect 18800 4146 18828 4694
rect 18984 4214 19012 4762
rect 19168 4622 19196 5034
rect 19156 4616 19208 4622
rect 19156 4558 19208 4564
rect 19168 4282 19196 4558
rect 19156 4276 19208 4282
rect 19156 4218 19208 4224
rect 18972 4208 19024 4214
rect 18972 4150 19024 4156
rect 18788 4140 18840 4146
rect 18788 4082 18840 4088
rect 5906 1728 5962 1737
rect 5906 1663 5962 1672
rect 17406 1728 17462 1737
rect 17406 1663 17462 1672
rect 19996 480 20024 5510
rect 20272 5370 20300 6598
rect 20548 6118 20576 6598
rect 20956 6556 21252 6576
rect 21012 6554 21036 6556
rect 21092 6554 21116 6556
rect 21172 6554 21196 6556
rect 21034 6502 21036 6554
rect 21098 6502 21110 6554
rect 21172 6502 21174 6554
rect 21012 6500 21036 6502
rect 21092 6500 21116 6502
rect 21172 6500 21196 6502
rect 20956 6480 21252 6500
rect 21284 6458 21312 6870
rect 21376 6730 21404 7686
rect 21560 7546 21588 7890
rect 21652 7886 21680 8230
rect 21744 8090 21772 11494
rect 21836 11234 21864 11494
rect 21836 11206 21956 11234
rect 21822 11112 21878 11121
rect 21822 11047 21878 11056
rect 21836 10266 21864 11047
rect 21824 10260 21876 10266
rect 21824 10202 21876 10208
rect 21822 9480 21878 9489
rect 21822 9415 21878 9424
rect 21836 8401 21864 9415
rect 21928 9110 21956 11206
rect 22284 11076 22336 11082
rect 22284 11018 22336 11024
rect 22296 10713 22324 11018
rect 22282 10704 22338 10713
rect 22282 10639 22338 10648
rect 22008 10464 22060 10470
rect 22008 10406 22060 10412
rect 22020 10305 22048 10406
rect 22006 10296 22062 10305
rect 22006 10231 22062 10240
rect 22376 10192 22428 10198
rect 22376 10134 22428 10140
rect 22388 9586 22416 10134
rect 22376 9580 22428 9586
rect 22376 9522 22428 9528
rect 22388 9382 22416 9522
rect 22376 9376 22428 9382
rect 22374 9344 22376 9353
rect 22428 9344 22430 9353
rect 22374 9279 22430 9288
rect 21916 9104 21968 9110
rect 21916 9046 21968 9052
rect 21928 8430 21956 9046
rect 22008 8560 22060 8566
rect 22008 8502 22060 8508
rect 21916 8424 21968 8430
rect 21822 8392 21878 8401
rect 21916 8366 21968 8372
rect 21822 8327 21878 8336
rect 21916 8288 21968 8294
rect 21822 8256 21878 8265
rect 21916 8230 21968 8236
rect 21822 8191 21878 8200
rect 21732 8084 21784 8090
rect 21732 8026 21784 8032
rect 21640 7880 21692 7886
rect 21836 7857 21864 8191
rect 21928 8090 21956 8230
rect 21916 8084 21968 8090
rect 21916 8026 21968 8032
rect 21916 7880 21968 7886
rect 21640 7822 21692 7828
rect 21822 7848 21878 7857
rect 21916 7822 21968 7828
rect 21822 7783 21878 7792
rect 21548 7540 21600 7546
rect 21548 7482 21600 7488
rect 21548 6928 21600 6934
rect 21548 6870 21600 6876
rect 21364 6724 21416 6730
rect 21364 6666 21416 6672
rect 21560 6662 21588 6870
rect 21640 6792 21692 6798
rect 21640 6734 21692 6740
rect 21548 6656 21600 6662
rect 21548 6598 21600 6604
rect 20812 6452 20864 6458
rect 20812 6394 20864 6400
rect 21272 6452 21324 6458
rect 21272 6394 21324 6400
rect 20536 6112 20588 6118
rect 20536 6054 20588 6060
rect 20260 5364 20312 5370
rect 20260 5306 20312 5312
rect 20272 5098 20300 5306
rect 20548 5137 20576 6054
rect 20824 5409 20852 6394
rect 21652 6254 21680 6734
rect 21928 6662 21956 7822
rect 21916 6656 21968 6662
rect 21916 6598 21968 6604
rect 21088 6248 21140 6254
rect 21088 6190 21140 6196
rect 21640 6248 21692 6254
rect 21640 6190 21692 6196
rect 21100 5710 21128 6190
rect 21652 5914 21680 6190
rect 21730 5944 21786 5953
rect 21640 5908 21692 5914
rect 21730 5879 21786 5888
rect 21640 5850 21692 5856
rect 21088 5704 21140 5710
rect 21088 5646 21140 5652
rect 21456 5704 21508 5710
rect 21456 5646 21508 5652
rect 20956 5468 21252 5488
rect 21012 5466 21036 5468
rect 21092 5466 21116 5468
rect 21172 5466 21196 5468
rect 21034 5414 21036 5466
rect 21098 5414 21110 5466
rect 21172 5414 21174 5466
rect 21012 5412 21036 5414
rect 21092 5412 21116 5414
rect 21172 5412 21196 5414
rect 20810 5400 20866 5409
rect 20956 5392 21252 5412
rect 21468 5370 21496 5646
rect 20810 5335 20866 5344
rect 21456 5364 21508 5370
rect 21456 5306 21508 5312
rect 20534 5128 20590 5137
rect 20260 5092 20312 5098
rect 21744 5098 21772 5879
rect 21824 5840 21876 5846
rect 21824 5782 21876 5788
rect 21836 5234 21864 5782
rect 21824 5228 21876 5234
rect 21824 5170 21876 5176
rect 20534 5063 20590 5072
rect 21732 5092 21784 5098
rect 20260 5034 20312 5040
rect 21732 5034 21784 5040
rect 21836 4826 21864 5170
rect 22020 4842 22048 8502
rect 22100 8424 22152 8430
rect 22100 8366 22152 8372
rect 22112 8022 22140 8366
rect 22468 8356 22520 8362
rect 22468 8298 22520 8304
rect 22376 8288 22428 8294
rect 22376 8230 22428 8236
rect 22100 8016 22152 8022
rect 22100 7958 22152 7964
rect 22388 7546 22416 8230
rect 22376 7540 22428 7546
rect 22376 7482 22428 7488
rect 22100 6656 22152 6662
rect 22100 6598 22152 6604
rect 22112 5370 22140 6598
rect 22480 6458 22508 8298
rect 22560 7200 22612 7206
rect 22560 7142 22612 7148
rect 22572 6730 22600 7142
rect 22560 6724 22612 6730
rect 22560 6666 22612 6672
rect 22468 6452 22520 6458
rect 22468 6394 22520 6400
rect 22480 5846 22508 6394
rect 22468 5840 22520 5846
rect 22468 5782 22520 5788
rect 22100 5364 22152 5370
rect 22100 5306 22152 5312
rect 22376 5296 22428 5302
rect 22376 5238 22428 5244
rect 22020 4826 22140 4842
rect 21824 4820 21876 4826
rect 22020 4820 22152 4826
rect 22020 4814 22100 4820
rect 21824 4762 21876 4768
rect 22100 4762 22152 4768
rect 20956 4380 21252 4400
rect 21012 4378 21036 4380
rect 21092 4378 21116 4380
rect 21172 4378 21196 4380
rect 21034 4326 21036 4378
rect 21098 4326 21110 4378
rect 21172 4326 21174 4378
rect 21012 4324 21036 4326
rect 21092 4324 21116 4326
rect 21172 4324 21196 4326
rect 20956 4304 21252 4324
rect 22112 4282 22140 4762
rect 22388 4758 22416 5238
rect 22376 4752 22428 4758
rect 22376 4694 22428 4700
rect 22284 4616 22336 4622
rect 22284 4558 22336 4564
rect 22100 4276 22152 4282
rect 22100 4218 22152 4224
rect 22296 4146 22324 4558
rect 22388 4146 22416 4694
rect 22664 4486 22692 12582
rect 22940 11354 22968 12854
rect 23400 12646 23428 13330
rect 23480 12776 23532 12782
rect 23480 12718 23532 12724
rect 23388 12640 23440 12646
rect 23388 12582 23440 12588
rect 23296 11552 23348 11558
rect 23296 11494 23348 11500
rect 23308 11354 23336 11494
rect 22928 11348 22980 11354
rect 22928 11290 22980 11296
rect 23296 11348 23348 11354
rect 23296 11290 23348 11296
rect 22940 10470 22968 11290
rect 23492 11082 23520 12718
rect 24400 12164 24452 12170
rect 24400 12106 24452 12112
rect 23756 11824 23808 11830
rect 23756 11766 23808 11772
rect 23572 11552 23624 11558
rect 23572 11494 23624 11500
rect 23480 11076 23532 11082
rect 23480 11018 23532 11024
rect 23018 10976 23074 10985
rect 23018 10911 23074 10920
rect 23032 10674 23060 10911
rect 23584 10742 23612 11494
rect 23768 11218 23796 11766
rect 24412 11762 24440 12106
rect 24400 11756 24452 11762
rect 24400 11698 24452 11704
rect 24400 11552 24452 11558
rect 24400 11494 24452 11500
rect 23848 11348 23900 11354
rect 23848 11290 23900 11296
rect 23756 11212 23808 11218
rect 23756 11154 23808 11160
rect 23768 11121 23796 11154
rect 23754 11112 23810 11121
rect 23754 11047 23810 11056
rect 23860 10810 23888 11290
rect 24412 11286 24440 11494
rect 24596 11286 24624 15520
rect 26988 13394 27016 15520
rect 27622 13628 27918 13648
rect 27678 13626 27702 13628
rect 27758 13626 27782 13628
rect 27838 13626 27862 13628
rect 27700 13574 27702 13626
rect 27764 13574 27776 13626
rect 27838 13574 27840 13626
rect 27678 13572 27702 13574
rect 27758 13572 27782 13574
rect 27838 13572 27862 13574
rect 27622 13552 27918 13572
rect 26976 13388 27028 13394
rect 26976 13330 27028 13336
rect 24860 13184 24912 13190
rect 24860 13126 24912 13132
rect 24872 12850 24900 13126
rect 25504 12980 25556 12986
rect 25504 12922 25556 12928
rect 25228 12912 25280 12918
rect 25228 12854 25280 12860
rect 24860 12844 24912 12850
rect 24860 12786 24912 12792
rect 24768 12708 24820 12714
rect 24768 12650 24820 12656
rect 24780 12617 24808 12650
rect 25136 12640 25188 12646
rect 24766 12608 24822 12617
rect 25136 12582 25188 12588
rect 24766 12543 24822 12552
rect 25044 12368 25096 12374
rect 25044 12310 25096 12316
rect 24952 12232 25004 12238
rect 24952 12174 25004 12180
rect 24676 12096 24728 12102
rect 24676 12038 24728 12044
rect 24688 11762 24716 12038
rect 24676 11756 24728 11762
rect 24676 11698 24728 11704
rect 24688 11370 24716 11698
rect 24688 11342 24808 11370
rect 24400 11280 24452 11286
rect 24400 11222 24452 11228
rect 24584 11280 24636 11286
rect 24584 11222 24636 11228
rect 24674 11248 24730 11257
rect 24674 11183 24730 11192
rect 24032 11144 24084 11150
rect 24032 11086 24084 11092
rect 24306 11112 24362 11121
rect 23848 10804 23900 10810
rect 23848 10746 23900 10752
rect 23572 10736 23624 10742
rect 24044 10713 24072 11086
rect 24306 11047 24362 11056
rect 24320 11014 24348 11047
rect 24308 11008 24360 11014
rect 24308 10950 24360 10956
rect 23572 10678 23624 10684
rect 24030 10704 24086 10713
rect 23020 10668 23072 10674
rect 24030 10639 24032 10648
rect 23020 10610 23072 10616
rect 24084 10639 24086 10648
rect 24032 10610 24084 10616
rect 24044 10579 24072 10610
rect 24320 10538 24348 10950
rect 24400 10668 24452 10674
rect 24400 10610 24452 10616
rect 24308 10532 24360 10538
rect 24308 10474 24360 10480
rect 22928 10464 22980 10470
rect 22928 10406 22980 10412
rect 24412 10266 24440 10610
rect 24492 10532 24544 10538
rect 24492 10474 24544 10480
rect 24400 10260 24452 10266
rect 24400 10202 24452 10208
rect 24400 10124 24452 10130
rect 24400 10066 24452 10072
rect 23480 9920 23532 9926
rect 23480 9862 23532 9868
rect 23388 9512 23440 9518
rect 23388 9454 23440 9460
rect 23020 9444 23072 9450
rect 23020 9386 23072 9392
rect 23032 9178 23060 9386
rect 23020 9172 23072 9178
rect 23020 9114 23072 9120
rect 23400 8634 23428 9454
rect 23492 9178 23520 9862
rect 24032 9648 24084 9654
rect 24032 9590 24084 9596
rect 23938 9344 23994 9353
rect 23938 9279 23994 9288
rect 23480 9172 23532 9178
rect 23480 9114 23532 9120
rect 23756 8832 23808 8838
rect 23756 8774 23808 8780
rect 23388 8628 23440 8634
rect 23388 8570 23440 8576
rect 23664 8492 23716 8498
rect 23664 8434 23716 8440
rect 23388 7744 23440 7750
rect 23388 7686 23440 7692
rect 22744 7268 22796 7274
rect 22744 7210 22796 7216
rect 22756 6866 22784 7210
rect 23400 7206 23428 7686
rect 23676 7546 23704 8434
rect 23768 8362 23796 8774
rect 23756 8356 23808 8362
rect 23756 8298 23808 8304
rect 23664 7540 23716 7546
rect 23664 7482 23716 7488
rect 23388 7200 23440 7206
rect 23388 7142 23440 7148
rect 23112 6928 23164 6934
rect 23112 6870 23164 6876
rect 22744 6860 22796 6866
rect 22744 6802 22796 6808
rect 23124 6458 23152 6870
rect 23400 6798 23428 7142
rect 23848 6860 23900 6866
rect 23848 6802 23900 6808
rect 23388 6792 23440 6798
rect 23388 6734 23440 6740
rect 23112 6452 23164 6458
rect 23112 6394 23164 6400
rect 23124 5681 23152 6394
rect 23400 5914 23428 6734
rect 23480 6724 23532 6730
rect 23480 6666 23532 6672
rect 23492 6458 23520 6666
rect 23480 6452 23532 6458
rect 23480 6394 23532 6400
rect 23492 6089 23520 6394
rect 23478 6080 23534 6089
rect 23478 6015 23534 6024
rect 23860 5914 23888 6802
rect 23952 6458 23980 9279
rect 24044 9217 24072 9590
rect 24412 9382 24440 10066
rect 24504 9926 24532 10474
rect 24688 9994 24716 11183
rect 24780 10849 24808 11342
rect 24860 11212 24912 11218
rect 24860 11154 24912 11160
rect 24766 10840 24822 10849
rect 24766 10775 24822 10784
rect 24780 10674 24808 10775
rect 24768 10668 24820 10674
rect 24768 10610 24820 10616
rect 24872 10470 24900 11154
rect 24964 11082 24992 12174
rect 25056 12073 25084 12310
rect 25042 12064 25098 12073
rect 25042 11999 25098 12008
rect 25056 11898 25084 11999
rect 25044 11892 25096 11898
rect 25044 11834 25096 11840
rect 25056 11665 25084 11834
rect 25042 11656 25098 11665
rect 25042 11591 25098 11600
rect 25148 11529 25176 12582
rect 25134 11520 25190 11529
rect 25134 11455 25190 11464
rect 24952 11076 25004 11082
rect 25240 11064 25268 12854
rect 25516 12102 25544 12922
rect 29380 12850 29408 15520
rect 31208 13728 31260 13734
rect 31208 13670 31260 13676
rect 31116 12980 31168 12986
rect 31116 12922 31168 12928
rect 26516 12844 26568 12850
rect 26516 12786 26568 12792
rect 29368 12844 29420 12850
rect 29368 12786 29420 12792
rect 25872 12232 25924 12238
rect 25872 12174 25924 12180
rect 25504 12096 25556 12102
rect 25504 12038 25556 12044
rect 25594 11928 25650 11937
rect 25594 11863 25650 11872
rect 25608 11529 25636 11863
rect 25884 11626 25912 12174
rect 25964 12096 26016 12102
rect 25964 12038 26016 12044
rect 25872 11620 25924 11626
rect 25872 11562 25924 11568
rect 25594 11520 25650 11529
rect 25594 11455 25650 11464
rect 24952 11018 25004 11024
rect 25148 11036 25268 11064
rect 25320 11076 25372 11082
rect 25044 11008 25096 11014
rect 25042 10976 25044 10985
rect 25096 10976 25098 10985
rect 25042 10911 25098 10920
rect 25148 10577 25176 11036
rect 25320 11018 25372 11024
rect 25226 10976 25282 10985
rect 25226 10911 25282 10920
rect 25134 10568 25190 10577
rect 25134 10503 25190 10512
rect 24860 10464 24912 10470
rect 24780 10424 24860 10452
rect 24676 9988 24728 9994
rect 24676 9930 24728 9936
rect 24492 9920 24544 9926
rect 24492 9862 24544 9868
rect 24504 9518 24532 9862
rect 24492 9512 24544 9518
rect 24492 9454 24544 9460
rect 24124 9376 24176 9382
rect 24124 9318 24176 9324
rect 24400 9376 24452 9382
rect 24400 9318 24452 9324
rect 24030 9208 24086 9217
rect 24030 9143 24086 9152
rect 24136 7342 24164 9318
rect 24780 8838 24808 10424
rect 24860 10406 24912 10412
rect 24952 9104 25004 9110
rect 24952 9046 25004 9052
rect 24768 8832 24820 8838
rect 24768 8774 24820 8780
rect 24964 8362 24992 9046
rect 25044 8968 25096 8974
rect 25044 8910 25096 8916
rect 25056 8634 25084 8910
rect 25044 8628 25096 8634
rect 25044 8570 25096 8576
rect 24952 8356 25004 8362
rect 24952 8298 25004 8304
rect 24964 7818 24992 8298
rect 25056 8090 25084 8570
rect 25044 8084 25096 8090
rect 25044 8026 25096 8032
rect 24952 7812 25004 7818
rect 24952 7754 25004 7760
rect 24124 7336 24176 7342
rect 24124 7278 24176 7284
rect 24676 6928 24728 6934
rect 24490 6896 24546 6905
rect 24676 6870 24728 6876
rect 24490 6831 24546 6840
rect 24124 6792 24176 6798
rect 24030 6760 24086 6769
rect 24124 6734 24176 6740
rect 24030 6695 24032 6704
rect 24084 6695 24086 6704
rect 24032 6666 24084 6672
rect 23940 6452 23992 6458
rect 23940 6394 23992 6400
rect 24136 6118 24164 6734
rect 24216 6656 24268 6662
rect 24216 6598 24268 6604
rect 24124 6112 24176 6118
rect 24124 6054 24176 6060
rect 23388 5908 23440 5914
rect 23388 5850 23440 5856
rect 23848 5908 23900 5914
rect 23848 5850 23900 5856
rect 23940 5704 23992 5710
rect 23110 5672 23166 5681
rect 23940 5646 23992 5652
rect 23110 5607 23166 5616
rect 22836 5568 22888 5574
rect 22836 5510 22888 5516
rect 22848 5098 22876 5510
rect 23952 5370 23980 5646
rect 24136 5409 24164 6054
rect 24228 5953 24256 6598
rect 24504 6458 24532 6831
rect 24688 6730 24716 6870
rect 24676 6724 24728 6730
rect 24676 6666 24728 6672
rect 24492 6452 24544 6458
rect 24492 6394 24544 6400
rect 24688 6225 24716 6666
rect 24952 6656 25004 6662
rect 24952 6598 25004 6604
rect 24674 6216 24730 6225
rect 24674 6151 24730 6160
rect 24768 6180 24820 6186
rect 24768 6122 24820 6128
rect 24214 5944 24270 5953
rect 24214 5879 24270 5888
rect 24216 5772 24268 5778
rect 24216 5714 24268 5720
rect 24122 5400 24178 5409
rect 23940 5364 23992 5370
rect 24122 5335 24178 5344
rect 23940 5306 23992 5312
rect 22836 5092 22888 5098
rect 22836 5034 22888 5040
rect 22848 4622 22876 5034
rect 22836 4616 22888 4622
rect 22836 4558 22888 4564
rect 22652 4480 22704 4486
rect 24136 4457 24164 5335
rect 24228 5098 24256 5714
rect 24780 5370 24808 6122
rect 24964 6118 24992 6598
rect 25148 6322 25176 10503
rect 25240 10062 25268 10911
rect 25332 10674 25360 11018
rect 25320 10668 25372 10674
rect 25320 10610 25372 10616
rect 25412 10192 25464 10198
rect 25412 10134 25464 10140
rect 25228 10056 25280 10062
rect 25320 10056 25372 10062
rect 25228 9998 25280 10004
rect 25318 10024 25320 10033
rect 25372 10024 25374 10033
rect 25240 9722 25268 9998
rect 25318 9959 25374 9968
rect 25228 9716 25280 9722
rect 25228 9658 25280 9664
rect 25424 9450 25452 10134
rect 25412 9444 25464 9450
rect 25412 9386 25464 9392
rect 25424 9178 25452 9386
rect 25412 9172 25464 9178
rect 25412 9114 25464 9120
rect 25504 8288 25556 8294
rect 25504 8230 25556 8236
rect 25516 7993 25544 8230
rect 25502 7984 25558 7993
rect 25502 7919 25504 7928
rect 25556 7919 25558 7928
rect 25504 7890 25556 7896
rect 25412 7880 25464 7886
rect 25412 7822 25464 7828
rect 25424 7546 25452 7822
rect 25412 7540 25464 7546
rect 25412 7482 25464 7488
rect 25412 7200 25464 7206
rect 25412 7142 25464 7148
rect 25424 6934 25452 7142
rect 25516 7002 25544 7890
rect 25504 6996 25556 7002
rect 25504 6938 25556 6944
rect 25412 6928 25464 6934
rect 25412 6870 25464 6876
rect 25136 6316 25188 6322
rect 25136 6258 25188 6264
rect 24952 6112 25004 6118
rect 24952 6054 25004 6060
rect 24768 5364 24820 5370
rect 24768 5306 24820 5312
rect 24216 5092 24268 5098
rect 24216 5034 24268 5040
rect 24964 4593 24992 6054
rect 25608 5001 25636 11455
rect 25884 11014 25912 11562
rect 25976 11558 26004 12038
rect 26528 11898 26556 12786
rect 27622 12540 27918 12560
rect 27678 12538 27702 12540
rect 27758 12538 27782 12540
rect 27838 12538 27862 12540
rect 27700 12486 27702 12538
rect 27764 12486 27776 12538
rect 27838 12486 27840 12538
rect 27678 12484 27702 12486
rect 27758 12484 27782 12486
rect 27838 12484 27862 12486
rect 27622 12464 27918 12484
rect 31128 12442 31156 12922
rect 31116 12436 31168 12442
rect 31116 12378 31168 12384
rect 29550 12336 29606 12345
rect 29550 12271 29606 12280
rect 27250 12200 27306 12209
rect 27250 12135 27306 12144
rect 26516 11892 26568 11898
rect 26516 11834 26568 11840
rect 25964 11552 26016 11558
rect 25964 11494 26016 11500
rect 25872 11008 25924 11014
rect 25872 10950 25924 10956
rect 25884 10810 25912 10950
rect 25872 10804 25924 10810
rect 25872 10746 25924 10752
rect 25884 9722 25912 10746
rect 25872 9716 25924 9722
rect 25872 9658 25924 9664
rect 25976 8673 26004 11494
rect 26332 11280 26384 11286
rect 26238 11248 26294 11257
rect 26332 11222 26384 11228
rect 26238 11183 26240 11192
rect 26292 11183 26294 11192
rect 26240 11154 26292 11160
rect 26344 10266 26372 11222
rect 26148 10260 26200 10266
rect 26148 10202 26200 10208
rect 26332 10260 26384 10266
rect 26332 10202 26384 10208
rect 26160 10033 26188 10202
rect 26528 10198 26556 11834
rect 27160 11824 27212 11830
rect 27160 11766 27212 11772
rect 27172 11286 27200 11766
rect 27264 11762 27292 12135
rect 27436 12096 27488 12102
rect 27436 12038 27488 12044
rect 27252 11756 27304 11762
rect 27252 11698 27304 11704
rect 27448 11626 27476 12038
rect 29564 11898 29592 12271
rect 30196 12096 30248 12102
rect 30196 12038 30248 12044
rect 31024 12096 31076 12102
rect 31024 12038 31076 12044
rect 29552 11892 29604 11898
rect 29552 11834 29604 11840
rect 29366 11792 29422 11801
rect 29366 11727 29422 11736
rect 29380 11694 29408 11727
rect 30208 11694 30236 12038
rect 30380 11824 30432 11830
rect 30380 11766 30432 11772
rect 29368 11688 29420 11694
rect 29920 11688 29972 11694
rect 29368 11630 29420 11636
rect 29918 11656 29920 11665
rect 30196 11688 30248 11694
rect 29972 11656 29974 11665
rect 27436 11620 27488 11626
rect 30196 11630 30248 11636
rect 29918 11591 29974 11600
rect 27436 11562 27488 11568
rect 27160 11280 27212 11286
rect 27160 11222 27212 11228
rect 26700 11144 26752 11150
rect 26606 11112 26662 11121
rect 26700 11086 26752 11092
rect 26606 11047 26608 11056
rect 26660 11047 26662 11056
rect 26608 11018 26660 11024
rect 26712 10606 26740 11086
rect 27342 10704 27398 10713
rect 27342 10639 27398 10648
rect 26700 10600 26752 10606
rect 26700 10542 26752 10548
rect 26712 10266 26740 10542
rect 27068 10532 27120 10538
rect 27068 10474 27120 10480
rect 26700 10260 26752 10266
rect 26700 10202 26752 10208
rect 26516 10192 26568 10198
rect 26516 10134 26568 10140
rect 27080 10130 27108 10474
rect 27356 10198 27384 10639
rect 27344 10192 27396 10198
rect 27344 10134 27396 10140
rect 27068 10124 27120 10130
rect 27068 10066 27120 10072
rect 26146 10024 26202 10033
rect 26146 9959 26202 9968
rect 27356 9722 27384 10134
rect 27344 9716 27396 9722
rect 27344 9658 27396 9664
rect 26056 9648 26108 9654
rect 26056 9590 26108 9596
rect 26882 9616 26938 9625
rect 26068 9042 26096 9590
rect 26882 9551 26938 9560
rect 26514 9480 26570 9489
rect 26514 9415 26570 9424
rect 26056 9036 26108 9042
rect 26056 8978 26108 8984
rect 25962 8664 26018 8673
rect 26068 8634 26096 8978
rect 26528 8634 26556 9415
rect 25962 8599 26018 8608
rect 26056 8628 26108 8634
rect 26056 8570 26108 8576
rect 26516 8628 26568 8634
rect 26516 8570 26568 8576
rect 26896 8566 26924 9551
rect 27068 9512 27120 9518
rect 27448 9489 27476 11562
rect 28264 11552 28316 11558
rect 28264 11494 28316 11500
rect 27622 11452 27918 11472
rect 27678 11450 27702 11452
rect 27758 11450 27782 11452
rect 27838 11450 27862 11452
rect 27700 11398 27702 11450
rect 27764 11398 27776 11450
rect 27838 11398 27840 11450
rect 27678 11396 27702 11398
rect 27758 11396 27782 11398
rect 27838 11396 27862 11398
rect 27622 11376 27918 11396
rect 28172 11144 28224 11150
rect 28172 11086 28224 11092
rect 27802 10840 27858 10849
rect 27802 10775 27804 10784
rect 27856 10775 27858 10784
rect 27804 10746 27856 10752
rect 28184 10538 28212 11086
rect 28172 10532 28224 10538
rect 28172 10474 28224 10480
rect 27622 10364 27918 10384
rect 27678 10362 27702 10364
rect 27758 10362 27782 10364
rect 27838 10362 27862 10364
rect 27700 10310 27702 10362
rect 27764 10310 27776 10362
rect 27838 10310 27840 10362
rect 27678 10308 27702 10310
rect 27758 10308 27782 10310
rect 27838 10308 27862 10310
rect 27622 10288 27918 10308
rect 27068 9454 27120 9460
rect 27434 9480 27490 9489
rect 26976 9104 27028 9110
rect 26974 9072 26976 9081
rect 27028 9072 27030 9081
rect 27080 9042 27108 9454
rect 27434 9415 27490 9424
rect 28172 9444 28224 9450
rect 28172 9386 28224 9392
rect 27622 9276 27918 9296
rect 27678 9274 27702 9276
rect 27758 9274 27782 9276
rect 27838 9274 27862 9276
rect 27700 9222 27702 9274
rect 27764 9222 27776 9274
rect 27838 9222 27840 9274
rect 27678 9220 27702 9222
rect 27758 9220 27782 9222
rect 27838 9220 27862 9222
rect 27622 9200 27918 9220
rect 27712 9104 27764 9110
rect 27712 9046 27764 9052
rect 26974 9007 27030 9016
rect 27068 9036 27120 9042
rect 27068 8978 27120 8984
rect 26884 8560 26936 8566
rect 26884 8502 26936 8508
rect 27160 8560 27212 8566
rect 27160 8502 27212 8508
rect 26896 8362 26924 8502
rect 26884 8356 26936 8362
rect 26884 8298 26936 8304
rect 27172 8090 27200 8502
rect 27724 8498 27752 9046
rect 28080 9036 28132 9042
rect 28080 8978 28132 8984
rect 28092 8634 28120 8978
rect 28184 8838 28212 9386
rect 28172 8832 28224 8838
rect 28172 8774 28224 8780
rect 28080 8628 28132 8634
rect 28000 8588 28080 8616
rect 27712 8492 27764 8498
rect 27712 8434 27764 8440
rect 27712 8356 27764 8362
rect 27448 8316 27712 8344
rect 27448 8129 27476 8316
rect 27712 8298 27764 8304
rect 27622 8188 27918 8208
rect 27678 8186 27702 8188
rect 27758 8186 27782 8188
rect 27838 8186 27862 8188
rect 27700 8134 27702 8186
rect 27764 8134 27776 8186
rect 27838 8134 27840 8186
rect 27678 8132 27702 8134
rect 27758 8132 27782 8134
rect 27838 8132 27862 8134
rect 27434 8120 27490 8129
rect 27160 8084 27212 8090
rect 27622 8112 27918 8132
rect 27434 8055 27490 8064
rect 27160 8026 27212 8032
rect 26332 7948 26384 7954
rect 26332 7890 26384 7896
rect 27344 7948 27396 7954
rect 27344 7890 27396 7896
rect 26344 7857 26372 7890
rect 27160 7880 27212 7886
rect 26330 7848 26386 7857
rect 26330 7783 26386 7792
rect 27066 7848 27122 7857
rect 27160 7822 27212 7828
rect 27066 7783 27122 7792
rect 26344 7478 26372 7783
rect 26332 7472 26384 7478
rect 26332 7414 26384 7420
rect 27080 7410 27108 7783
rect 26056 7404 26108 7410
rect 26056 7346 26108 7352
rect 27068 7404 27120 7410
rect 27068 7346 27120 7352
rect 26068 7313 26096 7346
rect 26054 7304 26110 7313
rect 27172 7274 27200 7822
rect 26054 7239 26110 7248
rect 27160 7268 27212 7274
rect 27160 7210 27212 7216
rect 27068 7200 27120 7206
rect 25686 7168 25742 7177
rect 27068 7142 27120 7148
rect 25686 7103 25742 7112
rect 25700 6934 25728 7103
rect 27080 7041 27108 7142
rect 27066 7032 27122 7041
rect 27172 7002 27200 7210
rect 27066 6967 27122 6976
rect 27160 6996 27212 7002
rect 25688 6928 25740 6934
rect 25688 6870 25740 6876
rect 26608 6860 26660 6866
rect 26608 6802 26660 6808
rect 25778 6760 25834 6769
rect 25778 6695 25834 6704
rect 25792 6458 25820 6695
rect 25964 6656 26016 6662
rect 25964 6598 26016 6604
rect 25780 6452 25832 6458
rect 25780 6394 25832 6400
rect 25976 6118 26004 6598
rect 26422 6488 26478 6497
rect 26422 6423 26424 6432
rect 26476 6423 26478 6432
rect 26424 6394 26476 6400
rect 26332 6384 26384 6390
rect 26332 6326 26384 6332
rect 25964 6112 26016 6118
rect 25964 6054 26016 6060
rect 26344 5710 26372 6326
rect 26620 6186 26648 6802
rect 26700 6792 26752 6798
rect 26700 6734 26752 6740
rect 26608 6180 26660 6186
rect 26608 6122 26660 6128
rect 26332 5704 26384 5710
rect 26332 5646 26384 5652
rect 26620 5642 26648 6122
rect 26608 5636 26660 5642
rect 26608 5578 26660 5584
rect 26712 5574 26740 6734
rect 27080 6458 27108 6967
rect 27160 6938 27212 6944
rect 27356 6769 27384 7890
rect 27342 6760 27398 6769
rect 27342 6695 27398 6704
rect 27356 6458 27384 6695
rect 27068 6452 27120 6458
rect 27068 6394 27120 6400
rect 27344 6452 27396 6458
rect 27344 6394 27396 6400
rect 27356 6118 27384 6394
rect 27344 6112 27396 6118
rect 27344 6054 27396 6060
rect 27342 5808 27398 5817
rect 27342 5743 27398 5752
rect 25688 5568 25740 5574
rect 25688 5510 25740 5516
rect 26700 5568 26752 5574
rect 27160 5568 27212 5574
rect 26700 5510 26752 5516
rect 27158 5536 27160 5545
rect 27212 5536 27214 5545
rect 25700 5166 25728 5510
rect 26712 5370 26740 5510
rect 27158 5471 27214 5480
rect 27172 5370 27200 5471
rect 26700 5364 26752 5370
rect 26700 5306 26752 5312
rect 27160 5364 27212 5370
rect 27212 5324 27292 5352
rect 27160 5306 27212 5312
rect 25688 5160 25740 5166
rect 25688 5102 25740 5108
rect 25594 4992 25650 5001
rect 25594 4927 25650 4936
rect 25700 4826 25728 5102
rect 25688 4820 25740 4826
rect 25688 4762 25740 4768
rect 24950 4584 25006 4593
rect 24950 4519 25006 4528
rect 22652 4422 22704 4428
rect 24122 4448 24178 4457
rect 24122 4383 24178 4392
rect 22284 4140 22336 4146
rect 22284 4082 22336 4088
rect 22376 4140 22428 4146
rect 22376 4082 22428 4088
rect 27264 4010 27292 5324
rect 27252 4004 27304 4010
rect 27252 3946 27304 3952
rect 27264 3738 27292 3946
rect 27356 3942 27384 5743
rect 27448 4690 27476 8055
rect 28000 7546 28028 8588
rect 28080 8570 28132 8576
rect 28184 8265 28212 8774
rect 28170 8256 28226 8265
rect 28170 8191 28226 8200
rect 28080 7880 28132 7886
rect 28080 7822 28132 7828
rect 28170 7848 28226 7857
rect 27988 7540 28040 7546
rect 27988 7482 28040 7488
rect 28092 7342 28120 7822
rect 28170 7783 28226 7792
rect 28080 7336 28132 7342
rect 27526 7304 27582 7313
rect 28080 7278 28132 7284
rect 27526 7239 27582 7248
rect 27540 7206 27568 7239
rect 27528 7200 27580 7206
rect 27528 7142 27580 7148
rect 27988 7200 28040 7206
rect 27988 7142 28040 7148
rect 27622 7100 27918 7120
rect 27678 7098 27702 7100
rect 27758 7098 27782 7100
rect 27838 7098 27862 7100
rect 27700 7046 27702 7098
rect 27764 7046 27776 7098
rect 27838 7046 27840 7098
rect 27678 7044 27702 7046
rect 27758 7044 27782 7046
rect 27838 7044 27862 7046
rect 27622 7024 27918 7044
rect 27528 6180 27580 6186
rect 27528 6122 27580 6128
rect 27436 4684 27488 4690
rect 27436 4626 27488 4632
rect 27540 4554 27568 6122
rect 27622 6012 27918 6032
rect 27678 6010 27702 6012
rect 27758 6010 27782 6012
rect 27838 6010 27862 6012
rect 27700 5958 27702 6010
rect 27764 5958 27776 6010
rect 27838 5958 27840 6010
rect 27678 5956 27702 5958
rect 27758 5956 27782 5958
rect 27838 5956 27862 5958
rect 27622 5936 27918 5956
rect 27804 5840 27856 5846
rect 27804 5782 27856 5788
rect 27816 5370 27844 5782
rect 27804 5364 27856 5370
rect 27804 5306 27856 5312
rect 27622 4924 27918 4944
rect 27678 4922 27702 4924
rect 27758 4922 27782 4924
rect 27838 4922 27862 4924
rect 27700 4870 27702 4922
rect 27764 4870 27776 4922
rect 27838 4870 27840 4922
rect 27678 4868 27702 4870
rect 27758 4868 27782 4870
rect 27838 4868 27862 4870
rect 27622 4848 27918 4868
rect 27712 4752 27764 4758
rect 27712 4694 27764 4700
rect 27528 4548 27580 4554
rect 27528 4490 27580 4496
rect 27724 4282 27752 4694
rect 27896 4684 27948 4690
rect 27896 4626 27948 4632
rect 27908 4282 27936 4626
rect 27712 4276 27764 4282
rect 27712 4218 27764 4224
rect 27896 4276 27948 4282
rect 27896 4218 27948 4224
rect 27528 4072 27580 4078
rect 27526 4040 27528 4049
rect 27580 4040 27582 4049
rect 27526 3975 27582 3984
rect 27344 3936 27396 3942
rect 27908 3924 27936 4218
rect 28000 4146 28028 7142
rect 28184 6338 28212 7783
rect 28276 7585 28304 11494
rect 28448 11212 28500 11218
rect 28448 11154 28500 11160
rect 28460 10810 28488 11154
rect 29552 11076 29604 11082
rect 29552 11018 29604 11024
rect 28448 10804 28500 10810
rect 28448 10746 28500 10752
rect 29564 10713 29592 11018
rect 29550 10704 29606 10713
rect 29550 10639 29606 10648
rect 29092 10532 29144 10538
rect 29092 10474 29144 10480
rect 28908 10192 28960 10198
rect 29000 10192 29052 10198
rect 28960 10152 29000 10180
rect 28908 10134 28960 10140
rect 29000 10134 29052 10140
rect 28448 9920 28500 9926
rect 28448 9862 28500 9868
rect 28460 9110 28488 9862
rect 29104 9722 29132 10474
rect 30012 10464 30064 10470
rect 30012 10406 30064 10412
rect 30024 10198 30052 10406
rect 30012 10192 30064 10198
rect 30012 10134 30064 10140
rect 30208 9994 30236 11630
rect 30392 11218 30420 11766
rect 31036 11626 31064 12038
rect 31220 11642 31248 13670
rect 31680 12850 31708 15520
rect 33140 13932 33192 13938
rect 33140 13874 33192 13880
rect 32312 13320 32364 13326
rect 32312 13262 32364 13268
rect 31668 12844 31720 12850
rect 31668 12786 31720 12792
rect 32036 12708 32088 12714
rect 32036 12650 32088 12656
rect 31300 12300 31352 12306
rect 31300 12242 31352 12248
rect 31024 11620 31076 11626
rect 31024 11562 31076 11568
rect 31128 11614 31248 11642
rect 30930 11384 30986 11393
rect 30930 11319 30986 11328
rect 30944 11286 30972 11319
rect 30932 11280 30984 11286
rect 30932 11222 30984 11228
rect 30380 11212 30432 11218
rect 30380 11154 30432 11160
rect 30392 11098 30420 11154
rect 30300 11070 30420 11098
rect 30300 10810 30328 11070
rect 30840 11008 30892 11014
rect 30840 10950 30892 10956
rect 30288 10804 30340 10810
rect 30288 10746 30340 10752
rect 30852 10538 30880 10950
rect 30840 10532 30892 10538
rect 30840 10474 30892 10480
rect 30564 10124 30616 10130
rect 30564 10066 30616 10072
rect 30196 9988 30248 9994
rect 30196 9930 30248 9936
rect 29092 9716 29144 9722
rect 29092 9658 29144 9664
rect 30288 9716 30340 9722
rect 30288 9658 30340 9664
rect 28908 9580 28960 9586
rect 28908 9522 28960 9528
rect 28920 9382 28948 9522
rect 28540 9376 28592 9382
rect 28540 9318 28592 9324
rect 28908 9376 28960 9382
rect 28960 9336 29040 9364
rect 28908 9318 28960 9324
rect 28448 9104 28500 9110
rect 28448 9046 28500 9052
rect 28356 8560 28408 8566
rect 28356 8502 28408 8508
rect 28262 7576 28318 7585
rect 28262 7511 28318 7520
rect 28092 6310 28212 6338
rect 28092 4758 28120 6310
rect 28264 6180 28316 6186
rect 28264 6122 28316 6128
rect 28276 5710 28304 6122
rect 28368 5778 28396 8502
rect 28460 8090 28488 9046
rect 28552 8634 28580 9318
rect 28630 9208 28686 9217
rect 28630 9143 28686 9152
rect 28540 8628 28592 8634
rect 28540 8570 28592 8576
rect 28644 8514 28672 9143
rect 28552 8486 28672 8514
rect 28552 8430 28580 8486
rect 28540 8424 28592 8430
rect 28540 8366 28592 8372
rect 28448 8084 28500 8090
rect 28448 8026 28500 8032
rect 28446 7576 28502 7585
rect 28446 7511 28502 7520
rect 28356 5772 28408 5778
rect 28356 5714 28408 5720
rect 28264 5704 28316 5710
rect 28264 5646 28316 5652
rect 28276 5166 28304 5646
rect 28368 5370 28396 5714
rect 28460 5681 28488 7511
rect 28552 5846 28580 8366
rect 28908 7948 28960 7954
rect 28908 7890 28960 7896
rect 28920 7018 28948 7890
rect 29012 7546 29040 9336
rect 29104 7954 29132 9658
rect 29828 9648 29880 9654
rect 29826 9616 29828 9625
rect 29880 9616 29882 9625
rect 30300 9602 30328 9658
rect 30300 9586 30420 9602
rect 30300 9580 30432 9586
rect 30300 9574 30380 9580
rect 29826 9551 29882 9560
rect 30380 9522 30432 9528
rect 30288 9376 30340 9382
rect 30288 9318 30340 9324
rect 29184 8832 29236 8838
rect 29184 8774 29236 8780
rect 29196 8430 29224 8774
rect 30012 8492 30064 8498
rect 30012 8434 30064 8440
rect 29184 8424 29236 8430
rect 29184 8366 29236 8372
rect 29196 7954 29224 8366
rect 29092 7948 29144 7954
rect 29092 7890 29144 7896
rect 29184 7948 29236 7954
rect 29184 7890 29236 7896
rect 29090 7712 29146 7721
rect 29090 7647 29146 7656
rect 29000 7540 29052 7546
rect 29000 7482 29052 7488
rect 29104 7478 29132 7647
rect 29092 7472 29144 7478
rect 29092 7414 29144 7420
rect 29104 7274 29132 7414
rect 29196 7410 29224 7890
rect 30024 7449 30052 8434
rect 30010 7440 30066 7449
rect 29184 7404 29236 7410
rect 30010 7375 30066 7384
rect 29184 7346 29236 7352
rect 29092 7268 29144 7274
rect 29092 7210 29144 7216
rect 28920 6990 29040 7018
rect 29196 7002 29224 7346
rect 29828 7268 29880 7274
rect 29828 7210 29880 7216
rect 29840 7177 29868 7210
rect 29826 7168 29882 7177
rect 29826 7103 29882 7112
rect 28908 6928 28960 6934
rect 28908 6870 28960 6876
rect 28816 6656 28868 6662
rect 28920 6633 28948 6870
rect 29012 6798 29040 6990
rect 29184 6996 29236 7002
rect 29184 6938 29236 6944
rect 29920 6860 29972 6866
rect 29920 6802 29972 6808
rect 29000 6792 29052 6798
rect 29000 6734 29052 6740
rect 28816 6598 28868 6604
rect 28906 6624 28962 6633
rect 28828 6474 28856 6598
rect 28906 6559 28962 6568
rect 28828 6446 28948 6474
rect 29012 6458 29040 6734
rect 29932 6458 29960 6802
rect 28920 6361 28948 6446
rect 29000 6452 29052 6458
rect 29000 6394 29052 6400
rect 29920 6452 29972 6458
rect 29920 6394 29972 6400
rect 29552 6384 29604 6390
rect 28906 6352 28962 6361
rect 29552 6326 29604 6332
rect 29826 6352 29882 6361
rect 28906 6287 28962 6296
rect 29564 5846 29592 6326
rect 29826 6287 29882 6296
rect 29840 6186 29868 6287
rect 29828 6180 29880 6186
rect 29828 6122 29880 6128
rect 29644 5908 29696 5914
rect 29644 5850 29696 5856
rect 28540 5840 28592 5846
rect 28540 5782 28592 5788
rect 29552 5840 29604 5846
rect 29552 5782 29604 5788
rect 29276 5704 29328 5710
rect 28446 5672 28502 5681
rect 28446 5607 28502 5616
rect 28630 5672 28686 5681
rect 29182 5672 29238 5681
rect 28630 5607 28686 5616
rect 28816 5636 28868 5642
rect 28644 5409 28672 5607
rect 29276 5646 29328 5652
rect 29366 5672 29422 5681
rect 29182 5607 29238 5616
rect 28816 5578 28868 5584
rect 28630 5400 28686 5409
rect 28356 5364 28408 5370
rect 28630 5335 28686 5344
rect 28356 5306 28408 5312
rect 28264 5160 28316 5166
rect 28264 5102 28316 5108
rect 28276 4826 28304 5102
rect 28368 5001 28396 5306
rect 28828 5273 28856 5578
rect 28814 5264 28870 5273
rect 28814 5199 28870 5208
rect 29196 5030 29224 5607
rect 29288 5302 29316 5646
rect 29366 5607 29422 5616
rect 29380 5370 29408 5607
rect 29368 5364 29420 5370
rect 29368 5306 29420 5312
rect 29276 5296 29328 5302
rect 29276 5238 29328 5244
rect 29550 5264 29606 5273
rect 29288 5137 29316 5238
rect 29550 5199 29606 5208
rect 29564 5166 29592 5199
rect 29552 5160 29604 5166
rect 29274 5128 29330 5137
rect 29552 5102 29604 5108
rect 29274 5063 29330 5072
rect 29184 5024 29236 5030
rect 28354 4992 28410 5001
rect 29184 4966 29236 4972
rect 28354 4927 28410 4936
rect 29656 4826 29684 5850
rect 29828 5568 29880 5574
rect 29828 5510 29880 5516
rect 29840 5098 29868 5510
rect 29932 5234 29960 6394
rect 29920 5228 29972 5234
rect 29920 5170 29972 5176
rect 29828 5092 29880 5098
rect 29828 5034 29880 5040
rect 29840 4826 29868 5034
rect 28264 4820 28316 4826
rect 28264 4762 28316 4768
rect 29644 4820 29696 4826
rect 29644 4762 29696 4768
rect 29828 4820 29880 4826
rect 29828 4762 29880 4768
rect 28080 4752 28132 4758
rect 28080 4694 28132 4700
rect 28276 4282 28304 4762
rect 29932 4758 29960 5170
rect 29920 4752 29972 4758
rect 29920 4694 29972 4700
rect 28264 4276 28316 4282
rect 28264 4218 28316 4224
rect 27988 4140 28040 4146
rect 27988 4082 28040 4088
rect 27908 3896 28028 3924
rect 27344 3878 27396 3884
rect 27622 3836 27918 3856
rect 27678 3834 27702 3836
rect 27758 3834 27782 3836
rect 27838 3834 27862 3836
rect 27700 3782 27702 3834
rect 27764 3782 27776 3834
rect 27838 3782 27840 3834
rect 27678 3780 27702 3782
rect 27758 3780 27782 3782
rect 27838 3780 27862 3782
rect 27622 3760 27918 3780
rect 27252 3732 27304 3738
rect 27252 3674 27304 3680
rect 20956 3292 21252 3312
rect 21012 3290 21036 3292
rect 21092 3290 21116 3292
rect 21172 3290 21196 3292
rect 21034 3238 21036 3290
rect 21098 3238 21110 3290
rect 21172 3238 21174 3290
rect 21012 3236 21036 3238
rect 21092 3236 21116 3238
rect 21172 3236 21196 3238
rect 20956 3216 21252 3236
rect 27622 2748 27918 2768
rect 27678 2746 27702 2748
rect 27758 2746 27782 2748
rect 27838 2746 27862 2748
rect 27700 2694 27702 2746
rect 27764 2694 27776 2746
rect 27838 2694 27840 2746
rect 27678 2692 27702 2694
rect 27758 2692 27782 2694
rect 27838 2692 27862 2694
rect 27622 2672 27918 2692
rect 28000 2553 28028 3896
rect 30024 3777 30052 7375
rect 30300 6186 30328 9318
rect 30576 8906 30604 10066
rect 30852 10062 30880 10474
rect 30932 10192 30984 10198
rect 30932 10134 30984 10140
rect 30840 10056 30892 10062
rect 30840 9998 30892 10004
rect 30852 9874 30880 9998
rect 30760 9846 30880 9874
rect 30760 9722 30788 9846
rect 30748 9716 30800 9722
rect 30748 9658 30800 9664
rect 30748 9104 30800 9110
rect 30748 9046 30800 9052
rect 30838 9072 30894 9081
rect 30760 8945 30788 9046
rect 30838 9007 30840 9016
rect 30892 9007 30894 9016
rect 30840 8978 30892 8984
rect 30746 8936 30802 8945
rect 30564 8900 30616 8906
rect 30746 8871 30802 8880
rect 30564 8842 30616 8848
rect 30378 8528 30434 8537
rect 30378 8463 30434 8472
rect 30392 8294 30420 8463
rect 30656 8424 30708 8430
rect 30654 8392 30656 8401
rect 30708 8392 30710 8401
rect 30654 8327 30710 8336
rect 30380 8288 30432 8294
rect 30380 8230 30432 8236
rect 30470 8256 30526 8265
rect 30470 8191 30526 8200
rect 30484 8090 30512 8191
rect 30760 8090 30788 8871
rect 30852 8566 30880 8978
rect 30944 8634 30972 10134
rect 31024 9920 31076 9926
rect 31024 9862 31076 9868
rect 31036 9450 31064 9862
rect 31024 9444 31076 9450
rect 31024 9386 31076 9392
rect 31036 8974 31064 9386
rect 31024 8968 31076 8974
rect 31024 8910 31076 8916
rect 30932 8628 30984 8634
rect 30932 8570 30984 8576
rect 30840 8560 30892 8566
rect 30840 8502 30892 8508
rect 31128 8430 31156 11614
rect 31312 11558 31340 12242
rect 31942 11928 31998 11937
rect 31942 11863 31944 11872
rect 31996 11863 31998 11872
rect 31944 11834 31996 11840
rect 31956 11694 31984 11834
rect 31668 11688 31720 11694
rect 31668 11630 31720 11636
rect 31944 11688 31996 11694
rect 31944 11630 31996 11636
rect 31208 11552 31260 11558
rect 31208 11494 31260 11500
rect 31300 11552 31352 11558
rect 31300 11494 31352 11500
rect 31220 10810 31248 11494
rect 31208 10804 31260 10810
rect 31208 10746 31260 10752
rect 31116 8424 31168 8430
rect 31116 8366 31168 8372
rect 30472 8084 30524 8090
rect 30472 8026 30524 8032
rect 30748 8084 30800 8090
rect 30748 8026 30800 8032
rect 30760 7449 30788 8026
rect 30746 7440 30802 7449
rect 30746 7375 30802 7384
rect 30748 6792 30800 6798
rect 30748 6734 30800 6740
rect 30760 6254 30788 6734
rect 31312 6497 31340 11494
rect 31680 10962 31708 11630
rect 31680 10934 31800 10962
rect 31668 10804 31720 10810
rect 31668 10746 31720 10752
rect 31680 10198 31708 10746
rect 31668 10192 31720 10198
rect 31668 10134 31720 10140
rect 31668 10056 31720 10062
rect 31668 9998 31720 10004
rect 31680 9382 31708 9998
rect 31668 9376 31720 9382
rect 31668 9318 31720 9324
rect 31484 8968 31536 8974
rect 31484 8910 31536 8916
rect 31496 8537 31524 8910
rect 31772 8906 31800 10934
rect 31852 10192 31904 10198
rect 31852 10134 31904 10140
rect 31864 9110 31892 10134
rect 31944 9376 31996 9382
rect 31944 9318 31996 9324
rect 31852 9104 31904 9110
rect 31852 9046 31904 9052
rect 31956 9042 31984 9318
rect 31944 9036 31996 9042
rect 31944 8978 31996 8984
rect 31760 8900 31812 8906
rect 31760 8842 31812 8848
rect 31482 8528 31538 8537
rect 31482 8463 31484 8472
rect 31536 8463 31538 8472
rect 31484 8434 31536 8440
rect 31496 8090 31524 8434
rect 31956 8090 31984 8978
rect 31484 8084 31536 8090
rect 31484 8026 31536 8032
rect 31944 8084 31996 8090
rect 31944 8026 31996 8032
rect 31760 7472 31812 7478
rect 31760 7414 31812 7420
rect 31576 7404 31628 7410
rect 31576 7346 31628 7352
rect 31484 7268 31536 7274
rect 31484 7210 31536 7216
rect 31392 7200 31444 7206
rect 31392 7142 31444 7148
rect 31404 6905 31432 7142
rect 31496 7002 31524 7210
rect 31484 6996 31536 7002
rect 31484 6938 31536 6944
rect 31390 6896 31446 6905
rect 31390 6831 31446 6840
rect 31484 6656 31536 6662
rect 31588 6644 31616 7346
rect 31772 6866 31800 7414
rect 31760 6860 31812 6866
rect 31760 6802 31812 6808
rect 31536 6616 31616 6644
rect 31484 6598 31536 6604
rect 31298 6488 31354 6497
rect 31298 6423 31354 6432
rect 30748 6248 30800 6254
rect 30748 6190 30800 6196
rect 30288 6180 30340 6186
rect 30288 6122 30340 6128
rect 30760 5914 30788 6190
rect 30748 5908 30800 5914
rect 30748 5850 30800 5856
rect 30380 5840 30432 5846
rect 30380 5782 30432 5788
rect 30392 5370 30420 5782
rect 30380 5364 30432 5370
rect 30380 5306 30432 5312
rect 31496 4049 31524 6598
rect 31772 5914 31800 6802
rect 32048 6730 32076 12650
rect 32324 12442 32352 13262
rect 33152 12918 33180 13874
rect 33416 13388 33468 13394
rect 33416 13330 33468 13336
rect 33140 12912 33192 12918
rect 33140 12854 33192 12860
rect 32312 12436 32364 12442
rect 32312 12378 32364 12384
rect 32956 12300 33008 12306
rect 32956 12242 33008 12248
rect 33324 12300 33376 12306
rect 33324 12242 33376 12248
rect 32772 12096 32824 12102
rect 32772 12038 32824 12044
rect 32312 11552 32364 11558
rect 32310 11520 32312 11529
rect 32364 11520 32366 11529
rect 32310 11455 32366 11464
rect 32680 11280 32732 11286
rect 32680 11222 32732 11228
rect 32692 10810 32720 11222
rect 32680 10804 32732 10810
rect 32680 10746 32732 10752
rect 32784 10606 32812 12038
rect 32864 11824 32916 11830
rect 32864 11766 32916 11772
rect 32876 11150 32904 11766
rect 32968 11558 32996 12242
rect 33138 12064 33194 12073
rect 33138 11999 33194 12008
rect 33152 11558 33180 11999
rect 33336 11898 33364 12242
rect 33324 11892 33376 11898
rect 33324 11834 33376 11840
rect 32956 11552 33008 11558
rect 32956 11494 33008 11500
rect 33140 11552 33192 11558
rect 33140 11494 33192 11500
rect 32864 11144 32916 11150
rect 32864 11086 32916 11092
rect 32876 10810 32904 11086
rect 32864 10804 32916 10810
rect 32864 10746 32916 10752
rect 32772 10600 32824 10606
rect 32772 10542 32824 10548
rect 32876 10130 32904 10746
rect 32968 10577 32996 11494
rect 33048 11212 33100 11218
rect 33048 11154 33100 11160
rect 33060 11098 33088 11154
rect 33060 11070 33180 11098
rect 33152 10674 33180 11070
rect 33140 10668 33192 10674
rect 33140 10610 33192 10616
rect 32954 10568 33010 10577
rect 32954 10503 33010 10512
rect 32968 10146 32996 10503
rect 32864 10124 32916 10130
rect 32968 10118 33272 10146
rect 32864 10066 32916 10072
rect 32588 9920 32640 9926
rect 32588 9862 32640 9868
rect 32600 9058 32628 9862
rect 32876 9364 32904 10066
rect 32956 9376 33008 9382
rect 32876 9336 32956 9364
rect 32956 9318 33008 9324
rect 33140 9376 33192 9382
rect 33140 9318 33192 9324
rect 32678 9072 32734 9081
rect 32600 9030 32678 9058
rect 32678 9007 32734 9016
rect 32692 8974 32720 9007
rect 32680 8968 32732 8974
rect 32680 8910 32732 8916
rect 32494 8664 32550 8673
rect 32494 8599 32550 8608
rect 32508 8362 32536 8599
rect 32772 8560 32824 8566
rect 32770 8528 32772 8537
rect 32824 8528 32826 8537
rect 32770 8463 32826 8472
rect 32968 8430 32996 9318
rect 33152 9217 33180 9318
rect 33138 9208 33194 9217
rect 33138 9143 33194 9152
rect 33140 9036 33192 9042
rect 33140 8978 33192 8984
rect 33048 8560 33100 8566
rect 33048 8502 33100 8508
rect 32956 8424 33008 8430
rect 32956 8366 33008 8372
rect 32496 8356 32548 8362
rect 32496 8298 32548 8304
rect 32220 8288 32272 8294
rect 32220 8230 32272 8236
rect 32036 6724 32088 6730
rect 32036 6666 32088 6672
rect 31760 5908 31812 5914
rect 31760 5850 31812 5856
rect 32232 4049 32260 8230
rect 32770 7984 32826 7993
rect 32404 7948 32456 7954
rect 32770 7919 32826 7928
rect 32404 7890 32456 7896
rect 32416 7546 32444 7890
rect 32404 7540 32456 7546
rect 32404 7482 32456 7488
rect 32680 6928 32732 6934
rect 32680 6870 32732 6876
rect 32404 6792 32456 6798
rect 32404 6734 32456 6740
rect 32416 6458 32444 6734
rect 32404 6452 32456 6458
rect 32404 6394 32456 6400
rect 32586 5944 32642 5953
rect 32692 5914 32720 6870
rect 32586 5879 32642 5888
rect 32680 5908 32732 5914
rect 32600 5302 32628 5879
rect 32680 5850 32732 5856
rect 32692 5681 32720 5850
rect 32678 5672 32734 5681
rect 32784 5642 32812 7919
rect 32968 7886 32996 8366
rect 32956 7880 33008 7886
rect 32876 7828 32956 7834
rect 32876 7822 33008 7828
rect 32876 7806 32996 7822
rect 32876 7478 32904 7806
rect 32956 7744 33008 7750
rect 32956 7686 33008 7692
rect 32864 7472 32916 7478
rect 32864 7414 32916 7420
rect 32862 7032 32918 7041
rect 32862 6967 32918 6976
rect 32678 5607 32734 5616
rect 32772 5636 32824 5642
rect 32772 5578 32824 5584
rect 32588 5296 32640 5302
rect 32588 5238 32640 5244
rect 32876 5234 32904 6967
rect 32772 5228 32824 5234
rect 32772 5170 32824 5176
rect 32864 5228 32916 5234
rect 32864 5170 32916 5176
rect 32784 4826 32812 5170
rect 32772 4820 32824 4826
rect 32772 4762 32824 4768
rect 32876 4758 32904 5170
rect 32968 4826 32996 7686
rect 33060 5370 33088 8502
rect 33152 7750 33180 8978
rect 33140 7744 33192 7750
rect 33140 7686 33192 7692
rect 33244 7342 33272 10118
rect 33428 8498 33456 13330
rect 33968 13184 34020 13190
rect 33968 13126 34020 13132
rect 33508 12912 33560 12918
rect 33508 12854 33560 12860
rect 33520 12714 33548 12854
rect 33784 12844 33836 12850
rect 33784 12786 33836 12792
rect 33508 12708 33560 12714
rect 33508 12650 33560 12656
rect 33796 12170 33824 12786
rect 33980 12646 34008 13126
rect 33968 12640 34020 12646
rect 33968 12582 34020 12588
rect 33784 12164 33836 12170
rect 33784 12106 33836 12112
rect 33692 12096 33744 12102
rect 33692 12038 33744 12044
rect 33704 11778 33732 12038
rect 33782 11792 33838 11801
rect 33704 11750 33782 11778
rect 33782 11727 33784 11736
rect 33836 11727 33838 11736
rect 33784 11698 33836 11704
rect 33876 11688 33928 11694
rect 33876 11630 33928 11636
rect 33784 11552 33836 11558
rect 33784 11494 33836 11500
rect 33692 11008 33744 11014
rect 33692 10950 33744 10956
rect 33704 10742 33732 10950
rect 33692 10736 33744 10742
rect 33796 10713 33824 11494
rect 33888 11286 33916 11630
rect 33876 11280 33928 11286
rect 33876 11222 33928 11228
rect 33876 11008 33928 11014
rect 33876 10950 33928 10956
rect 33692 10678 33744 10684
rect 33782 10704 33838 10713
rect 33704 10538 33732 10678
rect 33782 10639 33838 10648
rect 33888 10606 33916 10950
rect 33980 10810 34008 12582
rect 34072 11393 34100 15520
rect 34532 13870 34560 15807
rect 36358 15520 36414 16000
rect 38750 15520 38806 16000
rect 34610 15464 34666 15473
rect 34610 15399 34666 15408
rect 34520 13864 34572 13870
rect 34520 13806 34572 13812
rect 34624 13530 34652 15399
rect 34702 14648 34758 14657
rect 34702 14583 34758 14592
rect 34612 13524 34664 13530
rect 34612 13466 34664 13472
rect 34152 13388 34204 13394
rect 34152 13330 34204 13336
rect 34164 12968 34192 13330
rect 34716 13258 34744 14583
rect 34794 14240 34850 14249
rect 34794 14175 34850 14184
rect 34808 13938 34836 14175
rect 34796 13932 34848 13938
rect 34796 13874 34848 13880
rect 36176 13728 36228 13734
rect 36176 13670 36228 13676
rect 35346 13424 35402 13433
rect 35256 13388 35308 13394
rect 35346 13359 35402 13368
rect 35256 13330 35308 13336
rect 34796 13320 34848 13326
rect 34796 13262 34848 13268
rect 34704 13252 34756 13258
rect 34704 13194 34756 13200
rect 34289 13084 34585 13104
rect 34345 13082 34369 13084
rect 34425 13082 34449 13084
rect 34505 13082 34529 13084
rect 34367 13030 34369 13082
rect 34431 13030 34443 13082
rect 34505 13030 34507 13082
rect 34345 13028 34369 13030
rect 34425 13028 34449 13030
rect 34505 13028 34529 13030
rect 34289 13008 34585 13028
rect 34808 13025 34836 13262
rect 34888 13184 34940 13190
rect 34888 13126 34940 13132
rect 34794 13016 34850 13025
rect 34612 12980 34664 12986
rect 34164 12940 34376 12968
rect 34348 12646 34376 12940
rect 34794 12951 34850 12960
rect 34612 12922 34664 12928
rect 34624 12753 34652 12922
rect 34796 12912 34848 12918
rect 34796 12854 34848 12860
rect 34610 12744 34666 12753
rect 34610 12679 34666 12688
rect 34336 12640 34388 12646
rect 34336 12582 34388 12588
rect 34348 12209 34376 12582
rect 34334 12200 34390 12209
rect 34334 12135 34390 12144
rect 34612 12164 34664 12170
rect 34612 12106 34664 12112
rect 34289 11996 34585 12016
rect 34345 11994 34369 11996
rect 34425 11994 34449 11996
rect 34505 11994 34529 11996
rect 34367 11942 34369 11994
rect 34431 11942 34443 11994
rect 34505 11942 34507 11994
rect 34345 11940 34369 11942
rect 34425 11940 34449 11942
rect 34505 11940 34529 11942
rect 34289 11920 34585 11940
rect 34624 11898 34652 12106
rect 34612 11892 34664 11898
rect 34612 11834 34664 11840
rect 34152 11824 34204 11830
rect 34152 11766 34204 11772
rect 34058 11384 34114 11393
rect 34058 11319 34114 11328
rect 33968 10804 34020 10810
rect 33968 10746 34020 10752
rect 34164 10674 34192 11766
rect 34610 11656 34666 11665
rect 34610 11591 34612 11600
rect 34664 11591 34666 11600
rect 34612 11562 34664 11568
rect 34518 11112 34574 11121
rect 34518 11047 34520 11056
rect 34572 11047 34574 11056
rect 34520 11018 34572 11024
rect 34289 10908 34585 10928
rect 34345 10906 34369 10908
rect 34425 10906 34449 10908
rect 34505 10906 34529 10908
rect 34367 10854 34369 10906
rect 34431 10854 34443 10906
rect 34505 10854 34507 10906
rect 34345 10852 34369 10854
rect 34425 10852 34449 10854
rect 34505 10852 34529 10854
rect 34289 10832 34585 10852
rect 34152 10668 34204 10674
rect 34152 10610 34204 10616
rect 33876 10600 33928 10606
rect 33876 10542 33928 10548
rect 33692 10532 33744 10538
rect 33692 10474 33744 10480
rect 34612 10464 34664 10470
rect 34612 10406 34664 10412
rect 34150 10160 34206 10169
rect 34150 10095 34206 10104
rect 33876 9920 33928 9926
rect 33876 9862 33928 9868
rect 33888 9450 33916 9862
rect 34164 9761 34192 10095
rect 34624 10033 34652 10406
rect 34610 10024 34666 10033
rect 34610 9959 34666 9968
rect 34289 9820 34585 9840
rect 34345 9818 34369 9820
rect 34425 9818 34449 9820
rect 34505 9818 34529 9820
rect 34367 9766 34369 9818
rect 34431 9766 34443 9818
rect 34505 9766 34507 9818
rect 34345 9764 34369 9766
rect 34425 9764 34449 9766
rect 34505 9764 34529 9766
rect 34150 9752 34206 9761
rect 34289 9744 34585 9764
rect 34150 9687 34206 9696
rect 34624 9466 34652 9959
rect 34704 9920 34756 9926
rect 34704 9862 34756 9868
rect 33692 9444 33744 9450
rect 33692 9386 33744 9392
rect 33876 9444 33928 9450
rect 33876 9386 33928 9392
rect 34532 9438 34652 9466
rect 34716 9450 34744 9862
rect 34704 9444 34756 9450
rect 33600 8968 33652 8974
rect 33600 8910 33652 8916
rect 33416 8492 33468 8498
rect 33416 8434 33468 8440
rect 33612 8362 33640 8910
rect 33704 8906 33732 9386
rect 33692 8900 33744 8906
rect 33692 8842 33744 8848
rect 33600 8356 33652 8362
rect 33600 8298 33652 8304
rect 33508 8288 33560 8294
rect 33508 8230 33560 8236
rect 33324 7472 33376 7478
rect 33324 7414 33376 7420
rect 33232 7336 33284 7342
rect 33232 7278 33284 7284
rect 33140 7200 33192 7206
rect 33140 7142 33192 7148
rect 33152 6662 33180 7142
rect 33140 6656 33192 6662
rect 33140 6598 33192 6604
rect 33152 6458 33180 6598
rect 33140 6452 33192 6458
rect 33140 6394 33192 6400
rect 33232 5772 33284 5778
rect 33232 5714 33284 5720
rect 33048 5364 33100 5370
rect 33048 5306 33100 5312
rect 33060 5098 33088 5306
rect 33244 5234 33272 5714
rect 33336 5710 33364 7414
rect 33416 5840 33468 5846
rect 33416 5782 33468 5788
rect 33324 5704 33376 5710
rect 33324 5646 33376 5652
rect 33232 5228 33284 5234
rect 33232 5170 33284 5176
rect 33048 5092 33100 5098
rect 33048 5034 33100 5040
rect 33336 4826 33364 5646
rect 33428 5166 33456 5782
rect 33416 5160 33468 5166
rect 33520 5137 33548 8230
rect 33612 8090 33640 8298
rect 33600 8084 33652 8090
rect 33600 8026 33652 8032
rect 33612 7478 33640 8026
rect 33600 7472 33652 7478
rect 33600 7414 33652 7420
rect 33704 7290 33732 8842
rect 33784 8832 33836 8838
rect 33784 8774 33836 8780
rect 33612 7262 33732 7290
rect 33416 5102 33468 5108
rect 33506 5128 33562 5137
rect 32956 4820 33008 4826
rect 32956 4762 33008 4768
rect 33324 4820 33376 4826
rect 33324 4762 33376 4768
rect 32864 4752 32916 4758
rect 32864 4694 32916 4700
rect 33428 4554 33456 5102
rect 33506 5063 33562 5072
rect 33612 5001 33640 7262
rect 33796 7041 33824 8774
rect 33888 8362 33916 9386
rect 34152 9104 34204 9110
rect 34152 9046 34204 9052
rect 34164 8956 34192 9046
rect 34072 8928 34192 8956
rect 33968 8900 34020 8906
rect 33968 8842 34020 8848
rect 33876 8356 33928 8362
rect 33876 8298 33928 8304
rect 33980 8242 34008 8842
rect 34072 8809 34100 8928
rect 34532 8906 34560 9438
rect 34704 9386 34756 9392
rect 34612 9376 34664 9382
rect 34612 9318 34664 9324
rect 34520 8900 34572 8906
rect 34520 8842 34572 8848
rect 34058 8800 34114 8809
rect 34058 8735 34114 8744
rect 34072 8430 34100 8735
rect 34289 8732 34585 8752
rect 34345 8730 34369 8732
rect 34425 8730 34449 8732
rect 34505 8730 34529 8732
rect 34367 8678 34369 8730
rect 34431 8678 34443 8730
rect 34505 8678 34507 8730
rect 34345 8676 34369 8678
rect 34425 8676 34449 8678
rect 34505 8676 34529 8678
rect 34289 8656 34585 8676
rect 34060 8424 34112 8430
rect 34060 8366 34112 8372
rect 33888 8214 34008 8242
rect 33782 7032 33838 7041
rect 33782 6967 33838 6976
rect 33784 6724 33836 6730
rect 33784 6666 33836 6672
rect 33692 6656 33744 6662
rect 33692 6598 33744 6604
rect 33704 6390 33732 6598
rect 33692 6384 33744 6390
rect 33692 6326 33744 6332
rect 33704 5914 33732 6326
rect 33796 6322 33824 6666
rect 33784 6316 33836 6322
rect 33784 6258 33836 6264
rect 33796 6089 33824 6258
rect 33782 6080 33838 6089
rect 33782 6015 33838 6024
rect 33692 5908 33744 5914
rect 33692 5850 33744 5856
rect 33598 4992 33654 5001
rect 33598 4927 33654 4936
rect 33416 4548 33468 4554
rect 33416 4490 33468 4496
rect 31482 4040 31538 4049
rect 31482 3975 31538 3984
rect 32218 4040 32274 4049
rect 32218 3975 32274 3984
rect 30010 3768 30066 3777
rect 30010 3703 30066 3712
rect 33796 2961 33824 6015
rect 33888 5794 33916 8214
rect 33968 7404 34020 7410
rect 33968 7346 34020 7352
rect 33980 7002 34008 7346
rect 33968 6996 34020 7002
rect 33968 6938 34020 6944
rect 34072 6769 34100 8366
rect 34336 8356 34388 8362
rect 34336 8298 34388 8304
rect 34348 8090 34376 8298
rect 34336 8084 34388 8090
rect 34336 8026 34388 8032
rect 34624 7834 34652 9318
rect 34716 8430 34744 9386
rect 34704 8424 34756 8430
rect 34704 8366 34756 8372
rect 34716 8294 34744 8366
rect 34704 8288 34756 8294
rect 34704 8230 34756 8236
rect 34164 7806 34744 7834
rect 34808 7818 34836 12854
rect 34900 12782 34928 13126
rect 34888 12776 34940 12782
rect 34888 12718 34940 12724
rect 35268 12646 35296 13330
rect 35256 12640 35308 12646
rect 35256 12582 35308 12588
rect 34888 11552 34940 11558
rect 34888 11494 34940 11500
rect 34900 11082 34928 11494
rect 34888 11076 34940 11082
rect 34888 11018 34940 11024
rect 34900 9602 34928 11018
rect 35164 10736 35216 10742
rect 35070 10704 35126 10713
rect 35164 10678 35216 10684
rect 35070 10639 35126 10648
rect 34900 9574 35020 9602
rect 34886 9480 34942 9489
rect 34886 9415 34888 9424
rect 34940 9415 34942 9424
rect 34888 9386 34940 9392
rect 34900 9110 34928 9386
rect 34888 9104 34940 9110
rect 34888 9046 34940 9052
rect 34164 7585 34192 7806
rect 34289 7644 34585 7664
rect 34345 7642 34369 7644
rect 34425 7642 34449 7644
rect 34505 7642 34529 7644
rect 34367 7590 34369 7642
rect 34431 7590 34443 7642
rect 34505 7590 34507 7642
rect 34345 7588 34369 7590
rect 34425 7588 34449 7590
rect 34505 7588 34529 7590
rect 34150 7576 34206 7585
rect 34289 7568 34585 7588
rect 34150 7511 34206 7520
rect 34612 7268 34664 7274
rect 34612 7210 34664 7216
rect 34520 6928 34572 6934
rect 34520 6870 34572 6876
rect 34532 6798 34560 6870
rect 34520 6792 34572 6798
rect 34058 6760 34114 6769
rect 34520 6734 34572 6740
rect 34058 6695 34114 6704
rect 34289 6556 34585 6576
rect 34345 6554 34369 6556
rect 34425 6554 34449 6556
rect 34505 6554 34529 6556
rect 34367 6502 34369 6554
rect 34431 6502 34443 6554
rect 34505 6502 34507 6554
rect 34345 6500 34369 6502
rect 34425 6500 34449 6502
rect 34505 6500 34529 6502
rect 34289 6480 34585 6500
rect 34244 5840 34296 5846
rect 33888 5788 34244 5794
rect 34624 5794 34652 7210
rect 33888 5782 34296 5788
rect 33888 5766 34284 5782
rect 34440 5778 34652 5794
rect 34428 5772 34652 5778
rect 34060 5636 34112 5642
rect 34060 5578 34112 5584
rect 34072 4758 34100 5578
rect 34164 5370 34192 5766
rect 34480 5766 34652 5772
rect 34428 5714 34480 5720
rect 34612 5704 34664 5710
rect 34612 5646 34664 5652
rect 34289 5468 34585 5488
rect 34345 5466 34369 5468
rect 34425 5466 34449 5468
rect 34505 5466 34529 5468
rect 34367 5414 34369 5466
rect 34431 5414 34443 5466
rect 34505 5414 34507 5466
rect 34345 5412 34369 5414
rect 34425 5412 34449 5414
rect 34505 5412 34529 5414
rect 34289 5392 34585 5412
rect 34152 5364 34204 5370
rect 34152 5306 34204 5312
rect 34624 5302 34652 5646
rect 34716 5370 34744 7806
rect 34796 7812 34848 7818
rect 34796 7754 34848 7760
rect 34796 6860 34848 6866
rect 34796 6802 34848 6808
rect 34704 5364 34756 5370
rect 34704 5306 34756 5312
rect 34612 5296 34664 5302
rect 34612 5238 34664 5244
rect 34060 4752 34112 4758
rect 34060 4694 34112 4700
rect 34072 4282 34100 4694
rect 34289 4380 34585 4400
rect 34345 4378 34369 4380
rect 34425 4378 34449 4380
rect 34505 4378 34529 4380
rect 34367 4326 34369 4378
rect 34431 4326 34443 4378
rect 34505 4326 34507 4378
rect 34345 4324 34369 4326
rect 34425 4324 34449 4326
rect 34505 4324 34529 4326
rect 34289 4304 34585 4324
rect 34060 4276 34112 4282
rect 34060 4218 34112 4224
rect 34624 4026 34652 5238
rect 34716 5030 34744 5306
rect 34704 5024 34756 5030
rect 34704 4966 34756 4972
rect 34808 4758 34836 6802
rect 34900 5166 34928 9046
rect 34992 7954 35020 9574
rect 34980 7948 35032 7954
rect 34980 7890 35032 7896
rect 34980 7744 35032 7750
rect 34980 7686 35032 7692
rect 34992 7274 35020 7686
rect 35084 7585 35112 10639
rect 35176 10470 35204 10678
rect 35164 10464 35216 10470
rect 35164 10406 35216 10412
rect 35164 8288 35216 8294
rect 35164 8230 35216 8236
rect 35070 7576 35126 7585
rect 35070 7511 35126 7520
rect 35176 7426 35204 8230
rect 35268 7857 35296 12582
rect 35254 7848 35310 7857
rect 35254 7783 35310 7792
rect 35256 7744 35308 7750
rect 35256 7686 35308 7692
rect 35084 7398 35204 7426
rect 35084 7342 35112 7398
rect 35072 7336 35124 7342
rect 35072 7278 35124 7284
rect 35162 7304 35218 7313
rect 34980 7268 35032 7274
rect 34980 7210 35032 7216
rect 35084 7206 35112 7278
rect 35162 7239 35218 7248
rect 35072 7200 35124 7206
rect 34992 7148 35072 7154
rect 34992 7142 35124 7148
rect 34992 7126 35112 7142
rect 34992 6934 35020 7126
rect 35176 7041 35204 7239
rect 35162 7032 35218 7041
rect 35162 6967 35218 6976
rect 34980 6928 35032 6934
rect 35268 6905 35296 7686
rect 34980 6870 35032 6876
rect 35254 6896 35310 6905
rect 34992 6254 35020 6870
rect 35254 6831 35310 6840
rect 35070 6488 35126 6497
rect 35070 6423 35126 6432
rect 34980 6248 35032 6254
rect 34980 6190 35032 6196
rect 34992 5710 35020 6190
rect 35084 5817 35112 6423
rect 35164 6180 35216 6186
rect 35164 6122 35216 6128
rect 35176 5914 35204 6122
rect 35164 5908 35216 5914
rect 35164 5850 35216 5856
rect 35070 5808 35126 5817
rect 35070 5743 35126 5752
rect 34980 5704 35032 5710
rect 34980 5646 35032 5652
rect 34980 5296 35032 5302
rect 34980 5238 35032 5244
rect 34888 5160 34940 5166
rect 34888 5102 34940 5108
rect 34796 4752 34848 4758
rect 34796 4694 34848 4700
rect 34808 4214 34836 4694
rect 34900 4690 34928 5102
rect 34992 4826 35020 5238
rect 35176 5234 35204 5850
rect 35164 5228 35216 5234
rect 35164 5170 35216 5176
rect 35070 4992 35126 5001
rect 35070 4927 35126 4936
rect 34980 4820 35032 4826
rect 34980 4762 35032 4768
rect 34888 4684 34940 4690
rect 34888 4626 34940 4632
rect 34796 4208 34848 4214
rect 34796 4150 34848 4156
rect 34900 4162 34928 4626
rect 34992 4282 35020 4762
rect 35084 4706 35112 4927
rect 35176 4826 35204 5170
rect 35164 4820 35216 4826
rect 35164 4762 35216 4768
rect 35084 4678 35204 4706
rect 34980 4276 35032 4282
rect 34980 4218 35032 4224
rect 34900 4134 35112 4162
rect 34624 3998 34928 4026
rect 34289 3292 34585 3312
rect 34345 3290 34369 3292
rect 34425 3290 34449 3292
rect 34505 3290 34529 3292
rect 34367 3238 34369 3290
rect 34431 3238 34443 3290
rect 34505 3238 34507 3290
rect 34345 3236 34369 3238
rect 34425 3236 34449 3238
rect 34505 3236 34529 3238
rect 34289 3216 34585 3236
rect 33782 2952 33838 2961
rect 33782 2887 33838 2896
rect 27986 2544 28042 2553
rect 27986 2479 28042 2488
rect 20956 2204 21252 2224
rect 21012 2202 21036 2204
rect 21092 2202 21116 2204
rect 21172 2202 21196 2204
rect 21034 2150 21036 2202
rect 21098 2150 21110 2202
rect 21172 2150 21174 2202
rect 21012 2148 21036 2150
rect 21092 2148 21116 2150
rect 21172 2148 21196 2150
rect 20956 2128 21252 2148
rect 34289 2204 34585 2224
rect 34345 2202 34369 2204
rect 34425 2202 34449 2204
rect 34505 2202 34529 2204
rect 34367 2150 34369 2202
rect 34431 2150 34443 2202
rect 34505 2150 34507 2202
rect 34345 2148 34369 2150
rect 34425 2148 34449 2150
rect 34505 2148 34529 2150
rect 34289 2128 34585 2148
rect 22006 1864 22062 1873
rect 22006 1799 22062 1808
rect 22020 1465 22048 1799
rect 22006 1456 22062 1465
rect 22006 1391 22062 1400
rect 34900 1329 34928 3998
rect 34886 1320 34942 1329
rect 34886 1255 34942 1264
rect 35084 513 35112 4134
rect 35070 504 35126 513
rect 3606 232 3662 241
rect 3606 167 3662 176
rect 19982 0 20038 480
rect 35070 439 35126 448
rect 35176 241 35204 4678
rect 35360 3942 35388 13359
rect 35440 13184 35492 13190
rect 35440 13126 35492 13132
rect 35808 13184 35860 13190
rect 35808 13126 35860 13132
rect 35452 10305 35480 13126
rect 35714 12200 35770 12209
rect 35714 12135 35770 12144
rect 35532 12096 35584 12102
rect 35532 12038 35584 12044
rect 35544 11082 35572 12038
rect 35728 11286 35756 12135
rect 35716 11280 35768 11286
rect 35716 11222 35768 11228
rect 35532 11076 35584 11082
rect 35532 11018 35584 11024
rect 35624 11008 35676 11014
rect 35624 10950 35676 10956
rect 35532 10532 35584 10538
rect 35532 10474 35584 10480
rect 35438 10296 35494 10305
rect 35544 10266 35572 10474
rect 35636 10470 35664 10950
rect 35728 10810 35756 11222
rect 35820 11121 35848 13126
rect 36188 12782 36216 13670
rect 36372 12850 36400 15520
rect 36450 15056 36506 15065
rect 36450 14991 36506 15000
rect 36464 12986 36492 14991
rect 36634 13832 36690 13841
rect 36634 13767 36690 13776
rect 36452 12980 36504 12986
rect 36452 12922 36504 12928
rect 36360 12844 36412 12850
rect 36360 12786 36412 12792
rect 36176 12776 36228 12782
rect 36176 12718 36228 12724
rect 36268 12708 36320 12714
rect 36268 12650 36320 12656
rect 36280 12442 36308 12650
rect 36268 12436 36320 12442
rect 36268 12378 36320 12384
rect 36268 12300 36320 12306
rect 36268 12242 36320 12248
rect 36280 11898 36308 12242
rect 36268 11892 36320 11898
rect 36268 11834 36320 11840
rect 35992 11688 36044 11694
rect 35992 11630 36044 11636
rect 35806 11112 35862 11121
rect 35806 11047 35862 11056
rect 35716 10804 35768 10810
rect 35716 10746 35768 10752
rect 36004 10742 36032 11630
rect 36084 11552 36136 11558
rect 36084 11494 36136 11500
rect 36096 11150 36124 11494
rect 36360 11280 36412 11286
rect 36360 11222 36412 11228
rect 36084 11144 36136 11150
rect 36084 11086 36136 11092
rect 35992 10736 36044 10742
rect 35714 10704 35770 10713
rect 35992 10678 36044 10684
rect 35714 10639 35770 10648
rect 35624 10464 35676 10470
rect 35624 10406 35676 10412
rect 35438 10231 35494 10240
rect 35532 10260 35584 10266
rect 35532 10202 35584 10208
rect 35532 10124 35584 10130
rect 35532 10066 35584 10072
rect 35438 9888 35494 9897
rect 35438 9823 35494 9832
rect 35452 7256 35480 9823
rect 35544 9586 35572 10066
rect 35636 9722 35664 10406
rect 35624 9716 35676 9722
rect 35624 9658 35676 9664
rect 35728 9625 35756 10639
rect 35992 10600 36044 10606
rect 35992 10542 36044 10548
rect 35808 9648 35860 9654
rect 35714 9616 35770 9625
rect 35532 9580 35584 9586
rect 35808 9590 35860 9596
rect 35714 9551 35770 9560
rect 35532 9522 35584 9528
rect 35820 9178 35848 9590
rect 35900 9376 35952 9382
rect 35900 9318 35952 9324
rect 35808 9172 35860 9178
rect 35808 9114 35860 9120
rect 35624 9036 35676 9042
rect 35624 8978 35676 8984
rect 35532 7948 35584 7954
rect 35532 7890 35584 7896
rect 35544 7392 35572 7890
rect 35636 7750 35664 8978
rect 35820 8673 35848 9114
rect 35912 8974 35940 9318
rect 36004 9042 36032 10542
rect 36096 10266 36124 11086
rect 36268 10668 36320 10674
rect 36268 10610 36320 10616
rect 36084 10260 36136 10266
rect 36084 10202 36136 10208
rect 36280 9654 36308 10610
rect 36372 10470 36400 11222
rect 36360 10464 36412 10470
rect 36360 10406 36412 10412
rect 36372 10169 36400 10406
rect 36358 10160 36414 10169
rect 36358 10095 36414 10104
rect 36268 9648 36320 9654
rect 36268 9590 36320 9596
rect 36280 9450 36308 9590
rect 36268 9444 36320 9450
rect 36268 9386 36320 9392
rect 35992 9036 36044 9042
rect 35992 8978 36044 8984
rect 35900 8968 35952 8974
rect 35900 8910 35952 8916
rect 36268 8968 36320 8974
rect 36268 8910 36320 8916
rect 35900 8832 35952 8838
rect 35900 8774 35952 8780
rect 35806 8664 35862 8673
rect 35806 8599 35862 8608
rect 35806 8392 35862 8401
rect 35806 8327 35862 8336
rect 35624 7744 35676 7750
rect 35624 7686 35676 7692
rect 35544 7364 35664 7392
rect 35452 7228 35572 7256
rect 35438 7168 35494 7177
rect 35438 7103 35494 7112
rect 35452 5681 35480 7103
rect 35438 5672 35494 5681
rect 35438 5607 35494 5616
rect 35544 4826 35572 7228
rect 35636 6610 35664 7364
rect 35716 7268 35768 7274
rect 35716 7210 35768 7216
rect 35728 7002 35756 7210
rect 35716 6996 35768 7002
rect 35716 6938 35768 6944
rect 35820 6905 35848 8327
rect 35912 7041 35940 8774
rect 36280 8566 36308 8910
rect 36268 8560 36320 8566
rect 36266 8528 36268 8537
rect 36320 8528 36322 8537
rect 36266 8463 36322 8472
rect 36280 8090 36308 8463
rect 36268 8084 36320 8090
rect 36268 8026 36320 8032
rect 35992 8016 36044 8022
rect 35990 7984 35992 7993
rect 36044 7984 36046 7993
rect 36046 7942 36124 7970
rect 35990 7919 36046 7928
rect 35992 7880 36044 7886
rect 35992 7822 36044 7828
rect 36004 7546 36032 7822
rect 35992 7540 36044 7546
rect 35992 7482 36044 7488
rect 36096 7342 36124 7942
rect 36084 7336 36136 7342
rect 36084 7278 36136 7284
rect 35898 7032 35954 7041
rect 35898 6967 35954 6976
rect 35806 6896 35862 6905
rect 35806 6831 35862 6840
rect 35912 6644 35940 6967
rect 36082 6896 36138 6905
rect 36082 6831 36138 6840
rect 36268 6860 36320 6866
rect 35820 6616 35940 6644
rect 35636 6582 35756 6610
rect 35728 5778 35756 6582
rect 35716 5772 35768 5778
rect 35716 5714 35768 5720
rect 35532 4820 35584 4826
rect 35532 4762 35584 4768
rect 35438 4720 35494 4729
rect 35438 4655 35440 4664
rect 35492 4655 35494 4664
rect 35440 4626 35492 4632
rect 35452 4214 35480 4626
rect 35440 4208 35492 4214
rect 35440 4150 35492 4156
rect 35440 4072 35492 4078
rect 35440 4014 35492 4020
rect 35348 3936 35400 3942
rect 35348 3878 35400 3884
rect 35452 3777 35480 4014
rect 35438 3768 35494 3777
rect 35438 3703 35494 3712
rect 35820 921 35848 6616
rect 36096 5914 36124 6831
rect 36268 6802 36320 6808
rect 36280 6458 36308 6802
rect 36268 6452 36320 6458
rect 36268 6394 36320 6400
rect 36084 5908 36136 5914
rect 36084 5850 36136 5856
rect 35900 5772 35952 5778
rect 35900 5714 35952 5720
rect 35912 5030 35940 5714
rect 35900 5024 35952 5030
rect 35900 4966 35952 4972
rect 36372 4457 36400 10095
rect 36544 9648 36596 9654
rect 36544 9590 36596 9596
rect 36556 9081 36584 9590
rect 36542 9072 36598 9081
rect 36542 9007 36598 9016
rect 36452 7948 36504 7954
rect 36452 7890 36504 7896
rect 36464 6662 36492 7890
rect 36452 6656 36504 6662
rect 36452 6598 36504 6604
rect 36464 5953 36492 6598
rect 36450 5944 36506 5953
rect 36450 5879 36506 5888
rect 36648 5370 36676 13767
rect 37096 13320 37148 13326
rect 37096 13262 37148 13268
rect 37108 12986 37136 13262
rect 37096 12980 37148 12986
rect 37096 12922 37148 12928
rect 37280 12776 37332 12782
rect 37280 12718 37332 12724
rect 36820 11552 36872 11558
rect 36820 11494 36872 11500
rect 36832 9217 36860 11494
rect 37292 10674 37320 12718
rect 38764 12714 38792 15520
rect 38752 12708 38804 12714
rect 38752 12650 38804 12656
rect 37464 12640 37516 12646
rect 37464 12582 37516 12588
rect 37476 11937 37504 12582
rect 37462 11928 37518 11937
rect 37462 11863 37518 11872
rect 37554 11792 37610 11801
rect 37554 11727 37556 11736
rect 37608 11727 37610 11736
rect 37556 11698 37608 11704
rect 37280 10668 37332 10674
rect 37280 10610 37332 10616
rect 36912 10464 36964 10470
rect 36912 10406 36964 10412
rect 36818 9208 36874 9217
rect 36818 9143 36874 9152
rect 36924 8809 36952 10406
rect 37646 9616 37702 9625
rect 37646 9551 37702 9560
rect 37004 9376 37056 9382
rect 37004 9318 37056 9324
rect 37016 8838 37044 9318
rect 37370 9072 37426 9081
rect 37370 9007 37426 9016
rect 37004 8832 37056 8838
rect 36910 8800 36966 8809
rect 37004 8774 37056 8780
rect 36910 8735 36966 8744
rect 37278 8664 37334 8673
rect 37278 8599 37280 8608
rect 37332 8599 37334 8608
rect 37280 8570 37332 8576
rect 37384 8430 37412 9007
rect 37556 8560 37608 8566
rect 37556 8502 37608 8508
rect 37372 8424 37424 8430
rect 37372 8366 37424 8372
rect 37568 7993 37596 8502
rect 37554 7984 37610 7993
rect 37554 7919 37610 7928
rect 37660 6458 37688 9551
rect 37648 6452 37700 6458
rect 37648 6394 37700 6400
rect 37372 6248 37424 6254
rect 37372 6190 37424 6196
rect 36636 5364 36688 5370
rect 36636 5306 36688 5312
rect 36358 4448 36414 4457
rect 36358 4383 36414 4392
rect 37384 3913 37412 6190
rect 37370 3904 37426 3913
rect 37370 3839 37426 3848
rect 35806 912 35862 921
rect 35806 847 35862 856
rect 35162 232 35218 241
rect 35162 167 35218 176
<< via2 >>
rect 3606 15816 3662 15872
rect 3238 15408 3294 15464
rect 3146 14592 3202 14648
rect 3054 14184 3110 14240
rect 2778 13368 2834 13424
rect 1306 10920 1362 10976
rect 1582 8880 1638 8936
rect 2410 11620 2466 11656
rect 2410 11600 2412 11620
rect 2412 11600 2464 11620
rect 2464 11600 2466 11620
rect 2502 11464 2558 11520
rect 2502 9968 2558 10024
rect 2594 9832 2650 9888
rect 2870 10104 2926 10160
rect 2778 9696 2834 9752
rect 2686 9036 2742 9072
rect 2686 9016 2688 9036
rect 2688 9016 2740 9036
rect 2740 9016 2742 9036
rect 2410 8472 2466 8528
rect 2594 7520 2650 7576
rect 2318 4120 2374 4176
rect 2778 6976 2834 7032
rect 2042 4004 2098 4040
rect 2042 3984 2044 4004
rect 2044 3984 2096 4004
rect 2096 3984 2098 4004
rect 570 3712 626 3768
rect 1398 3596 1454 3632
rect 1398 3576 1400 3596
rect 1400 3576 1452 3596
rect 1452 3576 1454 3596
rect 3514 15000 3570 15056
rect 34518 15816 34574 15872
rect 3422 13776 3478 13832
rect 3422 12552 3478 12608
rect 4066 12980 4122 13016
rect 4066 12960 4068 12980
rect 4068 12960 4120 12980
rect 4120 12960 4122 12980
rect 3514 12144 3570 12200
rect 3882 11736 3938 11792
rect 3606 11076 3662 11112
rect 3606 11056 3608 11076
rect 3608 11056 3660 11076
rect 3660 11056 3662 11076
rect 4066 11328 4122 11384
rect 3882 10512 3938 10568
rect 3146 7148 3148 7168
rect 3148 7148 3200 7168
rect 3200 7148 3202 7168
rect 3146 7112 3202 7148
rect 3146 6840 3202 6896
rect 3238 6024 3294 6080
rect 3606 6704 3662 6760
rect 3330 5072 3386 5128
rect 3422 1264 3478 1320
rect 3238 856 3294 912
rect 2962 448 3018 504
rect 3974 9832 4030 9888
rect 4066 9288 4122 9344
rect 3882 8336 3938 8392
rect 3974 6976 4030 7032
rect 3974 5752 4030 5808
rect 4618 10004 4620 10024
rect 4620 10004 4672 10024
rect 4672 10004 4674 10024
rect 4618 9968 4674 10004
rect 4250 8200 4306 8256
rect 4342 8064 4398 8120
rect 4342 7692 4344 7712
rect 4344 7692 4396 7712
rect 4396 7692 4398 7712
rect 4342 7656 4398 7692
rect 4066 5364 4122 5400
rect 4066 5344 4068 5364
rect 4068 5344 4120 5364
rect 4120 5344 4122 5364
rect 3974 4936 4030 4992
rect 4066 4800 4122 4856
rect 3790 4528 3846 4584
rect 4710 4972 4712 4992
rect 4712 4972 4764 4992
rect 4764 4972 4766 4992
rect 4710 4936 4766 4972
rect 4526 4256 4582 4312
rect 5630 10784 5686 10840
rect 5630 10512 5686 10568
rect 5262 9152 5318 9208
rect 5354 8916 5356 8936
rect 5356 8916 5408 8936
rect 5408 8916 5410 8936
rect 5354 8880 5410 8916
rect 5538 8336 5594 8392
rect 5814 8472 5870 8528
rect 5446 7384 5502 7440
rect 4986 6568 5042 6624
rect 6826 11636 6828 11656
rect 6828 11636 6880 11656
rect 6880 11636 6882 11656
rect 6826 11600 6882 11636
rect 6182 8200 6238 8256
rect 6182 6060 6184 6080
rect 6184 6060 6236 6080
rect 6236 6060 6238 6080
rect 6182 6024 6238 6060
rect 7622 13082 7678 13084
rect 7702 13082 7758 13084
rect 7782 13082 7838 13084
rect 7862 13082 7918 13084
rect 7622 13030 7648 13082
rect 7648 13030 7678 13082
rect 7702 13030 7712 13082
rect 7712 13030 7758 13082
rect 7782 13030 7828 13082
rect 7828 13030 7838 13082
rect 7862 13030 7892 13082
rect 7892 13030 7918 13082
rect 7622 13028 7678 13030
rect 7702 13028 7758 13030
rect 7782 13028 7838 13030
rect 7862 13028 7918 13030
rect 6366 7248 6422 7304
rect 6274 5752 6330 5808
rect 5998 4528 6054 4584
rect 5906 3848 5962 3904
rect 4894 3032 4950 3088
rect 4802 2760 4858 2816
rect 4894 2080 4950 2136
rect 6642 9968 6698 10024
rect 7622 11994 7678 11996
rect 7702 11994 7758 11996
rect 7782 11994 7838 11996
rect 7862 11994 7918 11996
rect 7622 11942 7648 11994
rect 7648 11942 7678 11994
rect 7702 11942 7712 11994
rect 7712 11942 7758 11994
rect 7782 11942 7828 11994
rect 7828 11942 7838 11994
rect 7862 11942 7892 11994
rect 7892 11942 7918 11994
rect 7622 11940 7678 11942
rect 7702 11940 7758 11942
rect 7782 11940 7838 11942
rect 7862 11940 7918 11942
rect 8022 11872 8078 11928
rect 7562 11192 7618 11248
rect 7622 10906 7678 10908
rect 7702 10906 7758 10908
rect 7782 10906 7838 10908
rect 7862 10906 7918 10908
rect 7622 10854 7648 10906
rect 7648 10854 7678 10906
rect 7702 10854 7712 10906
rect 7712 10854 7758 10906
rect 7782 10854 7828 10906
rect 7828 10854 7838 10906
rect 7862 10854 7892 10906
rect 7892 10854 7918 10906
rect 7622 10852 7678 10854
rect 7702 10852 7758 10854
rect 7782 10852 7838 10854
rect 7862 10852 7918 10854
rect 8022 10240 8078 10296
rect 7622 9818 7678 9820
rect 7702 9818 7758 9820
rect 7782 9818 7838 9820
rect 7862 9818 7918 9820
rect 7622 9766 7648 9818
rect 7648 9766 7678 9818
rect 7702 9766 7712 9818
rect 7712 9766 7758 9818
rect 7782 9766 7828 9818
rect 7828 9766 7838 9818
rect 7862 9766 7892 9818
rect 7892 9766 7918 9818
rect 7622 9764 7678 9766
rect 7702 9764 7758 9766
rect 7782 9764 7838 9766
rect 7862 9764 7918 9766
rect 7286 9288 7342 9344
rect 7378 9052 7380 9072
rect 7380 9052 7432 9072
rect 7432 9052 7434 9072
rect 7378 9016 7434 9052
rect 8298 11600 8354 11656
rect 8114 9424 8170 9480
rect 8022 8744 8078 8800
rect 7622 8730 7678 8732
rect 7702 8730 7758 8732
rect 7782 8730 7838 8732
rect 7862 8730 7918 8732
rect 7622 8678 7648 8730
rect 7648 8678 7678 8730
rect 7702 8678 7712 8730
rect 7712 8678 7758 8730
rect 7782 8678 7828 8730
rect 7828 8678 7838 8730
rect 7862 8678 7892 8730
rect 7892 8678 7918 8730
rect 7622 8676 7678 8678
rect 7702 8676 7758 8678
rect 7782 8676 7838 8678
rect 7862 8676 7918 8678
rect 7286 8200 7342 8256
rect 7562 8200 7618 8256
rect 6734 7656 6790 7712
rect 6826 7520 6882 7576
rect 6550 7112 6606 7168
rect 7010 5364 7066 5400
rect 8390 9968 8446 10024
rect 7562 7792 7618 7848
rect 7622 7642 7678 7644
rect 7702 7642 7758 7644
rect 7782 7642 7838 7644
rect 7862 7642 7918 7644
rect 7622 7590 7648 7642
rect 7648 7590 7678 7642
rect 7702 7590 7712 7642
rect 7712 7590 7758 7642
rect 7782 7590 7828 7642
rect 7828 7590 7838 7642
rect 7862 7590 7892 7642
rect 7892 7590 7918 7642
rect 7622 7588 7678 7590
rect 7702 7588 7758 7590
rect 7782 7588 7838 7590
rect 7862 7588 7918 7590
rect 8206 7812 8262 7848
rect 8206 7792 8208 7812
rect 8208 7792 8260 7812
rect 8260 7792 8262 7812
rect 8574 9560 8630 9616
rect 9494 10684 9496 10704
rect 9496 10684 9548 10704
rect 9548 10684 9550 10704
rect 9494 10648 9550 10684
rect 9126 10376 9182 10432
rect 10690 11892 10746 11928
rect 10690 11872 10692 11892
rect 10692 11872 10744 11892
rect 10744 11872 10746 11892
rect 11610 11600 11666 11656
rect 10322 10260 10378 10296
rect 10322 10240 10324 10260
rect 10324 10240 10376 10260
rect 10376 10240 10378 10260
rect 10506 9716 10562 9752
rect 10506 9696 10508 9716
rect 10508 9696 10560 9716
rect 10560 9696 10562 9716
rect 8482 8608 8538 8664
rect 9678 9152 9734 9208
rect 10230 8628 10286 8664
rect 10230 8608 10232 8628
rect 10232 8608 10284 8628
rect 10284 8608 10286 8628
rect 8298 7520 8354 7576
rect 7286 6024 7342 6080
rect 9770 7384 9826 7440
rect 10138 7148 10140 7168
rect 10140 7148 10192 7168
rect 10192 7148 10194 7168
rect 7010 5344 7012 5364
rect 7012 5344 7064 5364
rect 7064 5344 7066 5364
rect 7562 6704 7618 6760
rect 7622 6554 7678 6556
rect 7702 6554 7758 6556
rect 7782 6554 7838 6556
rect 7862 6554 7918 6556
rect 7622 6502 7648 6554
rect 7648 6502 7678 6554
rect 7702 6502 7712 6554
rect 7712 6502 7758 6554
rect 7782 6502 7828 6554
rect 7828 6502 7838 6554
rect 7862 6502 7892 6554
rect 7892 6502 7918 6554
rect 7622 6500 7678 6502
rect 7702 6500 7758 6502
rect 7782 6500 7838 6502
rect 7862 6500 7918 6502
rect 9678 6840 9734 6896
rect 7654 5908 7710 5944
rect 7654 5888 7656 5908
rect 7656 5888 7708 5908
rect 7708 5888 7710 5908
rect 7622 5466 7678 5468
rect 7702 5466 7758 5468
rect 7782 5466 7838 5468
rect 7862 5466 7918 5468
rect 7622 5414 7648 5466
rect 7648 5414 7678 5466
rect 7702 5414 7712 5466
rect 7712 5414 7758 5466
rect 7782 5414 7828 5466
rect 7828 5414 7838 5466
rect 7862 5414 7892 5466
rect 7892 5414 7918 5466
rect 7622 5412 7678 5414
rect 7702 5412 7758 5414
rect 7782 5412 7838 5414
rect 7862 5412 7918 5414
rect 8022 5344 8078 5400
rect 9678 6196 9680 6216
rect 9680 6196 9732 6216
rect 9732 6196 9734 6216
rect 9678 6160 9734 6196
rect 8206 5752 8262 5808
rect 8114 4936 8170 4992
rect 8298 5480 8354 5536
rect 6458 3984 6514 4040
rect 7622 4378 7678 4380
rect 7702 4378 7758 4380
rect 7782 4378 7838 4380
rect 7862 4378 7918 4380
rect 7622 4326 7648 4378
rect 7648 4326 7678 4378
rect 7702 4326 7712 4378
rect 7712 4326 7758 4378
rect 7782 4326 7828 4378
rect 7828 4326 7838 4378
rect 7862 4326 7892 4378
rect 7892 4326 7918 4378
rect 7622 4324 7678 4326
rect 7702 4324 7758 4326
rect 7782 4324 7838 4326
rect 7862 4324 7918 4326
rect 9954 5752 10010 5808
rect 10138 7112 10194 7148
rect 10046 5616 10102 5672
rect 10322 5480 10378 5536
rect 10046 5072 10102 5128
rect 10506 6704 10562 6760
rect 10598 6160 10654 6216
rect 10506 5908 10562 5944
rect 10506 5888 10508 5908
rect 10508 5888 10560 5908
rect 10560 5888 10562 5908
rect 10414 4800 10470 4856
rect 9310 4120 9366 4176
rect 10782 11056 10838 11112
rect 11150 10376 11206 10432
rect 11702 11092 11704 11112
rect 11704 11092 11756 11112
rect 11756 11092 11758 11112
rect 11702 11056 11758 11092
rect 11610 9968 11666 10024
rect 10874 8880 10930 8936
rect 11334 8880 11390 8936
rect 14289 13626 14345 13628
rect 14369 13626 14425 13628
rect 14449 13626 14505 13628
rect 14529 13626 14585 13628
rect 14289 13574 14315 13626
rect 14315 13574 14345 13626
rect 14369 13574 14379 13626
rect 14379 13574 14425 13626
rect 14449 13574 14495 13626
rect 14495 13574 14505 13626
rect 14529 13574 14559 13626
rect 14559 13574 14585 13626
rect 14289 13572 14345 13574
rect 14369 13572 14425 13574
rect 14449 13572 14505 13574
rect 14529 13572 14585 13574
rect 11702 8608 11758 8664
rect 11334 7656 11390 7712
rect 10874 5344 10930 5400
rect 10874 4936 10930 4992
rect 11058 6876 11060 6896
rect 11060 6876 11112 6896
rect 11112 6876 11114 6896
rect 11058 6840 11114 6876
rect 10966 4800 11022 4856
rect 7622 3290 7678 3292
rect 7702 3290 7758 3292
rect 7782 3290 7838 3292
rect 7862 3290 7918 3292
rect 7622 3238 7648 3290
rect 7648 3238 7678 3290
rect 7702 3238 7712 3290
rect 7712 3238 7758 3290
rect 7782 3238 7828 3290
rect 7828 3238 7838 3290
rect 7862 3238 7892 3290
rect 7892 3238 7918 3290
rect 7622 3236 7678 3238
rect 7702 3236 7758 3238
rect 7782 3236 7838 3238
rect 7862 3236 7918 3238
rect 11150 4392 11206 4448
rect 11058 3984 11114 4040
rect 10598 3576 10654 3632
rect 12622 9424 12678 9480
rect 12162 7520 12218 7576
rect 12806 6568 12862 6624
rect 11426 4256 11482 4312
rect 11702 3612 11704 3632
rect 11704 3612 11756 3632
rect 11756 3612 11758 3632
rect 11702 3576 11758 3612
rect 12070 4664 12126 4720
rect 12530 6296 12586 6352
rect 12806 4800 12862 4856
rect 12530 4120 12586 4176
rect 12162 3884 12164 3904
rect 12164 3884 12216 3904
rect 12216 3884 12218 3904
rect 12162 3848 12218 3884
rect 11978 3440 12034 3496
rect 7470 2896 7526 2952
rect 12346 3032 12402 3088
rect 11610 2760 11666 2816
rect 6366 2488 6422 2544
rect 7622 2202 7678 2204
rect 7702 2202 7758 2204
rect 7782 2202 7838 2204
rect 7862 2202 7918 2204
rect 7622 2150 7648 2202
rect 7648 2150 7678 2202
rect 7702 2150 7712 2202
rect 7712 2150 7758 2202
rect 7782 2150 7828 2202
rect 7828 2150 7838 2202
rect 7862 2150 7892 2202
rect 7892 2150 7918 2202
rect 7622 2148 7678 2150
rect 7702 2148 7758 2150
rect 7782 2148 7838 2150
rect 7862 2148 7918 2150
rect 14289 12538 14345 12540
rect 14369 12538 14425 12540
rect 14449 12538 14505 12540
rect 14529 12538 14585 12540
rect 14289 12486 14315 12538
rect 14315 12486 14345 12538
rect 14369 12486 14379 12538
rect 14379 12486 14425 12538
rect 14449 12486 14495 12538
rect 14495 12486 14505 12538
rect 14529 12486 14559 12538
rect 14559 12486 14585 12538
rect 14289 12484 14345 12486
rect 14369 12484 14425 12486
rect 14449 12484 14505 12486
rect 14529 12484 14585 12486
rect 12990 9560 13046 9616
rect 14289 11450 14345 11452
rect 14369 11450 14425 11452
rect 14449 11450 14505 11452
rect 14529 11450 14585 11452
rect 14289 11398 14315 11450
rect 14315 11398 14345 11450
rect 14369 11398 14379 11450
rect 14379 11398 14425 11450
rect 14449 11398 14495 11450
rect 14495 11398 14505 11450
rect 14529 11398 14559 11450
rect 14559 11398 14585 11450
rect 14289 11396 14345 11398
rect 14369 11396 14425 11398
rect 14449 11396 14505 11398
rect 14529 11396 14585 11398
rect 15106 11192 15162 11248
rect 15750 11192 15806 11248
rect 13910 11056 13966 11112
rect 13266 9016 13322 9072
rect 13634 9424 13690 9480
rect 13358 7520 13414 7576
rect 13726 7948 13782 7984
rect 13726 7928 13728 7948
rect 13728 7928 13780 7948
rect 13780 7928 13782 7948
rect 13542 6296 13598 6352
rect 13450 5480 13506 5536
rect 13174 5344 13230 5400
rect 13174 5072 13230 5128
rect 12990 3576 13046 3632
rect 13818 6860 13874 6896
rect 13818 6840 13820 6860
rect 13820 6840 13872 6860
rect 13872 6840 13874 6860
rect 16486 11328 16542 11384
rect 14289 10362 14345 10364
rect 14369 10362 14425 10364
rect 14449 10362 14505 10364
rect 14529 10362 14585 10364
rect 14289 10310 14315 10362
rect 14315 10310 14345 10362
rect 14369 10310 14379 10362
rect 14379 10310 14425 10362
rect 14449 10310 14495 10362
rect 14495 10310 14505 10362
rect 14529 10310 14559 10362
rect 14559 10310 14585 10362
rect 14289 10308 14345 10310
rect 14369 10308 14425 10310
rect 14449 10308 14505 10310
rect 14529 10308 14585 10310
rect 15290 9716 15346 9752
rect 15290 9696 15292 9716
rect 15292 9696 15344 9716
rect 15344 9696 15346 9716
rect 14186 9560 14242 9616
rect 14094 8200 14150 8256
rect 14094 8064 14150 8120
rect 14289 9274 14345 9276
rect 14369 9274 14425 9276
rect 14449 9274 14505 9276
rect 14529 9274 14585 9276
rect 14289 9222 14315 9274
rect 14315 9222 14345 9274
rect 14369 9222 14379 9274
rect 14379 9222 14425 9274
rect 14449 9222 14495 9274
rect 14495 9222 14505 9274
rect 14529 9222 14559 9274
rect 14559 9222 14585 9274
rect 14289 9220 14345 9222
rect 14369 9220 14425 9222
rect 14449 9220 14505 9222
rect 14529 9220 14585 9222
rect 15382 9016 15438 9072
rect 15290 8356 15346 8392
rect 15290 8336 15292 8356
rect 15292 8336 15344 8356
rect 15344 8336 15346 8356
rect 14289 8186 14345 8188
rect 14369 8186 14425 8188
rect 14449 8186 14505 8188
rect 14529 8186 14585 8188
rect 14289 8134 14315 8186
rect 14315 8134 14345 8186
rect 14369 8134 14379 8186
rect 14379 8134 14425 8186
rect 14449 8134 14495 8186
rect 14495 8134 14505 8186
rect 14529 8134 14559 8186
rect 14559 8134 14585 8186
rect 14289 8132 14345 8134
rect 14369 8132 14425 8134
rect 14449 8132 14505 8134
rect 14529 8132 14585 8134
rect 17130 11600 17186 11656
rect 16026 9696 16082 9752
rect 16946 8880 17002 8936
rect 15750 8508 15752 8528
rect 15752 8508 15804 8528
rect 15804 8508 15806 8528
rect 15750 8472 15806 8508
rect 16210 8064 16266 8120
rect 15658 7928 15714 7984
rect 14738 7404 14794 7440
rect 14738 7384 14740 7404
rect 14740 7384 14792 7404
rect 14792 7384 14794 7404
rect 14738 7148 14740 7168
rect 14740 7148 14792 7168
rect 14792 7148 14794 7168
rect 14738 7112 14794 7148
rect 14289 7098 14345 7100
rect 14369 7098 14425 7100
rect 14449 7098 14505 7100
rect 14529 7098 14585 7100
rect 14289 7046 14315 7098
rect 14315 7046 14345 7098
rect 14369 7046 14379 7098
rect 14379 7046 14425 7098
rect 14449 7046 14495 7098
rect 14495 7046 14505 7098
rect 14529 7046 14559 7098
rect 14559 7046 14585 7098
rect 14289 7044 14345 7046
rect 14369 7044 14425 7046
rect 14449 7044 14505 7046
rect 14529 7044 14585 7046
rect 14094 6976 14150 7032
rect 16210 6840 16266 6896
rect 14289 6010 14345 6012
rect 14369 6010 14425 6012
rect 14449 6010 14505 6012
rect 14529 6010 14585 6012
rect 14289 5958 14315 6010
rect 14315 5958 14345 6010
rect 14369 5958 14379 6010
rect 14379 5958 14425 6010
rect 14449 5958 14495 6010
rect 14495 5958 14505 6010
rect 14529 5958 14559 6010
rect 14559 5958 14585 6010
rect 14289 5956 14345 5958
rect 14369 5956 14425 5958
rect 14449 5956 14505 5958
rect 14529 5956 14585 5958
rect 14289 4922 14345 4924
rect 14369 4922 14425 4924
rect 14449 4922 14505 4924
rect 14529 4922 14585 4924
rect 14289 4870 14315 4922
rect 14315 4870 14345 4922
rect 14369 4870 14379 4922
rect 14379 4870 14425 4922
rect 14449 4870 14495 4922
rect 14495 4870 14505 4922
rect 14529 4870 14559 4922
rect 14559 4870 14585 4922
rect 14289 4868 14345 4870
rect 14369 4868 14425 4870
rect 14449 4868 14505 4870
rect 14529 4868 14585 4870
rect 16302 6568 16358 6624
rect 20956 13082 21012 13084
rect 21036 13082 21092 13084
rect 21116 13082 21172 13084
rect 21196 13082 21252 13084
rect 20956 13030 20982 13082
rect 20982 13030 21012 13082
rect 21036 13030 21046 13082
rect 21046 13030 21092 13082
rect 21116 13030 21162 13082
rect 21162 13030 21172 13082
rect 21196 13030 21226 13082
rect 21226 13030 21252 13082
rect 20956 13028 21012 13030
rect 21036 13028 21092 13030
rect 21116 13028 21172 13030
rect 21196 13028 21252 13030
rect 19062 11464 19118 11520
rect 18878 11328 18934 11384
rect 17590 9560 17646 9616
rect 16946 7112 17002 7168
rect 16578 5888 16634 5944
rect 16578 5616 16634 5672
rect 16854 5516 16856 5536
rect 16856 5516 16908 5536
rect 16908 5516 16910 5536
rect 16854 5480 16910 5516
rect 16210 5208 16266 5264
rect 16578 5228 16634 5264
rect 16578 5208 16580 5228
rect 16580 5208 16632 5228
rect 16632 5208 16634 5228
rect 15658 4936 15714 4992
rect 14738 4664 14794 4720
rect 14646 4004 14702 4040
rect 14646 3984 14648 4004
rect 14648 3984 14700 4004
rect 14700 3984 14702 4004
rect 14289 3834 14345 3836
rect 14369 3834 14425 3836
rect 14449 3834 14505 3836
rect 14529 3834 14585 3836
rect 14289 3782 14315 3834
rect 14315 3782 14345 3834
rect 14369 3782 14379 3834
rect 14379 3782 14425 3834
rect 14449 3782 14495 3834
rect 14495 3782 14505 3834
rect 14529 3782 14559 3834
rect 14559 3782 14585 3834
rect 14289 3780 14345 3782
rect 14369 3780 14425 3782
rect 14449 3780 14505 3782
rect 14529 3780 14585 3782
rect 15750 4256 15806 4312
rect 18050 9424 18106 9480
rect 17590 8336 17646 8392
rect 17314 6432 17370 6488
rect 17314 5616 17370 5672
rect 18234 8336 18290 8392
rect 19062 10648 19118 10704
rect 19982 11736 20038 11792
rect 19890 9288 19946 9344
rect 18418 8608 18474 8664
rect 18602 8200 18658 8256
rect 18326 7656 18382 7712
rect 18602 7520 18658 7576
rect 19522 8084 19578 8120
rect 19522 8064 19524 8084
rect 19524 8064 19576 8084
rect 19576 8064 19578 8084
rect 19246 7692 19248 7712
rect 19248 7692 19300 7712
rect 19300 7692 19302 7712
rect 19246 7656 19302 7692
rect 19338 7112 19394 7168
rect 19062 6976 19118 7032
rect 18050 5092 18106 5128
rect 18050 5072 18052 5092
rect 18052 5072 18104 5092
rect 18104 5072 18106 5092
rect 17130 4700 17132 4720
rect 17132 4700 17184 4720
rect 17184 4700 17186 4720
rect 17130 4664 17186 4700
rect 18786 5888 18842 5944
rect 18970 6196 18972 6216
rect 18972 6196 19024 6216
rect 19024 6196 19026 6216
rect 18970 6160 19026 6196
rect 18970 5616 19026 5672
rect 20534 9152 20590 9208
rect 20166 7656 20222 7712
rect 19798 7112 19854 7168
rect 20956 11994 21012 11996
rect 21036 11994 21092 11996
rect 21116 11994 21172 11996
rect 21196 11994 21252 11996
rect 20956 11942 20982 11994
rect 20982 11942 21012 11994
rect 21036 11942 21046 11994
rect 21046 11942 21092 11994
rect 21116 11942 21162 11994
rect 21162 11942 21172 11994
rect 21196 11942 21226 11994
rect 21226 11942 21252 11994
rect 20956 11940 21012 11942
rect 21036 11940 21092 11942
rect 21116 11940 21172 11942
rect 21196 11940 21252 11942
rect 20810 11500 20812 11520
rect 20812 11500 20864 11520
rect 20864 11500 20866 11520
rect 20810 11464 20866 11500
rect 20956 10906 21012 10908
rect 21036 10906 21092 10908
rect 21116 10906 21172 10908
rect 21196 10906 21252 10908
rect 20956 10854 20982 10906
rect 20982 10854 21012 10906
rect 21036 10854 21046 10906
rect 21046 10854 21092 10906
rect 21116 10854 21162 10906
rect 21162 10854 21172 10906
rect 21196 10854 21226 10906
rect 21226 10854 21252 10906
rect 20956 10852 21012 10854
rect 21036 10852 21092 10854
rect 21116 10852 21172 10854
rect 21196 10852 21252 10854
rect 20810 9832 20866 9888
rect 20956 9818 21012 9820
rect 21036 9818 21092 9820
rect 21116 9818 21172 9820
rect 21196 9818 21252 9820
rect 20956 9766 20982 9818
rect 20982 9766 21012 9818
rect 21036 9766 21046 9818
rect 21046 9766 21092 9818
rect 21116 9766 21162 9818
rect 21162 9766 21172 9818
rect 21196 9766 21226 9818
rect 21226 9766 21252 9818
rect 20956 9764 21012 9766
rect 21036 9764 21092 9766
rect 21116 9764 21172 9766
rect 21196 9764 21252 9766
rect 21638 11228 21640 11248
rect 21640 11228 21692 11248
rect 21692 11228 21694 11248
rect 21638 11192 21694 11228
rect 20810 9016 20866 9072
rect 21362 9016 21418 9072
rect 20956 8730 21012 8732
rect 21036 8730 21092 8732
rect 21116 8730 21172 8732
rect 21196 8730 21252 8732
rect 20956 8678 20982 8730
rect 20982 8678 21012 8730
rect 21036 8678 21046 8730
rect 21046 8678 21092 8730
rect 21116 8678 21162 8730
rect 21162 8678 21172 8730
rect 21196 8678 21226 8730
rect 21226 8678 21252 8730
rect 20956 8676 21012 8678
rect 21036 8676 21092 8678
rect 21116 8676 21172 8678
rect 21196 8676 21252 8678
rect 20810 7656 20866 7712
rect 20956 7642 21012 7644
rect 21036 7642 21092 7644
rect 21116 7642 21172 7644
rect 21196 7642 21252 7644
rect 20956 7590 20982 7642
rect 20982 7590 21012 7642
rect 21036 7590 21046 7642
rect 21046 7590 21092 7642
rect 21116 7590 21162 7642
rect 21162 7590 21172 7642
rect 21196 7590 21226 7642
rect 21226 7590 21252 7642
rect 20956 7588 21012 7590
rect 21036 7588 21092 7590
rect 21116 7588 21172 7590
rect 21196 7588 21252 7590
rect 20810 7520 20866 7576
rect 19522 5908 19578 5944
rect 19522 5888 19524 5908
rect 19524 5888 19576 5908
rect 19576 5888 19578 5908
rect 19430 5208 19486 5264
rect 17222 4528 17278 4584
rect 16946 2896 17002 2952
rect 14289 2746 14345 2748
rect 14369 2746 14425 2748
rect 14449 2746 14505 2748
rect 14529 2746 14585 2748
rect 14289 2694 14315 2746
rect 14315 2694 14345 2746
rect 14369 2694 14379 2746
rect 14379 2694 14425 2746
rect 14449 2694 14495 2746
rect 14495 2694 14505 2746
rect 14529 2694 14559 2746
rect 14559 2694 14585 2746
rect 14289 2692 14345 2694
rect 14369 2692 14425 2694
rect 14449 2692 14505 2694
rect 14529 2692 14585 2694
rect 12530 1808 12586 1864
rect 5906 1672 5962 1728
rect 17406 1672 17462 1728
rect 20956 6554 21012 6556
rect 21036 6554 21092 6556
rect 21116 6554 21172 6556
rect 21196 6554 21252 6556
rect 20956 6502 20982 6554
rect 20982 6502 21012 6554
rect 21036 6502 21046 6554
rect 21046 6502 21092 6554
rect 21116 6502 21162 6554
rect 21162 6502 21172 6554
rect 21196 6502 21226 6554
rect 21226 6502 21252 6554
rect 20956 6500 21012 6502
rect 21036 6500 21092 6502
rect 21116 6500 21172 6502
rect 21196 6500 21252 6502
rect 21822 11056 21878 11112
rect 21822 9424 21878 9480
rect 22282 10648 22338 10704
rect 22006 10240 22062 10296
rect 22374 9324 22376 9344
rect 22376 9324 22428 9344
rect 22428 9324 22430 9344
rect 22374 9288 22430 9324
rect 21822 8336 21878 8392
rect 21822 8200 21878 8256
rect 21822 7792 21878 7848
rect 21730 5888 21786 5944
rect 20956 5466 21012 5468
rect 21036 5466 21092 5468
rect 21116 5466 21172 5468
rect 21196 5466 21252 5468
rect 20956 5414 20982 5466
rect 20982 5414 21012 5466
rect 21036 5414 21046 5466
rect 21046 5414 21092 5466
rect 21116 5414 21162 5466
rect 21162 5414 21172 5466
rect 21196 5414 21226 5466
rect 21226 5414 21252 5466
rect 20956 5412 21012 5414
rect 21036 5412 21092 5414
rect 21116 5412 21172 5414
rect 21196 5412 21252 5414
rect 20810 5344 20866 5400
rect 20534 5072 20590 5128
rect 20956 4378 21012 4380
rect 21036 4378 21092 4380
rect 21116 4378 21172 4380
rect 21196 4378 21252 4380
rect 20956 4326 20982 4378
rect 20982 4326 21012 4378
rect 21036 4326 21046 4378
rect 21046 4326 21092 4378
rect 21116 4326 21162 4378
rect 21162 4326 21172 4378
rect 21196 4326 21226 4378
rect 21226 4326 21252 4378
rect 20956 4324 21012 4326
rect 21036 4324 21092 4326
rect 21116 4324 21172 4326
rect 21196 4324 21252 4326
rect 23018 10920 23074 10976
rect 23754 11056 23810 11112
rect 27622 13626 27678 13628
rect 27702 13626 27758 13628
rect 27782 13626 27838 13628
rect 27862 13626 27918 13628
rect 27622 13574 27648 13626
rect 27648 13574 27678 13626
rect 27702 13574 27712 13626
rect 27712 13574 27758 13626
rect 27782 13574 27828 13626
rect 27828 13574 27838 13626
rect 27862 13574 27892 13626
rect 27892 13574 27918 13626
rect 27622 13572 27678 13574
rect 27702 13572 27758 13574
rect 27782 13572 27838 13574
rect 27862 13572 27918 13574
rect 24766 12552 24822 12608
rect 24674 11192 24730 11248
rect 24306 11056 24362 11112
rect 24030 10668 24086 10704
rect 24030 10648 24032 10668
rect 24032 10648 24084 10668
rect 24084 10648 24086 10668
rect 23938 9288 23994 9344
rect 23478 6024 23534 6080
rect 24766 10784 24822 10840
rect 25042 12008 25098 12064
rect 25042 11600 25098 11656
rect 25134 11464 25190 11520
rect 25594 11872 25650 11928
rect 25594 11464 25650 11520
rect 25042 10956 25044 10976
rect 25044 10956 25096 10976
rect 25096 10956 25098 10976
rect 25042 10920 25098 10956
rect 25226 10920 25282 10976
rect 25134 10512 25190 10568
rect 24030 9152 24086 9208
rect 24490 6840 24546 6896
rect 24030 6724 24086 6760
rect 24030 6704 24032 6724
rect 24032 6704 24084 6724
rect 24084 6704 24086 6724
rect 23110 5616 23166 5672
rect 24674 6160 24730 6216
rect 24214 5888 24270 5944
rect 24122 5344 24178 5400
rect 25318 10004 25320 10024
rect 25320 10004 25372 10024
rect 25372 10004 25374 10024
rect 25318 9968 25374 10004
rect 25502 7948 25558 7984
rect 25502 7928 25504 7948
rect 25504 7928 25556 7948
rect 25556 7928 25558 7948
rect 27622 12538 27678 12540
rect 27702 12538 27758 12540
rect 27782 12538 27838 12540
rect 27862 12538 27918 12540
rect 27622 12486 27648 12538
rect 27648 12486 27678 12538
rect 27702 12486 27712 12538
rect 27712 12486 27758 12538
rect 27782 12486 27828 12538
rect 27828 12486 27838 12538
rect 27862 12486 27892 12538
rect 27892 12486 27918 12538
rect 27622 12484 27678 12486
rect 27702 12484 27758 12486
rect 27782 12484 27838 12486
rect 27862 12484 27918 12486
rect 29550 12280 29606 12336
rect 27250 12144 27306 12200
rect 26238 11212 26294 11248
rect 26238 11192 26240 11212
rect 26240 11192 26292 11212
rect 26292 11192 26294 11212
rect 29366 11736 29422 11792
rect 29918 11636 29920 11656
rect 29920 11636 29972 11656
rect 29972 11636 29974 11656
rect 29918 11600 29974 11636
rect 26606 11076 26662 11112
rect 26606 11056 26608 11076
rect 26608 11056 26660 11076
rect 26660 11056 26662 11076
rect 27342 10648 27398 10704
rect 26146 9968 26202 10024
rect 26882 9560 26938 9616
rect 26514 9424 26570 9480
rect 25962 8608 26018 8664
rect 27622 11450 27678 11452
rect 27702 11450 27758 11452
rect 27782 11450 27838 11452
rect 27862 11450 27918 11452
rect 27622 11398 27648 11450
rect 27648 11398 27678 11450
rect 27702 11398 27712 11450
rect 27712 11398 27758 11450
rect 27782 11398 27828 11450
rect 27828 11398 27838 11450
rect 27862 11398 27892 11450
rect 27892 11398 27918 11450
rect 27622 11396 27678 11398
rect 27702 11396 27758 11398
rect 27782 11396 27838 11398
rect 27862 11396 27918 11398
rect 27802 10804 27858 10840
rect 27802 10784 27804 10804
rect 27804 10784 27856 10804
rect 27856 10784 27858 10804
rect 27622 10362 27678 10364
rect 27702 10362 27758 10364
rect 27782 10362 27838 10364
rect 27862 10362 27918 10364
rect 27622 10310 27648 10362
rect 27648 10310 27678 10362
rect 27702 10310 27712 10362
rect 27712 10310 27758 10362
rect 27782 10310 27828 10362
rect 27828 10310 27838 10362
rect 27862 10310 27892 10362
rect 27892 10310 27918 10362
rect 27622 10308 27678 10310
rect 27702 10308 27758 10310
rect 27782 10308 27838 10310
rect 27862 10308 27918 10310
rect 26974 9052 26976 9072
rect 26976 9052 27028 9072
rect 27028 9052 27030 9072
rect 26974 9016 27030 9052
rect 27434 9424 27490 9480
rect 27622 9274 27678 9276
rect 27702 9274 27758 9276
rect 27782 9274 27838 9276
rect 27862 9274 27918 9276
rect 27622 9222 27648 9274
rect 27648 9222 27678 9274
rect 27702 9222 27712 9274
rect 27712 9222 27758 9274
rect 27782 9222 27828 9274
rect 27828 9222 27838 9274
rect 27862 9222 27892 9274
rect 27892 9222 27918 9274
rect 27622 9220 27678 9222
rect 27702 9220 27758 9222
rect 27782 9220 27838 9222
rect 27862 9220 27918 9222
rect 27622 8186 27678 8188
rect 27702 8186 27758 8188
rect 27782 8186 27838 8188
rect 27862 8186 27918 8188
rect 27622 8134 27648 8186
rect 27648 8134 27678 8186
rect 27702 8134 27712 8186
rect 27712 8134 27758 8186
rect 27782 8134 27828 8186
rect 27828 8134 27838 8186
rect 27862 8134 27892 8186
rect 27892 8134 27918 8186
rect 27622 8132 27678 8134
rect 27702 8132 27758 8134
rect 27782 8132 27838 8134
rect 27862 8132 27918 8134
rect 27434 8064 27490 8120
rect 26330 7792 26386 7848
rect 27066 7792 27122 7848
rect 26054 7248 26110 7304
rect 25686 7112 25742 7168
rect 27066 6976 27122 7032
rect 25778 6704 25834 6760
rect 26422 6452 26478 6488
rect 26422 6432 26424 6452
rect 26424 6432 26476 6452
rect 26476 6432 26478 6452
rect 27342 6704 27398 6760
rect 27342 5752 27398 5808
rect 27158 5516 27160 5536
rect 27160 5516 27212 5536
rect 27212 5516 27214 5536
rect 27158 5480 27214 5516
rect 25594 4936 25650 4992
rect 24950 4528 25006 4584
rect 24122 4392 24178 4448
rect 28170 8200 28226 8256
rect 28170 7792 28226 7848
rect 27526 7248 27582 7304
rect 27622 7098 27678 7100
rect 27702 7098 27758 7100
rect 27782 7098 27838 7100
rect 27862 7098 27918 7100
rect 27622 7046 27648 7098
rect 27648 7046 27678 7098
rect 27702 7046 27712 7098
rect 27712 7046 27758 7098
rect 27782 7046 27828 7098
rect 27828 7046 27838 7098
rect 27862 7046 27892 7098
rect 27892 7046 27918 7098
rect 27622 7044 27678 7046
rect 27702 7044 27758 7046
rect 27782 7044 27838 7046
rect 27862 7044 27918 7046
rect 27622 6010 27678 6012
rect 27702 6010 27758 6012
rect 27782 6010 27838 6012
rect 27862 6010 27918 6012
rect 27622 5958 27648 6010
rect 27648 5958 27678 6010
rect 27702 5958 27712 6010
rect 27712 5958 27758 6010
rect 27782 5958 27828 6010
rect 27828 5958 27838 6010
rect 27862 5958 27892 6010
rect 27892 5958 27918 6010
rect 27622 5956 27678 5958
rect 27702 5956 27758 5958
rect 27782 5956 27838 5958
rect 27862 5956 27918 5958
rect 27622 4922 27678 4924
rect 27702 4922 27758 4924
rect 27782 4922 27838 4924
rect 27862 4922 27918 4924
rect 27622 4870 27648 4922
rect 27648 4870 27678 4922
rect 27702 4870 27712 4922
rect 27712 4870 27758 4922
rect 27782 4870 27828 4922
rect 27828 4870 27838 4922
rect 27862 4870 27892 4922
rect 27892 4870 27918 4922
rect 27622 4868 27678 4870
rect 27702 4868 27758 4870
rect 27782 4868 27838 4870
rect 27862 4868 27918 4870
rect 27526 4020 27528 4040
rect 27528 4020 27580 4040
rect 27580 4020 27582 4040
rect 27526 3984 27582 4020
rect 29550 10648 29606 10704
rect 30930 11328 30986 11384
rect 28262 7520 28318 7576
rect 28630 9152 28686 9208
rect 28446 7520 28502 7576
rect 29826 9596 29828 9616
rect 29828 9596 29880 9616
rect 29880 9596 29882 9616
rect 29826 9560 29882 9596
rect 29090 7656 29146 7712
rect 30010 7384 30066 7440
rect 29826 7112 29882 7168
rect 28906 6568 28962 6624
rect 28906 6296 28962 6352
rect 29826 6296 29882 6352
rect 28446 5616 28502 5672
rect 28630 5616 28686 5672
rect 29182 5616 29238 5672
rect 28630 5344 28686 5400
rect 28814 5208 28870 5264
rect 29366 5616 29422 5672
rect 29550 5208 29606 5264
rect 29274 5072 29330 5128
rect 28354 4936 28410 4992
rect 27622 3834 27678 3836
rect 27702 3834 27758 3836
rect 27782 3834 27838 3836
rect 27862 3834 27918 3836
rect 27622 3782 27648 3834
rect 27648 3782 27678 3834
rect 27702 3782 27712 3834
rect 27712 3782 27758 3834
rect 27782 3782 27828 3834
rect 27828 3782 27838 3834
rect 27862 3782 27892 3834
rect 27892 3782 27918 3834
rect 27622 3780 27678 3782
rect 27702 3780 27758 3782
rect 27782 3780 27838 3782
rect 27862 3780 27918 3782
rect 20956 3290 21012 3292
rect 21036 3290 21092 3292
rect 21116 3290 21172 3292
rect 21196 3290 21252 3292
rect 20956 3238 20982 3290
rect 20982 3238 21012 3290
rect 21036 3238 21046 3290
rect 21046 3238 21092 3290
rect 21116 3238 21162 3290
rect 21162 3238 21172 3290
rect 21196 3238 21226 3290
rect 21226 3238 21252 3290
rect 20956 3236 21012 3238
rect 21036 3236 21092 3238
rect 21116 3236 21172 3238
rect 21196 3236 21252 3238
rect 27622 2746 27678 2748
rect 27702 2746 27758 2748
rect 27782 2746 27838 2748
rect 27862 2746 27918 2748
rect 27622 2694 27648 2746
rect 27648 2694 27678 2746
rect 27702 2694 27712 2746
rect 27712 2694 27758 2746
rect 27782 2694 27828 2746
rect 27828 2694 27838 2746
rect 27862 2694 27892 2746
rect 27892 2694 27918 2746
rect 27622 2692 27678 2694
rect 27702 2692 27758 2694
rect 27782 2692 27838 2694
rect 27862 2692 27918 2694
rect 30838 9036 30894 9072
rect 30838 9016 30840 9036
rect 30840 9016 30892 9036
rect 30892 9016 30894 9036
rect 30746 8880 30802 8936
rect 30378 8472 30434 8528
rect 30654 8372 30656 8392
rect 30656 8372 30708 8392
rect 30708 8372 30710 8392
rect 30654 8336 30710 8372
rect 30470 8200 30526 8256
rect 31942 11892 31998 11928
rect 31942 11872 31944 11892
rect 31944 11872 31996 11892
rect 31996 11872 31998 11892
rect 30746 7384 30802 7440
rect 31482 8492 31538 8528
rect 31482 8472 31484 8492
rect 31484 8472 31536 8492
rect 31536 8472 31538 8492
rect 31390 6840 31446 6896
rect 31298 6432 31354 6488
rect 32310 11500 32312 11520
rect 32312 11500 32364 11520
rect 32364 11500 32366 11520
rect 32310 11464 32366 11500
rect 33138 12008 33194 12064
rect 32954 10512 33010 10568
rect 32678 9016 32734 9072
rect 32494 8608 32550 8664
rect 32770 8508 32772 8528
rect 32772 8508 32824 8528
rect 32824 8508 32826 8528
rect 32770 8472 32826 8508
rect 33138 9152 33194 9208
rect 32770 7928 32826 7984
rect 32586 5888 32642 5944
rect 32678 5616 32734 5672
rect 32862 6976 32918 7032
rect 33782 11756 33838 11792
rect 33782 11736 33784 11756
rect 33784 11736 33836 11756
rect 33836 11736 33838 11756
rect 33782 10648 33838 10704
rect 34610 15408 34666 15464
rect 34702 14592 34758 14648
rect 34794 14184 34850 14240
rect 35346 13368 35402 13424
rect 34289 13082 34345 13084
rect 34369 13082 34425 13084
rect 34449 13082 34505 13084
rect 34529 13082 34585 13084
rect 34289 13030 34315 13082
rect 34315 13030 34345 13082
rect 34369 13030 34379 13082
rect 34379 13030 34425 13082
rect 34449 13030 34495 13082
rect 34495 13030 34505 13082
rect 34529 13030 34559 13082
rect 34559 13030 34585 13082
rect 34289 13028 34345 13030
rect 34369 13028 34425 13030
rect 34449 13028 34505 13030
rect 34529 13028 34585 13030
rect 34794 12960 34850 13016
rect 34610 12688 34666 12744
rect 34334 12144 34390 12200
rect 34289 11994 34345 11996
rect 34369 11994 34425 11996
rect 34449 11994 34505 11996
rect 34529 11994 34585 11996
rect 34289 11942 34315 11994
rect 34315 11942 34345 11994
rect 34369 11942 34379 11994
rect 34379 11942 34425 11994
rect 34449 11942 34495 11994
rect 34495 11942 34505 11994
rect 34529 11942 34559 11994
rect 34559 11942 34585 11994
rect 34289 11940 34345 11942
rect 34369 11940 34425 11942
rect 34449 11940 34505 11942
rect 34529 11940 34585 11942
rect 34058 11328 34114 11384
rect 34610 11620 34666 11656
rect 34610 11600 34612 11620
rect 34612 11600 34664 11620
rect 34664 11600 34666 11620
rect 34518 11076 34574 11112
rect 34518 11056 34520 11076
rect 34520 11056 34572 11076
rect 34572 11056 34574 11076
rect 34289 10906 34345 10908
rect 34369 10906 34425 10908
rect 34449 10906 34505 10908
rect 34529 10906 34585 10908
rect 34289 10854 34315 10906
rect 34315 10854 34345 10906
rect 34369 10854 34379 10906
rect 34379 10854 34425 10906
rect 34449 10854 34495 10906
rect 34495 10854 34505 10906
rect 34529 10854 34559 10906
rect 34559 10854 34585 10906
rect 34289 10852 34345 10854
rect 34369 10852 34425 10854
rect 34449 10852 34505 10854
rect 34529 10852 34585 10854
rect 34150 10104 34206 10160
rect 34610 9968 34666 10024
rect 34289 9818 34345 9820
rect 34369 9818 34425 9820
rect 34449 9818 34505 9820
rect 34529 9818 34585 9820
rect 34289 9766 34315 9818
rect 34315 9766 34345 9818
rect 34369 9766 34379 9818
rect 34379 9766 34425 9818
rect 34449 9766 34495 9818
rect 34495 9766 34505 9818
rect 34529 9766 34559 9818
rect 34559 9766 34585 9818
rect 34289 9764 34345 9766
rect 34369 9764 34425 9766
rect 34449 9764 34505 9766
rect 34529 9764 34585 9766
rect 34150 9696 34206 9752
rect 33506 5072 33562 5128
rect 34058 8744 34114 8800
rect 34289 8730 34345 8732
rect 34369 8730 34425 8732
rect 34449 8730 34505 8732
rect 34529 8730 34585 8732
rect 34289 8678 34315 8730
rect 34315 8678 34345 8730
rect 34369 8678 34379 8730
rect 34379 8678 34425 8730
rect 34449 8678 34495 8730
rect 34495 8678 34505 8730
rect 34529 8678 34559 8730
rect 34559 8678 34585 8730
rect 34289 8676 34345 8678
rect 34369 8676 34425 8678
rect 34449 8676 34505 8678
rect 34529 8676 34585 8678
rect 33782 6976 33838 7032
rect 33782 6024 33838 6080
rect 33598 4936 33654 4992
rect 31482 3984 31538 4040
rect 32218 3984 32274 4040
rect 30010 3712 30066 3768
rect 35070 10648 35126 10704
rect 34886 9444 34942 9480
rect 34886 9424 34888 9444
rect 34888 9424 34940 9444
rect 34940 9424 34942 9444
rect 34289 7642 34345 7644
rect 34369 7642 34425 7644
rect 34449 7642 34505 7644
rect 34529 7642 34585 7644
rect 34289 7590 34315 7642
rect 34315 7590 34345 7642
rect 34369 7590 34379 7642
rect 34379 7590 34425 7642
rect 34449 7590 34495 7642
rect 34495 7590 34505 7642
rect 34529 7590 34559 7642
rect 34559 7590 34585 7642
rect 34289 7588 34345 7590
rect 34369 7588 34425 7590
rect 34449 7588 34505 7590
rect 34529 7588 34585 7590
rect 34150 7520 34206 7576
rect 34058 6704 34114 6760
rect 34289 6554 34345 6556
rect 34369 6554 34425 6556
rect 34449 6554 34505 6556
rect 34529 6554 34585 6556
rect 34289 6502 34315 6554
rect 34315 6502 34345 6554
rect 34369 6502 34379 6554
rect 34379 6502 34425 6554
rect 34449 6502 34495 6554
rect 34495 6502 34505 6554
rect 34529 6502 34559 6554
rect 34559 6502 34585 6554
rect 34289 6500 34345 6502
rect 34369 6500 34425 6502
rect 34449 6500 34505 6502
rect 34529 6500 34585 6502
rect 34289 5466 34345 5468
rect 34369 5466 34425 5468
rect 34449 5466 34505 5468
rect 34529 5466 34585 5468
rect 34289 5414 34315 5466
rect 34315 5414 34345 5466
rect 34369 5414 34379 5466
rect 34379 5414 34425 5466
rect 34449 5414 34495 5466
rect 34495 5414 34505 5466
rect 34529 5414 34559 5466
rect 34559 5414 34585 5466
rect 34289 5412 34345 5414
rect 34369 5412 34425 5414
rect 34449 5412 34505 5414
rect 34529 5412 34585 5414
rect 34289 4378 34345 4380
rect 34369 4378 34425 4380
rect 34449 4378 34505 4380
rect 34529 4378 34585 4380
rect 34289 4326 34315 4378
rect 34315 4326 34345 4378
rect 34369 4326 34379 4378
rect 34379 4326 34425 4378
rect 34449 4326 34495 4378
rect 34495 4326 34505 4378
rect 34529 4326 34559 4378
rect 34559 4326 34585 4378
rect 34289 4324 34345 4326
rect 34369 4324 34425 4326
rect 34449 4324 34505 4326
rect 34529 4324 34585 4326
rect 35070 7520 35126 7576
rect 35254 7792 35310 7848
rect 35162 7248 35218 7304
rect 35162 6976 35218 7032
rect 35254 6840 35310 6896
rect 35070 6432 35126 6488
rect 35070 5752 35126 5808
rect 35070 4936 35126 4992
rect 34289 3290 34345 3292
rect 34369 3290 34425 3292
rect 34449 3290 34505 3292
rect 34529 3290 34585 3292
rect 34289 3238 34315 3290
rect 34315 3238 34345 3290
rect 34369 3238 34379 3290
rect 34379 3238 34425 3290
rect 34449 3238 34495 3290
rect 34495 3238 34505 3290
rect 34529 3238 34559 3290
rect 34559 3238 34585 3290
rect 34289 3236 34345 3238
rect 34369 3236 34425 3238
rect 34449 3236 34505 3238
rect 34529 3236 34585 3238
rect 33782 2896 33838 2952
rect 27986 2488 28042 2544
rect 20956 2202 21012 2204
rect 21036 2202 21092 2204
rect 21116 2202 21172 2204
rect 21196 2202 21252 2204
rect 20956 2150 20982 2202
rect 20982 2150 21012 2202
rect 21036 2150 21046 2202
rect 21046 2150 21092 2202
rect 21116 2150 21162 2202
rect 21162 2150 21172 2202
rect 21196 2150 21226 2202
rect 21226 2150 21252 2202
rect 20956 2148 21012 2150
rect 21036 2148 21092 2150
rect 21116 2148 21172 2150
rect 21196 2148 21252 2150
rect 34289 2202 34345 2204
rect 34369 2202 34425 2204
rect 34449 2202 34505 2204
rect 34529 2202 34585 2204
rect 34289 2150 34315 2202
rect 34315 2150 34345 2202
rect 34369 2150 34379 2202
rect 34379 2150 34425 2202
rect 34449 2150 34495 2202
rect 34495 2150 34505 2202
rect 34529 2150 34559 2202
rect 34559 2150 34585 2202
rect 34289 2148 34345 2150
rect 34369 2148 34425 2150
rect 34449 2148 34505 2150
rect 34529 2148 34585 2150
rect 22006 1808 22062 1864
rect 22006 1400 22062 1456
rect 34886 1264 34942 1320
rect 3606 176 3662 232
rect 35070 448 35126 504
rect 35714 12144 35770 12200
rect 35438 10240 35494 10296
rect 36450 15000 36506 15056
rect 36634 13776 36690 13832
rect 35806 11056 35862 11112
rect 35714 10648 35770 10704
rect 35438 9832 35494 9888
rect 35714 9560 35770 9616
rect 36358 10104 36414 10160
rect 35806 8608 35862 8664
rect 35806 8336 35862 8392
rect 35438 7112 35494 7168
rect 35438 5616 35494 5672
rect 36266 8508 36268 8528
rect 36268 8508 36320 8528
rect 36320 8508 36322 8528
rect 36266 8472 36322 8508
rect 35990 7964 35992 7984
rect 35992 7964 36044 7984
rect 36044 7964 36046 7984
rect 35990 7928 36046 7964
rect 35898 6976 35954 7032
rect 35806 6840 35862 6896
rect 36082 6840 36138 6896
rect 35438 4684 35494 4720
rect 35438 4664 35440 4684
rect 35440 4664 35492 4684
rect 35492 4664 35494 4684
rect 35438 3712 35494 3768
rect 36542 9016 36598 9072
rect 36450 5888 36506 5944
rect 37462 11872 37518 11928
rect 37554 11756 37610 11792
rect 37554 11736 37556 11756
rect 37556 11736 37608 11756
rect 37608 11736 37610 11756
rect 36818 9152 36874 9208
rect 37646 9560 37702 9616
rect 37370 9016 37426 9072
rect 36910 8744 36966 8800
rect 37278 8628 37334 8664
rect 37278 8608 37280 8628
rect 37280 8608 37332 8628
rect 37332 8608 37334 8628
rect 37554 7928 37610 7984
rect 36358 4392 36414 4448
rect 37370 3848 37426 3904
rect 35806 856 35862 912
rect 35162 176 35218 232
<< metal3 >>
rect 0 15874 480 15904
rect 3601 15874 3667 15877
rect 0 15872 3667 15874
rect 0 15816 3606 15872
rect 3662 15816 3667 15872
rect 0 15814 3667 15816
rect 0 15784 480 15814
rect 3601 15811 3667 15814
rect 34513 15874 34579 15877
rect 39520 15874 40000 15904
rect 34513 15872 40000 15874
rect 34513 15816 34518 15872
rect 34574 15816 40000 15872
rect 34513 15814 40000 15816
rect 34513 15811 34579 15814
rect 39520 15784 40000 15814
rect 0 15466 480 15496
rect 3233 15466 3299 15469
rect 0 15464 3299 15466
rect 0 15408 3238 15464
rect 3294 15408 3299 15464
rect 0 15406 3299 15408
rect 0 15376 480 15406
rect 3233 15403 3299 15406
rect 34605 15466 34671 15469
rect 39520 15466 40000 15496
rect 34605 15464 40000 15466
rect 34605 15408 34610 15464
rect 34666 15408 40000 15464
rect 34605 15406 40000 15408
rect 34605 15403 34671 15406
rect 39520 15376 40000 15406
rect 0 15058 480 15088
rect 3509 15058 3575 15061
rect 0 15056 3575 15058
rect 0 15000 3514 15056
rect 3570 15000 3575 15056
rect 0 14998 3575 15000
rect 0 14968 480 14998
rect 3509 14995 3575 14998
rect 36445 15058 36511 15061
rect 39520 15058 40000 15088
rect 36445 15056 40000 15058
rect 36445 15000 36450 15056
rect 36506 15000 40000 15056
rect 36445 14998 40000 15000
rect 36445 14995 36511 14998
rect 39520 14968 40000 14998
rect 0 14650 480 14680
rect 3141 14650 3207 14653
rect 0 14648 3207 14650
rect 0 14592 3146 14648
rect 3202 14592 3207 14648
rect 0 14590 3207 14592
rect 0 14560 480 14590
rect 3141 14587 3207 14590
rect 34697 14650 34763 14653
rect 39520 14650 40000 14680
rect 34697 14648 40000 14650
rect 34697 14592 34702 14648
rect 34758 14592 40000 14648
rect 34697 14590 40000 14592
rect 34697 14587 34763 14590
rect 39520 14560 40000 14590
rect 0 14242 480 14272
rect 3049 14242 3115 14245
rect 0 14240 3115 14242
rect 0 14184 3054 14240
rect 3110 14184 3115 14240
rect 0 14182 3115 14184
rect 0 14152 480 14182
rect 3049 14179 3115 14182
rect 34789 14242 34855 14245
rect 39520 14242 40000 14272
rect 34789 14240 40000 14242
rect 34789 14184 34794 14240
rect 34850 14184 40000 14240
rect 34789 14182 40000 14184
rect 34789 14179 34855 14182
rect 39520 14152 40000 14182
rect 0 13834 480 13864
rect 3417 13834 3483 13837
rect 0 13832 3483 13834
rect 0 13776 3422 13832
rect 3478 13776 3483 13832
rect 0 13774 3483 13776
rect 0 13744 480 13774
rect 3417 13771 3483 13774
rect 36629 13834 36695 13837
rect 39520 13834 40000 13864
rect 36629 13832 40000 13834
rect 36629 13776 36634 13832
rect 36690 13776 40000 13832
rect 36629 13774 40000 13776
rect 36629 13771 36695 13774
rect 39520 13744 40000 13774
rect 14277 13632 14597 13633
rect 14277 13568 14285 13632
rect 14349 13568 14365 13632
rect 14429 13568 14445 13632
rect 14509 13568 14525 13632
rect 14589 13568 14597 13632
rect 14277 13567 14597 13568
rect 27610 13632 27930 13633
rect 27610 13568 27618 13632
rect 27682 13568 27698 13632
rect 27762 13568 27778 13632
rect 27842 13568 27858 13632
rect 27922 13568 27930 13632
rect 27610 13567 27930 13568
rect 0 13426 480 13456
rect 2773 13426 2839 13429
rect 0 13424 2839 13426
rect 0 13368 2778 13424
rect 2834 13368 2839 13424
rect 0 13366 2839 13368
rect 0 13336 480 13366
rect 2773 13363 2839 13366
rect 35341 13426 35407 13429
rect 39520 13426 40000 13456
rect 35341 13424 40000 13426
rect 35341 13368 35346 13424
rect 35402 13368 40000 13424
rect 35341 13366 40000 13368
rect 35341 13363 35407 13366
rect 39520 13336 40000 13366
rect 7610 13088 7930 13089
rect 0 13018 480 13048
rect 7610 13024 7618 13088
rect 7682 13024 7698 13088
rect 7762 13024 7778 13088
rect 7842 13024 7858 13088
rect 7922 13024 7930 13088
rect 7610 13023 7930 13024
rect 20944 13088 21264 13089
rect 20944 13024 20952 13088
rect 21016 13024 21032 13088
rect 21096 13024 21112 13088
rect 21176 13024 21192 13088
rect 21256 13024 21264 13088
rect 20944 13023 21264 13024
rect 34277 13088 34597 13089
rect 34277 13024 34285 13088
rect 34349 13024 34365 13088
rect 34429 13024 34445 13088
rect 34509 13024 34525 13088
rect 34589 13024 34597 13088
rect 34277 13023 34597 13024
rect 4061 13018 4127 13021
rect 0 13016 4127 13018
rect 0 12960 4066 13016
rect 4122 12960 4127 13016
rect 0 12958 4127 12960
rect 0 12928 480 12958
rect 4061 12955 4127 12958
rect 34789 13018 34855 13021
rect 39520 13018 40000 13048
rect 34789 13016 40000 13018
rect 34789 12960 34794 13016
rect 34850 12960 40000 13016
rect 34789 12958 40000 12960
rect 34789 12955 34855 12958
rect 39520 12928 40000 12958
rect 34605 12746 34671 12749
rect 39520 12746 40000 12776
rect 34605 12744 40000 12746
rect 34605 12688 34610 12744
rect 34666 12688 40000 12744
rect 34605 12686 40000 12688
rect 34605 12683 34671 12686
rect 39520 12656 40000 12686
rect 0 12610 480 12640
rect 3417 12610 3483 12613
rect 24761 12612 24827 12613
rect 0 12608 3483 12610
rect 0 12552 3422 12608
rect 3478 12552 3483 12608
rect 0 12550 3483 12552
rect 0 12520 480 12550
rect 3417 12547 3483 12550
rect 24710 12548 24716 12612
rect 24780 12610 24827 12612
rect 24780 12608 24872 12610
rect 24822 12552 24872 12608
rect 24780 12550 24872 12552
rect 24780 12548 24827 12550
rect 24761 12547 24827 12548
rect 14277 12544 14597 12545
rect 14277 12480 14285 12544
rect 14349 12480 14365 12544
rect 14429 12480 14445 12544
rect 14509 12480 14525 12544
rect 14589 12480 14597 12544
rect 14277 12479 14597 12480
rect 27610 12544 27930 12545
rect 27610 12480 27618 12544
rect 27682 12480 27698 12544
rect 27762 12480 27778 12544
rect 27842 12480 27858 12544
rect 27922 12480 27930 12544
rect 27610 12479 27930 12480
rect 29545 12338 29611 12341
rect 39520 12338 40000 12368
rect 29545 12336 40000 12338
rect 29545 12280 29550 12336
rect 29606 12280 40000 12336
rect 29545 12278 40000 12280
rect 29545 12275 29611 12278
rect 39520 12248 40000 12278
rect 0 12202 480 12232
rect 3509 12202 3575 12205
rect 0 12200 3575 12202
rect 0 12144 3514 12200
rect 3570 12144 3575 12200
rect 0 12142 3575 12144
rect 0 12112 480 12142
rect 3509 12139 3575 12142
rect 27245 12202 27311 12205
rect 34329 12202 34395 12205
rect 35709 12202 35775 12205
rect 27245 12200 35775 12202
rect 27245 12144 27250 12200
rect 27306 12144 34334 12200
rect 34390 12144 35714 12200
rect 35770 12144 35775 12200
rect 27245 12142 35775 12144
rect 27245 12139 27311 12142
rect 34329 12139 34395 12142
rect 35709 12139 35775 12142
rect 25037 12066 25103 12069
rect 33133 12066 33199 12069
rect 25037 12064 33199 12066
rect 25037 12008 25042 12064
rect 25098 12008 33138 12064
rect 33194 12008 33199 12064
rect 25037 12006 33199 12008
rect 25037 12003 25103 12006
rect 33133 12003 33199 12006
rect 7610 12000 7930 12001
rect 7610 11936 7618 12000
rect 7682 11936 7698 12000
rect 7762 11936 7778 12000
rect 7842 11936 7858 12000
rect 7922 11936 7930 12000
rect 7610 11935 7930 11936
rect 20944 12000 21264 12001
rect 20944 11936 20952 12000
rect 21016 11936 21032 12000
rect 21096 11936 21112 12000
rect 21176 11936 21192 12000
rect 21256 11936 21264 12000
rect 20944 11935 21264 11936
rect 34277 12000 34597 12001
rect 34277 11936 34285 12000
rect 34349 11936 34365 12000
rect 34429 11936 34445 12000
rect 34509 11936 34525 12000
rect 34589 11936 34597 12000
rect 34277 11935 34597 11936
rect 8017 11930 8083 11933
rect 10685 11930 10751 11933
rect 8017 11928 10751 11930
rect 8017 11872 8022 11928
rect 8078 11872 10690 11928
rect 10746 11872 10751 11928
rect 8017 11870 10751 11872
rect 8017 11867 8083 11870
rect 10685 11867 10751 11870
rect 25589 11930 25655 11933
rect 31937 11930 32003 11933
rect 25589 11928 32003 11930
rect 25589 11872 25594 11928
rect 25650 11872 31942 11928
rect 31998 11872 32003 11928
rect 25589 11870 32003 11872
rect 25589 11867 25655 11870
rect 31937 11867 32003 11870
rect 37457 11930 37523 11933
rect 39520 11930 40000 11960
rect 37457 11928 40000 11930
rect 37457 11872 37462 11928
rect 37518 11872 40000 11928
rect 37457 11870 40000 11872
rect 37457 11867 37523 11870
rect 39520 11840 40000 11870
rect 0 11794 480 11824
rect 3877 11794 3943 11797
rect 0 11792 3943 11794
rect 0 11736 3882 11792
rect 3938 11736 3943 11792
rect 0 11734 3943 11736
rect 0 11704 480 11734
rect 3877 11731 3943 11734
rect 19977 11794 20043 11797
rect 29361 11794 29427 11797
rect 19977 11792 29427 11794
rect 19977 11736 19982 11792
rect 20038 11736 29366 11792
rect 29422 11736 29427 11792
rect 19977 11734 29427 11736
rect 19977 11731 20043 11734
rect 29361 11731 29427 11734
rect 33777 11794 33843 11797
rect 37549 11794 37615 11797
rect 33777 11792 37615 11794
rect 33777 11736 33782 11792
rect 33838 11736 37554 11792
rect 37610 11736 37615 11792
rect 33777 11734 37615 11736
rect 33777 11731 33843 11734
rect 37549 11731 37615 11734
rect 2405 11658 2471 11661
rect 6821 11658 6887 11661
rect 2405 11656 6887 11658
rect 2405 11600 2410 11656
rect 2466 11600 6826 11656
rect 6882 11600 6887 11656
rect 2405 11598 6887 11600
rect 2405 11595 2471 11598
rect 6821 11595 6887 11598
rect 8293 11658 8359 11661
rect 11605 11658 11671 11661
rect 8293 11656 11671 11658
rect 8293 11600 8298 11656
rect 8354 11600 11610 11656
rect 11666 11600 11671 11656
rect 8293 11598 11671 11600
rect 8293 11595 8359 11598
rect 11605 11595 11671 11598
rect 17125 11658 17191 11661
rect 25037 11658 25103 11661
rect 17125 11656 25103 11658
rect 17125 11600 17130 11656
rect 17186 11600 25042 11656
rect 25098 11600 25103 11656
rect 17125 11598 25103 11600
rect 17125 11595 17191 11598
rect 25037 11595 25103 11598
rect 29913 11658 29979 11661
rect 34605 11658 34671 11661
rect 29913 11656 34671 11658
rect 29913 11600 29918 11656
rect 29974 11600 34610 11656
rect 34666 11600 34671 11656
rect 29913 11598 34671 11600
rect 29913 11595 29979 11598
rect 34605 11595 34671 11598
rect 2497 11522 2563 11525
rect 2998 11522 3004 11524
rect 2497 11520 3004 11522
rect 2497 11464 2502 11520
rect 2558 11464 3004 11520
rect 2497 11462 3004 11464
rect 2497 11459 2563 11462
rect 2998 11460 3004 11462
rect 3068 11460 3074 11524
rect 19057 11522 19123 11525
rect 20805 11522 20871 11525
rect 19057 11520 20871 11522
rect 19057 11464 19062 11520
rect 19118 11464 20810 11520
rect 20866 11464 20871 11520
rect 19057 11462 20871 11464
rect 19057 11459 19123 11462
rect 20805 11459 20871 11462
rect 25129 11522 25195 11525
rect 25589 11522 25655 11525
rect 25129 11520 25655 11522
rect 25129 11464 25134 11520
rect 25190 11464 25594 11520
rect 25650 11464 25655 11520
rect 25129 11462 25655 11464
rect 25129 11459 25195 11462
rect 25589 11459 25655 11462
rect 32305 11522 32371 11525
rect 39520 11522 40000 11552
rect 32305 11520 40000 11522
rect 32305 11464 32310 11520
rect 32366 11464 40000 11520
rect 32305 11462 40000 11464
rect 32305 11459 32371 11462
rect 14277 11456 14597 11457
rect 0 11386 480 11416
rect 14277 11392 14285 11456
rect 14349 11392 14365 11456
rect 14429 11392 14445 11456
rect 14509 11392 14525 11456
rect 14589 11392 14597 11456
rect 14277 11391 14597 11392
rect 27610 11456 27930 11457
rect 27610 11392 27618 11456
rect 27682 11392 27698 11456
rect 27762 11392 27778 11456
rect 27842 11392 27858 11456
rect 27922 11392 27930 11456
rect 39520 11432 40000 11462
rect 27610 11391 27930 11392
rect 4061 11386 4127 11389
rect 0 11384 4127 11386
rect 0 11328 4066 11384
rect 4122 11328 4127 11384
rect 0 11326 4127 11328
rect 0 11296 480 11326
rect 4061 11323 4127 11326
rect 16481 11386 16547 11389
rect 18873 11386 18939 11389
rect 16481 11384 18939 11386
rect 16481 11328 16486 11384
rect 16542 11328 18878 11384
rect 18934 11328 18939 11384
rect 16481 11326 18939 11328
rect 16481 11323 16547 11326
rect 18873 11323 18939 11326
rect 30925 11386 30991 11389
rect 34053 11386 34119 11389
rect 30925 11384 34119 11386
rect 30925 11328 30930 11384
rect 30986 11328 34058 11384
rect 34114 11328 34119 11384
rect 30925 11326 34119 11328
rect 30925 11323 30991 11326
rect 34053 11323 34119 11326
rect 7557 11250 7623 11253
rect 15101 11250 15167 11253
rect 7557 11248 15167 11250
rect 7557 11192 7562 11248
rect 7618 11192 15106 11248
rect 15162 11192 15167 11248
rect 7557 11190 15167 11192
rect 7557 11187 7623 11190
rect 15101 11187 15167 11190
rect 15745 11250 15811 11253
rect 21633 11250 21699 11253
rect 15745 11248 21699 11250
rect 15745 11192 15750 11248
rect 15806 11192 21638 11248
rect 21694 11192 21699 11248
rect 15745 11190 21699 11192
rect 15745 11187 15811 11190
rect 21633 11187 21699 11190
rect 24669 11250 24735 11253
rect 26233 11250 26299 11253
rect 24669 11248 26299 11250
rect 24669 11192 24674 11248
rect 24730 11192 26238 11248
rect 26294 11192 26299 11248
rect 24669 11190 26299 11192
rect 24669 11187 24735 11190
rect 26233 11187 26299 11190
rect 3601 11114 3667 11117
rect 10777 11114 10843 11117
rect 3601 11112 10843 11114
rect 3601 11056 3606 11112
rect 3662 11056 10782 11112
rect 10838 11056 10843 11112
rect 3601 11054 10843 11056
rect 3601 11051 3667 11054
rect 10777 11051 10843 11054
rect 11697 11114 11763 11117
rect 13905 11114 13971 11117
rect 11697 11112 13971 11114
rect 11697 11056 11702 11112
rect 11758 11056 13910 11112
rect 13966 11056 13971 11112
rect 11697 11054 13971 11056
rect 11697 11051 11763 11054
rect 13905 11051 13971 11054
rect 21817 11114 21883 11117
rect 23749 11114 23815 11117
rect 21817 11112 23815 11114
rect 21817 11056 21822 11112
rect 21878 11056 23754 11112
rect 23810 11056 23815 11112
rect 21817 11054 23815 11056
rect 21817 11051 21883 11054
rect 23749 11051 23815 11054
rect 24301 11114 24367 11117
rect 26601 11114 26667 11117
rect 34513 11114 34579 11117
rect 24301 11112 26667 11114
rect 24301 11056 24306 11112
rect 24362 11056 26606 11112
rect 26662 11056 26667 11112
rect 24301 11054 26667 11056
rect 24301 11051 24367 11054
rect 26601 11051 26667 11054
rect 34102 11112 34579 11114
rect 34102 11056 34518 11112
rect 34574 11056 34579 11112
rect 34102 11054 34579 11056
rect 0 10978 480 11008
rect 1301 10978 1367 10981
rect 0 10976 1367 10978
rect 0 10920 1306 10976
rect 1362 10920 1367 10976
rect 0 10918 1367 10920
rect 0 10888 480 10918
rect 1301 10915 1367 10918
rect 23013 10978 23079 10981
rect 25037 10978 25103 10981
rect 23013 10976 25103 10978
rect 23013 10920 23018 10976
rect 23074 10920 25042 10976
rect 25098 10920 25103 10976
rect 23013 10918 25103 10920
rect 23013 10915 23079 10918
rect 25037 10915 25103 10918
rect 25221 10978 25287 10981
rect 34102 10978 34162 11054
rect 34513 11051 34579 11054
rect 35801 11114 35867 11117
rect 39520 11114 40000 11144
rect 35801 11112 40000 11114
rect 35801 11056 35806 11112
rect 35862 11056 40000 11112
rect 35801 11054 40000 11056
rect 35801 11051 35867 11054
rect 39520 11024 40000 11054
rect 25221 10976 34162 10978
rect 25221 10920 25226 10976
rect 25282 10920 34162 10976
rect 25221 10918 34162 10920
rect 25221 10915 25287 10918
rect 7610 10912 7930 10913
rect 7610 10848 7618 10912
rect 7682 10848 7698 10912
rect 7762 10848 7778 10912
rect 7842 10848 7858 10912
rect 7922 10848 7930 10912
rect 7610 10847 7930 10848
rect 20944 10912 21264 10913
rect 20944 10848 20952 10912
rect 21016 10848 21032 10912
rect 21096 10848 21112 10912
rect 21176 10848 21192 10912
rect 21256 10848 21264 10912
rect 20944 10847 21264 10848
rect 34277 10912 34597 10913
rect 34277 10848 34285 10912
rect 34349 10848 34365 10912
rect 34429 10848 34445 10912
rect 34509 10848 34525 10912
rect 34589 10848 34597 10912
rect 34277 10847 34597 10848
rect 5625 10842 5691 10845
rect 24761 10842 24827 10845
rect 27797 10842 27863 10845
rect 5625 10840 7298 10842
rect 5625 10784 5630 10840
rect 5686 10784 7298 10840
rect 5625 10782 7298 10784
rect 5625 10779 5691 10782
rect 7238 10706 7298 10782
rect 24761 10840 27863 10842
rect 24761 10784 24766 10840
rect 24822 10784 27802 10840
rect 27858 10784 27863 10840
rect 24761 10782 27863 10784
rect 24761 10779 24827 10782
rect 27797 10779 27863 10782
rect 9489 10706 9555 10709
rect 7238 10704 9555 10706
rect 7238 10648 9494 10704
rect 9550 10648 9555 10704
rect 7238 10646 9555 10648
rect 9489 10643 9555 10646
rect 19057 10706 19123 10709
rect 22277 10706 22343 10709
rect 19057 10704 22343 10706
rect 19057 10648 19062 10704
rect 19118 10648 22282 10704
rect 22338 10648 22343 10704
rect 19057 10646 22343 10648
rect 19057 10643 19123 10646
rect 22277 10643 22343 10646
rect 24025 10706 24091 10709
rect 27337 10706 27403 10709
rect 29545 10706 29611 10709
rect 24025 10704 29611 10706
rect 24025 10648 24030 10704
rect 24086 10648 27342 10704
rect 27398 10648 29550 10704
rect 29606 10648 29611 10704
rect 24025 10646 29611 10648
rect 24025 10643 24091 10646
rect 27337 10643 27403 10646
rect 29545 10643 29611 10646
rect 33777 10706 33843 10709
rect 35065 10706 35131 10709
rect 33777 10704 35131 10706
rect 33777 10648 33782 10704
rect 33838 10648 35070 10704
rect 35126 10648 35131 10704
rect 33777 10646 35131 10648
rect 33777 10643 33843 10646
rect 35065 10643 35131 10646
rect 35709 10706 35775 10709
rect 39520 10706 40000 10736
rect 35709 10704 40000 10706
rect 35709 10648 35714 10704
rect 35770 10648 40000 10704
rect 35709 10646 40000 10648
rect 35709 10643 35775 10646
rect 39520 10616 40000 10646
rect 0 10570 480 10600
rect 3877 10570 3943 10573
rect 0 10568 3943 10570
rect 0 10512 3882 10568
rect 3938 10512 3943 10568
rect 0 10510 3943 10512
rect 0 10480 480 10510
rect 3877 10507 3943 10510
rect 5625 10570 5691 10573
rect 25129 10570 25195 10573
rect 32949 10570 33015 10573
rect 5625 10568 25195 10570
rect 5625 10512 5630 10568
rect 5686 10512 25134 10568
rect 25190 10512 25195 10568
rect 5625 10510 25195 10512
rect 5625 10507 5691 10510
rect 25129 10507 25195 10510
rect 26926 10568 33015 10570
rect 26926 10512 32954 10568
rect 33010 10512 33015 10568
rect 26926 10510 33015 10512
rect 9121 10434 9187 10437
rect 11145 10434 11211 10437
rect 9121 10432 11211 10434
rect 9121 10376 9126 10432
rect 9182 10376 11150 10432
rect 11206 10376 11211 10432
rect 9121 10374 11211 10376
rect 9121 10371 9187 10374
rect 11145 10371 11211 10374
rect 14277 10368 14597 10369
rect 14277 10304 14285 10368
rect 14349 10304 14365 10368
rect 14429 10304 14445 10368
rect 14509 10304 14525 10368
rect 14589 10304 14597 10368
rect 14277 10303 14597 10304
rect 8017 10298 8083 10301
rect 10317 10298 10383 10301
rect 8017 10296 10383 10298
rect 8017 10240 8022 10296
rect 8078 10240 10322 10296
rect 10378 10240 10383 10296
rect 8017 10238 10383 10240
rect 8017 10235 8083 10238
rect 10317 10235 10383 10238
rect 20662 10236 20668 10300
rect 20732 10298 20738 10300
rect 22001 10298 22067 10301
rect 26926 10298 26986 10510
rect 32949 10507 33015 10510
rect 27610 10368 27930 10369
rect 27610 10304 27618 10368
rect 27682 10304 27698 10368
rect 27762 10304 27778 10368
rect 27842 10304 27858 10368
rect 27922 10304 27930 10368
rect 27610 10303 27930 10304
rect 20732 10296 26986 10298
rect 20732 10240 22006 10296
rect 22062 10240 26986 10296
rect 20732 10238 26986 10240
rect 35433 10298 35499 10301
rect 39520 10298 40000 10328
rect 35433 10296 40000 10298
rect 35433 10240 35438 10296
rect 35494 10240 40000 10296
rect 35433 10238 40000 10240
rect 20732 10236 20738 10238
rect 22001 10235 22067 10238
rect 35433 10235 35499 10238
rect 39520 10208 40000 10238
rect 0 10162 480 10192
rect 2865 10162 2931 10165
rect 0 10160 2931 10162
rect 0 10104 2870 10160
rect 2926 10104 2931 10160
rect 0 10102 2931 10104
rect 0 10072 480 10102
rect 2865 10099 2931 10102
rect 34145 10162 34211 10165
rect 36353 10162 36419 10165
rect 34145 10160 36419 10162
rect 34145 10104 34150 10160
rect 34206 10104 36358 10160
rect 36414 10104 36419 10160
rect 34145 10102 36419 10104
rect 34145 10099 34211 10102
rect 36353 10099 36419 10102
rect 2497 10026 2563 10029
rect 4613 10026 4679 10029
rect 2497 10024 4679 10026
rect 2497 9968 2502 10024
rect 2558 9968 4618 10024
rect 4674 9968 4679 10024
rect 2497 9966 4679 9968
rect 2497 9963 2563 9966
rect 4613 9963 4679 9966
rect 6637 10026 6703 10029
rect 8385 10026 8451 10029
rect 6637 10024 8451 10026
rect 6637 9968 6642 10024
rect 6698 9968 8390 10024
rect 8446 9968 8451 10024
rect 6637 9966 8451 9968
rect 6637 9963 6703 9966
rect 8385 9963 8451 9966
rect 11605 10026 11671 10029
rect 25313 10026 25379 10029
rect 11605 10024 25379 10026
rect 11605 9968 11610 10024
rect 11666 9968 25318 10024
rect 25374 9968 25379 10024
rect 11605 9966 25379 9968
rect 11605 9963 11671 9966
rect 25313 9963 25379 9966
rect 26141 10026 26207 10029
rect 34605 10026 34671 10029
rect 26141 10024 34671 10026
rect 26141 9968 26146 10024
rect 26202 9968 34610 10024
rect 34666 9968 34671 10024
rect 26141 9966 34671 9968
rect 26141 9963 26207 9966
rect 34605 9963 34671 9966
rect 2589 9890 2655 9893
rect 3969 9890 4035 9893
rect 20805 9890 20871 9893
rect 2589 9888 4035 9890
rect 2589 9832 2594 9888
rect 2650 9832 3974 9888
rect 4030 9832 4035 9888
rect 2589 9830 4035 9832
rect 2589 9827 2655 9830
rect 3969 9827 4035 9830
rect 15886 9888 20871 9890
rect 15886 9832 20810 9888
rect 20866 9832 20871 9888
rect 15886 9830 20871 9832
rect 7610 9824 7930 9825
rect 0 9754 480 9784
rect 7610 9760 7618 9824
rect 7682 9760 7698 9824
rect 7762 9760 7778 9824
rect 7842 9760 7858 9824
rect 7922 9760 7930 9824
rect 7610 9759 7930 9760
rect 2773 9754 2839 9757
rect 0 9752 2839 9754
rect 0 9696 2778 9752
rect 2834 9696 2839 9752
rect 0 9694 2839 9696
rect 0 9664 480 9694
rect 2773 9691 2839 9694
rect 10501 9754 10567 9757
rect 15285 9754 15351 9757
rect 15886 9754 15946 9830
rect 20805 9827 20871 9830
rect 35433 9890 35499 9893
rect 39520 9890 40000 9920
rect 35433 9888 40000 9890
rect 35433 9832 35438 9888
rect 35494 9832 40000 9888
rect 35433 9830 40000 9832
rect 35433 9827 35499 9830
rect 20944 9824 21264 9825
rect 20944 9760 20952 9824
rect 21016 9760 21032 9824
rect 21096 9760 21112 9824
rect 21176 9760 21192 9824
rect 21256 9760 21264 9824
rect 20944 9759 21264 9760
rect 34277 9824 34597 9825
rect 34277 9760 34285 9824
rect 34349 9760 34365 9824
rect 34429 9760 34445 9824
rect 34509 9760 34525 9824
rect 34589 9760 34597 9824
rect 39520 9800 40000 9830
rect 34277 9759 34597 9760
rect 10501 9752 15946 9754
rect 10501 9696 10506 9752
rect 10562 9696 15290 9752
rect 15346 9696 15946 9752
rect 10501 9694 15946 9696
rect 16021 9754 16087 9757
rect 34145 9754 34211 9757
rect 16021 9752 20730 9754
rect 16021 9696 16026 9752
rect 16082 9696 20730 9752
rect 16021 9694 20730 9696
rect 10501 9691 10567 9694
rect 15285 9691 15351 9694
rect 16021 9691 16087 9694
rect 8569 9618 8635 9621
rect 12985 9618 13051 9621
rect 14181 9618 14247 9621
rect 17585 9618 17651 9621
rect 8569 9616 17651 9618
rect 8569 9560 8574 9616
rect 8630 9560 12990 9616
rect 13046 9560 14186 9616
rect 14242 9560 17590 9616
rect 17646 9560 17651 9616
rect 8569 9558 17651 9560
rect 20670 9618 20730 9694
rect 21406 9752 34211 9754
rect 21406 9696 34150 9752
rect 34206 9696 34211 9752
rect 21406 9694 34211 9696
rect 21406 9618 21466 9694
rect 34145 9691 34211 9694
rect 26877 9618 26943 9621
rect 20670 9558 21466 9618
rect 21590 9616 26943 9618
rect 21590 9560 26882 9616
rect 26938 9560 26943 9616
rect 21590 9558 26943 9560
rect 8569 9555 8635 9558
rect 12985 9555 13051 9558
rect 14181 9555 14247 9558
rect 17585 9555 17651 9558
rect 8109 9482 8175 9485
rect 12617 9482 12683 9485
rect 13629 9482 13695 9485
rect 18045 9482 18111 9485
rect 21590 9482 21650 9558
rect 26877 9555 26943 9558
rect 29821 9618 29887 9621
rect 35709 9618 35775 9621
rect 29821 9616 35775 9618
rect 29821 9560 29826 9616
rect 29882 9560 35714 9616
rect 35770 9560 35775 9616
rect 29821 9558 35775 9560
rect 29821 9555 29887 9558
rect 35709 9555 35775 9558
rect 37641 9618 37707 9621
rect 39520 9618 40000 9648
rect 37641 9616 40000 9618
rect 37641 9560 37646 9616
rect 37702 9560 40000 9616
rect 37641 9558 40000 9560
rect 37641 9555 37707 9558
rect 39520 9528 40000 9558
rect 8109 9480 21650 9482
rect 8109 9424 8114 9480
rect 8170 9424 12622 9480
rect 12678 9424 13634 9480
rect 13690 9424 18050 9480
rect 18106 9424 21650 9480
rect 8109 9422 21650 9424
rect 21817 9482 21883 9485
rect 26509 9482 26575 9485
rect 27429 9482 27495 9485
rect 34881 9482 34947 9485
rect 21817 9480 26575 9482
rect 21817 9424 21822 9480
rect 21878 9424 26514 9480
rect 26570 9424 26575 9480
rect 21817 9422 26575 9424
rect 8109 9419 8175 9422
rect 12617 9419 12683 9422
rect 13629 9419 13695 9422
rect 18045 9419 18111 9422
rect 21817 9419 21883 9422
rect 26509 9419 26575 9422
rect 26742 9480 34947 9482
rect 26742 9424 27434 9480
rect 27490 9424 34886 9480
rect 34942 9424 34947 9480
rect 26742 9422 34947 9424
rect 0 9346 480 9376
rect 4061 9346 4127 9349
rect 0 9344 4127 9346
rect 0 9288 4066 9344
rect 4122 9288 4127 9344
rect 0 9286 4127 9288
rect 0 9256 480 9286
rect 4061 9283 4127 9286
rect 7281 9346 7347 9349
rect 8150 9346 8156 9348
rect 7281 9344 8156 9346
rect 7281 9288 7286 9344
rect 7342 9288 8156 9344
rect 7281 9286 8156 9288
rect 7281 9283 7347 9286
rect 8150 9284 8156 9286
rect 8220 9284 8226 9348
rect 19885 9346 19951 9349
rect 22369 9346 22435 9349
rect 19885 9344 22435 9346
rect 19885 9288 19890 9344
rect 19946 9288 22374 9344
rect 22430 9288 22435 9344
rect 19885 9286 22435 9288
rect 19885 9283 19951 9286
rect 22369 9283 22435 9286
rect 23933 9346 23999 9349
rect 26742 9346 26802 9422
rect 27429 9419 27495 9422
rect 34881 9419 34947 9422
rect 23933 9344 26802 9346
rect 23933 9288 23938 9344
rect 23994 9288 26802 9344
rect 23933 9286 26802 9288
rect 23933 9283 23999 9286
rect 14277 9280 14597 9281
rect 14277 9216 14285 9280
rect 14349 9216 14365 9280
rect 14429 9216 14445 9280
rect 14509 9216 14525 9280
rect 14589 9216 14597 9280
rect 14277 9215 14597 9216
rect 27610 9280 27930 9281
rect 27610 9216 27618 9280
rect 27682 9216 27698 9280
rect 27762 9216 27778 9280
rect 27842 9216 27858 9280
rect 27922 9216 27930 9280
rect 27610 9215 27930 9216
rect 5257 9210 5323 9213
rect 9673 9210 9739 9213
rect 5257 9208 9739 9210
rect 5257 9152 5262 9208
rect 5318 9152 9678 9208
rect 9734 9152 9739 9208
rect 5257 9150 9739 9152
rect 5257 9147 5323 9150
rect 9673 9147 9739 9150
rect 20529 9210 20595 9213
rect 24025 9210 24091 9213
rect 20529 9208 24091 9210
rect 20529 9152 20534 9208
rect 20590 9152 24030 9208
rect 24086 9152 24091 9208
rect 20529 9150 24091 9152
rect 20529 9147 20595 9150
rect 24025 9147 24091 9150
rect 28625 9210 28691 9213
rect 33133 9210 33199 9213
rect 36813 9210 36879 9213
rect 39520 9210 40000 9240
rect 28625 9208 36738 9210
rect 28625 9152 28630 9208
rect 28686 9152 33138 9208
rect 33194 9152 36738 9208
rect 28625 9150 36738 9152
rect 28625 9147 28691 9150
rect 33133 9147 33199 9150
rect 2681 9074 2747 9077
rect 7373 9074 7439 9077
rect 2681 9072 7439 9074
rect 2681 9016 2686 9072
rect 2742 9016 7378 9072
rect 7434 9016 7439 9072
rect 2681 9014 7439 9016
rect 2681 9011 2747 9014
rect 7373 9011 7439 9014
rect 13261 9074 13327 9077
rect 15377 9074 15443 9077
rect 13261 9072 15443 9074
rect 13261 9016 13266 9072
rect 13322 9016 15382 9072
rect 15438 9016 15443 9072
rect 13261 9014 15443 9016
rect 13261 9011 13327 9014
rect 15377 9011 15443 9014
rect 20805 9074 20871 9077
rect 21357 9074 21423 9077
rect 26969 9074 27035 9077
rect 30833 9074 30899 9077
rect 20805 9072 26802 9074
rect 20805 9016 20810 9072
rect 20866 9016 21362 9072
rect 21418 9016 26802 9072
rect 20805 9014 26802 9016
rect 20805 9011 20871 9014
rect 21357 9011 21423 9014
rect 0 8938 480 8968
rect 1577 8938 1643 8941
rect 0 8936 1643 8938
rect 0 8880 1582 8936
rect 1638 8880 1643 8936
rect 0 8878 1643 8880
rect 0 8848 480 8878
rect 1577 8875 1643 8878
rect 5349 8938 5415 8941
rect 10869 8938 10935 8941
rect 5349 8936 10935 8938
rect 5349 8880 5354 8936
rect 5410 8880 10874 8936
rect 10930 8880 10935 8936
rect 5349 8878 10935 8880
rect 5349 8875 5415 8878
rect 10869 8875 10935 8878
rect 11329 8938 11395 8941
rect 16941 8938 17007 8941
rect 26742 8938 26802 9014
rect 26969 9072 30899 9074
rect 26969 9016 26974 9072
rect 27030 9016 30838 9072
rect 30894 9016 30899 9072
rect 26969 9014 30899 9016
rect 26969 9011 27035 9014
rect 30833 9011 30899 9014
rect 32673 9074 32739 9077
rect 36537 9074 36603 9077
rect 32673 9072 36603 9074
rect 32673 9016 32678 9072
rect 32734 9016 36542 9072
rect 36598 9016 36603 9072
rect 32673 9014 36603 9016
rect 36678 9074 36738 9150
rect 36813 9208 40000 9210
rect 36813 9152 36818 9208
rect 36874 9152 40000 9208
rect 36813 9150 40000 9152
rect 36813 9147 36879 9150
rect 39520 9120 40000 9150
rect 37365 9074 37431 9077
rect 36678 9072 37431 9074
rect 36678 9016 37370 9072
rect 37426 9016 37431 9072
rect 36678 9014 37431 9016
rect 32673 9011 32739 9014
rect 36537 9011 36603 9014
rect 37365 9011 37431 9014
rect 30741 8938 30807 8941
rect 11329 8936 17007 8938
rect 11329 8880 11334 8936
rect 11390 8880 16946 8936
rect 17002 8880 17007 8936
rect 11329 8878 17007 8880
rect 11329 8875 11395 8878
rect 16941 8875 17007 8878
rect 17174 8878 22018 8938
rect 26742 8936 30807 8938
rect 26742 8880 30746 8936
rect 30802 8880 30807 8936
rect 26742 8878 30807 8880
rect 8017 8802 8083 8805
rect 17174 8802 17234 8878
rect 8017 8800 17234 8802
rect 8017 8744 8022 8800
rect 8078 8744 17234 8800
rect 8017 8742 17234 8744
rect 8017 8739 8083 8742
rect 7610 8736 7930 8737
rect 7610 8672 7618 8736
rect 7682 8672 7698 8736
rect 7762 8672 7778 8736
rect 7842 8672 7858 8736
rect 7922 8672 7930 8736
rect 7610 8671 7930 8672
rect 20944 8736 21264 8737
rect 20944 8672 20952 8736
rect 21016 8672 21032 8736
rect 21096 8672 21112 8736
rect 21176 8672 21192 8736
rect 21256 8672 21264 8736
rect 20944 8671 21264 8672
rect 8477 8666 8543 8669
rect 10225 8666 10291 8669
rect 8477 8664 10291 8666
rect 8477 8608 8482 8664
rect 8538 8608 10230 8664
rect 10286 8608 10291 8664
rect 8477 8606 10291 8608
rect 8477 8603 8543 8606
rect 10225 8603 10291 8606
rect 11697 8666 11763 8669
rect 18413 8666 18479 8669
rect 11697 8664 18479 8666
rect 11697 8608 11702 8664
rect 11758 8608 18418 8664
rect 18474 8608 18479 8664
rect 11697 8606 18479 8608
rect 21958 8666 22018 8878
rect 30741 8875 30807 8878
rect 34053 8802 34119 8805
rect 22142 8800 34119 8802
rect 22142 8744 34058 8800
rect 34114 8744 34119 8800
rect 22142 8742 34119 8744
rect 22142 8666 22202 8742
rect 34053 8739 34119 8742
rect 36905 8802 36971 8805
rect 39520 8802 40000 8832
rect 36905 8800 40000 8802
rect 36905 8744 36910 8800
rect 36966 8744 40000 8800
rect 36905 8742 40000 8744
rect 36905 8739 36971 8742
rect 34277 8736 34597 8737
rect 34277 8672 34285 8736
rect 34349 8672 34365 8736
rect 34429 8672 34445 8736
rect 34509 8672 34525 8736
rect 34589 8672 34597 8736
rect 39520 8712 40000 8742
rect 34277 8671 34597 8672
rect 21958 8606 22202 8666
rect 25957 8666 26023 8669
rect 32489 8666 32555 8669
rect 25957 8664 32555 8666
rect 25957 8608 25962 8664
rect 26018 8608 32494 8664
rect 32550 8608 32555 8664
rect 25957 8606 32555 8608
rect 11697 8603 11763 8606
rect 18413 8603 18479 8606
rect 25957 8603 26023 8606
rect 32489 8603 32555 8606
rect 35801 8666 35867 8669
rect 37273 8666 37339 8669
rect 35801 8664 37339 8666
rect 35801 8608 35806 8664
rect 35862 8608 37278 8664
rect 37334 8608 37339 8664
rect 35801 8606 37339 8608
rect 35801 8603 35867 8606
rect 37273 8603 37339 8606
rect 0 8530 480 8560
rect 2405 8530 2471 8533
rect 0 8528 2471 8530
rect 0 8472 2410 8528
rect 2466 8472 2471 8528
rect 0 8470 2471 8472
rect 0 8440 480 8470
rect 2405 8467 2471 8470
rect 5809 8530 5875 8533
rect 15745 8530 15811 8533
rect 30373 8530 30439 8533
rect 5809 8528 30439 8530
rect 5809 8472 5814 8528
rect 5870 8472 15750 8528
rect 15806 8472 30378 8528
rect 30434 8472 30439 8528
rect 5809 8470 30439 8472
rect 5809 8467 5875 8470
rect 15745 8467 15811 8470
rect 30373 8467 30439 8470
rect 31477 8530 31543 8533
rect 31477 8528 32506 8530
rect 31477 8472 31482 8528
rect 31538 8472 32506 8528
rect 31477 8470 32506 8472
rect 31477 8467 31543 8470
rect 3877 8394 3943 8397
rect 5533 8394 5599 8397
rect 3877 8392 5599 8394
rect 3877 8336 3882 8392
rect 3938 8336 5538 8392
rect 5594 8336 5599 8392
rect 3877 8334 5599 8336
rect 3877 8331 3943 8334
rect 5533 8331 5599 8334
rect 15142 8332 15148 8396
rect 15212 8394 15218 8396
rect 15285 8394 15351 8397
rect 15212 8392 15351 8394
rect 15212 8336 15290 8392
rect 15346 8336 15351 8392
rect 15212 8334 15351 8336
rect 15212 8332 15218 8334
rect 15285 8331 15351 8334
rect 17585 8394 17651 8397
rect 18229 8394 18295 8397
rect 21817 8394 21883 8397
rect 30649 8396 30715 8397
rect 17585 8392 21883 8394
rect 17585 8336 17590 8392
rect 17646 8336 18234 8392
rect 18290 8336 21822 8392
rect 21878 8336 21883 8392
rect 17585 8334 21883 8336
rect 17585 8331 17651 8334
rect 18229 8331 18295 8334
rect 21817 8331 21883 8334
rect 30598 8332 30604 8396
rect 30668 8394 30715 8396
rect 32446 8394 32506 8470
rect 32622 8468 32628 8532
rect 32692 8530 32698 8532
rect 32765 8530 32831 8533
rect 36261 8530 36327 8533
rect 32692 8528 32831 8530
rect 32692 8472 32770 8528
rect 32826 8472 32831 8528
rect 32692 8470 32831 8472
rect 32692 8468 32698 8470
rect 32765 8467 32831 8470
rect 35390 8528 36327 8530
rect 35390 8472 36266 8528
rect 36322 8472 36327 8528
rect 35390 8470 36327 8472
rect 35390 8394 35450 8470
rect 36261 8467 36327 8470
rect 30668 8392 30760 8394
rect 30710 8336 30760 8392
rect 30668 8334 30760 8336
rect 32446 8334 35450 8394
rect 35801 8394 35867 8397
rect 39520 8394 40000 8424
rect 35801 8392 40000 8394
rect 35801 8336 35806 8392
rect 35862 8336 40000 8392
rect 35801 8334 40000 8336
rect 30668 8332 30715 8334
rect 30649 8331 30715 8332
rect 35801 8331 35867 8334
rect 39520 8304 40000 8334
rect 0 8258 480 8288
rect 4245 8258 4311 8261
rect 0 8256 4311 8258
rect 0 8200 4250 8256
rect 4306 8200 4311 8256
rect 0 8198 4311 8200
rect 0 8168 480 8198
rect 4245 8195 4311 8198
rect 6177 8258 6243 8261
rect 7281 8258 7347 8261
rect 6177 8256 7347 8258
rect 6177 8200 6182 8256
rect 6238 8200 7286 8256
rect 7342 8200 7347 8256
rect 6177 8198 7347 8200
rect 6177 8195 6243 8198
rect 7281 8195 7347 8198
rect 7557 8258 7623 8261
rect 14089 8258 14155 8261
rect 7557 8256 14155 8258
rect 7557 8200 7562 8256
rect 7618 8200 14094 8256
rect 14150 8200 14155 8256
rect 7557 8198 14155 8200
rect 7557 8195 7623 8198
rect 14089 8195 14155 8198
rect 18597 8258 18663 8261
rect 21817 8258 21883 8261
rect 28165 8258 28231 8261
rect 30465 8258 30531 8261
rect 18597 8256 21883 8258
rect 18597 8200 18602 8256
rect 18658 8200 21822 8256
rect 21878 8200 21883 8256
rect 18597 8198 21883 8200
rect 18597 8195 18663 8198
rect 21817 8195 21883 8198
rect 28030 8256 30531 8258
rect 28030 8200 28170 8256
rect 28226 8200 30470 8256
rect 30526 8200 30531 8256
rect 28030 8198 30531 8200
rect 14277 8192 14597 8193
rect 14277 8128 14285 8192
rect 14349 8128 14365 8192
rect 14429 8128 14445 8192
rect 14509 8128 14525 8192
rect 14589 8128 14597 8192
rect 14277 8127 14597 8128
rect 27610 8192 27930 8193
rect 27610 8128 27618 8192
rect 27682 8128 27698 8192
rect 27762 8128 27778 8192
rect 27842 8128 27858 8192
rect 27922 8128 27930 8192
rect 27610 8127 27930 8128
rect 4337 8122 4403 8125
rect 14089 8122 14155 8125
rect 4337 8120 14155 8122
rect 4337 8064 4342 8120
rect 4398 8064 14094 8120
rect 14150 8064 14155 8120
rect 4337 8062 14155 8064
rect 4337 8059 4403 8062
rect 14089 8059 14155 8062
rect 16205 8122 16271 8125
rect 19517 8122 19583 8125
rect 27429 8122 27495 8125
rect 16205 8120 19583 8122
rect 16205 8064 16210 8120
rect 16266 8064 19522 8120
rect 19578 8064 19583 8120
rect 16205 8062 19583 8064
rect 16205 8059 16271 8062
rect 19517 8059 19583 8062
rect 22004 8120 27495 8122
rect 22004 8064 27434 8120
rect 27490 8064 27495 8120
rect 22004 8062 27495 8064
rect 13721 7986 13787 7989
rect 15653 7986 15719 7989
rect 22004 7986 22064 8062
rect 27429 8059 27495 8062
rect 13721 7984 15719 7986
rect 13721 7928 13726 7984
rect 13782 7928 15658 7984
rect 15714 7928 15719 7984
rect 13721 7926 15719 7928
rect 13721 7923 13787 7926
rect 15653 7923 15719 7926
rect 16990 7926 22064 7986
rect 25497 7986 25563 7989
rect 28030 7986 28090 8198
rect 28165 8195 28231 8198
rect 30465 8195 30531 8198
rect 25497 7984 28090 7986
rect 25497 7928 25502 7984
rect 25558 7928 28090 7984
rect 25497 7926 28090 7928
rect 32765 7986 32831 7989
rect 35985 7986 36051 7989
rect 32765 7984 36051 7986
rect 32765 7928 32770 7984
rect 32826 7928 35990 7984
rect 36046 7928 36051 7984
rect 32765 7926 36051 7928
rect 0 7850 480 7880
rect 7557 7850 7623 7853
rect 0 7848 7623 7850
rect 0 7792 7562 7848
rect 7618 7792 7623 7848
rect 0 7790 7623 7792
rect 0 7760 480 7790
rect 7557 7787 7623 7790
rect 8201 7850 8267 7853
rect 16990 7850 17050 7926
rect 25497 7923 25563 7926
rect 32765 7923 32831 7926
rect 35985 7923 36051 7926
rect 37549 7986 37615 7989
rect 39520 7986 40000 8016
rect 37549 7984 40000 7986
rect 37549 7928 37554 7984
rect 37610 7928 40000 7984
rect 37549 7926 40000 7928
rect 37549 7923 37615 7926
rect 39520 7896 40000 7926
rect 21817 7850 21883 7853
rect 26325 7850 26391 7853
rect 8201 7848 17050 7850
rect 8201 7792 8206 7848
rect 8262 7792 17050 7848
rect 8201 7790 17050 7792
rect 17174 7790 21466 7850
rect 8201 7787 8267 7790
rect 4337 7714 4403 7717
rect 6729 7714 6795 7717
rect 4337 7712 6795 7714
rect 4337 7656 4342 7712
rect 4398 7656 6734 7712
rect 6790 7656 6795 7712
rect 4337 7654 6795 7656
rect 4337 7651 4403 7654
rect 6729 7651 6795 7654
rect 11329 7714 11395 7717
rect 17174 7714 17234 7790
rect 11329 7712 17234 7714
rect 11329 7656 11334 7712
rect 11390 7656 17234 7712
rect 11329 7654 17234 7656
rect 18321 7714 18387 7717
rect 19241 7714 19307 7717
rect 20161 7714 20227 7717
rect 20805 7714 20871 7717
rect 18321 7712 19074 7714
rect 18321 7656 18326 7712
rect 18382 7656 19074 7712
rect 18321 7654 19074 7656
rect 11329 7651 11395 7654
rect 18321 7651 18387 7654
rect 7610 7648 7930 7649
rect 7610 7584 7618 7648
rect 7682 7584 7698 7648
rect 7762 7584 7778 7648
rect 7842 7584 7858 7648
rect 7922 7584 7930 7648
rect 7610 7583 7930 7584
rect 2589 7578 2655 7581
rect 6821 7578 6887 7581
rect 2589 7576 6887 7578
rect 2589 7520 2594 7576
rect 2650 7520 6826 7576
rect 6882 7520 6887 7576
rect 2589 7518 6887 7520
rect 2589 7515 2655 7518
rect 6821 7515 6887 7518
rect 8293 7578 8359 7581
rect 12157 7578 12223 7581
rect 8293 7576 12223 7578
rect 8293 7520 8298 7576
rect 8354 7520 12162 7576
rect 12218 7520 12223 7576
rect 8293 7518 12223 7520
rect 8293 7515 8359 7518
rect 12157 7515 12223 7518
rect 13353 7578 13419 7581
rect 18597 7578 18663 7581
rect 13353 7576 18663 7578
rect 13353 7520 13358 7576
rect 13414 7520 18602 7576
rect 18658 7520 18663 7576
rect 13353 7518 18663 7520
rect 19014 7578 19074 7654
rect 19241 7712 20871 7714
rect 19241 7656 19246 7712
rect 19302 7656 20166 7712
rect 20222 7656 20810 7712
rect 20866 7656 20871 7712
rect 19241 7654 20871 7656
rect 21406 7714 21466 7790
rect 21817 7848 26391 7850
rect 21817 7792 21822 7848
rect 21878 7792 26330 7848
rect 26386 7792 26391 7848
rect 21817 7790 26391 7792
rect 21817 7787 21883 7790
rect 26325 7787 26391 7790
rect 27061 7850 27127 7853
rect 28165 7850 28231 7853
rect 35249 7850 35315 7853
rect 27061 7848 35315 7850
rect 27061 7792 27066 7848
rect 27122 7792 28170 7848
rect 28226 7792 35254 7848
rect 35310 7792 35315 7848
rect 27061 7790 35315 7792
rect 27061 7787 27127 7790
rect 28165 7787 28231 7790
rect 35249 7787 35315 7790
rect 29085 7714 29151 7717
rect 21406 7712 29151 7714
rect 21406 7656 29090 7712
rect 29146 7656 29151 7712
rect 21406 7654 29151 7656
rect 19241 7651 19307 7654
rect 20161 7651 20227 7654
rect 20805 7651 20871 7654
rect 29085 7651 29151 7654
rect 20944 7648 21264 7649
rect 20944 7584 20952 7648
rect 21016 7584 21032 7648
rect 21096 7584 21112 7648
rect 21176 7584 21192 7648
rect 21256 7584 21264 7648
rect 20944 7583 21264 7584
rect 34277 7648 34597 7649
rect 34277 7584 34285 7648
rect 34349 7584 34365 7648
rect 34429 7584 34445 7648
rect 34509 7584 34525 7648
rect 34589 7584 34597 7648
rect 34277 7583 34597 7584
rect 20805 7578 20871 7581
rect 19014 7576 20871 7578
rect 19014 7520 20810 7576
rect 20866 7520 20871 7576
rect 19014 7518 20871 7520
rect 13353 7515 13419 7518
rect 18597 7515 18663 7518
rect 20805 7515 20871 7518
rect 28257 7578 28323 7581
rect 28441 7578 28507 7581
rect 34145 7578 34211 7581
rect 28257 7576 34211 7578
rect 28257 7520 28262 7576
rect 28318 7520 28446 7576
rect 28502 7520 34150 7576
rect 34206 7520 34211 7576
rect 28257 7518 34211 7520
rect 28257 7515 28323 7518
rect 28441 7515 28507 7518
rect 34145 7515 34211 7518
rect 35065 7578 35131 7581
rect 39520 7578 40000 7608
rect 35065 7576 40000 7578
rect 35065 7520 35070 7576
rect 35126 7520 40000 7576
rect 35065 7518 40000 7520
rect 35065 7515 35131 7518
rect 39520 7488 40000 7518
rect 0 7442 480 7472
rect 3918 7442 3924 7444
rect 0 7382 3924 7442
rect 0 7352 480 7382
rect 3918 7380 3924 7382
rect 3988 7380 3994 7444
rect 5441 7442 5507 7445
rect 9765 7442 9831 7445
rect 5441 7440 9831 7442
rect 5441 7384 5446 7440
rect 5502 7384 9770 7440
rect 9826 7384 9831 7440
rect 5441 7382 9831 7384
rect 5441 7379 5507 7382
rect 9765 7379 9831 7382
rect 14733 7442 14799 7445
rect 30005 7442 30071 7445
rect 14733 7440 30071 7442
rect 14733 7384 14738 7440
rect 14794 7384 30010 7440
rect 30066 7384 30071 7440
rect 14733 7382 30071 7384
rect 14733 7379 14799 7382
rect 30005 7379 30071 7382
rect 30741 7442 30807 7445
rect 30741 7440 35634 7442
rect 30741 7384 30746 7440
rect 30802 7384 35634 7440
rect 30741 7382 35634 7384
rect 30741 7379 30807 7382
rect 6361 7306 6427 7309
rect 26049 7306 26115 7309
rect 6361 7304 26115 7306
rect 6361 7248 6366 7304
rect 6422 7248 26054 7304
rect 26110 7248 26115 7304
rect 6361 7246 26115 7248
rect 6361 7243 6427 7246
rect 26049 7243 26115 7246
rect 27521 7306 27587 7309
rect 35157 7306 35223 7309
rect 27521 7304 35223 7306
rect 27521 7248 27526 7304
rect 27582 7248 35162 7304
rect 35218 7248 35223 7304
rect 27521 7246 35223 7248
rect 27521 7243 27587 7246
rect 35157 7243 35223 7246
rect 2998 7170 3004 7172
rect 1350 7110 3004 7170
rect 0 7034 480 7064
rect 1350 7034 1410 7110
rect 2998 7108 3004 7110
rect 3068 7108 3074 7172
rect 3141 7170 3207 7173
rect 6545 7170 6611 7173
rect 10133 7170 10199 7173
rect 3141 7168 10199 7170
rect 3141 7112 3146 7168
rect 3202 7112 6550 7168
rect 6606 7112 10138 7168
rect 10194 7112 10199 7168
rect 3141 7110 10199 7112
rect 3141 7107 3207 7110
rect 6545 7107 6611 7110
rect 10133 7107 10199 7110
rect 14733 7170 14799 7173
rect 16941 7170 17007 7173
rect 19333 7172 19399 7173
rect 19333 7170 19380 7172
rect 14733 7168 17007 7170
rect 14733 7112 14738 7168
rect 14794 7112 16946 7168
rect 17002 7112 17007 7168
rect 14733 7110 17007 7112
rect 19288 7168 19380 7170
rect 19288 7112 19338 7168
rect 19288 7110 19380 7112
rect 14733 7107 14799 7110
rect 16941 7107 17007 7110
rect 19333 7108 19380 7110
rect 19444 7108 19450 7172
rect 19793 7170 19859 7173
rect 25681 7170 25747 7173
rect 19793 7168 25747 7170
rect 19793 7112 19798 7168
rect 19854 7112 25686 7168
rect 25742 7112 25747 7168
rect 19793 7110 25747 7112
rect 19333 7107 19399 7108
rect 19793 7107 19859 7110
rect 25681 7107 25747 7110
rect 29821 7170 29887 7173
rect 35433 7170 35499 7173
rect 29821 7168 35499 7170
rect 29821 7112 29826 7168
rect 29882 7112 35438 7168
rect 35494 7112 35499 7168
rect 29821 7110 35499 7112
rect 35574 7170 35634 7382
rect 39520 7170 40000 7200
rect 35574 7110 40000 7170
rect 29821 7107 29887 7110
rect 35433 7107 35499 7110
rect 14277 7104 14597 7105
rect 14277 7040 14285 7104
rect 14349 7040 14365 7104
rect 14429 7040 14445 7104
rect 14509 7040 14525 7104
rect 14589 7040 14597 7104
rect 14277 7039 14597 7040
rect 27610 7104 27930 7105
rect 27610 7040 27618 7104
rect 27682 7040 27698 7104
rect 27762 7040 27778 7104
rect 27842 7040 27858 7104
rect 27922 7040 27930 7104
rect 39520 7080 40000 7110
rect 27610 7039 27930 7040
rect 0 6974 1410 7034
rect 2773 7034 2839 7037
rect 3969 7034 4035 7037
rect 14089 7034 14155 7037
rect 2773 7032 14155 7034
rect 2773 6976 2778 7032
rect 2834 6976 3974 7032
rect 4030 6976 14094 7032
rect 14150 6976 14155 7032
rect 2773 6974 14155 6976
rect 0 6944 480 6974
rect 2773 6971 2839 6974
rect 3969 6971 4035 6974
rect 14089 6971 14155 6974
rect 19057 7034 19123 7037
rect 27061 7034 27127 7037
rect 19057 7032 27127 7034
rect 19057 6976 19062 7032
rect 19118 6976 27066 7032
rect 27122 6976 27127 7032
rect 19057 6974 27127 6976
rect 19057 6971 19123 6974
rect 27061 6971 27127 6974
rect 32857 7034 32923 7037
rect 33777 7034 33843 7037
rect 32857 7032 33843 7034
rect 32857 6976 32862 7032
rect 32918 6976 33782 7032
rect 33838 6976 33843 7032
rect 32857 6974 33843 6976
rect 32857 6971 32923 6974
rect 33777 6971 33843 6974
rect 35157 7034 35223 7037
rect 35893 7034 35959 7037
rect 35157 7032 35959 7034
rect 35157 6976 35162 7032
rect 35218 6976 35898 7032
rect 35954 6976 35959 7032
rect 35157 6974 35959 6976
rect 35157 6971 35223 6974
rect 35893 6971 35959 6974
rect 3141 6898 3207 6901
rect 9673 6898 9739 6901
rect 11053 6898 11119 6901
rect 13813 6898 13879 6901
rect 3141 6896 9874 6898
rect 3141 6840 3146 6896
rect 3202 6840 9678 6896
rect 9734 6840 9874 6896
rect 3141 6838 9874 6840
rect 3141 6835 3207 6838
rect 9673 6835 9739 6838
rect 3601 6762 3667 6765
rect 7557 6762 7623 6765
rect 3601 6760 7623 6762
rect 3601 6704 3606 6760
rect 3662 6704 7562 6760
rect 7618 6704 7623 6760
rect 3601 6702 7623 6704
rect 3601 6699 3667 6702
rect 7557 6699 7623 6702
rect 0 6626 480 6656
rect 4981 6626 5047 6629
rect 0 6624 5047 6626
rect 0 6568 4986 6624
rect 5042 6568 5047 6624
rect 0 6566 5047 6568
rect 0 6536 480 6566
rect 4981 6563 5047 6566
rect 7610 6560 7930 6561
rect 7610 6496 7618 6560
rect 7682 6496 7698 6560
rect 7762 6496 7778 6560
rect 7842 6496 7858 6560
rect 7922 6496 7930 6560
rect 7610 6495 7930 6496
rect 9814 6490 9874 6838
rect 11053 6896 13879 6898
rect 11053 6840 11058 6896
rect 11114 6840 13818 6896
rect 13874 6840 13879 6896
rect 11053 6838 13879 6840
rect 11053 6835 11119 6838
rect 13813 6835 13879 6838
rect 16205 6898 16271 6901
rect 24485 6898 24551 6901
rect 31385 6898 31451 6901
rect 35249 6898 35315 6901
rect 16205 6896 24410 6898
rect 16205 6840 16210 6896
rect 16266 6840 24410 6896
rect 16205 6838 24410 6840
rect 16205 6835 16271 6838
rect 10501 6762 10567 6765
rect 24025 6762 24091 6765
rect 10501 6760 24091 6762
rect 10501 6704 10506 6760
rect 10562 6704 24030 6760
rect 24086 6704 24091 6760
rect 10501 6702 24091 6704
rect 24350 6762 24410 6838
rect 24485 6896 31451 6898
rect 24485 6840 24490 6896
rect 24546 6840 31390 6896
rect 31446 6840 31451 6896
rect 24485 6838 31451 6840
rect 24485 6835 24551 6838
rect 31385 6835 31451 6838
rect 33918 6896 35315 6898
rect 33918 6840 35254 6896
rect 35310 6840 35315 6896
rect 33918 6838 35315 6840
rect 25773 6762 25839 6765
rect 24350 6760 25839 6762
rect 24350 6704 25778 6760
rect 25834 6704 25839 6760
rect 24350 6702 25839 6704
rect 10501 6699 10567 6702
rect 24025 6699 24091 6702
rect 25773 6699 25839 6702
rect 27337 6762 27403 6765
rect 33918 6762 33978 6838
rect 35249 6835 35315 6838
rect 35801 6898 35867 6901
rect 36077 6898 36143 6901
rect 35801 6896 36143 6898
rect 35801 6840 35806 6896
rect 35862 6840 36082 6896
rect 36138 6840 36143 6896
rect 35801 6838 36143 6840
rect 35801 6835 35867 6838
rect 36077 6835 36143 6838
rect 27337 6760 33978 6762
rect 27337 6704 27342 6760
rect 27398 6704 33978 6760
rect 27337 6702 33978 6704
rect 34053 6762 34119 6765
rect 39520 6762 40000 6792
rect 34053 6760 40000 6762
rect 34053 6704 34058 6760
rect 34114 6704 40000 6760
rect 34053 6702 40000 6704
rect 27337 6699 27403 6702
rect 34053 6699 34119 6702
rect 39520 6672 40000 6702
rect 12801 6626 12867 6629
rect 16297 6626 16363 6629
rect 12801 6624 16363 6626
rect 12801 6568 12806 6624
rect 12862 6568 16302 6624
rect 16358 6568 16363 6624
rect 12801 6566 16363 6568
rect 12801 6563 12867 6566
rect 16297 6563 16363 6566
rect 28901 6626 28967 6629
rect 28901 6624 34162 6626
rect 28901 6568 28906 6624
rect 28962 6568 34162 6624
rect 28901 6566 34162 6568
rect 28901 6563 28967 6566
rect 20944 6560 21264 6561
rect 20944 6496 20952 6560
rect 21016 6496 21032 6560
rect 21096 6496 21112 6560
rect 21176 6496 21192 6560
rect 21256 6496 21264 6560
rect 20944 6495 21264 6496
rect 17309 6490 17375 6493
rect 9814 6488 17375 6490
rect 9814 6432 17314 6488
rect 17370 6432 17375 6488
rect 9814 6430 17375 6432
rect 17309 6427 17375 6430
rect 26417 6490 26483 6493
rect 31293 6490 31359 6493
rect 26417 6488 31359 6490
rect 26417 6432 26422 6488
rect 26478 6432 31298 6488
rect 31354 6432 31359 6488
rect 26417 6430 31359 6432
rect 26417 6427 26483 6430
rect 31293 6427 31359 6430
rect 12525 6354 12591 6357
rect 13537 6354 13603 6357
rect 12525 6352 13603 6354
rect 12525 6296 12530 6352
rect 12586 6296 13542 6352
rect 13598 6296 13603 6352
rect 12525 6294 13603 6296
rect 12525 6291 12591 6294
rect 13537 6291 13603 6294
rect 28901 6354 28967 6357
rect 29821 6354 29887 6357
rect 28901 6352 29887 6354
rect 28901 6296 28906 6352
rect 28962 6296 29826 6352
rect 29882 6296 29887 6352
rect 28901 6294 29887 6296
rect 28901 6291 28967 6294
rect 29821 6291 29887 6294
rect 0 6218 480 6248
rect 9673 6218 9739 6221
rect 0 6216 9739 6218
rect 0 6160 9678 6216
rect 9734 6160 9739 6216
rect 0 6158 9739 6160
rect 0 6128 480 6158
rect 9673 6155 9739 6158
rect 10593 6218 10659 6221
rect 18965 6218 19031 6221
rect 10593 6216 19031 6218
rect 10593 6160 10598 6216
rect 10654 6160 18970 6216
rect 19026 6160 19031 6216
rect 10593 6158 19031 6160
rect 10593 6155 10659 6158
rect 18965 6155 19031 6158
rect 24669 6218 24735 6221
rect 24669 6216 28090 6218
rect 24669 6160 24674 6216
rect 24730 6160 28090 6216
rect 24669 6158 28090 6160
rect 24669 6155 24735 6158
rect 3233 6082 3299 6085
rect 6177 6082 6243 6085
rect 3233 6080 6243 6082
rect 3233 6024 3238 6080
rect 3294 6024 6182 6080
rect 6238 6024 6243 6080
rect 3233 6022 6243 6024
rect 3233 6019 3299 6022
rect 6177 6019 6243 6022
rect 7281 6082 7347 6085
rect 23473 6082 23539 6085
rect 7281 6080 12266 6082
rect 7281 6024 7286 6080
rect 7342 6024 12266 6080
rect 7281 6022 12266 6024
rect 7281 6019 7347 6022
rect 7649 5946 7715 5949
rect 10501 5946 10567 5949
rect 7649 5944 10567 5946
rect 7649 5888 7654 5944
rect 7710 5888 10506 5944
rect 10562 5888 10567 5944
rect 7649 5886 10567 5888
rect 12206 5946 12266 6022
rect 18830 6080 23539 6082
rect 18830 6024 23478 6080
rect 23534 6024 23539 6080
rect 18830 6022 23539 6024
rect 28030 6082 28090 6158
rect 33777 6082 33843 6085
rect 28030 6080 33843 6082
rect 28030 6024 33782 6080
rect 33838 6024 33843 6080
rect 28030 6022 33843 6024
rect 34102 6082 34162 6566
rect 34277 6560 34597 6561
rect 34277 6496 34285 6560
rect 34349 6496 34365 6560
rect 34429 6496 34445 6560
rect 34509 6496 34525 6560
rect 34589 6496 34597 6560
rect 34277 6495 34597 6496
rect 35065 6490 35131 6493
rect 39520 6490 40000 6520
rect 35065 6488 40000 6490
rect 35065 6432 35070 6488
rect 35126 6432 40000 6488
rect 35065 6430 40000 6432
rect 35065 6427 35131 6430
rect 39520 6400 40000 6430
rect 39520 6082 40000 6112
rect 34102 6022 40000 6082
rect 14277 6016 14597 6017
rect 14277 5952 14285 6016
rect 14349 5952 14365 6016
rect 14429 5952 14445 6016
rect 14509 5952 14525 6016
rect 14589 5952 14597 6016
rect 14277 5951 14597 5952
rect 18830 5949 18890 6022
rect 23473 6019 23539 6022
rect 33777 6019 33843 6022
rect 27610 6016 27930 6017
rect 27610 5952 27618 6016
rect 27682 5952 27698 6016
rect 27762 5952 27778 6016
rect 27842 5952 27858 6016
rect 27922 5952 27930 6016
rect 39520 5992 40000 6022
rect 27610 5951 27930 5952
rect 16573 5946 16639 5949
rect 18781 5946 18890 5949
rect 12206 5886 12588 5946
rect 7649 5883 7715 5886
rect 10501 5883 10567 5886
rect 0 5810 480 5840
rect 3969 5810 4035 5813
rect 6269 5812 6335 5813
rect 6269 5810 6316 5812
rect 0 5808 4035 5810
rect 0 5752 3974 5808
rect 4030 5752 4035 5808
rect 0 5750 4035 5752
rect 6224 5808 6316 5810
rect 6224 5752 6274 5808
rect 6224 5750 6316 5752
rect 0 5720 480 5750
rect 3969 5747 4035 5750
rect 6269 5748 6316 5750
rect 6380 5748 6386 5812
rect 8201 5810 8267 5813
rect 9949 5810 10015 5813
rect 8201 5808 10015 5810
rect 8201 5752 8206 5808
rect 8262 5752 9954 5808
rect 10010 5752 10015 5808
rect 8201 5750 10015 5752
rect 12528 5810 12588 5886
rect 16573 5944 18890 5946
rect 16573 5888 16578 5944
rect 16634 5888 18786 5944
rect 18842 5888 18890 5944
rect 16573 5886 18890 5888
rect 16573 5883 16639 5886
rect 18781 5883 18847 5886
rect 19374 5884 19380 5948
rect 19444 5946 19450 5948
rect 19517 5946 19583 5949
rect 19444 5944 19583 5946
rect 19444 5888 19522 5944
rect 19578 5888 19583 5944
rect 19444 5886 19583 5888
rect 19444 5884 19450 5886
rect 19517 5883 19583 5886
rect 21725 5946 21791 5949
rect 24209 5946 24275 5949
rect 21725 5944 24275 5946
rect 21725 5888 21730 5944
rect 21786 5888 24214 5944
rect 24270 5888 24275 5944
rect 21725 5886 24275 5888
rect 21725 5883 21791 5886
rect 24209 5883 24275 5886
rect 32581 5946 32647 5949
rect 36445 5946 36511 5949
rect 32581 5944 36511 5946
rect 32581 5888 32586 5944
rect 32642 5888 36450 5944
rect 36506 5888 36511 5944
rect 32581 5886 36511 5888
rect 32581 5883 32647 5886
rect 36445 5883 36511 5886
rect 27337 5810 27403 5813
rect 35065 5810 35131 5813
rect 12528 5808 35131 5810
rect 12528 5752 27342 5808
rect 27398 5752 35070 5808
rect 35126 5752 35131 5808
rect 12528 5750 35131 5752
rect 6269 5747 6335 5748
rect 8201 5747 8267 5750
rect 9949 5747 10015 5750
rect 27337 5747 27403 5750
rect 35065 5747 35131 5750
rect 10041 5674 10107 5677
rect 16573 5674 16639 5677
rect 10041 5672 16639 5674
rect 10041 5616 10046 5672
rect 10102 5616 16578 5672
rect 16634 5616 16639 5672
rect 10041 5614 16639 5616
rect 10041 5611 10107 5614
rect 16573 5611 16639 5614
rect 17309 5674 17375 5677
rect 18965 5674 19031 5677
rect 23105 5674 23171 5677
rect 28441 5674 28507 5677
rect 17309 5672 28507 5674
rect 17309 5616 17314 5672
rect 17370 5616 18970 5672
rect 19026 5616 23110 5672
rect 23166 5616 28446 5672
rect 28502 5616 28507 5672
rect 17309 5614 28507 5616
rect 17309 5611 17375 5614
rect 18965 5611 19031 5614
rect 23105 5611 23171 5614
rect 28441 5611 28507 5614
rect 28625 5674 28691 5677
rect 29177 5674 29243 5677
rect 28625 5672 29243 5674
rect 28625 5616 28630 5672
rect 28686 5616 29182 5672
rect 29238 5616 29243 5672
rect 28625 5614 29243 5616
rect 28625 5611 28691 5614
rect 29177 5611 29243 5614
rect 29361 5674 29427 5677
rect 32673 5674 32739 5677
rect 29361 5672 32739 5674
rect 29361 5616 29366 5672
rect 29422 5616 32678 5672
rect 32734 5616 32739 5672
rect 29361 5614 32739 5616
rect 29361 5611 29427 5614
rect 32673 5611 32739 5614
rect 35433 5674 35499 5677
rect 39520 5674 40000 5704
rect 35433 5672 40000 5674
rect 35433 5616 35438 5672
rect 35494 5616 40000 5672
rect 35433 5614 40000 5616
rect 35433 5611 35499 5614
rect 39520 5584 40000 5614
rect 8293 5538 8359 5541
rect 10317 5538 10383 5541
rect 13445 5538 13511 5541
rect 16849 5538 16915 5541
rect 8293 5536 10383 5538
rect 8293 5480 8298 5536
rect 8354 5480 10322 5536
rect 10378 5480 10383 5536
rect 8293 5478 10383 5480
rect 8293 5475 8359 5478
rect 10317 5475 10383 5478
rect 10550 5478 13370 5538
rect 7610 5472 7930 5473
rect 0 5402 480 5432
rect 7610 5408 7618 5472
rect 7682 5408 7698 5472
rect 7762 5408 7778 5472
rect 7842 5408 7858 5472
rect 7922 5408 7930 5472
rect 7610 5407 7930 5408
rect 3918 5402 3924 5404
rect 0 5342 3924 5402
rect 0 5312 480 5342
rect 3918 5340 3924 5342
rect 3988 5340 3994 5404
rect 4061 5402 4127 5405
rect 7005 5402 7071 5405
rect 4061 5400 7071 5402
rect 4061 5344 4066 5400
rect 4122 5344 7010 5400
rect 7066 5344 7071 5400
rect 4061 5342 7071 5344
rect 4061 5339 4127 5342
rect 7005 5339 7071 5342
rect 8017 5402 8083 5405
rect 10550 5402 10610 5478
rect 8017 5400 10610 5402
rect 8017 5344 8022 5400
rect 8078 5344 10610 5400
rect 8017 5342 10610 5344
rect 10869 5402 10935 5405
rect 13169 5402 13235 5405
rect 10869 5400 13235 5402
rect 10869 5344 10874 5400
rect 10930 5344 13174 5400
rect 13230 5344 13235 5400
rect 10869 5342 13235 5344
rect 13310 5402 13370 5478
rect 13445 5536 16915 5538
rect 13445 5480 13450 5536
rect 13506 5480 16854 5536
rect 16910 5480 16915 5536
rect 13445 5478 16915 5480
rect 13445 5475 13511 5478
rect 16849 5475 16915 5478
rect 27153 5538 27219 5541
rect 28942 5538 28948 5540
rect 27153 5536 28948 5538
rect 27153 5480 27158 5536
rect 27214 5480 28948 5536
rect 27153 5478 28948 5480
rect 27153 5475 27219 5478
rect 28942 5476 28948 5478
rect 29012 5476 29018 5540
rect 20944 5472 21264 5473
rect 20944 5408 20952 5472
rect 21016 5408 21032 5472
rect 21096 5408 21112 5472
rect 21176 5408 21192 5472
rect 21256 5408 21264 5472
rect 20944 5407 21264 5408
rect 34277 5472 34597 5473
rect 34277 5408 34285 5472
rect 34349 5408 34365 5472
rect 34429 5408 34445 5472
rect 34509 5408 34525 5472
rect 34589 5408 34597 5472
rect 34277 5407 34597 5408
rect 20805 5402 20871 5405
rect 13310 5400 20871 5402
rect 13310 5344 20810 5400
rect 20866 5344 20871 5400
rect 13310 5342 20871 5344
rect 8017 5339 8083 5342
rect 10869 5339 10935 5342
rect 13169 5339 13235 5342
rect 20805 5339 20871 5342
rect 24117 5402 24183 5405
rect 28625 5402 28691 5405
rect 24117 5400 28691 5402
rect 24117 5344 24122 5400
rect 24178 5344 28630 5400
rect 28686 5344 28691 5400
rect 24117 5342 28691 5344
rect 24117 5339 24183 5342
rect 28625 5339 28691 5342
rect 16205 5266 16271 5269
rect 2776 5264 16271 5266
rect 2776 5208 16210 5264
rect 16266 5208 16271 5264
rect 2776 5206 16271 5208
rect 2776 5130 2836 5206
rect 16205 5203 16271 5206
rect 16573 5266 16639 5269
rect 19425 5266 19491 5269
rect 16573 5264 19491 5266
rect 16573 5208 16578 5264
rect 16634 5208 19430 5264
rect 19486 5208 19491 5264
rect 16573 5206 19491 5208
rect 16573 5203 16639 5206
rect 19425 5203 19491 5206
rect 28809 5266 28875 5269
rect 29545 5266 29611 5269
rect 39520 5266 40000 5296
rect 28809 5264 29611 5266
rect 28809 5208 28814 5264
rect 28870 5208 29550 5264
rect 29606 5208 29611 5264
rect 28809 5206 29611 5208
rect 28809 5203 28875 5206
rect 29545 5203 29611 5206
rect 36678 5206 40000 5266
rect 2684 5070 2836 5130
rect 3325 5130 3391 5133
rect 10041 5130 10107 5133
rect 3325 5128 10107 5130
rect 3325 5072 3330 5128
rect 3386 5072 10046 5128
rect 10102 5072 10107 5128
rect 3325 5070 10107 5072
rect 0 4994 480 5024
rect 2684 4994 2744 5070
rect 3325 5067 3391 5070
rect 10041 5067 10107 5070
rect 13169 5130 13235 5133
rect 18045 5130 18111 5133
rect 20529 5130 20595 5133
rect 13169 5128 20595 5130
rect 13169 5072 13174 5128
rect 13230 5072 18050 5128
rect 18106 5072 20534 5128
rect 20590 5072 20595 5128
rect 13169 5070 20595 5072
rect 13169 5067 13235 5070
rect 18045 5067 18111 5070
rect 20529 5067 20595 5070
rect 28942 5068 28948 5132
rect 29012 5130 29018 5132
rect 29269 5130 29335 5133
rect 29012 5128 29335 5130
rect 29012 5072 29274 5128
rect 29330 5072 29335 5128
rect 29012 5070 29335 5072
rect 29012 5068 29018 5070
rect 29269 5067 29335 5070
rect 33501 5130 33567 5133
rect 36678 5130 36738 5206
rect 39520 5176 40000 5206
rect 33501 5128 36738 5130
rect 33501 5072 33506 5128
rect 33562 5072 36738 5128
rect 33501 5070 36738 5072
rect 33501 5067 33567 5070
rect 0 4934 2744 4994
rect 3969 4994 4035 4997
rect 4705 4994 4771 4997
rect 8109 4994 8175 4997
rect 10869 4994 10935 4997
rect 3969 4992 10935 4994
rect 3969 4936 3974 4992
rect 4030 4936 4710 4992
rect 4766 4936 8114 4992
rect 8170 4936 10874 4992
rect 10930 4936 10935 4992
rect 3969 4934 10935 4936
rect 0 4904 480 4934
rect 3969 4931 4035 4934
rect 4705 4931 4771 4934
rect 8109 4931 8175 4934
rect 10869 4931 10935 4934
rect 15653 4994 15719 4997
rect 25589 4994 25655 4997
rect 15653 4992 25655 4994
rect 15653 4936 15658 4992
rect 15714 4936 25594 4992
rect 25650 4936 25655 4992
rect 15653 4934 25655 4936
rect 15653 4931 15719 4934
rect 25589 4931 25655 4934
rect 28349 4994 28415 4997
rect 33593 4994 33659 4997
rect 35065 4994 35131 4997
rect 28349 4992 35131 4994
rect 28349 4936 28354 4992
rect 28410 4936 33598 4992
rect 33654 4936 35070 4992
rect 35126 4936 35131 4992
rect 28349 4934 35131 4936
rect 28349 4931 28415 4934
rect 33593 4931 33659 4934
rect 35065 4931 35131 4934
rect 14277 4928 14597 4929
rect 14277 4864 14285 4928
rect 14349 4864 14365 4928
rect 14429 4864 14445 4928
rect 14509 4864 14525 4928
rect 14589 4864 14597 4928
rect 14277 4863 14597 4864
rect 27610 4928 27930 4929
rect 27610 4864 27618 4928
rect 27682 4864 27698 4928
rect 27762 4864 27778 4928
rect 27842 4864 27858 4928
rect 27922 4864 27930 4928
rect 27610 4863 27930 4864
rect 4061 4858 4127 4861
rect 10409 4858 10475 4861
rect 4061 4856 10475 4858
rect 4061 4800 4066 4856
rect 4122 4800 10414 4856
rect 10470 4800 10475 4856
rect 4061 4798 10475 4800
rect 4061 4795 4127 4798
rect 10409 4795 10475 4798
rect 10961 4858 11027 4861
rect 12801 4858 12867 4861
rect 39520 4858 40000 4888
rect 10961 4856 12867 4858
rect 10961 4800 10966 4856
rect 11022 4800 12806 4856
rect 12862 4800 12867 4856
rect 10961 4798 12867 4800
rect 10961 4795 11027 4798
rect 12801 4795 12867 4798
rect 35574 4798 40000 4858
rect 12065 4722 12131 4725
rect 14733 4722 14799 4725
rect 12065 4720 14799 4722
rect 12065 4664 12070 4720
rect 12126 4664 14738 4720
rect 14794 4664 14799 4720
rect 12065 4662 14799 4664
rect 12065 4659 12131 4662
rect 14733 4659 14799 4662
rect 17125 4722 17191 4725
rect 35433 4722 35499 4725
rect 17125 4720 35499 4722
rect 17125 4664 17130 4720
rect 17186 4664 35438 4720
rect 35494 4664 35499 4720
rect 17125 4662 35499 4664
rect 17125 4659 17191 4662
rect 35433 4659 35499 4662
rect 0 4586 480 4616
rect 3785 4586 3851 4589
rect 0 4584 3851 4586
rect 0 4528 3790 4584
rect 3846 4528 3851 4584
rect 0 4526 3851 4528
rect 0 4496 480 4526
rect 3785 4523 3851 4526
rect 5993 4586 6059 4589
rect 17217 4586 17283 4589
rect 5993 4584 17283 4586
rect 5993 4528 5998 4584
rect 6054 4528 17222 4584
rect 17278 4528 17283 4584
rect 5993 4526 17283 4528
rect 5993 4523 6059 4526
rect 17217 4523 17283 4526
rect 24945 4586 25011 4589
rect 35574 4586 35634 4798
rect 39520 4768 40000 4798
rect 24945 4584 35634 4586
rect 24945 4528 24950 4584
rect 25006 4528 35634 4584
rect 24945 4526 35634 4528
rect 24945 4523 25011 4526
rect 11145 4450 11211 4453
rect 11278 4450 11284 4452
rect 11145 4448 11284 4450
rect 11145 4392 11150 4448
rect 11206 4392 11284 4448
rect 11145 4390 11284 4392
rect 11145 4387 11211 4390
rect 11278 4388 11284 4390
rect 11348 4388 11354 4452
rect 23974 4388 23980 4452
rect 24044 4450 24050 4452
rect 24117 4450 24183 4453
rect 24044 4448 24183 4450
rect 24044 4392 24122 4448
rect 24178 4392 24183 4448
rect 24044 4390 24183 4392
rect 24044 4388 24050 4390
rect 24117 4387 24183 4390
rect 36353 4450 36419 4453
rect 39520 4450 40000 4480
rect 36353 4448 40000 4450
rect 36353 4392 36358 4448
rect 36414 4392 40000 4448
rect 36353 4390 40000 4392
rect 36353 4387 36419 4390
rect 7610 4384 7930 4385
rect 7610 4320 7618 4384
rect 7682 4320 7698 4384
rect 7762 4320 7778 4384
rect 7842 4320 7858 4384
rect 7922 4320 7930 4384
rect 7610 4319 7930 4320
rect 20944 4384 21264 4385
rect 20944 4320 20952 4384
rect 21016 4320 21032 4384
rect 21096 4320 21112 4384
rect 21176 4320 21192 4384
rect 21256 4320 21264 4384
rect 20944 4319 21264 4320
rect 34277 4384 34597 4385
rect 34277 4320 34285 4384
rect 34349 4320 34365 4384
rect 34429 4320 34445 4384
rect 34509 4320 34525 4384
rect 34589 4320 34597 4384
rect 39520 4360 40000 4390
rect 34277 4319 34597 4320
rect 4521 4314 4587 4317
rect 2086 4312 4587 4314
rect 2086 4256 4526 4312
rect 4582 4256 4587 4312
rect 2086 4254 4587 4256
rect 0 4178 480 4208
rect 2086 4178 2146 4254
rect 4521 4251 4587 4254
rect 8150 4252 8156 4316
rect 8220 4314 8226 4316
rect 11421 4314 11487 4317
rect 15745 4314 15811 4317
rect 8220 4254 9506 4314
rect 8220 4252 8226 4254
rect 0 4118 2146 4178
rect 2313 4178 2379 4181
rect 9305 4178 9371 4181
rect 2313 4176 9371 4178
rect 2313 4120 2318 4176
rect 2374 4120 9310 4176
rect 9366 4120 9371 4176
rect 2313 4118 9371 4120
rect 9446 4178 9506 4254
rect 11421 4312 15811 4314
rect 11421 4256 11426 4312
rect 11482 4256 15750 4312
rect 15806 4256 15811 4312
rect 11421 4254 15811 4256
rect 11421 4251 11487 4254
rect 15745 4251 15811 4254
rect 12525 4178 12591 4181
rect 9446 4176 12591 4178
rect 9446 4120 12530 4176
rect 12586 4120 12591 4176
rect 9446 4118 12591 4120
rect 0 4088 480 4118
rect 2313 4115 2379 4118
rect 9305 4115 9371 4118
rect 12525 4115 12591 4118
rect 2037 4042 2103 4045
rect 6453 4042 6519 4045
rect 2037 4040 6519 4042
rect 2037 3984 2042 4040
rect 2098 3984 6458 4040
rect 6514 3984 6519 4040
rect 2037 3982 6519 3984
rect 2037 3979 2103 3982
rect 6453 3979 6519 3982
rect 11053 4042 11119 4045
rect 14641 4042 14707 4045
rect 11053 4040 14707 4042
rect 11053 3984 11058 4040
rect 11114 3984 14646 4040
rect 14702 3984 14707 4040
rect 11053 3982 14707 3984
rect 11053 3979 11119 3982
rect 14641 3979 14707 3982
rect 27521 4042 27587 4045
rect 31477 4042 31543 4045
rect 27521 4040 31543 4042
rect 27521 3984 27526 4040
rect 27582 3984 31482 4040
rect 31538 3984 31543 4040
rect 27521 3982 31543 3984
rect 27521 3979 27587 3982
rect 31477 3979 31543 3982
rect 32213 4042 32279 4045
rect 39520 4042 40000 4072
rect 32213 4040 40000 4042
rect 32213 3984 32218 4040
rect 32274 3984 40000 4040
rect 32213 3982 40000 3984
rect 32213 3979 32279 3982
rect 39520 3952 40000 3982
rect 5901 3906 5967 3909
rect 12157 3906 12223 3909
rect 37365 3906 37431 3909
rect 5901 3904 12223 3906
rect 5901 3848 5906 3904
rect 5962 3848 12162 3904
rect 12218 3848 12223 3904
rect 5901 3846 12223 3848
rect 5901 3843 5967 3846
rect 12157 3843 12223 3846
rect 28030 3904 37431 3906
rect 28030 3848 37370 3904
rect 37426 3848 37431 3904
rect 28030 3846 37431 3848
rect 14277 3840 14597 3841
rect 0 3770 480 3800
rect 14277 3776 14285 3840
rect 14349 3776 14365 3840
rect 14429 3776 14445 3840
rect 14509 3776 14525 3840
rect 14589 3776 14597 3840
rect 14277 3775 14597 3776
rect 27610 3840 27930 3841
rect 27610 3776 27618 3840
rect 27682 3776 27698 3840
rect 27762 3776 27778 3840
rect 27842 3776 27858 3840
rect 27922 3776 27930 3840
rect 27610 3775 27930 3776
rect 565 3770 631 3773
rect 0 3768 631 3770
rect 0 3712 570 3768
rect 626 3712 631 3768
rect 0 3710 631 3712
rect 0 3680 480 3710
rect 565 3707 631 3710
rect 1393 3634 1459 3637
rect 10593 3634 10659 3637
rect 1393 3632 10659 3634
rect 1393 3576 1398 3632
rect 1454 3576 10598 3632
rect 10654 3576 10659 3632
rect 1393 3574 10659 3576
rect 1393 3571 1459 3574
rect 10593 3571 10659 3574
rect 11697 3634 11763 3637
rect 11830 3634 11836 3636
rect 11697 3632 11836 3634
rect 11697 3576 11702 3632
rect 11758 3576 11836 3632
rect 11697 3574 11836 3576
rect 11697 3571 11763 3574
rect 11830 3572 11836 3574
rect 11900 3572 11906 3636
rect 12985 3634 13051 3637
rect 28030 3634 28090 3846
rect 37365 3843 37431 3846
rect 30005 3770 30071 3773
rect 35433 3770 35499 3773
rect 30005 3768 35499 3770
rect 30005 3712 30010 3768
rect 30066 3712 35438 3768
rect 35494 3712 35499 3768
rect 30005 3710 35499 3712
rect 30005 3707 30071 3710
rect 35433 3707 35499 3710
rect 12985 3632 28090 3634
rect 12985 3576 12990 3632
rect 13046 3576 28090 3632
rect 12985 3574 28090 3576
rect 12985 3571 13051 3574
rect 35566 3572 35572 3636
rect 35636 3634 35642 3636
rect 39520 3634 40000 3664
rect 35636 3574 40000 3634
rect 35636 3572 35642 3574
rect 39520 3544 40000 3574
rect 11973 3498 12039 3501
rect 4846 3496 12039 3498
rect 4846 3440 11978 3496
rect 12034 3440 12039 3496
rect 4846 3438 12039 3440
rect 0 3362 480 3392
rect 0 3302 2698 3362
rect 0 3272 480 3302
rect 2638 3226 2698 3302
rect 4846 3226 4906 3438
rect 11973 3435 12039 3438
rect 39520 3362 40000 3392
rect 35390 3302 40000 3362
rect 7610 3296 7930 3297
rect 7610 3232 7618 3296
rect 7682 3232 7698 3296
rect 7762 3232 7778 3296
rect 7842 3232 7858 3296
rect 7922 3232 7930 3296
rect 7610 3231 7930 3232
rect 20944 3296 21264 3297
rect 20944 3232 20952 3296
rect 21016 3232 21032 3296
rect 21096 3232 21112 3296
rect 21176 3232 21192 3296
rect 21256 3232 21264 3296
rect 20944 3231 21264 3232
rect 34277 3296 34597 3297
rect 34277 3232 34285 3296
rect 34349 3232 34365 3296
rect 34429 3232 34445 3296
rect 34509 3232 34525 3296
rect 34589 3232 34597 3296
rect 34277 3231 34597 3232
rect 2638 3166 4906 3226
rect 21958 3166 22202 3226
rect 4889 3090 4955 3093
rect 12341 3090 12407 3093
rect 4889 3088 12407 3090
rect 4889 3032 4894 3088
rect 4950 3032 12346 3088
rect 12402 3032 12407 3088
rect 4889 3030 12407 3032
rect 4889 3027 4955 3030
rect 12341 3027 12407 3030
rect 0 2954 480 2984
rect 7465 2954 7531 2957
rect 0 2952 7531 2954
rect 0 2896 7470 2952
rect 7526 2896 7531 2952
rect 0 2894 7531 2896
rect 0 2864 480 2894
rect 7465 2891 7531 2894
rect 16941 2954 17007 2957
rect 21958 2954 22018 3166
rect 22142 3090 22202 3166
rect 35390 3090 35450 3302
rect 39520 3272 40000 3302
rect 22142 3030 35450 3090
rect 16941 2952 22018 2954
rect 16941 2896 16946 2952
rect 17002 2896 22018 2952
rect 16941 2894 22018 2896
rect 33777 2954 33843 2957
rect 39520 2954 40000 2984
rect 33777 2952 40000 2954
rect 33777 2896 33782 2952
rect 33838 2896 40000 2952
rect 33777 2894 40000 2896
rect 16941 2891 17007 2894
rect 33777 2891 33843 2894
rect 39520 2864 40000 2894
rect 4797 2818 4863 2821
rect 11605 2818 11671 2821
rect 4797 2816 11671 2818
rect 4797 2760 4802 2816
rect 4858 2760 11610 2816
rect 11666 2760 11671 2816
rect 4797 2758 11671 2760
rect 4797 2755 4863 2758
rect 11605 2755 11671 2758
rect 14277 2752 14597 2753
rect 14277 2688 14285 2752
rect 14349 2688 14365 2752
rect 14429 2688 14445 2752
rect 14509 2688 14525 2752
rect 14589 2688 14597 2752
rect 14277 2687 14597 2688
rect 27610 2752 27930 2753
rect 27610 2688 27618 2752
rect 27682 2688 27698 2752
rect 27762 2688 27778 2752
rect 27842 2688 27858 2752
rect 27922 2688 27930 2752
rect 27610 2687 27930 2688
rect 0 2546 480 2576
rect 6361 2546 6427 2549
rect 0 2544 6427 2546
rect 0 2488 6366 2544
rect 6422 2488 6427 2544
rect 0 2486 6427 2488
rect 0 2456 480 2486
rect 6361 2483 6427 2486
rect 27981 2546 28047 2549
rect 39520 2546 40000 2576
rect 27981 2544 40000 2546
rect 27981 2488 27986 2544
rect 28042 2488 40000 2544
rect 27981 2486 40000 2488
rect 27981 2483 28047 2486
rect 39520 2456 40000 2486
rect 7610 2208 7930 2209
rect 0 2138 480 2168
rect 7610 2144 7618 2208
rect 7682 2144 7698 2208
rect 7762 2144 7778 2208
rect 7842 2144 7858 2208
rect 7922 2144 7930 2208
rect 7610 2143 7930 2144
rect 20944 2208 21264 2209
rect 20944 2144 20952 2208
rect 21016 2144 21032 2208
rect 21096 2144 21112 2208
rect 21176 2144 21192 2208
rect 21256 2144 21264 2208
rect 20944 2143 21264 2144
rect 34277 2208 34597 2209
rect 34277 2144 34285 2208
rect 34349 2144 34365 2208
rect 34429 2144 34445 2208
rect 34509 2144 34525 2208
rect 34589 2144 34597 2208
rect 34277 2143 34597 2144
rect 4889 2138 4955 2141
rect 39520 2138 40000 2168
rect 0 2136 4955 2138
rect 0 2080 4894 2136
rect 4950 2080 4955 2136
rect 0 2078 4955 2080
rect 0 2048 480 2078
rect 4889 2075 4955 2078
rect 35574 2078 40000 2138
rect 12525 1866 12591 1869
rect 22001 1866 22067 1869
rect 35574 1866 35634 2078
rect 39520 2048 40000 2078
rect 12525 1864 22067 1866
rect 12525 1808 12530 1864
rect 12586 1808 22006 1864
rect 22062 1808 22067 1864
rect 12525 1806 22067 1808
rect 12525 1803 12591 1806
rect 22001 1803 22067 1806
rect 22142 1806 35634 1866
rect 0 1730 480 1760
rect 5901 1730 5967 1733
rect 0 1728 5967 1730
rect 0 1672 5906 1728
rect 5962 1672 5967 1728
rect 0 1670 5967 1672
rect 0 1640 480 1670
rect 5901 1667 5967 1670
rect 17401 1730 17467 1733
rect 22142 1730 22202 1806
rect 39520 1730 40000 1760
rect 17401 1728 22202 1730
rect 17401 1672 17406 1728
rect 17462 1672 22202 1728
rect 17401 1670 22202 1672
rect 35574 1670 40000 1730
rect 17401 1667 17467 1670
rect 22001 1458 22067 1461
rect 35574 1458 35634 1670
rect 39520 1640 40000 1670
rect 22001 1456 35634 1458
rect 22001 1400 22006 1456
rect 22062 1400 35634 1456
rect 22001 1398 35634 1400
rect 22001 1395 22067 1398
rect 0 1322 480 1352
rect 3417 1322 3483 1325
rect 0 1320 3483 1322
rect 0 1264 3422 1320
rect 3478 1264 3483 1320
rect 0 1262 3483 1264
rect 0 1232 480 1262
rect 3417 1259 3483 1262
rect 34881 1322 34947 1325
rect 39520 1322 40000 1352
rect 34881 1320 40000 1322
rect 34881 1264 34886 1320
rect 34942 1264 40000 1320
rect 34881 1262 40000 1264
rect 34881 1259 34947 1262
rect 39520 1232 40000 1262
rect 0 914 480 944
rect 3233 914 3299 917
rect 0 912 3299 914
rect 0 856 3238 912
rect 3294 856 3299 912
rect 0 854 3299 856
rect 0 824 480 854
rect 3233 851 3299 854
rect 35801 914 35867 917
rect 39520 914 40000 944
rect 35801 912 40000 914
rect 35801 856 35806 912
rect 35862 856 40000 912
rect 35801 854 40000 856
rect 35801 851 35867 854
rect 39520 824 40000 854
rect 0 506 480 536
rect 2957 506 3023 509
rect 0 504 3023 506
rect 0 448 2962 504
rect 3018 448 3023 504
rect 0 446 3023 448
rect 0 416 480 446
rect 2957 443 3023 446
rect 35065 506 35131 509
rect 39520 506 40000 536
rect 35065 504 40000 506
rect 35065 448 35070 504
rect 35126 448 40000 504
rect 35065 446 40000 448
rect 35065 443 35131 446
rect 39520 416 40000 446
rect 0 234 480 264
rect 3601 234 3667 237
rect 0 232 3667 234
rect 0 176 3606 232
rect 3662 176 3667 232
rect 0 174 3667 176
rect 0 144 480 174
rect 3601 171 3667 174
rect 35157 234 35223 237
rect 39520 234 40000 264
rect 35157 232 40000 234
rect 35157 176 35162 232
rect 35218 176 40000 232
rect 35157 174 40000 176
rect 35157 171 35223 174
rect 39520 144 40000 174
<< via3 >>
rect 14285 13628 14349 13632
rect 14285 13572 14289 13628
rect 14289 13572 14345 13628
rect 14345 13572 14349 13628
rect 14285 13568 14349 13572
rect 14365 13628 14429 13632
rect 14365 13572 14369 13628
rect 14369 13572 14425 13628
rect 14425 13572 14429 13628
rect 14365 13568 14429 13572
rect 14445 13628 14509 13632
rect 14445 13572 14449 13628
rect 14449 13572 14505 13628
rect 14505 13572 14509 13628
rect 14445 13568 14509 13572
rect 14525 13628 14589 13632
rect 14525 13572 14529 13628
rect 14529 13572 14585 13628
rect 14585 13572 14589 13628
rect 14525 13568 14589 13572
rect 27618 13628 27682 13632
rect 27618 13572 27622 13628
rect 27622 13572 27678 13628
rect 27678 13572 27682 13628
rect 27618 13568 27682 13572
rect 27698 13628 27762 13632
rect 27698 13572 27702 13628
rect 27702 13572 27758 13628
rect 27758 13572 27762 13628
rect 27698 13568 27762 13572
rect 27778 13628 27842 13632
rect 27778 13572 27782 13628
rect 27782 13572 27838 13628
rect 27838 13572 27842 13628
rect 27778 13568 27842 13572
rect 27858 13628 27922 13632
rect 27858 13572 27862 13628
rect 27862 13572 27918 13628
rect 27918 13572 27922 13628
rect 27858 13568 27922 13572
rect 7618 13084 7682 13088
rect 7618 13028 7622 13084
rect 7622 13028 7678 13084
rect 7678 13028 7682 13084
rect 7618 13024 7682 13028
rect 7698 13084 7762 13088
rect 7698 13028 7702 13084
rect 7702 13028 7758 13084
rect 7758 13028 7762 13084
rect 7698 13024 7762 13028
rect 7778 13084 7842 13088
rect 7778 13028 7782 13084
rect 7782 13028 7838 13084
rect 7838 13028 7842 13084
rect 7778 13024 7842 13028
rect 7858 13084 7922 13088
rect 7858 13028 7862 13084
rect 7862 13028 7918 13084
rect 7918 13028 7922 13084
rect 7858 13024 7922 13028
rect 20952 13084 21016 13088
rect 20952 13028 20956 13084
rect 20956 13028 21012 13084
rect 21012 13028 21016 13084
rect 20952 13024 21016 13028
rect 21032 13084 21096 13088
rect 21032 13028 21036 13084
rect 21036 13028 21092 13084
rect 21092 13028 21096 13084
rect 21032 13024 21096 13028
rect 21112 13084 21176 13088
rect 21112 13028 21116 13084
rect 21116 13028 21172 13084
rect 21172 13028 21176 13084
rect 21112 13024 21176 13028
rect 21192 13084 21256 13088
rect 21192 13028 21196 13084
rect 21196 13028 21252 13084
rect 21252 13028 21256 13084
rect 21192 13024 21256 13028
rect 34285 13084 34349 13088
rect 34285 13028 34289 13084
rect 34289 13028 34345 13084
rect 34345 13028 34349 13084
rect 34285 13024 34349 13028
rect 34365 13084 34429 13088
rect 34365 13028 34369 13084
rect 34369 13028 34425 13084
rect 34425 13028 34429 13084
rect 34365 13024 34429 13028
rect 34445 13084 34509 13088
rect 34445 13028 34449 13084
rect 34449 13028 34505 13084
rect 34505 13028 34509 13084
rect 34445 13024 34509 13028
rect 34525 13084 34589 13088
rect 34525 13028 34529 13084
rect 34529 13028 34585 13084
rect 34585 13028 34589 13084
rect 34525 13024 34589 13028
rect 24716 12608 24780 12612
rect 24716 12552 24766 12608
rect 24766 12552 24780 12608
rect 24716 12548 24780 12552
rect 14285 12540 14349 12544
rect 14285 12484 14289 12540
rect 14289 12484 14345 12540
rect 14345 12484 14349 12540
rect 14285 12480 14349 12484
rect 14365 12540 14429 12544
rect 14365 12484 14369 12540
rect 14369 12484 14425 12540
rect 14425 12484 14429 12540
rect 14365 12480 14429 12484
rect 14445 12540 14509 12544
rect 14445 12484 14449 12540
rect 14449 12484 14505 12540
rect 14505 12484 14509 12540
rect 14445 12480 14509 12484
rect 14525 12540 14589 12544
rect 14525 12484 14529 12540
rect 14529 12484 14585 12540
rect 14585 12484 14589 12540
rect 14525 12480 14589 12484
rect 27618 12540 27682 12544
rect 27618 12484 27622 12540
rect 27622 12484 27678 12540
rect 27678 12484 27682 12540
rect 27618 12480 27682 12484
rect 27698 12540 27762 12544
rect 27698 12484 27702 12540
rect 27702 12484 27758 12540
rect 27758 12484 27762 12540
rect 27698 12480 27762 12484
rect 27778 12540 27842 12544
rect 27778 12484 27782 12540
rect 27782 12484 27838 12540
rect 27838 12484 27842 12540
rect 27778 12480 27842 12484
rect 27858 12540 27922 12544
rect 27858 12484 27862 12540
rect 27862 12484 27918 12540
rect 27918 12484 27922 12540
rect 27858 12480 27922 12484
rect 7618 11996 7682 12000
rect 7618 11940 7622 11996
rect 7622 11940 7678 11996
rect 7678 11940 7682 11996
rect 7618 11936 7682 11940
rect 7698 11996 7762 12000
rect 7698 11940 7702 11996
rect 7702 11940 7758 11996
rect 7758 11940 7762 11996
rect 7698 11936 7762 11940
rect 7778 11996 7842 12000
rect 7778 11940 7782 11996
rect 7782 11940 7838 11996
rect 7838 11940 7842 11996
rect 7778 11936 7842 11940
rect 7858 11996 7922 12000
rect 7858 11940 7862 11996
rect 7862 11940 7918 11996
rect 7918 11940 7922 11996
rect 7858 11936 7922 11940
rect 20952 11996 21016 12000
rect 20952 11940 20956 11996
rect 20956 11940 21012 11996
rect 21012 11940 21016 11996
rect 20952 11936 21016 11940
rect 21032 11996 21096 12000
rect 21032 11940 21036 11996
rect 21036 11940 21092 11996
rect 21092 11940 21096 11996
rect 21032 11936 21096 11940
rect 21112 11996 21176 12000
rect 21112 11940 21116 11996
rect 21116 11940 21172 11996
rect 21172 11940 21176 11996
rect 21112 11936 21176 11940
rect 21192 11996 21256 12000
rect 21192 11940 21196 11996
rect 21196 11940 21252 11996
rect 21252 11940 21256 11996
rect 21192 11936 21256 11940
rect 34285 11996 34349 12000
rect 34285 11940 34289 11996
rect 34289 11940 34345 11996
rect 34345 11940 34349 11996
rect 34285 11936 34349 11940
rect 34365 11996 34429 12000
rect 34365 11940 34369 11996
rect 34369 11940 34425 11996
rect 34425 11940 34429 11996
rect 34365 11936 34429 11940
rect 34445 11996 34509 12000
rect 34445 11940 34449 11996
rect 34449 11940 34505 11996
rect 34505 11940 34509 11996
rect 34445 11936 34509 11940
rect 34525 11996 34589 12000
rect 34525 11940 34529 11996
rect 34529 11940 34585 11996
rect 34585 11940 34589 11996
rect 34525 11936 34589 11940
rect 3004 11460 3068 11524
rect 14285 11452 14349 11456
rect 14285 11396 14289 11452
rect 14289 11396 14345 11452
rect 14345 11396 14349 11452
rect 14285 11392 14349 11396
rect 14365 11452 14429 11456
rect 14365 11396 14369 11452
rect 14369 11396 14425 11452
rect 14425 11396 14429 11452
rect 14365 11392 14429 11396
rect 14445 11452 14509 11456
rect 14445 11396 14449 11452
rect 14449 11396 14505 11452
rect 14505 11396 14509 11452
rect 14445 11392 14509 11396
rect 14525 11452 14589 11456
rect 14525 11396 14529 11452
rect 14529 11396 14585 11452
rect 14585 11396 14589 11452
rect 14525 11392 14589 11396
rect 27618 11452 27682 11456
rect 27618 11396 27622 11452
rect 27622 11396 27678 11452
rect 27678 11396 27682 11452
rect 27618 11392 27682 11396
rect 27698 11452 27762 11456
rect 27698 11396 27702 11452
rect 27702 11396 27758 11452
rect 27758 11396 27762 11452
rect 27698 11392 27762 11396
rect 27778 11452 27842 11456
rect 27778 11396 27782 11452
rect 27782 11396 27838 11452
rect 27838 11396 27842 11452
rect 27778 11392 27842 11396
rect 27858 11452 27922 11456
rect 27858 11396 27862 11452
rect 27862 11396 27918 11452
rect 27918 11396 27922 11452
rect 27858 11392 27922 11396
rect 7618 10908 7682 10912
rect 7618 10852 7622 10908
rect 7622 10852 7678 10908
rect 7678 10852 7682 10908
rect 7618 10848 7682 10852
rect 7698 10908 7762 10912
rect 7698 10852 7702 10908
rect 7702 10852 7758 10908
rect 7758 10852 7762 10908
rect 7698 10848 7762 10852
rect 7778 10908 7842 10912
rect 7778 10852 7782 10908
rect 7782 10852 7838 10908
rect 7838 10852 7842 10908
rect 7778 10848 7842 10852
rect 7858 10908 7922 10912
rect 7858 10852 7862 10908
rect 7862 10852 7918 10908
rect 7918 10852 7922 10908
rect 7858 10848 7922 10852
rect 20952 10908 21016 10912
rect 20952 10852 20956 10908
rect 20956 10852 21012 10908
rect 21012 10852 21016 10908
rect 20952 10848 21016 10852
rect 21032 10908 21096 10912
rect 21032 10852 21036 10908
rect 21036 10852 21092 10908
rect 21092 10852 21096 10908
rect 21032 10848 21096 10852
rect 21112 10908 21176 10912
rect 21112 10852 21116 10908
rect 21116 10852 21172 10908
rect 21172 10852 21176 10908
rect 21112 10848 21176 10852
rect 21192 10908 21256 10912
rect 21192 10852 21196 10908
rect 21196 10852 21252 10908
rect 21252 10852 21256 10908
rect 21192 10848 21256 10852
rect 34285 10908 34349 10912
rect 34285 10852 34289 10908
rect 34289 10852 34345 10908
rect 34345 10852 34349 10908
rect 34285 10848 34349 10852
rect 34365 10908 34429 10912
rect 34365 10852 34369 10908
rect 34369 10852 34425 10908
rect 34425 10852 34429 10908
rect 34365 10848 34429 10852
rect 34445 10908 34509 10912
rect 34445 10852 34449 10908
rect 34449 10852 34505 10908
rect 34505 10852 34509 10908
rect 34445 10848 34509 10852
rect 34525 10908 34589 10912
rect 34525 10852 34529 10908
rect 34529 10852 34585 10908
rect 34585 10852 34589 10908
rect 34525 10848 34589 10852
rect 14285 10364 14349 10368
rect 14285 10308 14289 10364
rect 14289 10308 14345 10364
rect 14345 10308 14349 10364
rect 14285 10304 14349 10308
rect 14365 10364 14429 10368
rect 14365 10308 14369 10364
rect 14369 10308 14425 10364
rect 14425 10308 14429 10364
rect 14365 10304 14429 10308
rect 14445 10364 14509 10368
rect 14445 10308 14449 10364
rect 14449 10308 14505 10364
rect 14505 10308 14509 10364
rect 14445 10304 14509 10308
rect 14525 10364 14589 10368
rect 14525 10308 14529 10364
rect 14529 10308 14585 10364
rect 14585 10308 14589 10364
rect 14525 10304 14589 10308
rect 20668 10236 20732 10300
rect 27618 10364 27682 10368
rect 27618 10308 27622 10364
rect 27622 10308 27678 10364
rect 27678 10308 27682 10364
rect 27618 10304 27682 10308
rect 27698 10364 27762 10368
rect 27698 10308 27702 10364
rect 27702 10308 27758 10364
rect 27758 10308 27762 10364
rect 27698 10304 27762 10308
rect 27778 10364 27842 10368
rect 27778 10308 27782 10364
rect 27782 10308 27838 10364
rect 27838 10308 27842 10364
rect 27778 10304 27842 10308
rect 27858 10364 27922 10368
rect 27858 10308 27862 10364
rect 27862 10308 27918 10364
rect 27918 10308 27922 10364
rect 27858 10304 27922 10308
rect 7618 9820 7682 9824
rect 7618 9764 7622 9820
rect 7622 9764 7678 9820
rect 7678 9764 7682 9820
rect 7618 9760 7682 9764
rect 7698 9820 7762 9824
rect 7698 9764 7702 9820
rect 7702 9764 7758 9820
rect 7758 9764 7762 9820
rect 7698 9760 7762 9764
rect 7778 9820 7842 9824
rect 7778 9764 7782 9820
rect 7782 9764 7838 9820
rect 7838 9764 7842 9820
rect 7778 9760 7842 9764
rect 7858 9820 7922 9824
rect 7858 9764 7862 9820
rect 7862 9764 7918 9820
rect 7918 9764 7922 9820
rect 7858 9760 7922 9764
rect 20952 9820 21016 9824
rect 20952 9764 20956 9820
rect 20956 9764 21012 9820
rect 21012 9764 21016 9820
rect 20952 9760 21016 9764
rect 21032 9820 21096 9824
rect 21032 9764 21036 9820
rect 21036 9764 21092 9820
rect 21092 9764 21096 9820
rect 21032 9760 21096 9764
rect 21112 9820 21176 9824
rect 21112 9764 21116 9820
rect 21116 9764 21172 9820
rect 21172 9764 21176 9820
rect 21112 9760 21176 9764
rect 21192 9820 21256 9824
rect 21192 9764 21196 9820
rect 21196 9764 21252 9820
rect 21252 9764 21256 9820
rect 21192 9760 21256 9764
rect 34285 9820 34349 9824
rect 34285 9764 34289 9820
rect 34289 9764 34345 9820
rect 34345 9764 34349 9820
rect 34285 9760 34349 9764
rect 34365 9820 34429 9824
rect 34365 9764 34369 9820
rect 34369 9764 34425 9820
rect 34425 9764 34429 9820
rect 34365 9760 34429 9764
rect 34445 9820 34509 9824
rect 34445 9764 34449 9820
rect 34449 9764 34505 9820
rect 34505 9764 34509 9820
rect 34445 9760 34509 9764
rect 34525 9820 34589 9824
rect 34525 9764 34529 9820
rect 34529 9764 34585 9820
rect 34585 9764 34589 9820
rect 34525 9760 34589 9764
rect 8156 9284 8220 9348
rect 14285 9276 14349 9280
rect 14285 9220 14289 9276
rect 14289 9220 14345 9276
rect 14345 9220 14349 9276
rect 14285 9216 14349 9220
rect 14365 9276 14429 9280
rect 14365 9220 14369 9276
rect 14369 9220 14425 9276
rect 14425 9220 14429 9276
rect 14365 9216 14429 9220
rect 14445 9276 14509 9280
rect 14445 9220 14449 9276
rect 14449 9220 14505 9276
rect 14505 9220 14509 9276
rect 14445 9216 14509 9220
rect 14525 9276 14589 9280
rect 14525 9220 14529 9276
rect 14529 9220 14585 9276
rect 14585 9220 14589 9276
rect 14525 9216 14589 9220
rect 27618 9276 27682 9280
rect 27618 9220 27622 9276
rect 27622 9220 27678 9276
rect 27678 9220 27682 9276
rect 27618 9216 27682 9220
rect 27698 9276 27762 9280
rect 27698 9220 27702 9276
rect 27702 9220 27758 9276
rect 27758 9220 27762 9276
rect 27698 9216 27762 9220
rect 27778 9276 27842 9280
rect 27778 9220 27782 9276
rect 27782 9220 27838 9276
rect 27838 9220 27842 9276
rect 27778 9216 27842 9220
rect 27858 9276 27922 9280
rect 27858 9220 27862 9276
rect 27862 9220 27918 9276
rect 27918 9220 27922 9276
rect 27858 9216 27922 9220
rect 7618 8732 7682 8736
rect 7618 8676 7622 8732
rect 7622 8676 7678 8732
rect 7678 8676 7682 8732
rect 7618 8672 7682 8676
rect 7698 8732 7762 8736
rect 7698 8676 7702 8732
rect 7702 8676 7758 8732
rect 7758 8676 7762 8732
rect 7698 8672 7762 8676
rect 7778 8732 7842 8736
rect 7778 8676 7782 8732
rect 7782 8676 7838 8732
rect 7838 8676 7842 8732
rect 7778 8672 7842 8676
rect 7858 8732 7922 8736
rect 7858 8676 7862 8732
rect 7862 8676 7918 8732
rect 7918 8676 7922 8732
rect 7858 8672 7922 8676
rect 20952 8732 21016 8736
rect 20952 8676 20956 8732
rect 20956 8676 21012 8732
rect 21012 8676 21016 8732
rect 20952 8672 21016 8676
rect 21032 8732 21096 8736
rect 21032 8676 21036 8732
rect 21036 8676 21092 8732
rect 21092 8676 21096 8732
rect 21032 8672 21096 8676
rect 21112 8732 21176 8736
rect 21112 8676 21116 8732
rect 21116 8676 21172 8732
rect 21172 8676 21176 8732
rect 21112 8672 21176 8676
rect 21192 8732 21256 8736
rect 21192 8676 21196 8732
rect 21196 8676 21252 8732
rect 21252 8676 21256 8732
rect 21192 8672 21256 8676
rect 34285 8732 34349 8736
rect 34285 8676 34289 8732
rect 34289 8676 34345 8732
rect 34345 8676 34349 8732
rect 34285 8672 34349 8676
rect 34365 8732 34429 8736
rect 34365 8676 34369 8732
rect 34369 8676 34425 8732
rect 34425 8676 34429 8732
rect 34365 8672 34429 8676
rect 34445 8732 34509 8736
rect 34445 8676 34449 8732
rect 34449 8676 34505 8732
rect 34505 8676 34509 8732
rect 34445 8672 34509 8676
rect 34525 8732 34589 8736
rect 34525 8676 34529 8732
rect 34529 8676 34585 8732
rect 34585 8676 34589 8732
rect 34525 8672 34589 8676
rect 15148 8332 15212 8396
rect 30604 8392 30668 8396
rect 32628 8468 32692 8532
rect 30604 8336 30654 8392
rect 30654 8336 30668 8392
rect 30604 8332 30668 8336
rect 14285 8188 14349 8192
rect 14285 8132 14289 8188
rect 14289 8132 14345 8188
rect 14345 8132 14349 8188
rect 14285 8128 14349 8132
rect 14365 8188 14429 8192
rect 14365 8132 14369 8188
rect 14369 8132 14425 8188
rect 14425 8132 14429 8188
rect 14365 8128 14429 8132
rect 14445 8188 14509 8192
rect 14445 8132 14449 8188
rect 14449 8132 14505 8188
rect 14505 8132 14509 8188
rect 14445 8128 14509 8132
rect 14525 8188 14589 8192
rect 14525 8132 14529 8188
rect 14529 8132 14585 8188
rect 14585 8132 14589 8188
rect 14525 8128 14589 8132
rect 27618 8188 27682 8192
rect 27618 8132 27622 8188
rect 27622 8132 27678 8188
rect 27678 8132 27682 8188
rect 27618 8128 27682 8132
rect 27698 8188 27762 8192
rect 27698 8132 27702 8188
rect 27702 8132 27758 8188
rect 27758 8132 27762 8188
rect 27698 8128 27762 8132
rect 27778 8188 27842 8192
rect 27778 8132 27782 8188
rect 27782 8132 27838 8188
rect 27838 8132 27842 8188
rect 27778 8128 27842 8132
rect 27858 8188 27922 8192
rect 27858 8132 27862 8188
rect 27862 8132 27918 8188
rect 27918 8132 27922 8188
rect 27858 8128 27922 8132
rect 7618 7644 7682 7648
rect 7618 7588 7622 7644
rect 7622 7588 7678 7644
rect 7678 7588 7682 7644
rect 7618 7584 7682 7588
rect 7698 7644 7762 7648
rect 7698 7588 7702 7644
rect 7702 7588 7758 7644
rect 7758 7588 7762 7644
rect 7698 7584 7762 7588
rect 7778 7644 7842 7648
rect 7778 7588 7782 7644
rect 7782 7588 7838 7644
rect 7838 7588 7842 7644
rect 7778 7584 7842 7588
rect 7858 7644 7922 7648
rect 7858 7588 7862 7644
rect 7862 7588 7918 7644
rect 7918 7588 7922 7644
rect 7858 7584 7922 7588
rect 20952 7644 21016 7648
rect 20952 7588 20956 7644
rect 20956 7588 21012 7644
rect 21012 7588 21016 7644
rect 20952 7584 21016 7588
rect 21032 7644 21096 7648
rect 21032 7588 21036 7644
rect 21036 7588 21092 7644
rect 21092 7588 21096 7644
rect 21032 7584 21096 7588
rect 21112 7644 21176 7648
rect 21112 7588 21116 7644
rect 21116 7588 21172 7644
rect 21172 7588 21176 7644
rect 21112 7584 21176 7588
rect 21192 7644 21256 7648
rect 21192 7588 21196 7644
rect 21196 7588 21252 7644
rect 21252 7588 21256 7644
rect 21192 7584 21256 7588
rect 34285 7644 34349 7648
rect 34285 7588 34289 7644
rect 34289 7588 34345 7644
rect 34345 7588 34349 7644
rect 34285 7584 34349 7588
rect 34365 7644 34429 7648
rect 34365 7588 34369 7644
rect 34369 7588 34425 7644
rect 34425 7588 34429 7644
rect 34365 7584 34429 7588
rect 34445 7644 34509 7648
rect 34445 7588 34449 7644
rect 34449 7588 34505 7644
rect 34505 7588 34509 7644
rect 34445 7584 34509 7588
rect 34525 7644 34589 7648
rect 34525 7588 34529 7644
rect 34529 7588 34585 7644
rect 34585 7588 34589 7644
rect 34525 7584 34589 7588
rect 3924 7380 3988 7444
rect 3004 7108 3068 7172
rect 19380 7168 19444 7172
rect 19380 7112 19394 7168
rect 19394 7112 19444 7168
rect 19380 7108 19444 7112
rect 14285 7100 14349 7104
rect 14285 7044 14289 7100
rect 14289 7044 14345 7100
rect 14345 7044 14349 7100
rect 14285 7040 14349 7044
rect 14365 7100 14429 7104
rect 14365 7044 14369 7100
rect 14369 7044 14425 7100
rect 14425 7044 14429 7100
rect 14365 7040 14429 7044
rect 14445 7100 14509 7104
rect 14445 7044 14449 7100
rect 14449 7044 14505 7100
rect 14505 7044 14509 7100
rect 14445 7040 14509 7044
rect 14525 7100 14589 7104
rect 14525 7044 14529 7100
rect 14529 7044 14585 7100
rect 14585 7044 14589 7100
rect 14525 7040 14589 7044
rect 27618 7100 27682 7104
rect 27618 7044 27622 7100
rect 27622 7044 27678 7100
rect 27678 7044 27682 7100
rect 27618 7040 27682 7044
rect 27698 7100 27762 7104
rect 27698 7044 27702 7100
rect 27702 7044 27758 7100
rect 27758 7044 27762 7100
rect 27698 7040 27762 7044
rect 27778 7100 27842 7104
rect 27778 7044 27782 7100
rect 27782 7044 27838 7100
rect 27838 7044 27842 7100
rect 27778 7040 27842 7044
rect 27858 7100 27922 7104
rect 27858 7044 27862 7100
rect 27862 7044 27918 7100
rect 27918 7044 27922 7100
rect 27858 7040 27922 7044
rect 7618 6556 7682 6560
rect 7618 6500 7622 6556
rect 7622 6500 7678 6556
rect 7678 6500 7682 6556
rect 7618 6496 7682 6500
rect 7698 6556 7762 6560
rect 7698 6500 7702 6556
rect 7702 6500 7758 6556
rect 7758 6500 7762 6556
rect 7698 6496 7762 6500
rect 7778 6556 7842 6560
rect 7778 6500 7782 6556
rect 7782 6500 7838 6556
rect 7838 6500 7842 6556
rect 7778 6496 7842 6500
rect 7858 6556 7922 6560
rect 7858 6500 7862 6556
rect 7862 6500 7918 6556
rect 7918 6500 7922 6556
rect 7858 6496 7922 6500
rect 20952 6556 21016 6560
rect 20952 6500 20956 6556
rect 20956 6500 21012 6556
rect 21012 6500 21016 6556
rect 20952 6496 21016 6500
rect 21032 6556 21096 6560
rect 21032 6500 21036 6556
rect 21036 6500 21092 6556
rect 21092 6500 21096 6556
rect 21032 6496 21096 6500
rect 21112 6556 21176 6560
rect 21112 6500 21116 6556
rect 21116 6500 21172 6556
rect 21172 6500 21176 6556
rect 21112 6496 21176 6500
rect 21192 6556 21256 6560
rect 21192 6500 21196 6556
rect 21196 6500 21252 6556
rect 21252 6500 21256 6556
rect 21192 6496 21256 6500
rect 34285 6556 34349 6560
rect 34285 6500 34289 6556
rect 34289 6500 34345 6556
rect 34345 6500 34349 6556
rect 34285 6496 34349 6500
rect 34365 6556 34429 6560
rect 34365 6500 34369 6556
rect 34369 6500 34425 6556
rect 34425 6500 34429 6556
rect 34365 6496 34429 6500
rect 34445 6556 34509 6560
rect 34445 6500 34449 6556
rect 34449 6500 34505 6556
rect 34505 6500 34509 6556
rect 34445 6496 34509 6500
rect 34525 6556 34589 6560
rect 34525 6500 34529 6556
rect 34529 6500 34585 6556
rect 34585 6500 34589 6556
rect 34525 6496 34589 6500
rect 14285 6012 14349 6016
rect 14285 5956 14289 6012
rect 14289 5956 14345 6012
rect 14345 5956 14349 6012
rect 14285 5952 14349 5956
rect 14365 6012 14429 6016
rect 14365 5956 14369 6012
rect 14369 5956 14425 6012
rect 14425 5956 14429 6012
rect 14365 5952 14429 5956
rect 14445 6012 14509 6016
rect 14445 5956 14449 6012
rect 14449 5956 14505 6012
rect 14505 5956 14509 6012
rect 14445 5952 14509 5956
rect 14525 6012 14589 6016
rect 14525 5956 14529 6012
rect 14529 5956 14585 6012
rect 14585 5956 14589 6012
rect 14525 5952 14589 5956
rect 27618 6012 27682 6016
rect 27618 5956 27622 6012
rect 27622 5956 27678 6012
rect 27678 5956 27682 6012
rect 27618 5952 27682 5956
rect 27698 6012 27762 6016
rect 27698 5956 27702 6012
rect 27702 5956 27758 6012
rect 27758 5956 27762 6012
rect 27698 5952 27762 5956
rect 27778 6012 27842 6016
rect 27778 5956 27782 6012
rect 27782 5956 27838 6012
rect 27838 5956 27842 6012
rect 27778 5952 27842 5956
rect 27858 6012 27922 6016
rect 27858 5956 27862 6012
rect 27862 5956 27918 6012
rect 27918 5956 27922 6012
rect 27858 5952 27922 5956
rect 6316 5808 6380 5812
rect 6316 5752 6330 5808
rect 6330 5752 6380 5808
rect 6316 5748 6380 5752
rect 19380 5884 19444 5948
rect 7618 5468 7682 5472
rect 7618 5412 7622 5468
rect 7622 5412 7678 5468
rect 7678 5412 7682 5468
rect 7618 5408 7682 5412
rect 7698 5468 7762 5472
rect 7698 5412 7702 5468
rect 7702 5412 7758 5468
rect 7758 5412 7762 5468
rect 7698 5408 7762 5412
rect 7778 5468 7842 5472
rect 7778 5412 7782 5468
rect 7782 5412 7838 5468
rect 7838 5412 7842 5468
rect 7778 5408 7842 5412
rect 7858 5468 7922 5472
rect 7858 5412 7862 5468
rect 7862 5412 7918 5468
rect 7918 5412 7922 5468
rect 7858 5408 7922 5412
rect 3924 5340 3988 5404
rect 28948 5476 29012 5540
rect 20952 5468 21016 5472
rect 20952 5412 20956 5468
rect 20956 5412 21012 5468
rect 21012 5412 21016 5468
rect 20952 5408 21016 5412
rect 21032 5468 21096 5472
rect 21032 5412 21036 5468
rect 21036 5412 21092 5468
rect 21092 5412 21096 5468
rect 21032 5408 21096 5412
rect 21112 5468 21176 5472
rect 21112 5412 21116 5468
rect 21116 5412 21172 5468
rect 21172 5412 21176 5468
rect 21112 5408 21176 5412
rect 21192 5468 21256 5472
rect 21192 5412 21196 5468
rect 21196 5412 21252 5468
rect 21252 5412 21256 5468
rect 21192 5408 21256 5412
rect 34285 5468 34349 5472
rect 34285 5412 34289 5468
rect 34289 5412 34345 5468
rect 34345 5412 34349 5468
rect 34285 5408 34349 5412
rect 34365 5468 34429 5472
rect 34365 5412 34369 5468
rect 34369 5412 34425 5468
rect 34425 5412 34429 5468
rect 34365 5408 34429 5412
rect 34445 5468 34509 5472
rect 34445 5412 34449 5468
rect 34449 5412 34505 5468
rect 34505 5412 34509 5468
rect 34445 5408 34509 5412
rect 34525 5468 34589 5472
rect 34525 5412 34529 5468
rect 34529 5412 34585 5468
rect 34585 5412 34589 5468
rect 34525 5408 34589 5412
rect 28948 5068 29012 5132
rect 14285 4924 14349 4928
rect 14285 4868 14289 4924
rect 14289 4868 14345 4924
rect 14345 4868 14349 4924
rect 14285 4864 14349 4868
rect 14365 4924 14429 4928
rect 14365 4868 14369 4924
rect 14369 4868 14425 4924
rect 14425 4868 14429 4924
rect 14365 4864 14429 4868
rect 14445 4924 14509 4928
rect 14445 4868 14449 4924
rect 14449 4868 14505 4924
rect 14505 4868 14509 4924
rect 14445 4864 14509 4868
rect 14525 4924 14589 4928
rect 14525 4868 14529 4924
rect 14529 4868 14585 4924
rect 14585 4868 14589 4924
rect 14525 4864 14589 4868
rect 27618 4924 27682 4928
rect 27618 4868 27622 4924
rect 27622 4868 27678 4924
rect 27678 4868 27682 4924
rect 27618 4864 27682 4868
rect 27698 4924 27762 4928
rect 27698 4868 27702 4924
rect 27702 4868 27758 4924
rect 27758 4868 27762 4924
rect 27698 4864 27762 4868
rect 27778 4924 27842 4928
rect 27778 4868 27782 4924
rect 27782 4868 27838 4924
rect 27838 4868 27842 4924
rect 27778 4864 27842 4868
rect 27858 4924 27922 4928
rect 27858 4868 27862 4924
rect 27862 4868 27918 4924
rect 27918 4868 27922 4924
rect 27858 4864 27922 4868
rect 11284 4388 11348 4452
rect 23980 4388 24044 4452
rect 7618 4380 7682 4384
rect 7618 4324 7622 4380
rect 7622 4324 7678 4380
rect 7678 4324 7682 4380
rect 7618 4320 7682 4324
rect 7698 4380 7762 4384
rect 7698 4324 7702 4380
rect 7702 4324 7758 4380
rect 7758 4324 7762 4380
rect 7698 4320 7762 4324
rect 7778 4380 7842 4384
rect 7778 4324 7782 4380
rect 7782 4324 7838 4380
rect 7838 4324 7842 4380
rect 7778 4320 7842 4324
rect 7858 4380 7922 4384
rect 7858 4324 7862 4380
rect 7862 4324 7918 4380
rect 7918 4324 7922 4380
rect 7858 4320 7922 4324
rect 20952 4380 21016 4384
rect 20952 4324 20956 4380
rect 20956 4324 21012 4380
rect 21012 4324 21016 4380
rect 20952 4320 21016 4324
rect 21032 4380 21096 4384
rect 21032 4324 21036 4380
rect 21036 4324 21092 4380
rect 21092 4324 21096 4380
rect 21032 4320 21096 4324
rect 21112 4380 21176 4384
rect 21112 4324 21116 4380
rect 21116 4324 21172 4380
rect 21172 4324 21176 4380
rect 21112 4320 21176 4324
rect 21192 4380 21256 4384
rect 21192 4324 21196 4380
rect 21196 4324 21252 4380
rect 21252 4324 21256 4380
rect 21192 4320 21256 4324
rect 34285 4380 34349 4384
rect 34285 4324 34289 4380
rect 34289 4324 34345 4380
rect 34345 4324 34349 4380
rect 34285 4320 34349 4324
rect 34365 4380 34429 4384
rect 34365 4324 34369 4380
rect 34369 4324 34425 4380
rect 34425 4324 34429 4380
rect 34365 4320 34429 4324
rect 34445 4380 34509 4384
rect 34445 4324 34449 4380
rect 34449 4324 34505 4380
rect 34505 4324 34509 4380
rect 34445 4320 34509 4324
rect 34525 4380 34589 4384
rect 34525 4324 34529 4380
rect 34529 4324 34585 4380
rect 34585 4324 34589 4380
rect 34525 4320 34589 4324
rect 8156 4252 8220 4316
rect 14285 3836 14349 3840
rect 14285 3780 14289 3836
rect 14289 3780 14345 3836
rect 14345 3780 14349 3836
rect 14285 3776 14349 3780
rect 14365 3836 14429 3840
rect 14365 3780 14369 3836
rect 14369 3780 14425 3836
rect 14425 3780 14429 3836
rect 14365 3776 14429 3780
rect 14445 3836 14509 3840
rect 14445 3780 14449 3836
rect 14449 3780 14505 3836
rect 14505 3780 14509 3836
rect 14445 3776 14509 3780
rect 14525 3836 14589 3840
rect 14525 3780 14529 3836
rect 14529 3780 14585 3836
rect 14585 3780 14589 3836
rect 14525 3776 14589 3780
rect 27618 3836 27682 3840
rect 27618 3780 27622 3836
rect 27622 3780 27678 3836
rect 27678 3780 27682 3836
rect 27618 3776 27682 3780
rect 27698 3836 27762 3840
rect 27698 3780 27702 3836
rect 27702 3780 27758 3836
rect 27758 3780 27762 3836
rect 27698 3776 27762 3780
rect 27778 3836 27842 3840
rect 27778 3780 27782 3836
rect 27782 3780 27838 3836
rect 27838 3780 27842 3836
rect 27778 3776 27842 3780
rect 27858 3836 27922 3840
rect 27858 3780 27862 3836
rect 27862 3780 27918 3836
rect 27918 3780 27922 3836
rect 27858 3776 27922 3780
rect 11836 3572 11900 3636
rect 35572 3572 35636 3636
rect 7618 3292 7682 3296
rect 7618 3236 7622 3292
rect 7622 3236 7678 3292
rect 7678 3236 7682 3292
rect 7618 3232 7682 3236
rect 7698 3292 7762 3296
rect 7698 3236 7702 3292
rect 7702 3236 7758 3292
rect 7758 3236 7762 3292
rect 7698 3232 7762 3236
rect 7778 3292 7842 3296
rect 7778 3236 7782 3292
rect 7782 3236 7838 3292
rect 7838 3236 7842 3292
rect 7778 3232 7842 3236
rect 7858 3292 7922 3296
rect 7858 3236 7862 3292
rect 7862 3236 7918 3292
rect 7918 3236 7922 3292
rect 7858 3232 7922 3236
rect 20952 3292 21016 3296
rect 20952 3236 20956 3292
rect 20956 3236 21012 3292
rect 21012 3236 21016 3292
rect 20952 3232 21016 3236
rect 21032 3292 21096 3296
rect 21032 3236 21036 3292
rect 21036 3236 21092 3292
rect 21092 3236 21096 3292
rect 21032 3232 21096 3236
rect 21112 3292 21176 3296
rect 21112 3236 21116 3292
rect 21116 3236 21172 3292
rect 21172 3236 21176 3292
rect 21112 3232 21176 3236
rect 21192 3292 21256 3296
rect 21192 3236 21196 3292
rect 21196 3236 21252 3292
rect 21252 3236 21256 3292
rect 21192 3232 21256 3236
rect 34285 3292 34349 3296
rect 34285 3236 34289 3292
rect 34289 3236 34345 3292
rect 34345 3236 34349 3292
rect 34285 3232 34349 3236
rect 34365 3292 34429 3296
rect 34365 3236 34369 3292
rect 34369 3236 34425 3292
rect 34425 3236 34429 3292
rect 34365 3232 34429 3236
rect 34445 3292 34509 3296
rect 34445 3236 34449 3292
rect 34449 3236 34505 3292
rect 34505 3236 34509 3292
rect 34445 3232 34509 3236
rect 34525 3292 34589 3296
rect 34525 3236 34529 3292
rect 34529 3236 34585 3292
rect 34585 3236 34589 3292
rect 34525 3232 34589 3236
rect 14285 2748 14349 2752
rect 14285 2692 14289 2748
rect 14289 2692 14345 2748
rect 14345 2692 14349 2748
rect 14285 2688 14349 2692
rect 14365 2748 14429 2752
rect 14365 2692 14369 2748
rect 14369 2692 14425 2748
rect 14425 2692 14429 2748
rect 14365 2688 14429 2692
rect 14445 2748 14509 2752
rect 14445 2692 14449 2748
rect 14449 2692 14505 2748
rect 14505 2692 14509 2748
rect 14445 2688 14509 2692
rect 14525 2748 14589 2752
rect 14525 2692 14529 2748
rect 14529 2692 14585 2748
rect 14585 2692 14589 2748
rect 14525 2688 14589 2692
rect 27618 2748 27682 2752
rect 27618 2692 27622 2748
rect 27622 2692 27678 2748
rect 27678 2692 27682 2748
rect 27618 2688 27682 2692
rect 27698 2748 27762 2752
rect 27698 2692 27702 2748
rect 27702 2692 27758 2748
rect 27758 2692 27762 2748
rect 27698 2688 27762 2692
rect 27778 2748 27842 2752
rect 27778 2692 27782 2748
rect 27782 2692 27838 2748
rect 27838 2692 27842 2748
rect 27778 2688 27842 2692
rect 27858 2748 27922 2752
rect 27858 2692 27862 2748
rect 27862 2692 27918 2748
rect 27918 2692 27922 2748
rect 27858 2688 27922 2692
rect 7618 2204 7682 2208
rect 7618 2148 7622 2204
rect 7622 2148 7678 2204
rect 7678 2148 7682 2204
rect 7618 2144 7682 2148
rect 7698 2204 7762 2208
rect 7698 2148 7702 2204
rect 7702 2148 7758 2204
rect 7758 2148 7762 2204
rect 7698 2144 7762 2148
rect 7778 2204 7842 2208
rect 7778 2148 7782 2204
rect 7782 2148 7838 2204
rect 7838 2148 7842 2204
rect 7778 2144 7842 2148
rect 7858 2204 7922 2208
rect 7858 2148 7862 2204
rect 7862 2148 7918 2204
rect 7918 2148 7922 2204
rect 7858 2144 7922 2148
rect 20952 2204 21016 2208
rect 20952 2148 20956 2204
rect 20956 2148 21012 2204
rect 21012 2148 21016 2204
rect 20952 2144 21016 2148
rect 21032 2204 21096 2208
rect 21032 2148 21036 2204
rect 21036 2148 21092 2204
rect 21092 2148 21096 2204
rect 21032 2144 21096 2148
rect 21112 2204 21176 2208
rect 21112 2148 21116 2204
rect 21116 2148 21172 2204
rect 21172 2148 21176 2204
rect 21112 2144 21176 2148
rect 21192 2204 21256 2208
rect 21192 2148 21196 2204
rect 21196 2148 21252 2204
rect 21252 2148 21256 2204
rect 21192 2144 21256 2148
rect 34285 2204 34349 2208
rect 34285 2148 34289 2204
rect 34289 2148 34345 2204
rect 34345 2148 34349 2204
rect 34285 2144 34349 2148
rect 34365 2204 34429 2208
rect 34365 2148 34369 2204
rect 34369 2148 34425 2204
rect 34425 2148 34429 2204
rect 34365 2144 34429 2148
rect 34445 2204 34509 2208
rect 34445 2148 34449 2204
rect 34449 2148 34505 2204
rect 34505 2148 34509 2204
rect 34445 2144 34509 2148
rect 34525 2204 34589 2208
rect 34525 2148 34529 2204
rect 34529 2148 34585 2204
rect 34585 2148 34589 2204
rect 34525 2144 34589 2148
<< metal4 >>
rect 7610 13088 7931 13648
rect 7610 13024 7618 13088
rect 7682 13024 7698 13088
rect 7762 13024 7778 13088
rect 7842 13024 7858 13088
rect 7922 13024 7931 13088
rect 7610 12000 7931 13024
rect 7610 11936 7618 12000
rect 7682 11936 7698 12000
rect 7762 11936 7778 12000
rect 7842 11936 7858 12000
rect 7922 11936 7931 12000
rect 3003 11524 3069 11525
rect 3003 11460 3004 11524
rect 3068 11460 3069 11524
rect 3003 11459 3069 11460
rect 3006 8618 3066 11459
rect 7610 10912 7931 11936
rect 7610 10848 7618 10912
rect 7682 10848 7698 10912
rect 7762 10848 7778 10912
rect 7842 10848 7858 10912
rect 7922 10848 7931 10912
rect 7610 9824 7931 10848
rect 7610 9760 7618 9824
rect 7682 9760 7698 9824
rect 7762 9760 7778 9824
rect 7842 9760 7858 9824
rect 7922 9760 7931 9824
rect 7610 8736 7931 9760
rect 14277 13632 14597 13648
rect 14277 13568 14285 13632
rect 14349 13568 14365 13632
rect 14429 13568 14445 13632
rect 14509 13568 14525 13632
rect 14589 13568 14597 13632
rect 14277 12544 14597 13568
rect 14277 12480 14285 12544
rect 14349 12480 14365 12544
rect 14429 12480 14445 12544
rect 14509 12480 14525 12544
rect 14589 12480 14597 12544
rect 14277 11456 14597 12480
rect 14277 11392 14285 11456
rect 14349 11392 14365 11456
rect 14429 11392 14445 11456
rect 14509 11392 14525 11456
rect 14589 11392 14597 11456
rect 14277 10368 14597 11392
rect 14277 10304 14285 10368
rect 14349 10304 14365 10368
rect 14429 10304 14445 10368
rect 14509 10304 14525 10368
rect 14589 10304 14597 10368
rect 8155 9348 8221 9349
rect 8155 9284 8156 9348
rect 8220 9284 8221 9348
rect 8155 9283 8221 9284
rect 7610 8672 7618 8736
rect 7682 8672 7698 8736
rect 7762 8672 7778 8736
rect 7842 8672 7858 8736
rect 7922 8672 7931 8736
rect 3006 7173 3066 8382
rect 3926 7445 3986 7702
rect 7610 7648 7931 8672
rect 7610 7584 7618 7648
rect 7682 7584 7698 7648
rect 7762 7584 7778 7648
rect 7842 7584 7858 7648
rect 7922 7584 7931 7648
rect 3923 7444 3989 7445
rect 3923 7380 3924 7444
rect 3988 7380 3989 7444
rect 3923 7379 3989 7380
rect 3003 7172 3069 7173
rect 3003 7108 3004 7172
rect 3068 7108 3069 7172
rect 3003 7107 3069 7108
rect 7610 6560 7931 7584
rect 7610 6496 7618 6560
rect 7682 6496 7698 6560
rect 7762 6496 7778 6560
rect 7842 6496 7858 6560
rect 7922 6496 7931 6560
rect 7610 5472 7931 6496
rect 7610 5408 7618 5472
rect 7682 5408 7698 5472
rect 7762 5408 7778 5472
rect 7842 5408 7858 5472
rect 7922 5408 7931 5472
rect 3923 5404 3989 5405
rect 3923 5340 3924 5404
rect 3988 5340 3989 5404
rect 3923 5339 3989 5340
rect 3926 5218 3986 5339
rect 7610 4384 7931 5408
rect 7610 4320 7618 4384
rect 7682 4320 7698 4384
rect 7762 4320 7778 4384
rect 7842 4320 7858 4384
rect 7922 4320 7931 4384
rect 7610 3296 7931 4320
rect 8158 4317 8218 9283
rect 14277 9280 14597 10304
rect 20944 13088 21264 13648
rect 20944 13024 20952 13088
rect 21016 13024 21032 13088
rect 21096 13024 21112 13088
rect 21176 13024 21192 13088
rect 21256 13024 21264 13088
rect 20944 12000 21264 13024
rect 27610 13632 27930 13648
rect 27610 13568 27618 13632
rect 27682 13568 27698 13632
rect 27762 13568 27778 13632
rect 27842 13568 27858 13632
rect 27922 13568 27930 13632
rect 24715 12612 24781 12613
rect 24715 12548 24716 12612
rect 24780 12548 24781 12612
rect 24715 12547 24781 12548
rect 20944 11936 20952 12000
rect 21016 11936 21032 12000
rect 21096 11936 21112 12000
rect 21176 11936 21192 12000
rect 21256 11936 21264 12000
rect 20944 10912 21264 11936
rect 20944 10848 20952 10912
rect 21016 10848 21032 10912
rect 21096 10848 21112 10912
rect 21176 10848 21192 10912
rect 21256 10848 21264 10912
rect 20667 10300 20733 10301
rect 20667 10236 20668 10300
rect 20732 10236 20733 10300
rect 20667 10235 20733 10236
rect 14277 9216 14285 9280
rect 14349 9216 14365 9280
rect 14429 9216 14445 9280
rect 14509 9216 14525 9280
rect 14589 9216 14597 9280
rect 14277 8192 14597 9216
rect 15147 8396 15213 8397
rect 15147 8332 15148 8396
rect 15212 8332 15213 8396
rect 15147 8331 15213 8332
rect 14277 8128 14285 8192
rect 14349 8128 14365 8192
rect 14429 8128 14445 8192
rect 14509 8128 14525 8192
rect 14589 8128 14597 8192
rect 14277 7104 14597 8128
rect 15150 7938 15210 8331
rect 19382 7173 19442 7702
rect 19379 7172 19445 7173
rect 19379 7108 19380 7172
rect 19444 7108 19445 7172
rect 19379 7107 19445 7108
rect 14277 7040 14285 7104
rect 14349 7040 14365 7104
rect 14429 7040 14445 7104
rect 14509 7040 14525 7104
rect 14589 7040 14597 7104
rect 14277 6016 14597 7040
rect 14277 5952 14285 6016
rect 14349 5952 14365 6016
rect 14429 5952 14445 6016
rect 14509 5952 14525 6016
rect 14589 5952 14597 6016
rect 14277 4928 14597 5952
rect 19379 5948 19445 5949
rect 19379 5898 19380 5948
rect 19444 5898 19445 5948
rect 20670 5218 20730 10235
rect 20944 9824 21264 10848
rect 20944 9760 20952 9824
rect 21016 9760 21032 9824
rect 21096 9760 21112 9824
rect 21176 9760 21192 9824
rect 21256 9760 21264 9824
rect 20944 8736 21264 9760
rect 20944 8672 20952 8736
rect 21016 8672 21032 8736
rect 21096 8672 21112 8736
rect 21176 8672 21192 8736
rect 21256 8672 21264 8736
rect 20944 7648 21264 8672
rect 20944 7584 20952 7648
rect 21016 7584 21032 7648
rect 21096 7584 21112 7648
rect 21176 7584 21192 7648
rect 21256 7584 21264 7648
rect 20944 6560 21264 7584
rect 20944 6496 20952 6560
rect 21016 6496 21032 6560
rect 21096 6496 21112 6560
rect 21176 6496 21192 6560
rect 21256 6496 21264 6560
rect 20944 5472 21264 6496
rect 20944 5408 20952 5472
rect 21016 5408 21032 5472
rect 21096 5408 21112 5472
rect 21176 5408 21192 5472
rect 21256 5408 21264 5472
rect 14277 4864 14285 4928
rect 14349 4864 14365 4928
rect 14429 4864 14445 4928
rect 14509 4864 14525 4928
rect 14589 4864 14597 4928
rect 8155 4316 8221 4317
rect 8155 4252 8156 4316
rect 8220 4252 8221 4316
rect 8155 4251 8221 4252
rect 14277 3840 14597 4864
rect 14277 3776 14285 3840
rect 14349 3776 14365 3840
rect 14429 3776 14445 3840
rect 14509 3776 14525 3840
rect 14589 3776 14597 3840
rect 11835 3572 11836 3622
rect 11900 3572 11901 3622
rect 11835 3571 11901 3572
rect 7610 3232 7618 3296
rect 7682 3232 7698 3296
rect 7762 3232 7778 3296
rect 7842 3232 7858 3296
rect 7922 3232 7931 3296
rect 7610 2208 7931 3232
rect 7610 2144 7618 2208
rect 7682 2144 7698 2208
rect 7762 2144 7778 2208
rect 7842 2144 7858 2208
rect 7922 2144 7931 2208
rect 7610 2128 7931 2144
rect 14277 2752 14597 3776
rect 14277 2688 14285 2752
rect 14349 2688 14365 2752
rect 14429 2688 14445 2752
rect 14509 2688 14525 2752
rect 14589 2688 14597 2752
rect 14277 2128 14597 2688
rect 20944 4384 21264 5408
rect 20944 4320 20952 4384
rect 21016 4320 21032 4384
rect 21096 4320 21112 4384
rect 21176 4320 21192 4384
rect 21256 4320 21264 4384
rect 20944 3296 21264 4320
rect 24718 3858 24778 12547
rect 27610 12544 27930 13568
rect 27610 12480 27618 12544
rect 27682 12480 27698 12544
rect 27762 12480 27778 12544
rect 27842 12480 27858 12544
rect 27922 12480 27930 12544
rect 27610 11456 27930 12480
rect 27610 11392 27618 11456
rect 27682 11392 27698 11456
rect 27762 11392 27778 11456
rect 27842 11392 27858 11456
rect 27922 11392 27930 11456
rect 27610 10368 27930 11392
rect 27610 10304 27618 10368
rect 27682 10304 27698 10368
rect 27762 10304 27778 10368
rect 27842 10304 27858 10368
rect 27922 10304 27930 10368
rect 27610 9280 27930 10304
rect 27610 9216 27618 9280
rect 27682 9216 27698 9280
rect 27762 9216 27778 9280
rect 27842 9216 27858 9280
rect 27922 9216 27930 9280
rect 27610 8192 27930 9216
rect 34277 13088 34597 13648
rect 34277 13024 34285 13088
rect 34349 13024 34365 13088
rect 34429 13024 34445 13088
rect 34509 13024 34525 13088
rect 34589 13024 34597 13088
rect 34277 12000 34597 13024
rect 34277 11936 34285 12000
rect 34349 11936 34365 12000
rect 34429 11936 34445 12000
rect 34509 11936 34525 12000
rect 34589 11936 34597 12000
rect 34277 10912 34597 11936
rect 34277 10848 34285 10912
rect 34349 10848 34365 10912
rect 34429 10848 34445 10912
rect 34509 10848 34525 10912
rect 34589 10848 34597 10912
rect 34277 9824 34597 10848
rect 34277 9760 34285 9824
rect 34349 9760 34365 9824
rect 34429 9760 34445 9824
rect 34509 9760 34525 9824
rect 34589 9760 34597 9824
rect 34277 8736 34597 9760
rect 34277 8672 34285 8736
rect 34349 8672 34365 8736
rect 34429 8672 34445 8736
rect 34509 8672 34525 8736
rect 34589 8672 34597 8736
rect 30603 8396 30669 8397
rect 30603 8332 30604 8396
rect 30668 8332 30669 8396
rect 30603 8331 30669 8332
rect 27610 8128 27618 8192
rect 27682 8128 27698 8192
rect 27762 8128 27778 8192
rect 27842 8128 27858 8192
rect 27922 8128 27930 8192
rect 27610 7104 27930 8128
rect 30606 7938 30666 8331
rect 27610 7040 27618 7104
rect 27682 7040 27698 7104
rect 27762 7040 27778 7104
rect 27842 7040 27858 7104
rect 27922 7040 27930 7104
rect 27610 6016 27930 7040
rect 27610 5952 27618 6016
rect 27682 5952 27698 6016
rect 27762 5952 27778 6016
rect 27842 5952 27858 6016
rect 27922 5952 27930 6016
rect 27610 4928 27930 5952
rect 34277 7648 34597 8672
rect 34277 7584 34285 7648
rect 34349 7584 34365 7648
rect 34429 7584 34445 7648
rect 34509 7584 34525 7648
rect 34589 7584 34597 7648
rect 34277 6560 34597 7584
rect 34277 6496 34285 6560
rect 34349 6496 34365 6560
rect 34429 6496 34445 6560
rect 34509 6496 34525 6560
rect 34589 6496 34597 6560
rect 28947 5540 29013 5541
rect 28947 5476 28948 5540
rect 29012 5476 29013 5540
rect 28947 5475 29013 5476
rect 28950 5133 29010 5475
rect 34277 5472 34597 6496
rect 34277 5408 34285 5472
rect 34349 5408 34365 5472
rect 34429 5408 34445 5472
rect 34509 5408 34525 5472
rect 34589 5408 34597 5472
rect 28947 5132 29013 5133
rect 28947 5068 28948 5132
rect 29012 5068 29013 5132
rect 28947 5067 29013 5068
rect 27610 4864 27618 4928
rect 27682 4864 27698 4928
rect 27762 4864 27778 4928
rect 27842 4864 27858 4928
rect 27922 4864 27930 4928
rect 27610 3840 27930 4864
rect 27610 3776 27618 3840
rect 27682 3776 27698 3840
rect 27762 3776 27778 3840
rect 27842 3776 27858 3840
rect 27922 3776 27930 3840
rect 20944 3232 20952 3296
rect 21016 3232 21032 3296
rect 21096 3232 21112 3296
rect 21176 3232 21192 3296
rect 21256 3232 21264 3296
rect 20944 2208 21264 3232
rect 20944 2144 20952 2208
rect 21016 2144 21032 2208
rect 21096 2144 21112 2208
rect 21176 2144 21192 2208
rect 21256 2144 21264 2208
rect 20944 2128 21264 2144
rect 27610 2752 27930 3776
rect 27610 2688 27618 2752
rect 27682 2688 27698 2752
rect 27762 2688 27778 2752
rect 27842 2688 27858 2752
rect 27922 2688 27930 2752
rect 27610 2128 27930 2688
rect 34277 4384 34597 5408
rect 34277 4320 34285 4384
rect 34349 4320 34365 4384
rect 34429 4320 34445 4384
rect 34509 4320 34525 4384
rect 34589 4320 34597 4384
rect 34277 3296 34597 4320
rect 35571 3572 35572 3622
rect 35636 3572 35637 3622
rect 35571 3571 35637 3572
rect 34277 3232 34285 3296
rect 34349 3232 34365 3296
rect 34429 3232 34445 3296
rect 34509 3232 34525 3296
rect 34589 3232 34597 3296
rect 34277 2208 34597 3232
rect 34277 2144 34285 2208
rect 34349 2144 34365 2208
rect 34429 2144 34445 2208
rect 34509 2144 34525 2208
rect 34589 2144 34597 2208
rect 34277 2128 34597 2144
<< via4 >>
rect 2918 8382 3154 8618
rect 3838 7702 4074 7938
rect 6230 5812 6466 5898
rect 6230 5748 6316 5812
rect 6316 5748 6380 5812
rect 6380 5748 6466 5812
rect 6230 5662 6466 5748
rect 3838 4982 4074 5218
rect 15062 7702 15298 7938
rect 19294 7702 19530 7938
rect 19294 5884 19380 5898
rect 19380 5884 19444 5898
rect 19444 5884 19530 5898
rect 19294 5662 19530 5884
rect 20582 4982 20818 5218
rect 11198 4452 11434 4538
rect 11198 4388 11284 4452
rect 11284 4388 11348 4452
rect 11348 4388 11434 4452
rect 11198 4302 11434 4388
rect 11750 3636 11986 3858
rect 11750 3622 11836 3636
rect 11836 3622 11900 3636
rect 11900 3622 11986 3636
rect 23894 4452 24130 4538
rect 23894 4388 23980 4452
rect 23980 4388 24044 4452
rect 24044 4388 24130 4452
rect 23894 4302 24130 4388
rect 32542 8532 32778 8618
rect 32542 8468 32628 8532
rect 32628 8468 32692 8532
rect 32692 8468 32778 8532
rect 32542 8382 32778 8468
rect 30518 7702 30754 7938
rect 24630 3622 24866 3858
rect 35486 3636 35722 3858
rect 35486 3622 35572 3636
rect 35572 3622 35636 3636
rect 35636 3622 35722 3636
<< metal5 >>
rect 2876 8618 32820 8660
rect 2876 8382 2918 8618
rect 3154 8382 32542 8618
rect 32778 8382 32820 8618
rect 2876 8340 32820 8382
rect 3796 7938 30796 7980
rect 3796 7702 3838 7938
rect 4074 7702 15062 7938
rect 15298 7702 19294 7938
rect 19530 7702 30518 7938
rect 30754 7702 30796 7938
rect 3796 7660 30796 7702
rect 6188 5898 19572 5940
rect 6188 5662 6230 5898
rect 6466 5662 19294 5898
rect 19530 5662 19572 5898
rect 6188 5620 19572 5662
rect 3796 5218 20860 5260
rect 3796 4982 3838 5218
rect 4074 4982 20582 5218
rect 20818 4982 20860 5218
rect 3796 4940 20860 4982
rect 11156 4538 24172 4580
rect 11156 4302 11198 4538
rect 11434 4302 23894 4538
rect 24130 4302 24172 4538
rect 11156 4260 24172 4302
rect 11708 3858 35764 3900
rect 11708 3622 11750 3858
rect 11986 3622 24630 3858
rect 24866 3622 35486 3858
rect 35722 3622 35764 3858
rect 11708 3580 35764 3622
use scs8hd_decap_3  PHY_0 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1104 0 -1 2720
box -38 -48 314 592
use scs8hd_decap_3  PHY_2
timestamp 1586364061
transform 1 0 1104 0 1 2720
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__36__A tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1564 0 1 2720
box -38 -48 222 592
use scs8hd_decap_12  FILLER_0_3 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1380 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_15
timestamp 1586364061
transform 1 0 2484 0 -1 2720
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_1_3 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1380 0 1 2720
box -38 -48 222 592
use scs8hd_decap_12  FILLER_1_7
timestamp 1586364061
transform 1 0 1748 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_19
timestamp 1586364061
transform 1 0 2852 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_42 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 3956 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_4  FILLER_0_27 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 3588 0 -1 2720
box -38 -48 406 592
use scs8hd_decap_12  FILLER_0_32
timestamp 1586364061
transform 1 0 4048 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_31
timestamp 1586364061
transform 1 0 3956 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_44
timestamp 1586364061
transform 1 0 5152 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_0_56 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 6256 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_1_43
timestamp 1586364061
transform 1 0 5060 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_1_55
timestamp 1586364061
transform 1 0 6164 0 1 2720
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_43
timestamp 1586364061
transform 1 0 6808 0 -1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_55
timestamp 1586364061
transform 1 0 6716 0 1 2720
box -38 -48 130 592
use scs8hd_decap_12  FILLER_0_63
timestamp 1586364061
transform 1 0 6900 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_75
timestamp 1586364061
transform 1 0 8004 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_62
timestamp 1586364061
transform 1 0 6808 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_74
timestamp 1586364061
transform 1 0 7912 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_44
timestamp 1586364061
transform 1 0 9660 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_87
timestamp 1586364061
transform 1 0 9108 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_0_94
timestamp 1586364061
transform 1 0 9752 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_86
timestamp 1586364061
transform 1 0 9016 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_1_98 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 10120 0 1 2720
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_5.mux_l2_in_2__A0
timestamp 1586364061
transform 1 0 11224 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_5.mux_l2_in_2__A1
timestamp 1586364061
transform 1 0 11592 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_5.mux_l2_in_2__S
timestamp 1586364061
transform 1 0 10856 0 1 2720
box -38 -48 222 592
use scs8hd_decap_12  FILLER_0_106
timestamp 1586364061
transform 1 0 10856 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_0_118
timestamp 1586364061
transform 1 0 11960 0 -1 2720
box -38 -48 590 592
use scs8hd_fill_2  FILLER_1_108
timestamp 1586364061
transform 1 0 11040 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_112
timestamp 1586364061
transform 1 0 11408 0 1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_1_116
timestamp 1586364061
transform 1 0 11776 0 1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_0_125
timestamp 1586364061
transform 1 0 12604 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_4.mux_l3_in_1__A1
timestamp 1586364061
transform 1 0 12788 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_4.mux_l3_in_1__S
timestamp 1586364061
transform 1 0 12144 0 1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_56
timestamp 1586364061
transform 1 0 12328 0 1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_45
timestamp 1586364061
transform 1 0 12512 0 -1 2720
box -38 -48 130 592
use scs8hd_mux2_2  mux_bottom_ipin_4.mux_l3_in_1_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 12420 0 1 2720
box -38 -48 866 592
use scs8hd_fill_2  FILLER_1_136
timestamp 1586364061
transform 1 0 13616 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_132
timestamp 1586364061
transform 1 0 13248 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_133
timestamp 1586364061
transform 1 0 13340 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_129
timestamp 1586364061
transform 1 0 12972 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_4.mux_l4_in_0__A0
timestamp 1586364061
transform 1 0 13524 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_4.mux_l4_in_0__A1
timestamp 1586364061
transform 1 0 13800 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_4.mux_l3_in_1__A0
timestamp 1586364061
transform 1 0 13156 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_4.mux_l4_in_0__S
timestamp 1586364061
transform 1 0 13432 0 1 2720
box -38 -48 222 592
use scs8hd_decap_12  FILLER_0_137
timestamp 1586364061
transform 1 0 13708 0 -1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_46
timestamp 1586364061
transform 1 0 15364 0 -1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_5.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 14168 0 1 2720
box -38 -48 222 592
use scs8hd_decap_6  FILLER_0_149
timestamp 1586364061
transform 1 0 14812 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_0_156
timestamp 1586364061
transform 1 0 15456 0 -1 2720
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_1_140
timestamp 1586364061
transform 1 0 13984 0 1 2720
box -38 -48 222 592
use scs8hd_decap_12  FILLER_1_144
timestamp 1586364061
transform 1 0 14352 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_156
timestamp 1586364061
transform 1 0 15456 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_168
timestamp 1586364061
transform 1 0 16560 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_168
timestamp 1586364061
transform 1 0 16560 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_47
timestamp 1586364061
transform 1 0 18216 0 -1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_57
timestamp 1586364061
transform 1 0 17940 0 1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_180
timestamp 1586364061
transform 1 0 17664 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_0_187
timestamp 1586364061
transform 1 0 18308 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_1_180
timestamp 1586364061
transform 1 0 17664 0 1 2720
box -38 -48 314 592
use scs8hd_decap_12  FILLER_1_184
timestamp 1586364061
transform 1 0 18032 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_196
timestamp 1586364061
transform 1 0 19136 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_48
timestamp 1586364061
transform 1 0 21068 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_12  FILLER_0_199
timestamp 1586364061
transform 1 0 19412 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_0_211
timestamp 1586364061
transform 1 0 20516 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_0_218
timestamp 1586364061
transform 1 0 21160 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_208
timestamp 1586364061
transform 1 0 20240 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_230
timestamp 1586364061
transform 1 0 22264 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_220
timestamp 1586364061
transform 1 0 21344 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_232
timestamp 1586364061
transform 1 0 22448 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_49
timestamp 1586364061
transform 1 0 23920 0 -1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_58
timestamp 1586364061
transform 1 0 23552 0 1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_242
timestamp 1586364061
transform 1 0 23368 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_0_249
timestamp 1586364061
transform 1 0 24012 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_245
timestamp 1586364061
transform 1 0 23644 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_257
timestamp 1586364061
transform 1 0 24748 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_261
timestamp 1586364061
transform 1 0 25116 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_0_273
timestamp 1586364061
transform 1 0 26220 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_1_269
timestamp 1586364061
transform 1 0 25852 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_50
timestamp 1586364061
transform 1 0 26772 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_12  FILLER_0_280
timestamp 1586364061
transform 1 0 26864 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_292
timestamp 1586364061
transform 1 0 27968 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_281
timestamp 1586364061
transform 1 0 26956 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_293
timestamp 1586364061
transform 1 0 28060 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_51
timestamp 1586364061
transform 1 0 29624 0 -1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_59
timestamp 1586364061
transform 1 0 29164 0 1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_304
timestamp 1586364061
transform 1 0 29072 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_0_311
timestamp 1586364061
transform 1 0 29716 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_306
timestamp 1586364061
transform 1 0 29256 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_323
timestamp 1586364061
transform 1 0 30820 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_0_335
timestamp 1586364061
transform 1 0 31924 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_1_318
timestamp 1586364061
transform 1 0 30360 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_330
timestamp 1586364061
transform 1 0 31464 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_52
timestamp 1586364061
transform 1 0 32476 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_12  FILLER_0_342
timestamp 1586364061
transform 1 0 32568 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_354
timestamp 1586364061
transform 1 0 33672 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_342
timestamp 1586364061
transform 1 0 32568 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_354
timestamp 1586364061
transform 1 0 33672 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_53
timestamp 1586364061
transform 1 0 35328 0 -1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_60
timestamp 1586364061
transform 1 0 34776 0 1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_366
timestamp 1586364061
transform 1 0 34776 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_0_373
timestamp 1586364061
transform 1 0 35420 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_367
timestamp 1586364061
transform 1 0 34868 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_385
timestamp 1586364061
transform 1 0 36524 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_379
timestamp 1586364061
transform 1 0 35972 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_391
timestamp 1586364061
transform 1 0 37076 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_3  PHY_1
timestamp 1586364061
transform -1 0 38824 0 -1 2720
box -38 -48 314 592
use scs8hd_decap_3  PHY_3
timestamp 1586364061
transform -1 0 38824 0 1 2720
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_54
timestamp 1586364061
transform 1 0 38180 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_397
timestamp 1586364061
transform 1 0 37628 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_3  FILLER_0_404
timestamp 1586364061
transform 1 0 38272 0 -1 2720
box -38 -48 314 592
use scs8hd_decap_4  FILLER_1_403
timestamp 1586364061
transform 1 0 38180 0 1 2720
box -38 -48 406 592
use scs8hd_buf_2  _36_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1380 0 -1 3808
box -38 -48 406 592
use scs8hd_decap_3  PHY_4
timestamp 1586364061
transform 1 0 1104 0 -1 3808
box -38 -48 314 592
use scs8hd_decap_12  FILLER_2_7
timestamp 1586364061
transform 1 0 1748 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_19
timestamp 1586364061
transform 1 0 2852 0 -1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_61
timestamp 1586364061
transform 1 0 3956 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_2_32
timestamp 1586364061
transform 1 0 4048 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_44
timestamp 1586364061
transform 1 0 5152 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_56
timestamp 1586364061
transform 1 0 6256 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_68
timestamp 1586364061
transform 1 0 7360 0 -1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_62
timestamp 1586364061
transform 1 0 9568 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_2_80
timestamp 1586364061
transform 1 0 8464 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_2_93
timestamp 1586364061
transform 1 0 9660 0 -1 3808
box -38 -48 774 592
use scs8hd_mux2_2  mux_bottom_ipin_5.mux_l2_in_2_
timestamp 1586364061
transform 1 0 11224 0 -1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_5.mux_l2_in_3__A0
timestamp 1586364061
transform 1 0 10764 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_5.mux_l3_in_1__S
timestamp 1586364061
transform 1 0 10396 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_103
timestamp 1586364061
transform 1 0 10580 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_3  FILLER_2_107
timestamp 1586364061
transform 1 0 10948 0 -1 3808
box -38 -48 314 592
use scs8hd_decap_4  FILLER_2_119
timestamp 1586364061
transform 1 0 12052 0 -1 3808
box -38 -48 406 592
use scs8hd_mux2_2  mux_bottom_ipin_4.mux_l4_in_0_
timestamp 1586364061
transform 1 0 12788 0 -1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_4.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 13800 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_4.mux_l1_in_2__A0
timestamp 1586364061
transform 1 0 12420 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_125
timestamp 1586364061
transform 1 0 12604 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_136
timestamp 1586364061
transform 1 0 13616 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_2_148
timestamp 1586364061
transform 1 0 14720 0 -1 3808
box -38 -48 406 592
use scs8hd_fill_2  FILLER_2_144
timestamp 1586364061
transform 1 0 14352 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_140
timestamp 1586364061
transform 1 0 13984 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_5.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 14536 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_4.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 14168 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_154
timestamp 1586364061
transform 1 0 15272 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_1  FILLER_2_152 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 15088 0 -1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_5.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 15456 0 -1 3808
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_63
timestamp 1586364061
transform 1 0 15180 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_2_158
timestamp 1586364061
transform 1 0 15640 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_170
timestamp 1586364061
transform 1 0 16744 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_182
timestamp 1586364061
transform 1 0 17848 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_194
timestamp 1586364061
transform 1 0 18952 0 -1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_64
timestamp 1586364061
transform 1 0 20792 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_8  FILLER_2_206
timestamp 1586364061
transform 1 0 20056 0 -1 3808
box -38 -48 774 592
use scs8hd_decap_12  FILLER_2_215
timestamp 1586364061
transform 1 0 20884 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_227
timestamp 1586364061
transform 1 0 21988 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_239
timestamp 1586364061
transform 1 0 23092 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_251
timestamp 1586364061
transform 1 0 24196 0 -1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_65
timestamp 1586364061
transform 1 0 26404 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_2_263
timestamp 1586364061
transform 1 0 25300 0 -1 3808
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_2_276
timestamp 1586364061
transform 1 0 26496 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_12.mux_l2_in_3__S
timestamp 1586364061
transform 1 0 26680 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_12  FILLER_2_280
timestamp 1586364061
transform 1 0 26864 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_292
timestamp 1586364061
transform 1 0 27968 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_304
timestamp 1586364061
transform 1 0 29072 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_316
timestamp 1586364061
transform 1 0 30176 0 -1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_66
timestamp 1586364061
transform 1 0 32016 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_8  FILLER_2_328
timestamp 1586364061
transform 1 0 31280 0 -1 3808
box -38 -48 774 592
use scs8hd_decap_12  FILLER_2_337
timestamp 1586364061
transform 1 0 32108 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_349
timestamp 1586364061
transform 1 0 33212 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_361
timestamp 1586364061
transform 1 0 34316 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_373
timestamp 1586364061
transform 1 0 35420 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_385
timestamp 1586364061
transform 1 0 36524 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_3  PHY_5
timestamp 1586364061
transform -1 0 38824 0 -1 3808
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_67
timestamp 1586364061
transform 1 0 37628 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_8  FILLER_2_398
timestamp 1586364061
transform 1 0 37720 0 -1 3808
box -38 -48 774 592
use scs8hd_fill_1  FILLER_2_406
timestamp 1586364061
transform 1 0 38456 0 -1 3808
box -38 -48 130 592
use scs8hd_conb_1  _27_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 2484 0 1 3808
box -38 -48 314 592
use scs8hd_buf_2  _49_
timestamp 1586364061
transform 1 0 1380 0 1 3808
box -38 -48 406 592
use scs8hd_decap_3  PHY_6
timestamp 1586364061
transform 1 0 1104 0 1 3808
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__49__A
timestamp 1586364061
transform 1 0 1932 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__44__A
timestamp 1586364061
transform 1 0 2300 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_7
timestamp 1586364061
transform 1 0 1748 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_11
timestamp 1586364061
transform 1 0 2116 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_18
timestamp 1586364061
transform 1 0 2760 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__50__A
timestamp 1586364061
transform 1 0 2944 0 1 3808
box -38 -48 222 592
use scs8hd_decap_12  FILLER_3_22
timestamp 1586364061
transform 1 0 3128 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_34
timestamp 1586364061
transform 1 0 4232 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_46
timestamp 1586364061
transform 1 0 5336 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_3_58
timestamp 1586364061
transform 1 0 6440 0 1 3808
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_68
timestamp 1586364061
transform 1 0 6716 0 1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_3.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 7544 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_3.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 7912 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_3.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 8280 0 1 3808
box -38 -48 222 592
use scs8hd_decap_8  FILLER_3_62
timestamp 1586364061
transform 1 0 6808 0 1 3808
box -38 -48 774 592
use scs8hd_fill_2  FILLER_3_72
timestamp 1586364061
transform 1 0 7728 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_76
timestamp 1586364061
transform 1 0 8096 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_5.mux_l2_in_3__S
timestamp 1586364061
transform 1 0 10212 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_5.mux_l3_in_1__A1
timestamp 1586364061
transform 1 0 9844 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_5.mux_l3_in_1__A0
timestamp 1586364061
transform 1 0 9476 0 1 3808
box -38 -48 222 592
use scs8hd_decap_8  FILLER_3_80
timestamp 1586364061
transform 1 0 8464 0 1 3808
box -38 -48 774 592
use scs8hd_decap_3  FILLER_3_88
timestamp 1586364061
transform 1 0 9200 0 1 3808
box -38 -48 314 592
use scs8hd_fill_2  FILLER_3_93
timestamp 1586364061
transform 1 0 9660 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_97
timestamp 1586364061
transform 1 0 10028 0 1 3808
box -38 -48 222 592
use scs8hd_mux2_2  mux_bottom_ipin_5.mux_l2_in_3_
timestamp 1586364061
transform 1 0 10764 0 1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_5.mux_l2_in_3__A1
timestamp 1586364061
transform 1 0 10580 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_4.mux_l1_in_2__S
timestamp 1586364061
transform 1 0 11776 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_101
timestamp 1586364061
transform 1 0 10396 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_114
timestamp 1586364061
transform 1 0 11592 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_118
timestamp 1586364061
transform 1 0 11960 0 1 3808
box -38 -48 222 592
use scs8hd_mux2_2  mux_bottom_ipin_4.mux_l1_in_2_
timestamp 1586364061
transform 1 0 12420 0 1 3808
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_69
timestamp 1586364061
transform 1 0 12328 0 1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_4.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 13524 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_4.mux_l1_in_2__A1
timestamp 1586364061
transform 1 0 12144 0 1 3808
box -38 -48 222 592
use scs8hd_decap_3  FILLER_3_132
timestamp 1586364061
transform 1 0 13248 0 1 3808
box -38 -48 314 592
use scs8hd_decap_3  FILLER_3_137
timestamp 1586364061
transform 1 0 13708 0 1 3808
box -38 -48 314 592
use scs8hd_mux2_2  mux_bottom_ipin_5.mux_l3_in_0_
timestamp 1586364061
transform 1 0 13984 0 1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_5.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 15272 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_5.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 15640 0 1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_3_149
timestamp 1586364061
transform 1 0 14812 0 1 3808
box -38 -48 406 592
use scs8hd_fill_1  FILLER_3_153
timestamp 1586364061
transform 1 0 15180 0 1 3808
box -38 -48 130 592
use scs8hd_fill_2  FILLER_3_156
timestamp 1586364061
transform 1 0 15456 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_5.mux_l1_in_2__A1
timestamp 1586364061
transform 1 0 16836 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_5.mux_l1_in_2__A0
timestamp 1586364061
transform 1 0 17204 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_5.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 16008 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_160
timestamp 1586364061
transform 1 0 15824 0 1 3808
box -38 -48 222 592
use scs8hd_decap_6  FILLER_3_164
timestamp 1586364061
transform 1 0 16192 0 1 3808
box -38 -48 590 592
use scs8hd_fill_1  FILLER_3_170
timestamp 1586364061
transform 1 0 16744 0 1 3808
box -38 -48 130 592
use scs8hd_fill_2  FILLER_3_173
timestamp 1586364061
transform 1 0 17020 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_177
timestamp 1586364061
transform 1 0 17388 0 1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_3_184
timestamp 1586364061
transform 1 0 18032 0 1 3808
box -38 -48 406 592
use scs8hd_fill_2  FILLER_3_181
timestamp 1586364061
transform 1 0 17756 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_5.mux_l1_in_2__S
timestamp 1586364061
transform 1 0 17572 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_5.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 18400 0 1 3808
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_70
timestamp 1586364061
transform 1 0 17940 0 1 3808
box -38 -48 130 592
use scs8hd_fill_2  FILLER_3_194
timestamp 1586364061
transform 1 0 18952 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_190
timestamp 1586364061
transform 1 0 18584 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_5.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 19136 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_5.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 18768 0 1 3808
box -38 -48 222 592
use scs8hd_decap_12  FILLER_3_198
timestamp 1586364061
transform 1 0 19320 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_210
timestamp 1586364061
transform 1 0 20424 0 1 3808
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_11.mux_l4_in_0__S
timestamp 1586364061
transform 1 0 21988 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_11.mux_l4_in_0__A1
timestamp 1586364061
transform 1 0 22356 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_11.mux_l4_in_0__A0
timestamp 1586364061
transform 1 0 22724 0 1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_3_222
timestamp 1586364061
transform 1 0 21528 0 1 3808
box -38 -48 406 592
use scs8hd_fill_1  FILLER_3_226
timestamp 1586364061
transform 1 0 21896 0 1 3808
box -38 -48 130 592
use scs8hd_fill_2  FILLER_3_229
timestamp 1586364061
transform 1 0 22172 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_233
timestamp 1586364061
transform 1 0 22540 0 1 3808
box -38 -48 222 592
use scs8hd_decap_6  FILLER_3_237
timestamp 1586364061
transform 1 0 22908 0 1 3808
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_71
timestamp 1586364061
transform 1 0 23552 0 1 3808
box -38 -48 130 592
use scs8hd_fill_1  FILLER_3_243
timestamp 1586364061
transform 1 0 23460 0 1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_3_245
timestamp 1586364061
transform 1 0 23644 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_257
timestamp 1586364061
transform 1 0 24748 0 1 3808
box -38 -48 1142 592
use scs8hd_mux2_2  mux_bottom_ipin_12.mux_l2_in_3_
timestamp 1586364061
transform 1 0 26588 0 1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_12.mux_l2_in_3__A1
timestamp 1586364061
transform 1 0 26404 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_12.mux_l2_in_3__A0
timestamp 1586364061
transform 1 0 26036 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_269
timestamp 1586364061
transform 1 0 25852 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_273
timestamp 1586364061
transform 1 0 26220 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_12.mux_l1_in_2__A1
timestamp 1586364061
transform 1 0 27600 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_12.mux_l1_in_2__A0
timestamp 1586364061
transform 1 0 27968 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_12.mux_l1_in_2__S
timestamp 1586364061
transform 1 0 28336 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_286
timestamp 1586364061
transform 1 0 27416 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_290
timestamp 1586364061
transform 1 0 27784 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_294
timestamp 1586364061
transform 1 0 28152 0 1 3808
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_72
timestamp 1586364061
transform 1 0 29164 0 1 3808
box -38 -48 130 592
use scs8hd_decap_6  FILLER_3_298
timestamp 1586364061
transform 1 0 28520 0 1 3808
box -38 -48 590 592
use scs8hd_fill_1  FILLER_3_304
timestamp 1586364061
transform 1 0 29072 0 1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_3_306
timestamp 1586364061
transform 1 0 29256 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_318
timestamp 1586364061
transform 1 0 30360 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_330
timestamp 1586364061
transform 1 0 31464 0 1 3808
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_13.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 33948 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_13.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 33580 0 1 3808
box -38 -48 222 592
use scs8hd_decap_8  FILLER_3_342
timestamp 1586364061
transform 1 0 32568 0 1 3808
box -38 -48 774 592
use scs8hd_decap_3  FILLER_3_350
timestamp 1586364061
transform 1 0 33304 0 1 3808
box -38 -48 314 592
use scs8hd_fill_2  FILLER_3_355
timestamp 1586364061
transform 1 0 33764 0 1 3808
box -38 -48 222 592
use scs8hd_buf_2  _57_
timestamp 1586364061
transform 1 0 35420 0 1 3808
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_73
timestamp 1586364061
transform 1 0 34776 0 1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_13.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 34316 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_359
timestamp 1586364061
transform 1 0 34132 0 1 3808
box -38 -48 222 592
use scs8hd_decap_3  FILLER_3_363
timestamp 1586364061
transform 1 0 34500 0 1 3808
box -38 -48 314 592
use scs8hd_decap_6  FILLER_3_367
timestamp 1586364061
transform 1 0 34868 0 1 3808
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA__57__A
timestamp 1586364061
transform 1 0 35972 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__66__A
timestamp 1586364061
transform 1 0 36340 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_377
timestamp 1586364061
transform 1 0 35788 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_381
timestamp 1586364061
transform 1 0 36156 0 1 3808
box -38 -48 222 592
use scs8hd_decap_12  FILLER_3_385
timestamp 1586364061
transform 1 0 36524 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_3  PHY_7
timestamp 1586364061
transform -1 0 38824 0 1 3808
box -38 -48 314 592
use scs8hd_decap_8  FILLER_3_397
timestamp 1586364061
transform 1 0 37628 0 1 3808
box -38 -48 774 592
use scs8hd_fill_2  FILLER_3_405
timestamp 1586364061
transform 1 0 38364 0 1 3808
box -38 -48 222 592
use scs8hd_buf_2  _44_
timestamp 1586364061
transform 1 0 1380 0 -1 4896
box -38 -48 406 592
use scs8hd_buf_2  _50_
timestamp 1586364061
transform 1 0 2484 0 -1 4896
box -38 -48 406 592
use scs8hd_decap_3  PHY_8
timestamp 1586364061
transform 1 0 1104 0 -1 4896
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_3.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 2024 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_3  FILLER_4_7
timestamp 1586364061
transform 1 0 1748 0 -1 4896
box -38 -48 314 592
use scs8hd_decap_3  FILLER_4_12
timestamp 1586364061
transform 1 0 2208 0 -1 4896
box -38 -48 314 592
use scs8hd_fill_2  FILLER_4_19
timestamp 1586364061
transform 1 0 2852 0 -1 4896
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_74
timestamp 1586364061
transform 1 0 3956 0 -1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_3.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 3036 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_3.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 3404 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_3.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 3772 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_3.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 4232 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_23
timestamp 1586364061
transform 1 0 3220 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_27
timestamp 1586364061
transform 1 0 3588 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_32
timestamp 1586364061
transform 1 0 4048 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_12  FILLER_4_36
timestamp 1586364061
transform 1 0 4416 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_48
timestamp 1586364061
transform 1 0 5520 0 -1 4896
box -38 -48 1142 592
use scs8hd_mux2_2  mux_bottom_ipin_3.mux_l2_in_1_
timestamp 1586364061
transform 1 0 7544 0 -1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_3.mux_l4_in_0__A0
timestamp 1586364061
transform 1 0 7360 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_8  FILLER_4_60
timestamp 1586364061
transform 1 0 6624 0 -1 4896
box -38 -48 774 592
use scs8hd_fill_2  FILLER_4_79
timestamp 1586364061
transform 1 0 8372 0 -1 4896
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_75
timestamp 1586364061
transform 1 0 9568 0 -1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_3.mux_l2_in_3__A0
timestamp 1586364061
transform 1 0 9844 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_4.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 8556 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_8  FILLER_4_83
timestamp 1586364061
transform 1 0 8740 0 -1 4896
box -38 -48 774 592
use scs8hd_fill_1  FILLER_4_91
timestamp 1586364061
transform 1 0 9476 0 -1 4896
box -38 -48 130 592
use scs8hd_fill_2  FILLER_4_93
timestamp 1586364061
transform 1 0 9660 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_4_97
timestamp 1586364061
transform 1 0 10028 0 -1 4896
box -38 -48 406 592
use scs8hd_mux2_2  mux_bottom_ipin_4.mux_l2_in_0_
timestamp 1586364061
transform 1 0 11960 0 -1 4896
box -38 -48 866 592
use scs8hd_mux2_2  mux_bottom_ipin_5.mux_l3_in_1_
timestamp 1586364061
transform 1 0 10396 0 -1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_4.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 11776 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_4.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 11408 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_110
timestamp 1586364061
transform 1 0 11224 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_114
timestamp 1586364061
transform 1 0 11592 0 -1 4896
box -38 -48 222 592
use scs8hd_mux2_2  mux_bottom_ipin_4.mux_l1_in_0_
timestamp 1586364061
transform 1 0 13524 0 -1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_4.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 12972 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_4.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 13340 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_127
timestamp 1586364061
transform 1 0 12788 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_131
timestamp 1586364061
transform 1 0 13156 0 -1 4896
box -38 -48 222 592
use scs8hd_mux2_2  mux_bottom_ipin_5.mux_l2_in_1_
timestamp 1586364061
transform 1 0 15272 0 -1 4896
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_76
timestamp 1586364061
transform 1 0 15180 0 -1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_5.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 14536 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_144
timestamp 1586364061
transform 1 0 14352 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_4_148
timestamp 1586364061
transform 1 0 14720 0 -1 4896
box -38 -48 406 592
use scs8hd_fill_1  FILLER_4_152
timestamp 1586364061
transform 1 0 15088 0 -1 4896
box -38 -48 130 592
use scs8hd_mux2_2  mux_bottom_ipin_5.mux_l1_in_2_
timestamp 1586364061
transform 1 0 16836 0 -1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_5.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 16284 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_5.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 16652 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_163
timestamp 1586364061
transform 1 0 16100 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_167
timestamp 1586364061
transform 1 0 16468 0 -1 4896
box -38 -48 222 592
use scs8hd_mux2_2  mux_bottom_ipin_5.mux_l1_in_0_
timestamp 1586364061
transform 1 0 18400 0 -1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_5.mux_l1_in_1__A0
timestamp 1586364061
transform 1 0 18032 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_4_180
timestamp 1586364061
transform 1 0 17664 0 -1 4896
box -38 -48 406 592
use scs8hd_fill_2  FILLER_4_186
timestamp 1586364061
transform 1 0 18216 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_12  FILLER_4_197
timestamp 1586364061
transform 1 0 19228 0 -1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_77
timestamp 1586364061
transform 1 0 20792 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_4  FILLER_4_209
timestamp 1586364061
transform 1 0 20332 0 -1 4896
box -38 -48 406 592
use scs8hd_fill_1  FILLER_4_213
timestamp 1586364061
transform 1 0 20700 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_6  FILLER_4_215
timestamp 1586364061
transform 1 0 20884 0 -1 4896
box -38 -48 590 592
use scs8hd_mux2_2  mux_bottom_ipin_11.mux_l4_in_0_
timestamp 1586364061
transform 1 0 21988 0 -1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_11.scs8hd_dfxbp_1_3__D
timestamp 1586364061
transform 1 0 21436 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_4_223
timestamp 1586364061
transform 1 0 21620 0 -1 4896
box -38 -48 406 592
use scs8hd_decap_12  FILLER_4_236
timestamp 1586364061
transform 1 0 22816 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_248
timestamp 1586364061
transform 1 0 23920 0 -1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_78
timestamp 1586364061
transform 1 0 26404 0 -1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_12.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 25576 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_6  FILLER_4_260
timestamp 1586364061
transform 1 0 25024 0 -1 4896
box -38 -48 590 592
use scs8hd_decap_6  FILLER_4_268
timestamp 1586364061
transform 1 0 25760 0 -1 4896
box -38 -48 590 592
use scs8hd_fill_1  FILLER_4_274
timestamp 1586364061
transform 1 0 26312 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_8  FILLER_4_276
timestamp 1586364061
transform 1 0 26496 0 -1 4896
box -38 -48 774 592
use scs8hd_mux2_2  mux_bottom_ipin_12.mux_l1_in_2_
timestamp 1586364061
transform 1 0 27508 0 -1 4896
box -38 -48 866 592
use scs8hd_decap_3  FILLER_4_284
timestamp 1586364061
transform 1 0 27232 0 -1 4896
box -38 -48 314 592
use scs8hd_decap_8  FILLER_4_296
timestamp 1586364061
transform 1 0 28336 0 -1 4896
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_12.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 29256 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_12.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 29624 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_12.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 29992 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_304
timestamp 1586364061
transform 1 0 29072 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_308
timestamp 1586364061
transform 1 0 29440 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_312
timestamp 1586364061
transform 1 0 29808 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_12  FILLER_4_316
timestamp 1586364061
transform 1 0 30176 0 -1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_79
timestamp 1586364061
transform 1 0 32016 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_8  FILLER_4_328
timestamp 1586364061
transform 1 0 31280 0 -1 4896
box -38 -48 774 592
use scs8hd_decap_3  FILLER_4_337
timestamp 1586364061
transform 1 0 32108 0 -1 4896
box -38 -48 314 592
use scs8hd_conb_1  _24_
timestamp 1586364061
transform 1 0 32936 0 -1 4896
box -38 -48 314 592
use scs8hd_mux2_2  mux_bottom_ipin_13.mux_l2_in_0_
timestamp 1586364061
transform 1 0 33948 0 -1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_13.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 32752 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_13.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 33396 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_13.mux_l3_in_1__A0
timestamp 1586364061
transform 1 0 32384 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_342
timestamp 1586364061
transform 1 0 32568 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_349
timestamp 1586364061
transform 1 0 33212 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_4_353
timestamp 1586364061
transform 1 0 33580 0 -1 4896
box -38 -48 406 592
use scs8hd_buf_2  _66_
timestamp 1586364061
transform 1 0 35512 0 -1 4896
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_13.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 34960 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_13.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 35328 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_366
timestamp 1586364061
transform 1 0 34776 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_370
timestamp 1586364061
transform 1 0 35144 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_12  FILLER_4_378
timestamp 1586364061
transform 1 0 35880 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_4_390
timestamp 1586364061
transform 1 0 36984 0 -1 4896
box -38 -48 590 592
use scs8hd_fill_1  FILLER_4_396
timestamp 1586364061
transform 1 0 37536 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_3  PHY_9
timestamp 1586364061
transform -1 0 38824 0 -1 4896
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_80
timestamp 1586364061
transform 1 0 37628 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_8  FILLER_4_398
timestamp 1586364061
transform 1 0 37720 0 -1 4896
box -38 -48 774 592
use scs8hd_fill_1  FILLER_4_406
timestamp 1586364061
transform 1 0 38456 0 -1 4896
box -38 -48 130 592
use scs8hd_mux2_2  mux_bottom_ipin_3.mux_l1_in_0_
timestamp 1586364061
transform 1 0 2024 0 1 4896
box -38 -48 866 592
use scs8hd_decap_3  PHY_10
timestamp 1586364061
transform 1 0 1104 0 1 4896
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_3.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 1840 0 1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_5_3
timestamp 1586364061
transform 1 0 1380 0 1 4896
box -38 -48 406 592
use scs8hd_fill_1  FILLER_5_7
timestamp 1586364061
transform 1 0 1748 0 1 4896
box -38 -48 130 592
use scs8hd_fill_2  FILLER_5_19
timestamp 1586364061
transform 1 0 2852 0 1 4896
box -38 -48 222 592
use scs8hd_mux2_2  mux_bottom_ipin_3.mux_l2_in_0_
timestamp 1586364061
transform 1 0 3588 0 1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_3.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 3404 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__48__A
timestamp 1586364061
transform 1 0 4600 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_3.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 3036 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_23
timestamp 1586364061
transform 1 0 3220 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_36
timestamp 1586364061
transform 1 0 4416 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_3.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 5244 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_3.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 5612 0 1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_5_40
timestamp 1586364061
transform 1 0 4784 0 1 4896
box -38 -48 406 592
use scs8hd_fill_1  FILLER_5_44
timestamp 1586364061
transform 1 0 5152 0 1 4896
box -38 -48 130 592
use scs8hd_fill_2  FILLER_5_47
timestamp 1586364061
transform 1 0 5428 0 1 4896
box -38 -48 222 592
use scs8hd_decap_8  FILLER_5_51
timestamp 1586364061
transform 1 0 5796 0 1 4896
box -38 -48 774 592
use scs8hd_fill_2  FILLER_5_59
timestamp 1586364061
transform 1 0 6532 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_66
timestamp 1586364061
transform 1 0 7176 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_62
timestamp 1586364061
transform 1 0 6808 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_3.mux_l4_in_0__A1
timestamp 1586364061
transform 1 0 7360 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_3.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 6992 0 1 4896
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_81
timestamp 1586364061
transform 1 0 6716 0 1 4896
box -38 -48 130 592
use scs8hd_decap_3  FILLER_5_74
timestamp 1586364061
transform 1 0 7912 0 1 4896
box -38 -48 314 592
use scs8hd_fill_2  FILLER_5_70
timestamp 1586364061
transform 1 0 7544 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_3.mux_l4_in_0__S
timestamp 1586364061
transform 1 0 7728 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_4.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 8188 0 1 4896
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_bottom_ipin_4.scs8hd_dfxbp_1_0_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 8372 0 1 4896
box -38 -48 1786 592
use scs8hd_fill_2  FILLER_5_98
timestamp 1586364061
transform 1 0 10120 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_102
timestamp 1586364061
transform 1 0 10488 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_3.mux_l2_in_3__S
timestamp 1586364061
transform 1 0 10672 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_3.mux_l2_in_3__A1
timestamp 1586364061
transform 1 0 10304 0 1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_5_106
timestamp 1586364061
transform 1 0 10856 0 1 4896
box -38 -48 406 592
use scs8hd_fill_2  FILLER_5_113
timestamp 1586364061
transform 1 0 11500 0 1 4896
box -38 -48 222 592
use scs8hd_fill_1  FILLER_5_110
timestamp 1586364061
transform 1 0 11224 0 1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_4.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 11316 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_117
timestamp 1586364061
transform 1 0 11868 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_4.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 11684 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_4.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 12052 0 1 4896
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_bottom_ipin_4.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 12420 0 1 4896
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_82
timestamp 1586364061
transform 1 0 12328 0 1 4896
box -38 -48 130 592
use scs8hd_fill_1  FILLER_5_121
timestamp 1586364061
transform 1 0 12236 0 1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_4.scs8hd_dfxbp_1_3__CLK
timestamp 1586364061
transform 1 0 15456 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_4.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 14352 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_4.scs8hd_dfxbp_1_3__D
timestamp 1586364061
transform 1 0 15088 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_4.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 14720 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_142
timestamp 1586364061
transform 1 0 14168 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_146
timestamp 1586364061
transform 1 0 14536 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_150
timestamp 1586364061
transform 1 0 14904 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_154
timestamp 1586364061
transform 1 0 15272 0 1 4896
box -38 -48 222 592
use scs8hd_decap_3  FILLER_5_158
timestamp 1586364061
transform 1 0 15640 0 1 4896
box -38 -48 314 592
use scs8hd_mux2_2  mux_bottom_ipin_5.mux_l2_in_0_
timestamp 1586364061
transform 1 0 15916 0 1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_5.mux_l1_in_1__S
timestamp 1586364061
transform 1 0 17388 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_8.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 17020 0 1 4896
box -38 -48 222 592
use scs8hd_decap_3  FILLER_5_170
timestamp 1586364061
transform 1 0 16744 0 1 4896
box -38 -48 314 592
use scs8hd_fill_2  FILLER_5_175
timestamp 1586364061
transform 1 0 17204 0 1 4896
box -38 -48 222 592
use scs8hd_mux2_2  mux_bottom_ipin_5.mux_l1_in_1_
timestamp 1586364061
transform 1 0 18032 0 1 4896
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_83
timestamp 1586364061
transform 1 0 17940 0 1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_5.mux_l1_in_1__A1
timestamp 1586364061
transform 1 0 17756 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_8.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 19044 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_179
timestamp 1586364061
transform 1 0 17572 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_193
timestamp 1586364061
transform 1 0 18860 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_197
timestamp 1586364061
transform 1 0 19228 0 1 4896
box -38 -48 222 592
use scs8hd_mux2_2  mux_bottom_ipin_11.mux_l3_in_1_
timestamp 1586364061
transform 1 0 21160 0 1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_11.mux_l3_in_1__S
timestamp 1586364061
transform 1 0 20976 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_11.mux_l3_in_1__A1
timestamp 1586364061
transform 1 0 20608 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_11.mux_l3_in_1__A0
timestamp 1586364061
transform 1 0 20240 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_8.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 19412 0 1 4896
box -38 -48 222 592
use scs8hd_decap_6  FILLER_5_201
timestamp 1586364061
transform 1 0 19596 0 1 4896
box -38 -48 590 592
use scs8hd_fill_1  FILLER_5_207
timestamp 1586364061
transform 1 0 20148 0 1 4896
box -38 -48 130 592
use scs8hd_fill_2  FILLER_5_210
timestamp 1586364061
transform 1 0 20424 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_214
timestamp 1586364061
transform 1 0 20792 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_11.scs8hd_dfxbp_1_3__CLK
timestamp 1586364061
transform 1 0 22172 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_227
timestamp 1586364061
transform 1 0 21988 0 1 4896
box -38 -48 222 592
use scs8hd_decap_12  FILLER_5_231
timestamp 1586364061
transform 1 0 22356 0 1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_84
timestamp 1586364061
transform 1 0 23552 0 1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_12.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 23920 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_12.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 24288 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_12.mux_l2_in_2__S
timestamp 1586364061
transform 1 0 24656 0 1 4896
box -38 -48 222 592
use scs8hd_fill_1  FILLER_5_243
timestamp 1586364061
transform 1 0 23460 0 1 4896
box -38 -48 130 592
use scs8hd_decap_3  FILLER_5_245
timestamp 1586364061
transform 1 0 23644 0 1 4896
box -38 -48 314 592
use scs8hd_fill_2  FILLER_5_250
timestamp 1586364061
transform 1 0 24104 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_254
timestamp 1586364061
transform 1 0 24472 0 1 4896
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_bottom_ipin_12.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 25576 0 1 4896
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_12.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 25392 0 1 4896
box -38 -48 222 592
use scs8hd_decap_6  FILLER_5_258
timestamp 1586364061
transform 1 0 24840 0 1 4896
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_12.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 27600 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_12.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 27968 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_12.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 28336 0 1 4896
box -38 -48 222 592
use scs8hd_decap_3  FILLER_5_285
timestamp 1586364061
transform 1 0 27324 0 1 4896
box -38 -48 314 592
use scs8hd_fill_2  FILLER_5_290
timestamp 1586364061
transform 1 0 27784 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_294
timestamp 1586364061
transform 1 0 28152 0 1 4896
box -38 -48 222 592
use scs8hd_mux2_2  mux_bottom_ipin_12.mux_l3_in_0_
timestamp 1586364061
transform 1 0 29256 0 1 4896
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_85
timestamp 1586364061
transform 1 0 29164 0 1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_12.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 28980 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_12.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 30268 0 1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_5_298
timestamp 1586364061
transform 1 0 28520 0 1 4896
box -38 -48 406 592
use scs8hd_fill_1  FILLER_5_302
timestamp 1586364061
transform 1 0 28888 0 1 4896
box -38 -48 130 592
use scs8hd_fill_2  FILLER_5_315
timestamp 1586364061
transform 1 0 30084 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_12.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 30636 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_13.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 32016 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_13.mux_l3_in_1__A1
timestamp 1586364061
transform 1 0 31648 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_319
timestamp 1586364061
transform 1 0 30452 0 1 4896
box -38 -48 222 592
use scs8hd_decap_8  FILLER_5_323
timestamp 1586364061
transform 1 0 30820 0 1 4896
box -38 -48 774 592
use scs8hd_fill_1  FILLER_5_331
timestamp 1586364061
transform 1 0 31556 0 1 4896
box -38 -48 130 592
use scs8hd_fill_2  FILLER_5_334
timestamp 1586364061
transform 1 0 31832 0 1 4896
box -38 -48 222 592
use scs8hd_mux2_2  mux_bottom_ipin_13.mux_l3_in_1_
timestamp 1586364061
transform 1 0 32568 0 1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_13.mux_l1_in_1__A0
timestamp 1586364061
transform 1 0 33856 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_13.mux_l3_in_1__S
timestamp 1586364061
transform 1 0 32384 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_338
timestamp 1586364061
transform 1 0 32200 0 1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_5_351
timestamp 1586364061
transform 1 0 33396 0 1 4896
box -38 -48 406 592
use scs8hd_fill_1  FILLER_5_355
timestamp 1586364061
transform 1 0 33764 0 1 4896
box -38 -48 130 592
use scs8hd_mux2_2  mux_bottom_ipin_13.mux_l1_in_0_
timestamp 1586364061
transform 1 0 34868 0 1 4896
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_86
timestamp 1586364061
transform 1 0 34776 0 1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_13.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 34592 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_13.mux_l1_in_1__A1
timestamp 1586364061
transform 1 0 34224 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_358
timestamp 1586364061
transform 1 0 34040 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_362
timestamp 1586364061
transform 1 0 34408 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_376
timestamp 1586364061
transform 1 0 35696 0 1 4896
box -38 -48 222 592
use scs8hd_buf_2  _56_
timestamp 1586364061
transform 1 0 36432 0 1 4896
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__56__A
timestamp 1586364061
transform 1 0 36984 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__70__A
timestamp 1586364061
transform 1 0 35880 0 1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_5_380
timestamp 1586364061
transform 1 0 36064 0 1 4896
box -38 -48 406 592
use scs8hd_fill_2  FILLER_5_388
timestamp 1586364061
transform 1 0 36800 0 1 4896
box -38 -48 222 592
use scs8hd_decap_12  FILLER_5_392
timestamp 1586364061
transform 1 0 37168 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_3  PHY_11
timestamp 1586364061
transform -1 0 38824 0 1 4896
box -38 -48 314 592
use scs8hd_decap_3  FILLER_5_404
timestamp 1586364061
transform 1 0 38272 0 1 4896
box -38 -48 314 592
use scs8hd_dfxbp_1  mem_bottom_ipin_2.scs8hd_dfxbp_1_3_
timestamp 1586364061
transform 1 0 1748 0 1 5984
box -38 -48 1786 592
use scs8hd_dfxbp_1  mem_bottom_ipin_3.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 1472 0 -1 5984
box -38 -48 1786 592
use scs8hd_decap_3  PHY_12
timestamp 1586364061
transform 1 0 1104 0 -1 5984
box -38 -48 314 592
use scs8hd_decap_3  PHY_14
timestamp 1586364061
transform 1 0 1104 0 1 5984
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_2.scs8hd_dfxbp_1_3__CLK
timestamp 1586364061
transform 1 0 1564 0 1 5984
box -38 -48 222 592
use scs8hd_fill_1  FILLER_6_3
timestamp 1586364061
transform 1 0 1380 0 -1 5984
box -38 -48 130 592
use scs8hd_fill_2  FILLER_7_3
timestamp 1586364061
transform 1 0 1380 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_26
timestamp 1586364061
transform 1 0 3496 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_27
timestamp 1586364061
transform 1 0 3588 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_23
timestamp 1586364061
transform 1 0 3220 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l3_in_1__A0
timestamp 1586364061
transform 1 0 3772 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_2.scs8hd_dfxbp_1_3__D
timestamp 1586364061
transform 1 0 3404 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_3.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 3680 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_30
timestamp 1586364061
transform 1 0 3864 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_36
timestamp 1586364061
transform 1 0 4416 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_3.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 4600 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__51__A
timestamp 1586364061
transform 1 0 4048 0 1 5984
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_87
timestamp 1586364061
transform 1 0 3956 0 -1 5984
box -38 -48 130 592
use scs8hd_buf_2  _48_
timestamp 1586364061
transform 1 0 4048 0 -1 5984
box -38 -48 406 592
use scs8hd_dfxbp_1  mem_bottom_ipin_3.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 4232 0 1 5984
box -38 -48 1786 592
use scs8hd_dfxbp_1  mem_bottom_ipin_3.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 5244 0 -1 5984
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 6164 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 6532 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 5060 0 -1 5984
box -38 -48 222 592
use scs8hd_decap_3  FILLER_6_40
timestamp 1586364061
transform 1 0 4784 0 -1 5984
box -38 -48 314 592
use scs8hd_fill_2  FILLER_7_53
timestamp 1586364061
transform 1 0 5980 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_57
timestamp 1586364061
transform 1 0 6348 0 1 5984
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_bottom_ipin_3.scs8hd_dfxbp_1_3_
timestamp 1586364061
transform 1 0 7360 0 1 5984
box -38 -48 1786 592
use scs8hd_mux2_2  mux_bottom_ipin_3.mux_l4_in_0_
timestamp 1586364061
transform 1 0 7728 0 -1 5984
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_94
timestamp 1586364061
transform 1 0 6716 0 1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_3.scs8hd_dfxbp_1_3__CLK
timestamp 1586364061
transform 1 0 7176 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_3.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 7176 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_3.scs8hd_dfxbp_1_3__D
timestamp 1586364061
transform 1 0 7544 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_64
timestamp 1586364061
transform 1 0 6992 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_68
timestamp 1586364061
transform 1 0 7360 0 -1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_7_62
timestamp 1586364061
transform 1 0 6808 0 1 5984
box -38 -48 406 592
use scs8hd_fill_2  FILLER_7_87
timestamp 1586364061
transform 1 0 9108 0 1 5984
box -38 -48 222 592
use scs8hd_fill_1  FILLER_6_89
timestamp 1586364061
transform 1 0 9292 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_8  FILLER_6_81
timestamp 1586364061
transform 1 0 8556 0 -1 5984
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_3.mux_l2_in_2__A1
timestamp 1586364061
transform 1 0 9292 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_91
timestamp 1586364061
transform 1 0 9476 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_3.mux_l3_in_1__A1
timestamp 1586364061
transform 1 0 9384 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_3.mux_l2_in_2__A0
timestamp 1586364061
transform 1 0 9660 0 1 5984
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_88
timestamp 1586364061
transform 1 0 9568 0 -1 5984
box -38 -48 130 592
use scs8hd_mux2_2  mux_bottom_ipin_3.mux_l3_in_1_
timestamp 1586364061
transform 1 0 9844 0 1 5984
box -38 -48 866 592
use scs8hd_mux2_2  mux_bottom_ipin_3.mux_l2_in_3_
timestamp 1586364061
transform 1 0 9660 0 -1 5984
box -38 -48 866 592
use scs8hd_decap_3  FILLER_7_108
timestamp 1586364061
transform 1 0 11040 0 1 5984
box -38 -48 314 592
use scs8hd_fill_2  FILLER_7_104
timestamp 1586364061
transform 1 0 10672 0 1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_6_106
timestamp 1586364061
transform 1 0 10856 0 -1 5984
box -38 -48 406 592
use scs8hd_fill_2  FILLER_6_102
timestamp 1586364061
transform 1 0 10488 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_3.mux_l3_in_1__S
timestamp 1586364061
transform 1 0 10672 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_3.mux_l2_in_2__S
timestamp 1586364061
transform 1 0 10856 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_118
timestamp 1586364061
transform 1 0 11960 0 1 5984
box -38 -48 222 592
use scs8hd_decap_3  FILLER_7_113
timestamp 1586364061
transform 1 0 11500 0 1 5984
box -38 -48 314 592
use scs8hd_fill_2  FILLER_6_117
timestamp 1586364061
transform 1 0 11868 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_113
timestamp 1586364061
transform 1 0 11500 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_1  FILLER_6_110
timestamp 1586364061
transform 1 0 11224 0 -1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_5.scs8hd_dfxbp_1_3__D
timestamp 1586364061
transform 1 0 11684 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_5.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 11316 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_5.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 11316 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_4.mux_l1_in_1__A0
timestamp 1586364061
transform 1 0 11776 0 1 5984
box -38 -48 222 592
use scs8hd_mux2_2  mux_bottom_ipin_4.mux_l2_in_1_
timestamp 1586364061
transform 1 0 12052 0 -1 5984
box -38 -48 866 592
use scs8hd_fill_2  FILLER_6_128
timestamp 1586364061
transform 1 0 12880 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_4.mux_l1_in_1__A1
timestamp 1586364061
transform 1 0 12144 0 1 5984
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_95
timestamp 1586364061
transform 1 0 12328 0 1 5984
box -38 -48 130 592
use scs8hd_mux2_2  mux_bottom_ipin_4.mux_l1_in_1_
timestamp 1586364061
transform 1 0 12420 0 1 5984
box -38 -48 866 592
use scs8hd_decap_6  FILLER_7_136
timestamp 1586364061
transform 1 0 13616 0 1 5984
box -38 -48 590 592
use scs8hd_fill_2  FILLER_7_132
timestamp 1586364061
transform 1 0 13248 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_132
timestamp 1586364061
transform 1 0 13248 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_4.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 13432 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_4.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 13064 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_4.mux_l1_in_1__S
timestamp 1586364061
transform 1 0 13432 0 1 5984
box -38 -48 222 592
use scs8hd_mux2_2  mux_bottom_ipin_4.mux_l3_in_0_
timestamp 1586364061
transform 1 0 13616 0 -1 5984
box -38 -48 866 592
use scs8hd_dfxbp_1  mem_bottom_ipin_4.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 14352 0 1 5984
box -38 -48 1786 592
use scs8hd_dfxbp_1  mem_bottom_ipin_4.scs8hd_dfxbp_1_3_
timestamp 1586364061
transform 1 0 15456 0 -1 5984
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_89
timestamp 1586364061
transform 1 0 15180 0 -1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_4.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 14168 0 1 5984
box -38 -48 222 592
use scs8hd_decap_8  FILLER_6_145
timestamp 1586364061
transform 1 0 14444 0 -1 5984
box -38 -48 774 592
use scs8hd_fill_2  FILLER_6_154
timestamp 1586364061
transform 1 0 15272 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_5.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 16744 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_5.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 17112 0 1 5984
box -38 -48 222 592
use scs8hd_decap_8  FILLER_6_175
timestamp 1586364061
transform 1 0 17204 0 -1 5984
box -38 -48 774 592
use scs8hd_decap_6  FILLER_7_163
timestamp 1586364061
transform 1 0 16100 0 1 5984
box -38 -48 590 592
use scs8hd_fill_1  FILLER_7_169
timestamp 1586364061
transform 1 0 16652 0 1 5984
box -38 -48 130 592
use scs8hd_fill_2  FILLER_7_172
timestamp 1586364061
transform 1 0 16928 0 1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_7_176
timestamp 1586364061
transform 1 0 17296 0 1 5984
box -38 -48 406 592
use scs8hd_fill_2  FILLER_7_188
timestamp 1586364061
transform 1 0 18400 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_184
timestamp 1586364061
transform 1 0 18032 0 1 5984
box -38 -48 222 592
use scs8hd_fill_1  FILLER_7_182
timestamp 1586364061
transform 1 0 17848 0 1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_8.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 17664 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_5.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 18216 0 1 5984
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_96
timestamp 1586364061
transform 1 0 17940 0 1 5984
box -38 -48 130 592
use scs8hd_mux2_2  mux_bottom_ipin_8.mux_l2_in_0_
timestamp 1586364061
transform 1 0 17940 0 -1 5984
box -38 -48 866 592
use scs8hd_fill_2  FILLER_7_196
timestamp 1586364061
transform 1 0 19136 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_192
timestamp 1586364061
transform 1 0 18768 0 1 5984
box -38 -48 222 592
use scs8hd_decap_8  FILLER_6_192
timestamp 1586364061
transform 1 0 18768 0 -1 5984
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_11.mux_l2_in_3__A0
timestamp 1586364061
transform 1 0 18584 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_11.mux_l2_in_3__A1
timestamp 1586364061
transform 1 0 18952 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_8.mux_l2_in_2__A0
timestamp 1586364061
transform 1 0 19320 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_206
timestamp 1586364061
transform 1 0 20056 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_202
timestamp 1586364061
transform 1 0 19688 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_8.mux_l2_in_2__S
timestamp 1586364061
transform 1 0 20240 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_11.mux_l2_in_3__S
timestamp 1586364061
transform 1 0 19872 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_8.mux_l2_in_2__A1
timestamp 1586364061
transform 1 0 19504 0 -1 5984
box -38 -48 222 592
use scs8hd_mux2_2  mux_bottom_ipin_8.mux_l2_in_2_
timestamp 1586364061
transform 1 0 19504 0 1 5984
box -38 -48 866 592
use scs8hd_fill_2  FILLER_7_213
timestamp 1586364061
transform 1 0 20700 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_209
timestamp 1586364061
transform 1 0 20332 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_215
timestamp 1586364061
transform 1 0 20884 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_210
timestamp 1586364061
transform 1 0 20424 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_11.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 20608 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_11.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 21068 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_11.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 20516 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_11.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 20884 0 1 5984
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_90
timestamp 1586364061
transform 1 0 20792 0 -1 5984
box -38 -48 130 592
use scs8hd_dfxbp_1  mem_bottom_ipin_11.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 21068 0 1 5984
box -38 -48 1786 592
use scs8hd_dfxbp_1  mem_bottom_ipin_11.scs8hd_dfxbp_1_3_
timestamp 1586364061
transform 1 0 21436 0 -1 5984
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_11.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 23000 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_219
timestamp 1586364061
transform 1 0 21252 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_236
timestamp 1586364061
transform 1 0 22816 0 1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_7_245
timestamp 1586364061
transform 1 0 23644 0 1 5984
box -38 -48 406 592
use scs8hd_fill_2  FILLER_7_240
timestamp 1586364061
transform 1 0 23184 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_244
timestamp 1586364061
transform 1 0 23552 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_240
timestamp 1586364061
transform 1 0 23184 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_11.mux_l2_in_2__S
timestamp 1586364061
transform 1 0 23736 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_11.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 23368 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_11.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 23368 0 1 5984
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_97
timestamp 1586364061
transform 1 0 23552 0 1 5984
box -38 -48 130 592
use scs8hd_fill_1  FILLER_7_252
timestamp 1586364061
transform 1 0 24288 0 1 5984
box -38 -48 130 592
use scs8hd_fill_1  FILLER_7_249
timestamp 1586364061
transform 1 0 24012 0 1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_11.mux_l2_in_2__A0
timestamp 1586364061
transform 1 0 24104 0 1 5984
box -38 -48 222 592
use scs8hd_mux2_2  mux_bottom_ipin_12.mux_l2_in_2_
timestamp 1586364061
transform 1 0 24380 0 1 5984
box -38 -48 866 592
use scs8hd_dfxbp_1  mem_bottom_ipin_12.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 23920 0 -1 5984
box -38 -48 1786 592
use scs8hd_fill_2  FILLER_7_266
timestamp 1586364061
transform 1 0 25576 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_262
timestamp 1586364061
transform 1 0 25208 0 1 5984
box -38 -48 222 592
use scs8hd_decap_3  FILLER_6_267
timestamp 1586364061
transform 1 0 25668 0 -1 5984
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_12.mux_l2_in_2__A0
timestamp 1586364061
transform 1 0 25392 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_276
timestamp 1586364061
transform 1 0 26496 0 -1 5984
box -38 -48 222 592
use scs8hd_decap_3  FILLER_6_272
timestamp 1586364061
transform 1 0 26128 0 -1 5984
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_12.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 25944 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_12.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 25760 0 1 5984
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_91
timestamp 1586364061
transform 1 0 26404 0 -1 5984
box -38 -48 130 592
use scs8hd_mux2_2  mux_bottom_ipin_12.mux_l2_in_1_
timestamp 1586364061
transform 1 0 25944 0 1 5984
box -38 -48 866 592
use scs8hd_fill_2  FILLER_7_283
timestamp 1586364061
transform 1 0 27140 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_279
timestamp 1586364061
transform 1 0 26772 0 1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_6_284
timestamp 1586364061
transform 1 0 27232 0 -1 5984
box -38 -48 406 592
use scs8hd_fill_2  FILLER_6_280
timestamp 1586364061
transform 1 0 26864 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_12.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 27048 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_12.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 26680 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_12.mux_l1_in_1__A0
timestamp 1586364061
transform 1 0 26956 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_12.mux_l1_in_1__A1
timestamp 1586364061
transform 1 0 27324 0 1 5984
box -38 -48 222 592
use scs8hd_mux2_2  mux_bottom_ipin_12.mux_l1_in_1_
timestamp 1586364061
transform 1 0 27508 0 1 5984
box -38 -48 866 592
use scs8hd_fill_2  FILLER_7_296
timestamp 1586364061
transform 1 0 28336 0 1 5984
box -38 -48 222 592
use scs8hd_decap_8  FILLER_6_297
timestamp 1586364061
transform 1 0 28428 0 -1 5984
box -38 -48 774 592
use scs8hd_mux2_2  mux_bottom_ipin_12.mux_l1_in_0_
timestamp 1586364061
transform 1 0 27600 0 -1 5984
box -38 -48 866 592
use scs8hd_fill_2  FILLER_7_306
timestamp 1586364061
transform 1 0 29256 0 1 5984
box -38 -48 222 592
use scs8hd_fill_1  FILLER_7_304
timestamp 1586364061
transform 1 0 29072 0 1 5984
box -38 -48 130 592
use scs8hd_decap_4  FILLER_7_300
timestamp 1586364061
transform 1 0 28704 0 1 5984
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_12.mux_l1_in_1__S
timestamp 1586364061
transform 1 0 28520 0 1 5984
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_98
timestamp 1586364061
transform 1 0 29164 0 1 5984
box -38 -48 130 592
use scs8hd_mux2_2  mux_bottom_ipin_12.mux_l2_in_0_
timestamp 1586364061
transform 1 0 29164 0 -1 5984
box -38 -48 866 592
use scs8hd_decap_3  FILLER_7_314
timestamp 1586364061
transform 1 0 29992 0 1 5984
box -38 -48 314 592
use scs8hd_fill_2  FILLER_7_310
timestamp 1586364061
transform 1 0 29624 0 1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_6_314
timestamp 1586364061
transform 1 0 29992 0 -1 5984
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_12.scs8hd_dfxbp_1_3__D
timestamp 1586364061
transform 1 0 29808 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_12.scs8hd_dfxbp_1_3__CLK
timestamp 1586364061
transform 1 0 29440 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_13.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 30268 0 1 5984
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_bottom_ipin_13.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 30452 0 1 5984
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_92
timestamp 1586364061
transform 1 0 32016 0 -1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_13.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 30452 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_12.mux_l4_in_0__A0
timestamp 1586364061
transform 1 0 31832 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_1  FILLER_6_318
timestamp 1586364061
transform 1 0 30360 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_321
timestamp 1586364061
transform 1 0 30636 0 -1 5984
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_6_333
timestamp 1586364061
transform 1 0 31740 0 -1 5984
box -38 -48 130 592
use scs8hd_fill_2  FILLER_6_337
timestamp 1586364061
transform 1 0 32108 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_1  FILLER_7_346
timestamp 1586364061
transform 1 0 32936 0 1 5984
box -38 -48 130 592
use scs8hd_decap_4  FILLER_7_342
timestamp 1586364061
transform 1 0 32568 0 1 5984
box -38 -48 406 592
use scs8hd_fill_2  FILLER_7_338
timestamp 1586364061
transform 1 0 32200 0 1 5984
box -38 -48 222 592
use scs8hd_decap_3  FILLER_6_341
timestamp 1586364061
transform 1 0 32476 0 -1 5984
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_12.mux_l4_in_0__A1
timestamp 1586364061
transform 1 0 32292 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_12.mux_l4_in_0__S
timestamp 1586364061
transform 1 0 32384 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_13.mux_l1_in_2__A1
timestamp 1586364061
transform 1 0 33028 0 1 5984
box -38 -48 222 592
use scs8hd_mux2_2  mux_bottom_ipin_13.mux_l3_in_0_
timestamp 1586364061
transform 1 0 32752 0 -1 5984
box -38 -48 866 592
use scs8hd_decap_6  FILLER_6_353
timestamp 1586364061
transform 1 0 33580 0 -1 5984
box -38 -48 590 592
use scs8hd_mux2_2  mux_bottom_ipin_13.mux_l1_in_2_
timestamp 1586364061
transform 1 0 33212 0 1 5984
box -38 -48 866 592
use scs8hd_fill_1  FILLER_7_365
timestamp 1586364061
transform 1 0 34684 0 1 5984
box -38 -48 130 592
use scs8hd_fill_1  FILLER_7_362
timestamp 1586364061
transform 1 0 34408 0 1 5984
box -38 -48 130 592
use scs8hd_decap_4  FILLER_7_358
timestamp 1586364061
transform 1 0 34040 0 1 5984
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_13.mux_l1_in_1__S
timestamp 1586364061
transform 1 0 34132 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_13.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 34500 0 1 5984
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_99
timestamp 1586364061
transform 1 0 34776 0 1 5984
box -38 -48 130 592
use scs8hd_mux2_2  mux_bottom_ipin_13.mux_l1_in_1_
timestamp 1586364061
transform 1 0 34316 0 -1 5984
box -38 -48 866 592
use scs8hd_fill_2  FILLER_6_374
timestamp 1586364061
transform 1 0 35512 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_370
timestamp 1586364061
transform 1 0 35144 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_13.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 35696 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_13.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 35328 0 -1 5984
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_bottom_ipin_13.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 34868 0 1 5984
box -38 -48 1786 592
use scs8hd_buf_2  _67_
timestamp 1586364061
transform 1 0 37352 0 1 5984
box -38 -48 406 592
use scs8hd_buf_2  _70_
timestamp 1586364061
transform 1 0 35880 0 -1 5984
box -38 -48 406 592
use scs8hd_decap_12  FILLER_6_382
timestamp 1586364061
transform 1 0 36248 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_6_394
timestamp 1586364061
transform 1 0 37352 0 -1 5984
box -38 -48 314 592
use scs8hd_decap_8  FILLER_7_386
timestamp 1586364061
transform 1 0 36616 0 1 5984
box -38 -48 774 592
use scs8hd_decap_3  PHY_13
timestamp 1586364061
transform -1 0 38824 0 -1 5984
box -38 -48 314 592
use scs8hd_decap_3  PHY_15
timestamp 1586364061
transform -1 0 38824 0 1 5984
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_93
timestamp 1586364061
transform 1 0 37628 0 -1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__67__A
timestamp 1586364061
transform 1 0 37904 0 1 5984
box -38 -48 222 592
use scs8hd_decap_8  FILLER_6_398
timestamp 1586364061
transform 1 0 37720 0 -1 5984
box -38 -48 774 592
use scs8hd_fill_1  FILLER_6_406
timestamp 1586364061
transform 1 0 38456 0 -1 5984
box -38 -48 130 592
use scs8hd_fill_2  FILLER_7_398
timestamp 1586364061
transform 1 0 37720 0 1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_7_402
timestamp 1586364061
transform 1 0 38088 0 1 5984
box -38 -48 406 592
use scs8hd_fill_1  FILLER_7_406
timestamp 1586364061
transform 1 0 38456 0 1 5984
box -38 -48 130 592
use scs8hd_mux2_2  mux_bottom_ipin_2.mux_l3_in_1_
timestamp 1586364061
transform 1 0 1564 0 -1 7072
box -38 -48 866 592
use scs8hd_decap_3  PHY_16
timestamp 1586364061
transform 1 0 1104 0 -1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l2_in_2__A1
timestamp 1586364061
transform 1 0 2576 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_3
timestamp 1586364061
transform 1 0 1380 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_14
timestamp 1586364061
transform 1 0 2392 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_18
timestamp 1586364061
transform 1 0 2760 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_22
timestamp 1586364061
transform 1 0 3128 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l3_in_1__S
timestamp 1586364061
transform 1 0 3312 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l2_in_2__S
timestamp 1586364061
transform 1 0 2944 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_26
timestamp 1586364061
transform 1 0 3496 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l3_in_1__A1
timestamp 1586364061
transform 1 0 3680 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_1  FILLER_8_30
timestamp 1586364061
transform 1 0 3864 0 -1 7072
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_100
timestamp 1586364061
transform 1 0 3956 0 -1 7072
box -38 -48 130 592
use scs8hd_buf_2  _51_
timestamp 1586364061
transform 1 0 4048 0 -1 7072
box -38 -48 406 592
use scs8hd_decap_3  FILLER_8_36
timestamp 1586364061
transform 1 0 4416 0 -1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_2.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 4692 0 -1 7072
box -38 -48 222 592
use scs8hd_mux2_2  mux_bottom_ipin_2.mux_l2_in_0_
timestamp 1586364061
transform 1 0 5428 0 -1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_2.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 5060 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_3.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 6440 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_41
timestamp 1586364061
transform 1 0 4876 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_45
timestamp 1586364061
transform 1 0 5244 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_56
timestamp 1586364061
transform 1 0 6256 0 -1 7072
box -38 -48 222 592
use scs8hd_mux2_2  mux_bottom_ipin_3.mux_l3_in_0_
timestamp 1586364061
transform 1 0 6992 0 -1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_2.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 8004 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 6808 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_60
timestamp 1586364061
transform 1 0 6624 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_73
timestamp 1586364061
transform 1 0 7820 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_8_77
timestamp 1586364061
transform 1 0 8188 0 -1 7072
box -38 -48 406 592
use scs8hd_conb_1  _28_
timestamp 1586364061
transform 1 0 8556 0 -1 7072
box -38 -48 314 592
use scs8hd_mux2_2  mux_bottom_ipin_3.mux_l2_in_2_
timestamp 1586364061
transform 1 0 9660 0 -1 7072
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_101
timestamp 1586364061
transform 1 0 9568 0 -1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_3.mux_l3_in_1__A0
timestamp 1586364061
transform 1 0 9384 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_6  FILLER_8_84
timestamp 1586364061
transform 1 0 8832 0 -1 7072
box -38 -48 590 592
use scs8hd_dfxbp_1  mem_bottom_ipin_5.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 11316 0 -1 7072
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_4.mux_l2_in_3__A0
timestamp 1586364061
transform 1 0 10764 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_4.mux_l2_in_3__S
timestamp 1586364061
transform 1 0 11132 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_3  FILLER_8_102
timestamp 1586364061
transform 1 0 10488 0 -1 7072
box -38 -48 314 592
use scs8hd_fill_2  FILLER_8_107
timestamp 1586364061
transform 1 0 10948 0 -1 7072
box -38 -48 222 592
use scs8hd_conb_1  _29_
timestamp 1586364061
transform 1 0 13800 0 -1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_6.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 13248 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_6.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 13616 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_130
timestamp 1586364061
transform 1 0 13064 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_134
timestamp 1586364061
transform 1 0 13432 0 -1 7072
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_102
timestamp 1586364061
transform 1 0 15180 0 -1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_4.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 14352 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_3  FILLER_8_141
timestamp 1586364061
transform 1 0 14076 0 -1 7072
box -38 -48 314 592
use scs8hd_decap_6  FILLER_8_146
timestamp 1586364061
transform 1 0 14536 0 -1 7072
box -38 -48 590 592
use scs8hd_fill_1  FILLER_8_152
timestamp 1586364061
transform 1 0 15088 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_8  FILLER_8_154
timestamp 1586364061
transform 1 0 15272 0 -1 7072
box -38 -48 774 592
use scs8hd_dfxbp_1  mem_bottom_ipin_5.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 16744 0 -1 7072
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_8.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 16376 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_8.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 16008 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_164
timestamp 1586364061
transform 1 0 16192 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_168
timestamp 1586364061
transform 1 0 16560 0 -1 7072
box -38 -48 222 592
use scs8hd_mux2_2  mux_bottom_ipin_11.mux_l2_in_3_
timestamp 1586364061
transform 1 0 19228 0 -1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_5.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 18676 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_189
timestamp 1586364061
transform 1 0 18492 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_8_193
timestamp 1586364061
transform 1 0 18860 0 -1 7072
box -38 -48 406 592
use scs8hd_mux2_2  mux_bottom_ipin_11.mux_l2_in_1_
timestamp 1586364061
transform 1 0 20976 0 -1 7072
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_103
timestamp 1586364061
transform 1 0 20792 0 -1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_11.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 20608 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_6  FILLER_8_206
timestamp 1586364061
transform 1 0 20056 0 -1 7072
box -38 -48 590 592
use scs8hd_fill_1  FILLER_8_215
timestamp 1586364061
transform 1 0 20884 0 -1 7072
box -38 -48 130 592
use scs8hd_mux2_2  mux_bottom_ipin_11.mux_l1_in_0_
timestamp 1586364061
transform 1 0 22540 0 -1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_11.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 21988 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_11.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 22356 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_225
timestamp 1586364061
transform 1 0 21804 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_229
timestamp 1586364061
transform 1 0 22172 0 -1 7072
box -38 -48 222 592
use scs8hd_mux2_2  mux_bottom_ipin_11.mux_l2_in_2_
timestamp 1586364061
transform 1 0 24104 0 -1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_11.mux_l2_in_2__A1
timestamp 1586364061
transform 1 0 23920 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_6  FILLER_8_242
timestamp 1586364061
transform 1 0 23368 0 -1 7072
box -38 -48 590 592
use scs8hd_fill_2  FILLER_8_259
timestamp 1586364061
transform 1 0 24932 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_263
timestamp 1586364061
transform 1 0 25300 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_12.mux_l2_in_2__A1
timestamp 1586364061
transform 1 0 25116 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_10.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 25484 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_267
timestamp 1586364061
transform 1 0 25668 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_12.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 25852 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_271
timestamp 1586364061
transform 1 0 26036 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_10.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 26220 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_276
timestamp 1586364061
transform 1 0 26496 0 -1 7072
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_104
timestamp 1586364061
transform 1 0 26404 0 -1 7072
box -38 -48 130 592
use scs8hd_dfxbp_1  mem_bottom_ipin_12.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 26680 0 -1 7072
box -38 -48 1786 592
use scs8hd_decap_6  FILLER_8_297
timestamp 1586364061
transform 1 0 28428 0 -1 7072
box -38 -48 590 592
use scs8hd_dfxbp_1  mem_bottom_ipin_12.scs8hd_dfxbp_1_3_
timestamp 1586364061
transform 1 0 29164 0 -1 7072
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_10.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 28980 0 -1 7072
box -38 -48 222 592
use scs8hd_mux2_2  mux_bottom_ipin_12.mux_l4_in_0_
timestamp 1586364061
transform 1 0 32108 0 -1 7072
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_105
timestamp 1586364061
transform 1 0 32016 0 -1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_12.mux_l3_in_1__S
timestamp 1586364061
transform 1 0 31096 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_12.mux_l3_in_1__A0
timestamp 1586364061
transform 1 0 31464 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_13.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 31832 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_324
timestamp 1586364061
transform 1 0 30912 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_328
timestamp 1586364061
transform 1 0 31280 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_332
timestamp 1586364061
transform 1 0 31648 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_13.mux_l1_in_2__A0
timestamp 1586364061
transform 1 0 33212 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_13.mux_l1_in_2__S
timestamp 1586364061
transform 1 0 33580 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_13.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 33948 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_3  FILLER_8_346
timestamp 1586364061
transform 1 0 32936 0 -1 7072
box -38 -48 314 592
use scs8hd_fill_2  FILLER_8_351
timestamp 1586364061
transform 1 0 33396 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_355
timestamp 1586364061
transform 1 0 33764 0 -1 7072
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_bottom_ipin_13.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 34500 0 -1 7072
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_13.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 34316 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_359
timestamp 1586364061
transform 1 0 34132 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_13.mux_l4_in_0__A0
timestamp 1586364061
transform 1 0 36432 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_382
timestamp 1586364061
transform 1 0 36248 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_8  FILLER_8_386
timestamp 1586364061
transform 1 0 36616 0 -1 7072
box -38 -48 774 592
use scs8hd_decap_3  FILLER_8_394
timestamp 1586364061
transform 1 0 37352 0 -1 7072
box -38 -48 314 592
use scs8hd_decap_3  PHY_17
timestamp 1586364061
transform -1 0 38824 0 -1 7072
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_106
timestamp 1586364061
transform 1 0 37628 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_8  FILLER_8_398
timestamp 1586364061
transform 1 0 37720 0 -1 7072
box -38 -48 774 592
use scs8hd_fill_1  FILLER_8_406
timestamp 1586364061
transform 1 0 38456 0 -1 7072
box -38 -48 130 592
use scs8hd_mux2_2  mux_bottom_ipin_2.mux_l2_in_2_
timestamp 1586364061
transform 1 0 1840 0 1 7072
box -38 -48 866 592
use scs8hd_decap_3  PHY_18
timestamp 1586364061
transform 1 0 1104 0 1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l2_in_2__A0
timestamp 1586364061
transform 1 0 1656 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l2_in_3__A1
timestamp 1586364061
transform 1 0 2852 0 1 7072
box -38 -48 222 592
use scs8hd_decap_3  FILLER_9_3
timestamp 1586364061
transform 1 0 1380 0 1 7072
box -38 -48 314 592
use scs8hd_fill_2  FILLER_9_17
timestamp 1586364061
transform 1 0 2668 0 1 7072
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_bottom_ipin_2.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 4048 0 1 7072
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_2.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 3864 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l2_in_3__A0
timestamp 1586364061
transform 1 0 3220 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_21
timestamp 1586364061
transform 1 0 3036 0 1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_9_25
timestamp 1586364061
transform 1 0 3404 0 1 7072
box -38 -48 406 592
use scs8hd_fill_1  FILLER_9_29
timestamp 1586364061
transform 1 0 3772 0 1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 6532 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_2.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 6164 0 1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_9_51
timestamp 1586364061
transform 1 0 5796 0 1 7072
box -38 -48 406 592
use scs8hd_fill_2  FILLER_9_57
timestamp 1586364061
transform 1 0 6348 0 1 7072
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_bottom_ipin_2.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 7360 0 1 7072
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_107
timestamp 1586364061
transform 1 0 6716 0 1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 7176 0 1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_9_62
timestamp 1586364061
transform 1 0 6808 0 1 7072
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 9660 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 10028 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 9292 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_87
timestamp 1586364061
transform 1 0 9108 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_91
timestamp 1586364061
transform 1 0 9476 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_95
timestamp 1586364061
transform 1 0 9844 0 1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_9_99
timestamp 1586364061
transform 1 0 10212 0 1 7072
box -38 -48 406 592
use scs8hd_mux2_2  mux_bottom_ipin_4.mux_l2_in_3_
timestamp 1586364061
transform 1 0 10764 0 1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_4.mux_l2_in_3__A1
timestamp 1586364061
transform 1 0 10580 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_5.scs8hd_dfxbp_1_3__CLK
timestamp 1586364061
transform 1 0 11776 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_114
timestamp 1586364061
transform 1 0 11592 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_118
timestamp 1586364061
transform 1 0 11960 0 1 7072
box -38 -48 222 592
use scs8hd_mux2_2  mux_bottom_ipin_6.mux_l2_in_0_
timestamp 1586364061
transform 1 0 12604 0 1 7072
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_108
timestamp 1586364061
transform 1 0 12328 0 1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_6.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 12144 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_4.mux_l2_in_2__S
timestamp 1586364061
transform 1 0 13616 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_123
timestamp 1586364061
transform 1 0 12420 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_134
timestamp 1586364061
transform 1 0 13432 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_138
timestamp 1586364061
transform 1 0 13800 0 1 7072
box -38 -48 222 592
use scs8hd_mux2_2  mux_bottom_ipin_4.mux_l2_in_2_
timestamp 1586364061
transform 1 0 14168 0 1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_4.mux_l2_in_2__A0
timestamp 1586364061
transform 1 0 13984 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_8.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 15456 0 1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_9_151
timestamp 1586364061
transform 1 0 14996 0 1 7072
box -38 -48 406 592
use scs8hd_fill_1  FILLER_9_155
timestamp 1586364061
transform 1 0 15364 0 1 7072
box -38 -48 130 592
use scs8hd_fill_2  FILLER_9_158
timestamp 1586364061
transform 1 0 15640 0 1 7072
box -38 -48 222 592
use scs8hd_mux2_2  mux_bottom_ipin_8.mux_l2_in_1_
timestamp 1586364061
transform 1 0 16376 0 1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_8.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 16192 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_8.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 15824 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_162
timestamp 1586364061
transform 1 0 16008 0 1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_9_175
timestamp 1586364061
transform 1 0 17204 0 1 7072
box -38 -48 406 592
use scs8hd_dfxbp_1  mem_bottom_ipin_5.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 18032 0 1 7072
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_109
timestamp 1586364061
transform 1 0 17940 0 1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_8.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 17664 0 1 7072
box -38 -48 222 592
use scs8hd_fill_1  FILLER_9_179
timestamp 1586364061
transform 1 0 17572 0 1 7072
box -38 -48 130 592
use scs8hd_fill_1  FILLER_9_182
timestamp 1586364061
transform 1 0 17848 0 1 7072
box -38 -48 130 592
use scs8hd_conb_1  _22_
timestamp 1586364061
transform 1 0 20884 0 1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_8.mux_l4_in_0__A0
timestamp 1586364061
transform 1 0 19964 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_203
timestamp 1586364061
transform 1 0 19780 0 1 7072
box -38 -48 222 592
use scs8hd_decap_8  FILLER_9_207
timestamp 1586364061
transform 1 0 20148 0 1 7072
box -38 -48 774 592
use scs8hd_decap_3  FILLER_9_218
timestamp 1586364061
transform 1 0 21160 0 1 7072
box -38 -48 314 592
use scs8hd_mux2_2  mux_bottom_ipin_11.mux_l2_in_0_
timestamp 1586364061
transform 1 0 21988 0 1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_11.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 21804 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_11.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 21436 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_11.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 23000 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_223
timestamp 1586364061
transform 1 0 21620 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_236
timestamp 1586364061
transform 1 0 22816 0 1 7072
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_bottom_ipin_11.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 24012 0 1 7072
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_110
timestamp 1586364061
transform 1 0 23552 0 1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_11.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 23828 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_11.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 23368 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_240
timestamp 1586364061
transform 1 0 23184 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_245
timestamp 1586364061
transform 1 0 23644 0 1 7072
box -38 -48 222 592
use scs8hd_mux2_2  mux_bottom_ipin_10.mux_l2_in_1_
timestamp 1586364061
transform 1 0 26496 0 1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_10.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 26312 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_10.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 25944 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_268
timestamp 1586364061
transform 1 0 25760 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_272
timestamp 1586364061
transform 1 0 26128 0 1 7072
box -38 -48 222 592
use scs8hd_conb_1  _23_
timestamp 1586364061
transform 1 0 28060 0 1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_10.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 27508 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_10.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 27876 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_285
timestamp 1586364061
transform 1 0 27324 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_289
timestamp 1586364061
transform 1 0 27692 0 1 7072
box -38 -48 222 592
use scs8hd_decap_3  FILLER_9_296
timestamp 1586364061
transform 1 0 28336 0 1 7072
box -38 -48 314 592
use scs8hd_mux2_2  mux_bottom_ipin_10.mux_l2_in_3_
timestamp 1586364061
transform 1 0 29256 0 1 7072
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_111
timestamp 1586364061
transform 1 0 29164 0 1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_10.mux_l2_in_3__A1
timestamp 1586364061
transform 1 0 28980 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_10.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 28612 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_10.mux_l2_in_3__A0
timestamp 1586364061
transform 1 0 30268 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_301
timestamp 1586364061
transform 1 0 28796 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_315
timestamp 1586364061
transform 1 0 30084 0 1 7072
box -38 -48 222 592
use scs8hd_mux2_2  mux_bottom_ipin_12.mux_l3_in_1_
timestamp 1586364061
transform 1 0 30820 0 1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_10.mux_l2_in_3__S
timestamp 1586364061
transform 1 0 30636 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_12.mux_l3_in_1__A1
timestamp 1586364061
transform 1 0 31832 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_319
timestamp 1586364061
transform 1 0 30452 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_332
timestamp 1586364061
transform 1 0 31648 0 1 7072
box -38 -48 222 592
use scs8hd_decap_3  FILLER_9_336
timestamp 1586364061
transform 1 0 32016 0 1 7072
box -38 -48 314 592
use scs8hd_mux2_2  mux_bottom_ipin_13.mux_l2_in_1_
timestamp 1586364061
transform 1 0 33212 0 1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_13.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 33028 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_14.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 32660 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_14.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 32292 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_341
timestamp 1586364061
transform 1 0 32476 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_345
timestamp 1586364061
transform 1 0 32844 0 1 7072
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_bottom_ipin_13.scs8hd_dfxbp_1_3_
timestamp 1586364061
transform 1 0 35236 0 1 7072
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_112
timestamp 1586364061
transform 1 0 34776 0 1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_13.scs8hd_dfxbp_1_3__CLK
timestamp 1586364061
transform 1 0 35052 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_13.mux_l4_in_0__S
timestamp 1586364061
transform 1 0 34592 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_13.mux_l2_in_3__S
timestamp 1586364061
transform 1 0 34224 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_358
timestamp 1586364061
transform 1 0 34040 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_362
timestamp 1586364061
transform 1 0 34408 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_367
timestamp 1586364061
transform 1 0 34868 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_13.mux_l4_in_0__A1
timestamp 1586364061
transform 1 0 37168 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_390
timestamp 1586364061
transform 1 0 36984 0 1 7072
box -38 -48 222 592
use scs8hd_decap_12  FILLER_9_394
timestamp 1586364061
transform 1 0 37352 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_3  PHY_19
timestamp 1586364061
transform -1 0 38824 0 1 7072
box -38 -48 314 592
use scs8hd_fill_1  FILLER_9_406
timestamp 1586364061
transform 1 0 38456 0 1 7072
box -38 -48 130 592
use scs8hd_mux2_2  mux_bottom_ipin_2.mux_l2_in_3_
timestamp 1586364061
transform 1 0 1748 0 -1 8160
box -38 -48 866 592
use scs8hd_decap_3  PHY_20
timestamp 1586364061
transform 1 0 1104 0 -1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l4_in_0__S
timestamp 1586364061
transform 1 0 2760 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l2_in_3__S
timestamp 1586364061
transform 1 0 1564 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_3
timestamp 1586364061
transform 1 0 1380 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_16
timestamp 1586364061
transform 1 0 2576 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_1  FILLER_10_28
timestamp 1586364061
transform 1 0 3680 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_4  FILLER_10_24
timestamp 1586364061
transform 1 0 3312 0 -1 8160
box -38 -48 406 592
use scs8hd_fill_2  FILLER_10_20
timestamp 1586364061
transform 1 0 2944 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 3772 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.mux_l4_in_0__A0
timestamp 1586364061
transform 1 0 3128 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_3  FILLER_10_36
timestamp 1586364061
transform 1 0 4416 0 -1 8160
box -38 -48 314 592
use scs8hd_fill_2  FILLER_10_32
timestamp 1586364061
transform 1 0 4048 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_2.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 4232 0 -1 8160
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_113
timestamp 1586364061
transform 1 0 3956 0 -1 8160
box -38 -48 130 592
use scs8hd_dfxbp_1  mem_bottom_ipin_2.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 4692 0 -1 8160
box -38 -48 1786 592
use scs8hd_fill_2  FILLER_10_58
timestamp 1586364061
transform 1 0 6440 0 -1 8160
box -38 -48 222 592
use scs8hd_mux2_2  mux_bottom_ipin_2.mux_l1_in_0_
timestamp 1586364061
transform 1 0 7176 0 -1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 6624 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__45__A
timestamp 1586364061
transform 1 0 6992 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_1.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 8280 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_62
timestamp 1586364061
transform 1 0 6808 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_3  FILLER_10_75
timestamp 1586364061
transform 1 0 8004 0 -1 8160
box -38 -48 314 592
use scs8hd_mux2_2  mux_bottom_ipin_1.mux_l1_in_0_
timestamp 1586364061
transform 1 0 9660 0 -1 8160
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_114
timestamp 1586364061
transform 1 0 9568 0 -1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 8648 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_1.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 9016 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_80
timestamp 1586364061
transform 1 0 8464 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_84
timestamp 1586364061
transform 1 0 8832 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_10_88
timestamp 1586364061
transform 1 0 9200 0 -1 8160
box -38 -48 406 592
use scs8hd_dfxbp_1  mem_bottom_ipin_5.scs8hd_dfxbp_1_3_
timestamp 1586364061
transform 1 0 11224 0 -1 8160
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.mux_l1_in_1__A0
timestamp 1586364061
transform 1 0 10764 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_3  FILLER_10_102
timestamp 1586364061
transform 1 0 10488 0 -1 8160
box -38 -48 314 592
use scs8hd_decap_3  FILLER_10_107
timestamp 1586364061
transform 1 0 10948 0 -1 8160
box -38 -48 314 592
use scs8hd_conb_1  _31_
timestamp 1586364061
transform 1 0 13708 0 -1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_6.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 13156 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_6.mux_l3_in_1__S
timestamp 1586364061
transform 1 0 13524 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_129
timestamp 1586364061
transform 1 0 12972 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_133
timestamp 1586364061
transform 1 0 13340 0 -1 8160
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_115
timestamp 1586364061
transform 1 0 15180 0 -1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_4.mux_l2_in_2__A1
timestamp 1586364061
transform 1 0 14168 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_140
timestamp 1586364061
transform 1 0 13984 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_8  FILLER_10_144
timestamp 1586364061
transform 1 0 14352 0 -1 8160
box -38 -48 774 592
use scs8hd_fill_1  FILLER_10_152
timestamp 1586364061
transform 1 0 15088 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_6  FILLER_10_154
timestamp 1586364061
transform 1 0 15272 0 -1 8160
box -38 -48 590 592
use scs8hd_mux2_2  mux_bottom_ipin_8.mux_l3_in_0_
timestamp 1586364061
transform 1 0 16100 0 -1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_8.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 17480 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_8.mux_l1_in_2__S
timestamp 1586364061
transform 1 0 17112 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_8.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 15916 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_1  FILLER_10_160
timestamp 1586364061
transform 1 0 15824 0 -1 8160
box -38 -48 130 592
use scs8hd_fill_2  FILLER_10_172
timestamp 1586364061
transform 1 0 16928 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_176
timestamp 1586364061
transform 1 0 17296 0 -1 8160
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_bottom_ipin_8.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 17664 0 -1 8160
box -38 -48 1786 592
use scs8hd_decap_4  FILLER_10_203
timestamp 1586364061
transform 1 0 19780 0 -1 8160
box -38 -48 406 592
use scs8hd_fill_2  FILLER_10_199
timestamp 1586364061
transform 1 0 19412 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_8.mux_l4_in_0__A1
timestamp 1586364061
transform 1 0 19596 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_8.mux_l3_in_1__S
timestamp 1586364061
transform 1 0 20148 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_209
timestamp 1586364061
transform 1 0 20332 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_8.mux_l3_in_1__A0
timestamp 1586364061
transform 1 0 20516 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_1  FILLER_10_215
timestamp 1586364061
transform 1 0 20884 0 -1 8160
box -38 -48 130 592
use scs8hd_fill_1  FILLER_10_213
timestamp 1586364061
transform 1 0 20700 0 -1 8160
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_116
timestamp 1586364061
transform 1 0 20792 0 -1 8160
box -38 -48 130 592
use scs8hd_conb_1  _17_
timestamp 1586364061
transform 1 0 20976 0 -1 8160
box -38 -48 314 592
use scs8hd_dfxbp_1  mem_bottom_ipin_11.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 21988 0 -1 8160
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_11.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 21804 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_11.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 21436 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_219
timestamp 1586364061
transform 1 0 21252 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_223
timestamp 1586364061
transform 1 0 21620 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_10.mux_l4_in_0__S
timestamp 1586364061
transform 1 0 24288 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_10.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 24656 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_10.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 23920 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_246
timestamp 1586364061
transform 1 0 23736 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_250
timestamp 1586364061
transform 1 0 24104 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_254
timestamp 1586364061
transform 1 0 24472 0 -1 8160
box -38 -48 222 592
use scs8hd_mux2_2  mux_bottom_ipin_10.mux_l2_in_0_
timestamp 1586364061
transform 1 0 26496 0 -1 8160
box -38 -48 866 592
use scs8hd_mux2_2  mux_bottom_ipin_10.mux_l3_in_0_
timestamp 1586364061
transform 1 0 24840 0 -1 8160
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_117
timestamp 1586364061
transform 1 0 26404 0 -1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_10.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 26220 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_6  FILLER_10_267
timestamp 1586364061
transform 1 0 25668 0 -1 8160
box -38 -48 590 592
use scs8hd_conb_1  _21_
timestamp 1586364061
transform 1 0 28060 0 -1 8160
box -38 -48 314 592
use scs8hd_decap_8  FILLER_10_285
timestamp 1586364061
transform 1 0 27324 0 -1 8160
box -38 -48 774 592
use scs8hd_fill_2  FILLER_10_296
timestamp 1586364061
transform 1 0 28336 0 -1 8160
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_bottom_ipin_10.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 29072 0 -1 8160
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_10.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 28520 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_10_300
timestamp 1586364061
transform 1 0 28704 0 -1 8160
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_118
timestamp 1586364061
transform 1 0 32016 0 -1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_14.mux_l2_in_3__A1
timestamp 1586364061
transform 1 0 31004 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_14.mux_l2_in_2__S
timestamp 1586364061
transform 1 0 31372 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_14.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 31832 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_323
timestamp 1586364061
transform 1 0 30820 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_327
timestamp 1586364061
transform 1 0 31188 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_3  FILLER_10_331
timestamp 1586364061
transform 1 0 31556 0 -1 8160
box -38 -48 314 592
use scs8hd_decap_3  FILLER_10_337
timestamp 1586364061
transform 1 0 32108 0 -1 8160
box -38 -48 314 592
use scs8hd_dfxbp_1  mem_bottom_ipin_14.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 32936 0 -1 8160
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_13.mux_l2_in_3__A0
timestamp 1586364061
transform 1 0 32752 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_13.mux_l2_in_2__S
timestamp 1586364061
transform 1 0 32384 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_342
timestamp 1586364061
transform 1 0 32568 0 -1 8160
box -38 -48 222 592
use scs8hd_mux2_2  mux_bottom_ipin_13.mux_l4_in_0_
timestamp 1586364061
transform 1 0 35420 0 -1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_14.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 35236 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_13.scs8hd_dfxbp_1_3__D
timestamp 1586364061
transform 1 0 34868 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_365
timestamp 1586364061
transform 1 0 34684 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_369
timestamp 1586364061
transform 1 0 35052 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_14.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 36432 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_382
timestamp 1586364061
transform 1 0 36248 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_8  FILLER_10_386
timestamp 1586364061
transform 1 0 36616 0 -1 8160
box -38 -48 774 592
use scs8hd_decap_3  FILLER_10_394
timestamp 1586364061
transform 1 0 37352 0 -1 8160
box -38 -48 314 592
use scs8hd_decap_3  PHY_21
timestamp 1586364061
transform -1 0 38824 0 -1 8160
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_119
timestamp 1586364061
transform 1 0 37628 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_8  FILLER_10_398
timestamp 1586364061
transform 1 0 37720 0 -1 8160
box -38 -48 774 592
use scs8hd_fill_1  FILLER_10_406
timestamp 1586364061
transform 1 0 38456 0 -1 8160
box -38 -48 130 592
use scs8hd_dfxbp_1  mem_bottom_ipin_1.scs8hd_dfxbp_1_3_
timestamp 1586364061
transform 1 0 2116 0 1 8160
box -38 -48 1786 592
use scs8hd_decap_3  PHY_22
timestamp 1586364061
transform 1 0 1104 0 1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_1.scs8hd_dfxbp_1_3__CLK
timestamp 1586364061
transform 1 0 1932 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_1.scs8hd_dfxbp_1_3__D
timestamp 1586364061
transform 1 0 1564 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_3
timestamp 1586364061
transform 1 0 1380 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_7
timestamp 1586364061
transform 1 0 1748 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 4416 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 4048 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_30
timestamp 1586364061
transform 1 0 3864 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_34
timestamp 1586364061
transform 1 0 4232 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_38
timestamp 1586364061
transform 1 0 4600 0 1 8160
box -38 -48 222 592
use scs8hd_mux2_2  mux_bottom_ipin_2.mux_l3_in_0_
timestamp 1586364061
transform 1 0 5152 0 1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 6348 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 4784 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_42
timestamp 1586364061
transform 1 0 4968 0 1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_11_53
timestamp 1586364061
transform 1 0 5980 0 1 8160
box -38 -48 406 592
use scs8hd_fill_2  FILLER_11_59
timestamp 1586364061
transform 1 0 6532 0 1 8160
box -38 -48 222 592
use scs8hd_buf_2  _45_
timestamp 1586364061
transform 1 0 6808 0 1 8160
box -38 -48 406 592
use scs8hd_dfxbp_1  mem_bottom_ipin_1.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 8280 0 1 8160
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_120
timestamp 1586364061
transform 1 0 6716 0 1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 8004 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 7636 0 1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_11_66
timestamp 1586364061
transform 1 0 7176 0 1 8160
box -38 -48 406 592
use scs8hd_fill_1  FILLER_11_70
timestamp 1586364061
transform 1 0 7544 0 1 8160
box -38 -48 130 592
use scs8hd_fill_2  FILLER_11_73
timestamp 1586364061
transform 1 0 7820 0 1 8160
box -38 -48 222 592
use scs8hd_fill_1  FILLER_11_77
timestamp 1586364061
transform 1 0 8188 0 1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_6.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 10212 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_97
timestamp 1586364061
transform 1 0 10028 0 1 8160
box -38 -48 222 592
use scs8hd_mux2_2  mux_bottom_ipin_1.mux_l1_in_1_
timestamp 1586364061
transform 1 0 10764 0 1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_6.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 11776 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.mux_l1_in_1__A1
timestamp 1586364061
transform 1 0 10580 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_101
timestamp 1586364061
transform 1 0 10396 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_114
timestamp 1586364061
transform 1 0 11592 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_118
timestamp 1586364061
transform 1 0 11960 0 1 8160
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_bottom_ipin_6.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 12604 0 1 8160
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_121
timestamp 1586364061
transform 1 0 12328 0 1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_6.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 12144 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_123
timestamp 1586364061
transform 1 0 12420 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_6.mux_l2_in_2__A0
timestamp 1586364061
transform 1 0 15272 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_6.mux_l2_in_2__A1
timestamp 1586364061
transform 1 0 15640 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_6.mux_l2_in_2__S
timestamp 1586364061
transform 1 0 14904 0 1 8160
box -38 -48 222 592
use scs8hd_decap_6  FILLER_11_144
timestamp 1586364061
transform 1 0 14352 0 1 8160
box -38 -48 590 592
use scs8hd_fill_2  FILLER_11_152
timestamp 1586364061
transform 1 0 15088 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_156
timestamp 1586364061
transform 1 0 15456 0 1 8160
box -38 -48 222 592
use scs8hd_mux2_2  mux_bottom_ipin_8.mux_l1_in_2_
timestamp 1586364061
transform 1 0 16376 0 1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_8.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 17480 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_8.mux_l1_in_2__A1
timestamp 1586364061
transform 1 0 16192 0 1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_11_160
timestamp 1586364061
transform 1 0 15824 0 1 8160
box -38 -48 406 592
use scs8hd_decap_3  FILLER_11_175
timestamp 1586364061
transform 1 0 17204 0 1 8160
box -38 -48 314 592
use scs8hd_mux2_2  mux_bottom_ipin_8.mux_l1_in_1_
timestamp 1586364061
transform 1 0 18032 0 1 8160
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_122
timestamp 1586364061
transform 1 0 17940 0 1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_8.mux_l1_in_1__A0
timestamp 1586364061
transform 1 0 19044 0 1 8160
box -38 -48 222 592
use scs8hd_decap_3  FILLER_11_180
timestamp 1586364061
transform 1 0 17664 0 1 8160
box -38 -48 314 592
use scs8hd_fill_2  FILLER_11_193
timestamp 1586364061
transform 1 0 18860 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_197
timestamp 1586364061
transform 1 0 19228 0 1 8160
box -38 -48 222 592
use scs8hd_mux2_2  mux_bottom_ipin_8.mux_l3_in_1_
timestamp 1586364061
transform 1 0 20148 0 1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_8.mux_l4_in_0__S
timestamp 1586364061
transform 1 0 19412 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_8.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 19780 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_201
timestamp 1586364061
transform 1 0 19596 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_205
timestamp 1586364061
transform 1 0 19964 0 1 8160
box -38 -48 222 592
use scs8hd_decap_3  FILLER_11_216
timestamp 1586364061
transform 1 0 20976 0 1 8160
box -38 -48 314 592
use scs8hd_mux2_2  mux_bottom_ipin_11.mux_l3_in_0_
timestamp 1586364061
transform 1 0 21804 0 1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_8.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 21620 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_8.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 21252 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_11.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 22816 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_221
timestamp 1586364061
transform 1 0 21436 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_234
timestamp 1586364061
transform 1 0 22632 0 1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_11_238
timestamp 1586364061
transform 1 0 23000 0 1 8160
box -38 -48 406 592
use scs8hd_dfxbp_1  mem_bottom_ipin_10.scs8hd_dfxbp_1_3_
timestamp 1586364061
transform 1 0 23644 0 1 8160
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_123
timestamp 1586364061
transform 1 0 23552 0 1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_10.scs8hd_dfxbp_1_3__CLK
timestamp 1586364061
transform 1 0 23368 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_10.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 26496 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_10.mux_l4_in_0__A1
timestamp 1586364061
transform 1 0 25576 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_10.mux_l4_in_0__A0
timestamp 1586364061
transform 1 0 25944 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_264
timestamp 1586364061
transform 1 0 25392 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_268
timestamp 1586364061
transform 1 0 25760 0 1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_11_272
timestamp 1586364061
transform 1 0 26128 0 1 8160
box -38 -48 406 592
use scs8hd_mux2_2  mux_bottom_ipin_10.mux_l1_in_0_
timestamp 1586364061
transform 1 0 27048 0 1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_10.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 26864 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_10.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 28060 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_278
timestamp 1586364061
transform 1 0 26680 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_291
timestamp 1586364061
transform 1 0 27876 0 1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_11_295
timestamp 1586364061
transform 1 0 28244 0 1 8160
box -38 -48 406 592
use scs8hd_mux2_2  mux_bottom_ipin_10.mux_l2_in_2_
timestamp 1586364061
transform 1 0 29256 0 1 8160
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_124
timestamp 1586364061
transform 1 0 29164 0 1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_10.mux_l2_in_2__A0
timestamp 1586364061
transform 1 0 28980 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_14.mux_l2_in_2__A1
timestamp 1586364061
transform 1 0 30268 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_10.mux_l2_in_2__A1
timestamp 1586364061
transform 1 0 28612 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_301
timestamp 1586364061
transform 1 0 28796 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_315
timestamp 1586364061
transform 1 0 30084 0 1 8160
box -38 -48 222 592
use scs8hd_mux2_2  mux_bottom_ipin_14.mux_l2_in_2_
timestamp 1586364061
transform 1 0 30820 0 1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_14.mux_l2_in_2__A0
timestamp 1586364061
transform 1 0 30636 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_14.mux_l2_in_3__A0
timestamp 1586364061
transform 1 0 31832 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_319
timestamp 1586364061
transform 1 0 30452 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_332
timestamp 1586364061
transform 1 0 31648 0 1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_11_336
timestamp 1586364061
transform 1 0 32016 0 1 8160
box -38 -48 406 592
use scs8hd_mux2_2  mux_bottom_ipin_13.mux_l2_in_2_
timestamp 1586364061
transform 1 0 32936 0 1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_13.mux_l2_in_2__A0
timestamp 1586364061
transform 1 0 32752 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_13.mux_l2_in_2__A1
timestamp 1586364061
transform 1 0 32384 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_13.mux_l2_in_3__A1
timestamp 1586364061
transform 1 0 33948 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_342
timestamp 1586364061
transform 1 0 32568 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_355
timestamp 1586364061
transform 1 0 33764 0 1 8160
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_bottom_ipin_14.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 34868 0 1 8160
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_125
timestamp 1586364061
transform 1 0 34776 0 1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_14.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 34592 0 1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_11_359
timestamp 1586364061
transform 1 0 34132 0 1 8160
box -38 -48 406 592
use scs8hd_fill_1  FILLER_11_363
timestamp 1586364061
transform 1 0 34500 0 1 8160
box -38 -48 130 592
use scs8hd_buf_2  _71_
timestamp 1586364061
transform 1 0 37352 0 1 8160
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_14.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 36800 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_14.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 37168 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_386
timestamp 1586364061
transform 1 0 36616 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_390
timestamp 1586364061
transform 1 0 36984 0 1 8160
box -38 -48 222 592
use scs8hd_decap_3  PHY_23
timestamp 1586364061
transform -1 0 38824 0 1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__71__A
timestamp 1586364061
transform 1 0 37904 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_398
timestamp 1586364061
transform 1 0 37720 0 1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_11_402
timestamp 1586364061
transform 1 0 38088 0 1 8160
box -38 -48 406 592
use scs8hd_fill_1  FILLER_11_406
timestamp 1586364061
transform 1 0 38456 0 1 8160
box -38 -48 130 592
use scs8hd_mux2_2  mux_bottom_ipin_2.mux_l4_in_0_
timestamp 1586364061
transform 1 0 2208 0 -1 9248
box -38 -48 866 592
use scs8hd_decap_3  PHY_24
timestamp 1586364061
transform 1 0 1104 0 -1 9248
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.mux_l3_in_1__S
timestamp 1586364061
transform 1 0 1932 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.mux_l3_in_1__A1
timestamp 1586364061
transform 1 0 1564 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_3
timestamp 1586364061
transform 1 0 1380 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_7
timestamp 1586364061
transform 1 0 1748 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_1  FILLER_12_11
timestamp 1586364061
transform 1 0 2116 0 -1 9248
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_126
timestamp 1586364061
transform 1 0 3956 0 -1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__43__A
timestamp 1586364061
transform 1 0 4232 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_1.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 3496 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 4600 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_12_21
timestamp 1586364061
transform 1 0 3036 0 -1 9248
box -38 -48 406 592
use scs8hd_fill_1  FILLER_12_25
timestamp 1586364061
transform 1 0 3404 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_3  FILLER_12_28
timestamp 1586364061
transform 1 0 3680 0 -1 9248
box -38 -48 314 592
use scs8hd_fill_2  FILLER_12_32
timestamp 1586364061
transform 1 0 4048 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_36
timestamp 1586364061
transform 1 0 4416 0 -1 9248
box -38 -48 222 592
use scs8hd_mux2_2  mux_bottom_ipin_1.mux_l2_in_0_
timestamp 1586364061
transform 1 0 4784 0 -1 9248
box -38 -48 866 592
use scs8hd_mux2_2  mux_bottom_ipin_2.mux_l2_in_1_
timestamp 1586364061
transform 1 0 6348 0 -1 9248
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 6164 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 5796 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_49
timestamp 1586364061
transform 1 0 5612 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_53
timestamp 1586364061
transform 1 0 5980 0 -1 9248
box -38 -48 222 592
use scs8hd_mux2_2  mux_bottom_ipin_0.mux_l1_in_0_
timestamp 1586364061
transform 1 0 8004 0 -1 9248
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l1_in_1__A0
timestamp 1586364061
transform 1 0 7820 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l4_in_0__A0
timestamp 1586364061
transform 1 0 7360 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_66
timestamp 1586364061
transform 1 0 7176 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_3  FILLER_12_70
timestamp 1586364061
transform 1 0 7544 0 -1 9248
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_127
timestamp 1586364061
transform 1 0 9568 0 -1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_0.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 9016 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_84
timestamp 1586364061
transform 1 0 8832 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_12_88
timestamp 1586364061
transform 1 0 9200 0 -1 9248
box -38 -48 406 592
use scs8hd_decap_8  FILLER_12_93
timestamp 1586364061
transform 1 0 9660 0 -1 9248
box -38 -48 774 592
use scs8hd_mux2_2  mux_bottom_ipin_6.mux_l2_in_1_
timestamp 1586364061
transform 1 0 11132 0 -1 9248
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.mux_l1_in_1__S
timestamp 1586364061
transform 1 0 10764 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_6.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 10396 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_103
timestamp 1586364061
transform 1 0 10580 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_107
timestamp 1586364061
transform 1 0 10948 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_118
timestamp 1586364061
transform 1 0 11960 0 -1 9248
box -38 -48 222 592
use scs8hd_mux2_2  mux_bottom_ipin_6.mux_l3_in_1_
timestamp 1586364061
transform 1 0 12696 0 -1 9248
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_6.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 13708 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_6.mux_l3_in_1__A1
timestamp 1586364061
transform 1 0 12512 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_6.mux_l3_in_1__A0
timestamp 1586364061
transform 1 0 12144 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_122
timestamp 1586364061
transform 1 0 12328 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_135
timestamp 1586364061
transform 1 0 13524 0 -1 9248
box -38 -48 222 592
use scs8hd_mux2_2  mux_bottom_ipin_6.mux_l2_in_2_
timestamp 1586364061
transform 1 0 15272 0 -1 9248
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_128
timestamp 1586364061
transform 1 0 15180 0 -1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_6.mux_l2_in_3__S
timestamp 1586364061
transform 1 0 14996 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_12  FILLER_12_139
timestamp 1586364061
transform 1 0 13892 0 -1 9248
box -38 -48 1142 592
use scs8hd_mux2_2  mux_bottom_ipin_8.mux_l1_in_0_
timestamp 1586364061
transform 1 0 17480 0 -1 9248
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_7.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 16376 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_8.mux_l1_in_2__A0
timestamp 1586364061
transform 1 0 16744 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_7.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 17112 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_3  FILLER_12_163
timestamp 1586364061
transform 1 0 16100 0 -1 9248
box -38 -48 314 592
use scs8hd_fill_2  FILLER_12_168
timestamp 1586364061
transform 1 0 16560 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_172
timestamp 1586364061
transform 1 0 16928 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_176
timestamp 1586364061
transform 1 0 17296 0 -1 9248
box -38 -48 222 592
use scs8hd_mux2_2  mux_bottom_ipin_8.mux_l4_in_0_
timestamp 1586364061
transform 1 0 19228 0 -1 9248
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_8.mux_l1_in_1__A1
timestamp 1586364061
transform 1 0 18492 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_8.mux_l1_in_1__S
timestamp 1586364061
transform 1 0 18860 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_187
timestamp 1586364061
transform 1 0 18308 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_191
timestamp 1586364061
transform 1 0 18676 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_195
timestamp 1586364061
transform 1 0 19044 0 -1 9248
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_129
timestamp 1586364061
transform 1 0 20792 0 -1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_8.mux_l3_in_1__A1
timestamp 1586364061
transform 1 0 20240 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_206
timestamp 1586364061
transform 1 0 20056 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_12_210
timestamp 1586364061
transform 1 0 20424 0 -1 9248
box -38 -48 406 592
use scs8hd_decap_8  FILLER_12_215
timestamp 1586364061
transform 1 0 20884 0 -1 9248
box -38 -48 774 592
use scs8hd_dfxbp_1  mem_bottom_ipin_8.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 21620 0 -1 9248
box -38 -48 1786 592
use scs8hd_mux2_2  mux_bottom_ipin_10.mux_l4_in_0_
timestamp 1586364061
transform 1 0 24288 0 -1 9248
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_10.scs8hd_dfxbp_1_3__D
timestamp 1586364061
transform 1 0 23644 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_9.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 24104 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_3  FILLER_12_242
timestamp 1586364061
transform 1 0 23368 0 -1 9248
box -38 -48 314 592
use scs8hd_decap_3  FILLER_12_247
timestamp 1586364061
transform 1 0 23828 0 -1 9248
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_130
timestamp 1586364061
transform 1 0 26404 0 -1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_9.mux_l1_in_1__S
timestamp 1586364061
transform 1 0 25300 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_261
timestamp 1586364061
transform 1 0 25116 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_8  FILLER_12_265
timestamp 1586364061
transform 1 0 25484 0 -1 9248
box -38 -48 774 592
use scs8hd_fill_2  FILLER_12_273
timestamp 1586364061
transform 1 0 26220 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_12_276
timestamp 1586364061
transform 1 0 26496 0 -1 9248
box -38 -48 406 592
use scs8hd_conb_1  _25_
timestamp 1586364061
transform 1 0 26956 0 -1 9248
box -38 -48 314 592
use scs8hd_dfxbp_1  mem_bottom_ipin_10.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 27968 0 -1 9248
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_10.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 27416 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_10.mux_l3_in_1__S
timestamp 1586364061
transform 1 0 27784 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_1  FILLER_12_280
timestamp 1586364061
transform 1 0 26864 0 -1 9248
box -38 -48 130 592
use scs8hd_fill_2  FILLER_12_284
timestamp 1586364061
transform 1 0 27232 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_288
timestamp 1586364061
transform 1 0 27600 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_10.mux_l2_in_2__S
timestamp 1586364061
transform 1 0 29900 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_14.mux_l2_in_3__S
timestamp 1586364061
transform 1 0 30268 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_311
timestamp 1586364061
transform 1 0 29716 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_315
timestamp 1586364061
transform 1 0 30084 0 -1 9248
box -38 -48 222 592
use scs8hd_mux2_2  mux_bottom_ipin_14.mux_l2_in_3_
timestamp 1586364061
transform 1 0 30452 0 -1 9248
box -38 -48 866 592
use scs8hd_mux2_2  mux_bottom_ipin_14.mux_l3_in_0_
timestamp 1586364061
transform 1 0 32108 0 -1 9248
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_131
timestamp 1586364061
transform 1 0 32016 0 -1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_15.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 31832 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_14.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 31464 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_328
timestamp 1586364061
transform 1 0 31280 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_332
timestamp 1586364061
transform 1 0 31648 0 -1 9248
box -38 -48 222 592
use scs8hd_mux2_2  mux_bottom_ipin_13.mux_l2_in_3_
timestamp 1586364061
transform 1 0 33672 0 -1 9248
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_14.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 33212 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_3  FILLER_12_346
timestamp 1586364061
transform 1 0 32936 0 -1 9248
box -38 -48 314 592
use scs8hd_decap_3  FILLER_12_351
timestamp 1586364061
transform 1 0 33396 0 -1 9248
box -38 -48 314 592
use scs8hd_mux2_2  mux_bottom_ipin_14.mux_l2_in_0_
timestamp 1586364061
transform 1 0 35236 0 -1 9248
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_15.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 34868 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_12_363
timestamp 1586364061
transform 1 0 34500 0 -1 9248
box -38 -48 406 592
use scs8hd_fill_2  FILLER_12_369
timestamp 1586364061
transform 1 0 35052 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_14.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 36432 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_12_380
timestamp 1586364061
transform 1 0 36064 0 -1 9248
box -38 -48 406 592
use scs8hd_decap_8  FILLER_12_386
timestamp 1586364061
transform 1 0 36616 0 -1 9248
box -38 -48 774 592
use scs8hd_decap_3  FILLER_12_394
timestamp 1586364061
transform 1 0 37352 0 -1 9248
box -38 -48 314 592
use scs8hd_decap_3  PHY_25
timestamp 1586364061
transform -1 0 38824 0 -1 9248
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_132
timestamp 1586364061
transform 1 0 37628 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_8  FILLER_12_398
timestamp 1586364061
transform 1 0 37720 0 -1 9248
box -38 -48 774 592
use scs8hd_fill_1  FILLER_12_406
timestamp 1586364061
transform 1 0 38456 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_4  FILLER_14_3
timestamp 1586364061
transform 1 0 1380 0 -1 10336
box -38 -48 406 592
use scs8hd_decap_4  FILLER_13_3
timestamp 1586364061
transform 1 0 1380 0 1 9248
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 1748 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.mux_l4_in_0__S
timestamp 1586364061
transform 1 0 1748 0 1 9248
box -38 -48 222 592
use scs8hd_decap_3  PHY_28
timestamp 1586364061
transform 1 0 1104 0 -1 10336
box -38 -48 314 592
use scs8hd_decap_3  PHY_26
timestamp 1586364061
transform 1 0 1104 0 1 9248
box -38 -48 314 592
use scs8hd_mux2_2  mux_bottom_ipin_1.mux_l4_in_0_
timestamp 1586364061
transform 1 0 1932 0 1 9248
box -38 -48 866 592
use scs8hd_mux2_2  mux_bottom_ipin_1.mux_l3_in_1_
timestamp 1586364061
transform 1 0 1932 0 -1 10336
box -38 -48 866 592
use scs8hd_fill_2  FILLER_14_18
timestamp 1586364061
transform 1 0 2760 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_18
timestamp 1586364061
transform 1 0 2760 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_26
timestamp 1586364061
transform 1 0 3496 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_22
timestamp 1586364061
transform 1 0 3128 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_22
timestamp 1586364061
transform 1 0 3128 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.mux_l3_in_1__A0
timestamp 1586364061
transform 1 0 3680 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 2944 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 3312 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.mux_l2_in_3__S
timestamp 1586364061
transform 1 0 2944 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_1.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 3312 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_36
timestamp 1586364061
transform 1 0 4416 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_1  FILLER_14_30
timestamp 1586364061
transform 1 0 3864 0 -1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.mux_l4_in_0__A1
timestamp 1586364061
transform 1 0 4600 0 -1 10336
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_139
timestamp 1586364061
transform 1 0 3956 0 -1 10336
box -38 -48 130 592
use scs8hd_buf_2  _43_
timestamp 1586364061
transform 1 0 4048 0 -1 10336
box -38 -48 406 592
use scs8hd_dfxbp_1  mem_bottom_ipin_1.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 3496 0 1 9248
box -38 -48 1786 592
use scs8hd_fill_1  FILLER_14_44
timestamp 1586364061
transform 1 0 5152 0 -1 10336
box -38 -48 130 592
use scs8hd_fill_2  FILLER_14_40
timestamp 1586364061
transform 1 0 4784 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_49
timestamp 1586364061
transform 1 0 5612 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_45
timestamp 1586364061
transform 1 0 5244 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l4_in_0__A1
timestamp 1586364061
transform 1 0 4968 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_1.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 5428 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_57
timestamp 1586364061
transform 1 0 6348 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_53
timestamp 1586364061
transform 1 0 5980 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_1.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 5796 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l1_in_2__A0
timestamp 1586364061
transform 1 0 6164 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l1_in_2__A1
timestamp 1586364061
transform 1 0 6532 0 1 9248
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_bottom_ipin_1.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 5244 0 -1 10336
box -38 -48 1786 592
use scs8hd_decap_4  FILLER_14_68
timestamp 1586364061
transform 1 0 7360 0 -1 10336
box -38 -48 406 592
use scs8hd_fill_2  FILLER_14_64
timestamp 1586364061
transform 1 0 6992 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_1  FILLER_13_62
timestamp 1586364061
transform 1 0 6808 0 1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l1_in_2__S
timestamp 1586364061
transform 1 0 7176 0 -1 10336
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_133
timestamp 1586364061
transform 1 0 6716 0 1 9248
box -38 -48 130 592
use scs8hd_mux2_2  mux_bottom_ipin_0.mux_l1_in_2_
timestamp 1586364061
transform 1 0 6900 0 1 9248
box -38 -48 866 592
use scs8hd_fill_1  FILLER_14_72
timestamp 1586364061
transform 1 0 7728 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_3  FILLER_13_77
timestamp 1586364061
transform 1 0 8188 0 1 9248
box -38 -48 314 592
use scs8hd_decap_3  FILLER_13_72
timestamp 1586364061
transform 1 0 7728 0 1 9248
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l1_in_1__S
timestamp 1586364061
transform 1 0 7820 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l1_in_1__A1
timestamp 1586364061
transform 1 0 8004 0 1 9248
box -38 -48 222 592
use scs8hd_mux2_2  mux_bottom_ipin_0.mux_l1_in_1_
timestamp 1586364061
transform 1 0 8004 0 -1 10336
box -38 -48 866 592
use scs8hd_buf_2  _33_
timestamp 1586364061
transform 1 0 9660 0 -1 10336
box -38 -48 406 592
use scs8hd_dfxbp_1  mem_bottom_ipin_0.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 8464 0 1 9248
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_140
timestamp 1586364061
transform 1 0 9568 0 -1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_0.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 9016 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_99
timestamp 1586364061
transform 1 0 10212 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_84
timestamp 1586364061
transform 1 0 8832 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_14_88
timestamp 1586364061
transform 1 0 9200 0 -1 10336
box -38 -48 406 592
use scs8hd_decap_3  FILLER_14_97
timestamp 1586364061
transform 1 0 10028 0 -1 10336
box -38 -48 314 592
use scs8hd_decap_3  FILLER_14_106
timestamp 1586364061
transform 1 0 10856 0 -1 10336
box -38 -48 314 592
use scs8hd_fill_2  FILLER_14_102
timestamp 1586364061
transform 1 0 10488 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_103
timestamp 1586364061
transform 1 0 10580 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_6.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 10764 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 10304 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 10672 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__33__A
timestamp 1586364061
transform 1 0 10396 0 1 9248
box -38 -48 222 592
use scs8hd_mux2_2  mux_bottom_ipin_6.mux_l3_in_0_
timestamp 1586364061
transform 1 0 11132 0 -1 10336
box -38 -48 866 592
use scs8hd_conb_1  _30_
timestamp 1586364061
transform 1 0 10948 0 1 9248
box -38 -48 314 592
use scs8hd_decap_4  FILLER_14_118
timestamp 1586364061
transform 1 0 11960 0 -1 10336
box -38 -48 406 592
use scs8hd_fill_2  FILLER_13_118
timestamp 1586364061
transform 1 0 11960 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_114
timestamp 1586364061
transform 1 0 11592 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_110
timestamp 1586364061
transform 1 0 11224 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_6.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 11776 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_6.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 11408 0 1 9248
box -38 -48 222 592
use scs8hd_fill_1  FILLER_14_125
timestamp 1586364061
transform 1 0 12604 0 -1 10336
box -38 -48 130 592
use scs8hd_fill_1  FILLER_14_122
timestamp 1586364061
transform 1 0 12328 0 -1 10336
box -38 -48 130 592
use scs8hd_fill_2  FILLER_13_128
timestamp 1586364061
transform 1 0 12880 0 1 9248
box -38 -48 222 592
use scs8hd_decap_3  FILLER_13_123
timestamp 1586364061
transform 1 0 12420 0 1 9248
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_6.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 12144 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_6.mux_l4_in_0__S
timestamp 1586364061
transform 1 0 12420 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_6.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 12696 0 1 9248
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_134
timestamp 1586364061
transform 1 0 12328 0 1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_6.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 13064 0 1 9248
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_bottom_ipin_6.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 12696 0 -1 10336
box -38 -48 1786 592
use scs8hd_dfxbp_1  mem_bottom_ipin_6.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 13248 0 1 9248
box -38 -48 1786 592
use scs8hd_mux2_2  mux_bottom_ipin_6.mux_l2_in_3_
timestamp 1586364061
transform 1 0 15272 0 -1 10336
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_141
timestamp 1586364061
transform 1 0 15180 0 -1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_6.mux_l2_in_3__A1
timestamp 1586364061
transform 1 0 15272 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_7.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 14996 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_6.mux_l2_in_3__A0
timestamp 1586364061
transform 1 0 15640 0 1 9248
box -38 -48 222 592
use scs8hd_decap_3  FILLER_13_151
timestamp 1586364061
transform 1 0 14996 0 1 9248
box -38 -48 314 592
use scs8hd_fill_2  FILLER_13_156
timestamp 1586364061
transform 1 0 15456 0 1 9248
box -38 -48 222 592
use scs8hd_decap_6  FILLER_14_145
timestamp 1586364061
transform 1 0 14444 0 -1 10336
box -38 -48 590 592
use scs8hd_dfxbp_1  mem_bottom_ipin_7.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 16836 0 -1 10336
box -38 -48 1786 592
use scs8hd_mux2_2  mux_bottom_ipin_7.mux_l1_in_0_
timestamp 1586364061
transform 1 0 16376 0 1 9248
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_7.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 16192 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_7.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 17388 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_7.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 16376 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_13_160
timestamp 1586364061
transform 1 0 15824 0 1 9248
box -38 -48 406 592
use scs8hd_fill_2  FILLER_13_175
timestamp 1586364061
transform 1 0 17204 0 1 9248
box -38 -48 222 592
use scs8hd_decap_3  FILLER_14_163
timestamp 1586364061
transform 1 0 16100 0 -1 10336
box -38 -48 314 592
use scs8hd_decap_3  FILLER_14_168
timestamp 1586364061
transform 1 0 16560 0 -1 10336
box -38 -48 314 592
use scs8hd_decap_3  FILLER_13_184
timestamp 1586364061
transform 1 0 18032 0 1 9248
box -38 -48 314 592
use scs8hd_fill_2  FILLER_13_179
timestamp 1586364061
transform 1 0 17572 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_8.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 17756 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_8.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 18308 0 1 9248
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_135
timestamp 1586364061
transform 1 0 17940 0 1 9248
box -38 -48 130 592
use scs8hd_decap_3  FILLER_14_198
timestamp 1586364061
transform 1 0 19320 0 -1 10336
box -38 -48 314 592
use scs8hd_fill_2  FILLER_14_194
timestamp 1586364061
transform 1 0 18952 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_190
timestamp 1586364061
transform 1 0 18584 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_7.mux_l3_in_1__A0
timestamp 1586364061
transform 1 0 19136 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_7.mux_l3_in_1__A1
timestamp 1586364061
transform 1 0 18768 0 -1 10336
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_bottom_ipin_8.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 18492 0 1 9248
box -38 -48 1786 592
use scs8hd_decap_8  FILLER_14_203
timestamp 1586364061
transform 1 0 19780 0 -1 10336
box -38 -48 774 592
use scs8hd_fill_2  FILLER_13_208
timestamp 1586364061
transform 1 0 20240 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_7.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 19596 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_8  FILLER_14_215
timestamp 1586364061
transform 1 0 20884 0 -1 10336
box -38 -48 774 592
use scs8hd_decap_3  FILLER_14_211
timestamp 1586364061
transform 1 0 20516 0 -1 10336
box -38 -48 314 592
use scs8hd_fill_2  FILLER_13_212
timestamp 1586364061
transform 1 0 20608 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_8.scs8hd_dfxbp_1_3__D
timestamp 1586364061
transform 1 0 20424 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_8.scs8hd_dfxbp_1_3__CLK
timestamp 1586364061
transform 1 0 20792 0 1 9248
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_142
timestamp 1586364061
transform 1 0 20792 0 -1 10336
box -38 -48 130 592
use scs8hd_dfxbp_1  mem_bottom_ipin_8.scs8hd_dfxbp_1_3_
timestamp 1586364061
transform 1 0 20976 0 1 9248
box -38 -48 1786 592
use scs8hd_dfxbp_1  mem_bottom_ipin_9.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 21896 0 -1 10336
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_9.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 22908 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_9.mux_l4_in_0__A0
timestamp 1586364061
transform 1 0 21712 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_235
timestamp 1586364061
transform 1 0 22724 0 1 9248
box -38 -48 222 592
use scs8hd_fill_1  FILLER_14_223
timestamp 1586364061
transform 1 0 21620 0 -1 10336
box -38 -48 130 592
use scs8hd_fill_2  FILLER_14_245
timestamp 1586364061
transform 1 0 23644 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_3  FILLER_13_245
timestamp 1586364061
transform 1 0 23644 0 1 9248
box -38 -48 314 592
use scs8hd_fill_1  FILLER_13_243
timestamp 1586364061
transform 1 0 23460 0 1 9248
box -38 -48 130 592
use scs8hd_fill_2  FILLER_13_239
timestamp 1586364061
transform 1 0 23092 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_9.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 23828 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_9.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 23276 0 1 9248
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_136
timestamp 1586364061
transform 1 0 23552 0 1 9248
box -38 -48 130 592
use scs8hd_fill_1  FILLER_14_253
timestamp 1586364061
transform 1 0 24380 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_4  FILLER_14_249
timestamp 1586364061
transform 1 0 24012 0 -1 10336
box -38 -48 406 592
use scs8hd_fill_2  FILLER_13_250
timestamp 1586364061
transform 1 0 24104 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_9.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 24472 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_9.mux_l1_in_1__A0
timestamp 1586364061
transform 1 0 23920 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_9.mux_l1_in_1__A1
timestamp 1586364061
transform 1 0 24288 0 1 9248
box -38 -48 222 592
use scs8hd_mux2_2  mux_bottom_ipin_9.mux_l1_in_1_
timestamp 1586364061
transform 1 0 24656 0 -1 10336
box -38 -48 866 592
use scs8hd_dfxbp_1  mem_bottom_ipin_9.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 24472 0 1 9248
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_143
timestamp 1586364061
transform 1 0 26404 0 -1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_9.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 26220 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_13_273
timestamp 1586364061
transform 1 0 26220 0 1 9248
box -38 -48 406 592
use scs8hd_fill_1  FILLER_13_277
timestamp 1586364061
transform 1 0 26588 0 1 9248
box -38 -48 130 592
use scs8hd_decap_8  FILLER_14_265
timestamp 1586364061
transform 1 0 25484 0 -1 10336
box -38 -48 774 592
use scs8hd_fill_2  FILLER_14_276
timestamp 1586364061
transform 1 0 26496 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_280
timestamp 1586364061
transform 1 0 26864 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_284
timestamp 1586364061
transform 1 0 27232 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_280
timestamp 1586364061
transform 1 0 26864 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_9.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 26680 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_10.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 26680 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_10.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 27048 0 1 9248
box -38 -48 222 592
use scs8hd_mux2_2  mux_bottom_ipin_10.mux_l3_in_1_
timestamp 1586364061
transform 1 0 27416 0 1 9248
box -38 -48 866 592
use scs8hd_fill_2  FILLER_13_295
timestamp 1586364061
transform 1 0 28244 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_10.mux_l3_in_1__A1
timestamp 1586364061
transform 1 0 28428 0 1 9248
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_bottom_ipin_10.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 27048 0 -1 10336
box -38 -48 1786 592
use scs8hd_decap_8  FILLER_14_301
timestamp 1586364061
transform 1 0 28796 0 -1 10336
box -38 -48 774 592
use scs8hd_fill_2  FILLER_13_306
timestamp 1586364061
transform 1 0 29256 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_303
timestamp 1586364061
transform 1 0 28980 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_299
timestamp 1586364061
transform 1 0 28612 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_10.mux_l3_in_1__A0
timestamp 1586364061
transform 1 0 28796 0 1 9248
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_137
timestamp 1586364061
transform 1 0 29164 0 1 9248
box -38 -48 130 592
use scs8hd_fill_2  FILLER_14_312
timestamp 1586364061
transform 1 0 29808 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_1  FILLER_14_309
timestamp 1586364061
transform 1 0 29532 0 -1 10336
box -38 -48 130 592
use scs8hd_fill_2  FILLER_13_314
timestamp 1586364061
transform 1 0 29992 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_14.mux_l3_in_1__A0
timestamp 1586364061
transform 1 0 29624 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_14.mux_l3_in_1__A1
timestamp 1586364061
transform 1 0 29992 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_14.mux_l3_in_1__S
timestamp 1586364061
transform 1 0 29440 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__64__A
timestamp 1586364061
transform 1 0 30176 0 1 9248
box -38 -48 222 592
use scs8hd_mux2_2  mux_bottom_ipin_14.mux_l3_in_1_
timestamp 1586364061
transform 1 0 30176 0 -1 10336
box -38 -48 866 592
use scs8hd_buf_2  _64_
timestamp 1586364061
transform 1 0 29624 0 1 9248
box -38 -48 406 592
use scs8hd_fill_2  FILLER_14_325
timestamp 1586364061
transform 1 0 31004 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_318
timestamp 1586364061
transform 1 0 30360 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_14.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 31188 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_14.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 30544 0 1 9248
box -38 -48 222 592
use scs8hd_fill_1  FILLER_14_337
timestamp 1586364061
transform 1 0 32108 0 -1 10336
box -38 -48 130 592
use scs8hd_fill_1  FILLER_14_333
timestamp 1586364061
transform 1 0 31740 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_4  FILLER_14_329
timestamp 1586364061
transform 1 0 31372 0 -1 10336
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_14.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 31832 0 -1 10336
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_144
timestamp 1586364061
transform 1 0 32016 0 -1 10336
box -38 -48 130 592
use scs8hd_dfxbp_1  mem_bottom_ipin_14.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 30728 0 1 9248
box -38 -48 1786 592
use scs8hd_dfxbp_1  mem_bottom_ipin_15.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 32200 0 -1 10336
box -38 -48 1786 592
use scs8hd_mux2_2  mux_bottom_ipin_14.mux_l1_in_0_
timestamp 1586364061
transform 1 0 33212 0 1 9248
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_14.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 33028 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_15.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 32660 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_341
timestamp 1586364061
transform 1 0 32476 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_345
timestamp 1586364061
transform 1 0 32844 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_357
timestamp 1586364061
transform 1 0 33948 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_1  FILLER_14_365
timestamp 1586364061
transform 1 0 34684 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_4  FILLER_14_361
timestamp 1586364061
transform 1 0 34316 0 -1 10336
box -38 -48 406 592
use scs8hd_fill_2  FILLER_13_362
timestamp 1586364061
transform 1 0 34408 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_358
timestamp 1586364061
transform 1 0 34040 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_15.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 34776 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_14.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 34132 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_15.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 34224 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_15.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 34592 0 1 9248
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_138
timestamp 1586364061
transform 1 0 34776 0 1 9248
box -38 -48 130 592
use scs8hd_fill_2  FILLER_13_376
timestamp 1586364061
transform 1 0 35696 0 1 9248
box -38 -48 222 592
use scs8hd_mux2_2  mux_bottom_ipin_15.mux_l1_in_0_
timestamp 1586364061
transform 1 0 34868 0 1 9248
box -38 -48 866 592
use scs8hd_dfxbp_1  mem_bottom_ipin_15.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 34960 0 -1 10336
box -38 -48 1786 592
use scs8hd_mux2_2  mux_bottom_ipin_14.mux_l2_in_1_
timestamp 1586364061
transform 1 0 36432 0 1 9248
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_14.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 36248 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_14.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 35880 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_15.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 37444 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_380
timestamp 1586364061
transform 1 0 36064 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_393
timestamp 1586364061
transform 1 0 37260 0 1 9248
box -38 -48 222 592
use scs8hd_decap_8  FILLER_14_387
timestamp 1586364061
transform 1 0 36708 0 -1 10336
box -38 -48 774 592
use scs8hd_fill_2  FILLER_14_395
timestamp 1586364061
transform 1 0 37444 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_3  PHY_27
timestamp 1586364061
transform -1 0 38824 0 1 9248
box -38 -48 314 592
use scs8hd_decap_3  PHY_29
timestamp 1586364061
transform -1 0 38824 0 -1 10336
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_145
timestamp 1586364061
transform 1 0 37628 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_8  FILLER_13_397
timestamp 1586364061
transform 1 0 37628 0 1 9248
box -38 -48 774 592
use scs8hd_fill_2  FILLER_13_405
timestamp 1586364061
transform 1 0 38364 0 1 9248
box -38 -48 222 592
use scs8hd_decap_8  FILLER_14_398
timestamp 1586364061
transform 1 0 37720 0 -1 10336
box -38 -48 774 592
use scs8hd_fill_1  FILLER_14_406
timestamp 1586364061
transform 1 0 38456 0 -1 10336
box -38 -48 130 592
use scs8hd_mux2_2  mux_bottom_ipin_1.mux_l2_in_3_
timestamp 1586364061
transform 1 0 2116 0 1 10336
box -38 -48 866 592
use scs8hd_decap_3  PHY_30
timestamp 1586364061
transform 1 0 1104 0 1 10336
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.mux_l2_in_3__A1
timestamp 1586364061
transform 1 0 1932 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.mux_l2_in_3__A0
timestamp 1586364061
transform 1 0 1564 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_3
timestamp 1586364061
transform 1 0 1380 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_7
timestamp 1586364061
transform 1 0 1748 0 1 10336
box -38 -48 222 592
use scs8hd_buf_2  _42_
timestamp 1586364061
transform 1 0 3680 0 1 10336
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l2_in_2__A1
timestamp 1586364061
transform 1 0 4600 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__42__A
timestamp 1586364061
transform 1 0 4232 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_0.scs8hd_dfxbp_1_3__CLK
timestamp 1586364061
transform 1 0 3496 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_0.scs8hd_dfxbp_1_3__D
timestamp 1586364061
transform 1 0 3128 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_20
timestamp 1586364061
transform 1 0 2944 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_24
timestamp 1586364061
transform 1 0 3312 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_32
timestamp 1586364061
transform 1 0 4048 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_36
timestamp 1586364061
transform 1 0 4416 0 1 10336
box -38 -48 222 592
use scs8hd_mux2_2  mux_bottom_ipin_0.mux_l2_in_2_
timestamp 1586364061
transform 1 0 5152 0 1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l2_in_2__A0
timestamp 1586364061
transform 1 0 4968 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l2_in_3__A1
timestamp 1586364061
transform 1 0 6532 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l2_in_3__A0
timestamp 1586364061
transform 1 0 6164 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_40
timestamp 1586364061
transform 1 0 4784 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_53
timestamp 1586364061
transform 1 0 5980 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_57
timestamp 1586364061
transform 1 0 6348 0 1 10336
box -38 -48 222 592
use scs8hd_buf_2  _37_
timestamp 1586364061
transform 1 0 6808 0 1 10336
box -38 -48 406 592
use scs8hd_dfxbp_1  mem_bottom_ipin_0.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 8188 0 1 10336
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_146
timestamp 1586364061
transform 1 0 6716 0 1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__37__A
timestamp 1586364061
transform 1 0 7360 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__34__A
timestamp 1586364061
transform 1 0 8004 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_66
timestamp 1586364061
transform 1 0 7176 0 1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_15_70
timestamp 1586364061
transform 1 0 7544 0 1 10336
box -38 -48 406 592
use scs8hd_fill_1  FILLER_15_74
timestamp 1586364061
transform 1 0 7912 0 1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_0.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 10120 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_96
timestamp 1586364061
transform 1 0 9936 0 1 10336
box -38 -48 222 592
use scs8hd_mux2_2  mux_bottom_ipin_0.mux_l3_in_0_
timestamp 1586364061
transform 1 0 10672 0 1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_0.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 10488 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_6.scs8hd_dfxbp_1_3__D
timestamp 1586364061
transform 1 0 11776 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_100
timestamp 1586364061
transform 1 0 10304 0 1 10336
box -38 -48 222 592
use scs8hd_decap_3  FILLER_15_113
timestamp 1586364061
transform 1 0 11500 0 1 10336
box -38 -48 314 592
use scs8hd_fill_2  FILLER_15_118
timestamp 1586364061
transform 1 0 11960 0 1 10336
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_bottom_ipin_6.scs8hd_dfxbp_1_3_
timestamp 1586364061
transform 1 0 12604 0 1 10336
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_147
timestamp 1586364061
transform 1 0 12328 0 1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_6.scs8hd_dfxbp_1_3__CLK
timestamp 1586364061
transform 1 0 12144 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_123
timestamp 1586364061
transform 1 0 12420 0 1 10336
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_bottom_ipin_7.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 15088 0 1 10336
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_7.mux_l2_in_2__A0
timestamp 1586364061
transform 1 0 14904 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_7.mux_l2_in_2__A1
timestamp 1586364061
transform 1 0 14536 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_144
timestamp 1586364061
transform 1 0 14352 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_148
timestamp 1586364061
transform 1 0 14720 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_7.mux_l4_in_0__S
timestamp 1586364061
transform 1 0 17020 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_7.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 17388 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_171
timestamp 1586364061
transform 1 0 16836 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_175
timestamp 1586364061
transform 1 0 17204 0 1 10336
box -38 -48 222 592
use scs8hd_mux2_2  mux_bottom_ipin_7.mux_l2_in_0_
timestamp 1586364061
transform 1 0 18032 0 1 10336
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_148
timestamp 1586364061
transform 1 0 17940 0 1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_7.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 17756 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_7.mux_l3_in_1__S
timestamp 1586364061
transform 1 0 19044 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_179
timestamp 1586364061
transform 1 0 17572 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_193
timestamp 1586364061
transform 1 0 18860 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_197
timestamp 1586364061
transform 1 0 19228 0 1 10336
box -38 -48 222 592
use scs8hd_mux2_2  mux_bottom_ipin_7.mux_l2_in_1_
timestamp 1586364061
transform 1 0 19596 0 1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_7.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 19412 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_7.scs8hd_dfxbp_1_3__CLK
timestamp 1586364061
transform 1 0 20884 0 1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_15_210
timestamp 1586364061
transform 1 0 20424 0 1 10336
box -38 -48 406 592
use scs8hd_fill_1  FILLER_15_214
timestamp 1586364061
transform 1 0 20792 0 1 10336
box -38 -48 130 592
use scs8hd_fill_2  FILLER_15_217
timestamp 1586364061
transform 1 0 21068 0 1 10336
box -38 -48 222 592
use scs8hd_mux2_2  mux_bottom_ipin_9.mux_l2_in_1_
timestamp 1586364061
transform 1 0 21988 0 1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_9.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 21804 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_7.scs8hd_dfxbp_1_3__D
timestamp 1586364061
transform 1 0 21252 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_9.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 23000 0 1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_15_221
timestamp 1586364061
transform 1 0 21436 0 1 10336
box -38 -48 406 592
use scs8hd_fill_2  FILLER_15_236
timestamp 1586364061
transform 1 0 22816 0 1 10336
box -38 -48 222 592
use scs8hd_mux2_2  mux_bottom_ipin_9.mux_l3_in_0_
timestamp 1586364061
transform 1 0 23736 0 1 10336
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_149
timestamp 1586364061
transform 1 0 23552 0 1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_9.mux_l4_in_0__S
timestamp 1586364061
transform 1 0 23368 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_240
timestamp 1586364061
transform 1 0 23184 0 1 10336
box -38 -48 222 592
use scs8hd_fill_1  FILLER_15_245
timestamp 1586364061
transform 1 0 23644 0 1 10336
box -38 -48 130 592
use scs8hd_decap_4  FILLER_15_255
timestamp 1586364061
transform 1 0 24564 0 1 10336
box -38 -48 406 592
use scs8hd_conb_1  _18_
timestamp 1586364061
transform 1 0 25300 0 1 10336
box -38 -48 314 592
use scs8hd_dfxbp_1  mem_bottom_ipin_9.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 26404 0 1 10336
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_9.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 26220 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_9.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 25852 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_10.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 24932 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_261
timestamp 1586364061
transform 1 0 25116 0 1 10336
box -38 -48 222 592
use scs8hd_decap_3  FILLER_15_266
timestamp 1586364061
transform 1 0 25576 0 1 10336
box -38 -48 314 592
use scs8hd_fill_2  FILLER_15_271
timestamp 1586364061
transform 1 0 26036 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_9.scs8hd_dfxbp_1_3__CLK
timestamp 1586364061
transform 1 0 28336 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_294
timestamp 1586364061
transform 1 0 28152 0 1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_15_306
timestamp 1586364061
transform 1 0 29256 0 1 10336
box -38 -48 406 592
use scs8hd_decap_3  FILLER_15_302
timestamp 1586364061
transform 1 0 28888 0 1 10336
box -38 -48 314 592
use scs8hd_fill_2  FILLER_15_298
timestamp 1586364061
transform 1 0 28520 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_9.scs8hd_dfxbp_1_3__D
timestamp 1586364061
transform 1 0 28704 0 1 10336
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_150
timestamp 1586364061
transform 1 0 29164 0 1 10336
box -38 -48 130 592
use scs8hd_fill_2  FILLER_15_313
timestamp 1586364061
transform 1 0 29900 0 1 10336
box -38 -48 222 592
use scs8hd_fill_1  FILLER_15_310
timestamp 1586364061
transform 1 0 29624 0 1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_14.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 29716 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_14.scs8hd_dfxbp_1_3__CLK
timestamp 1586364061
transform 1 0 30084 0 1 10336
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_bottom_ipin_14.scs8hd_dfxbp_1_3_
timestamp 1586364061
transform 1 0 30268 0 1 10336
box -38 -48 1786 592
use scs8hd_fill_2  FILLER_15_336
timestamp 1586364061
transform 1 0 32016 0 1 10336
box -38 -48 222 592
use scs8hd_mux2_2  mux_bottom_ipin_15.mux_l3_in_0_
timestamp 1586364061
transform 1 0 33212 0 1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_15.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 32936 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_15.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 32568 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_15.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 32200 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_340
timestamp 1586364061
transform 1 0 32384 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_344
timestamp 1586364061
transform 1 0 32752 0 1 10336
box -38 -48 222 592
use scs8hd_fill_1  FILLER_15_348
timestamp 1586364061
transform 1 0 33120 0 1 10336
box -38 -48 130 592
use scs8hd_mux2_2  mux_bottom_ipin_15.mux_l2_in_0_
timestamp 1586364061
transform 1 0 34868 0 1 10336
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_151
timestamp 1586364061
transform 1 0 34776 0 1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_15.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 34592 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_15.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 34224 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_358
timestamp 1586364061
transform 1 0 34040 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_362
timestamp 1586364061
transform 1 0 34408 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_376
timestamp 1586364061
transform 1 0 35696 0 1 10336
box -38 -48 222 592
use scs8hd_buf_2  _69_
timestamp 1586364061
transform 1 0 36432 0 1 10336
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_15.mux_l2_in_2__A0
timestamp 1586364061
transform 1 0 35880 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__69__A
timestamp 1586364061
transform 1 0 36984 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_15.mux_l2_in_2__A1
timestamp 1586364061
transform 1 0 36248 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_380
timestamp 1586364061
transform 1 0 36064 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_388
timestamp 1586364061
transform 1 0 36800 0 1 10336
box -38 -48 222 592
use scs8hd_decap_12  FILLER_15_392
timestamp 1586364061
transform 1 0 37168 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_3  PHY_31
timestamp 1586364061
transform -1 0 38824 0 1 10336
box -38 -48 314 592
use scs8hd_decap_3  FILLER_15_404
timestamp 1586364061
transform 1 0 38272 0 1 10336
box -38 -48 314 592
use scs8hd_conb_1  _20_
timestamp 1586364061
transform 1 0 1380 0 -1 11424
box -38 -48 314 592
use scs8hd_mux2_2  mux_bottom_ipin_1.mux_l3_in_0_
timestamp 1586364061
transform 1 0 2392 0 -1 11424
box -38 -48 866 592
use scs8hd_decap_3  PHY_32
timestamp 1586364061
transform 1 0 1104 0 -1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.mux_l2_in_2__A1
timestamp 1586364061
transform 1 0 1932 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_3  FILLER_16_6
timestamp 1586364061
transform 1 0 1656 0 -1 11424
box -38 -48 314 592
use scs8hd_decap_3  FILLER_16_11
timestamp 1586364061
transform 1 0 2116 0 -1 11424
box -38 -48 314 592
use scs8hd_dfxbp_1  mem_bottom_ipin_0.scs8hd_dfxbp_1_3_
timestamp 1586364061
transform 1 0 4048 0 -1 11424
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_152
timestamp 1586364061
transform 1 0 3956 0 -1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l4_in_0__A1
timestamp 1586364061
transform 1 0 3496 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_3  FILLER_16_23
timestamp 1586364061
transform 1 0 3220 0 -1 11424
box -38 -48 314 592
use scs8hd_decap_3  FILLER_16_28
timestamp 1586364061
transform 1 0 3680 0 -1 11424
box -38 -48 314 592
use scs8hd_mux2_2  mux_bottom_ipin_0.mux_l2_in_3_
timestamp 1586364061
transform 1 0 6532 0 -1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l2_in_3__S
timestamp 1586364061
transform 1 0 6348 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l2_in_2__S
timestamp 1586364061
transform 1 0 5980 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_51
timestamp 1586364061
transform 1 0 5796 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_55
timestamp 1586364061
transform 1 0 6164 0 -1 11424
box -38 -48 222 592
use scs8hd_buf_2  _34_
timestamp 1586364061
transform 1 0 8096 0 -1 11424
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 7912 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_6  FILLER_16_68
timestamp 1586364061
transform 1 0 7360 0 -1 11424
box -38 -48 590 592
use scs8hd_dfxbp_1  mem_bottom_ipin_0.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 9660 0 -1 11424
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_153
timestamp 1586364061
transform 1 0 9568 0 -1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_0.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 8648 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_0.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 9016 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_80
timestamp 1586364061
transform 1 0 8464 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_84
timestamp 1586364061
transform 1 0 8832 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_16_88
timestamp 1586364061
transform 1 0 9200 0 -1 11424
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_5.mux_l4_in_0__A1
timestamp 1586364061
transform 1 0 11592 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_5.mux_l4_in_0__A0
timestamp 1586364061
transform 1 0 11960 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_112
timestamp 1586364061
transform 1 0 11408 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_116
timestamp 1586364061
transform 1 0 11776 0 -1 11424
box -38 -48 222 592
use scs8hd_mux2_2  mux_bottom_ipin_6.mux_l4_in_0_
timestamp 1586364061
transform 1 0 12420 0 -1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_6.mux_l4_in_0__A1
timestamp 1586364061
transform 1 0 13432 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_6.mux_l4_in_0__A0
timestamp 1586364061
transform 1 0 13800 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_3  FILLER_16_120
timestamp 1586364061
transform 1 0 12144 0 -1 11424
box -38 -48 314 592
use scs8hd_fill_2  FILLER_16_132
timestamp 1586364061
transform 1 0 13248 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_136
timestamp 1586364061
transform 1 0 13616 0 -1 11424
box -38 -48 222 592
use scs8hd_mux2_2  mux_bottom_ipin_7.mux_l2_in_2_
timestamp 1586364061
transform 1 0 15272 0 -1 11424
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_154
timestamp 1586364061
transform 1 0 15180 0 -1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_7.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 14996 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_8  FILLER_16_140
timestamp 1586364061
transform 1 0 13984 0 -1 11424
box -38 -48 774 592
use scs8hd_decap_3  FILLER_16_148
timestamp 1586364061
transform 1 0 14720 0 -1 11424
box -38 -48 314 592
use scs8hd_mux2_2  mux_bottom_ipin_7.mux_l4_in_0_
timestamp 1586364061
transform 1 0 16836 0 -1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_7.mux_l2_in_3__A0
timestamp 1586364061
transform 1 0 16376 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_3  FILLER_16_163
timestamp 1586364061
transform 1 0 16100 0 -1 11424
box -38 -48 314 592
use scs8hd_decap_3  FILLER_16_168
timestamp 1586364061
transform 1 0 16560 0 -1 11424
box -38 -48 314 592
use scs8hd_mux2_2  mux_bottom_ipin_7.mux_l3_in_1_
timestamp 1586364061
transform 1 0 18400 0 -1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_7.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 18032 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_16_180
timestamp 1586364061
transform 1 0 17664 0 -1 11424
box -38 -48 406 592
use scs8hd_fill_2  FILLER_16_186
timestamp 1586364061
transform 1 0 18216 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_16_197
timestamp 1586364061
transform 1 0 19228 0 -1 11424
box -38 -48 406 592
use scs8hd_dfxbp_1  mem_bottom_ipin_7.scs8hd_dfxbp_1_3_
timestamp 1586364061
transform 1 0 20884 0 -1 11424
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_155
timestamp 1586364061
transform 1 0 20792 0 -1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_7.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 19596 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_8  FILLER_16_203
timestamp 1586364061
transform 1 0 19780 0 -1 11424
box -38 -48 774 592
use scs8hd_decap_3  FILLER_16_211
timestamp 1586364061
transform 1 0 20516 0 -1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_9.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 22816 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_234
timestamp 1586364061
transform 1 0 22632 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_238
timestamp 1586364061
transform 1 0 23000 0 -1 11424
box -38 -48 222 592
use scs8hd_mux2_2  mux_bottom_ipin_9.mux_l4_in_0_
timestamp 1586364061
transform 1 0 23368 0 -1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_9.mux_l2_in_3__A0
timestamp 1586364061
transform 1 0 24380 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_9.mux_l2_in_3__S
timestamp 1586364061
transform 1 0 24748 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_9.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 23184 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_251
timestamp 1586364061
transform 1 0 24196 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_255
timestamp 1586364061
transform 1 0 24564 0 -1 11424
box -38 -48 222 592
use scs8hd_buf_4  mux_bottom_ipin_10.scs8hd_buf_4_0_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 24932 0 -1 11424
box -38 -48 590 592
use scs8hd_mux2_2  mux_bottom_ipin_9.mux_l2_in_0_
timestamp 1586364061
transform 1 0 26496 0 -1 11424
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_156
timestamp 1586364061
transform 1 0 26404 0 -1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_9.mux_l2_in_2__S
timestamp 1586364061
transform 1 0 25668 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_9.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 26220 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_265
timestamp 1586364061
transform 1 0 25484 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_16_269
timestamp 1586364061
transform 1 0 25852 0 -1 11424
box -38 -48 406 592
use scs8hd_dfxbp_1  mem_bottom_ipin_9.scs8hd_dfxbp_1_3_
timestamp 1586364061
transform 1 0 28152 0 -1 11424
box -38 -48 1786 592
use scs8hd_decap_8  FILLER_16_285
timestamp 1586364061
transform 1 0 27324 0 -1 11424
box -38 -48 774 592
use scs8hd_fill_1  FILLER_16_293
timestamp 1586364061
transform 1 0 28060 0 -1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_14.scs8hd_dfxbp_1_3__D
timestamp 1586364061
transform 1 0 30268 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_16_313
timestamp 1586364061
transform 1 0 29900 0 -1 11424
box -38 -48 406 592
use scs8hd_buf_4  mux_bottom_ipin_14.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 30636 0 -1 11424
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_157
timestamp 1586364061
transform 1 0 32016 0 -1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_15.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 31832 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_319
timestamp 1586364061
transform 1 0 30452 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_6  FILLER_16_327
timestamp 1586364061
transform 1 0 31188 0 -1 11424
box -38 -48 590 592
use scs8hd_fill_1  FILLER_16_333
timestamp 1586364061
transform 1 0 31740 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_3  FILLER_16_337
timestamp 1586364061
transform 1 0 32108 0 -1 11424
box -38 -48 314 592
use scs8hd_dfxbp_1  mem_bottom_ipin_15.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 32936 0 -1 11424
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_15.mux_l2_in_3__S
timestamp 1586364061
transform 1 0 32752 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_15.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 32384 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_342
timestamp 1586364061
transform 1 0 32568 0 -1 11424
box -38 -48 222 592
use scs8hd_mux2_2  mux_bottom_ipin_15.mux_l2_in_2_
timestamp 1586364061
transform 1 0 35420 0 -1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_15.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 34868 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_15.mux_l2_in_2__S
timestamp 1586364061
transform 1 0 35236 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_365
timestamp 1586364061
transform 1 0 34684 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_369
timestamp 1586364061
transform 1 0 35052 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_15.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 36432 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_382
timestamp 1586364061
transform 1 0 36248 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_8  FILLER_16_386
timestamp 1586364061
transform 1 0 36616 0 -1 11424
box -38 -48 774 592
use scs8hd_decap_3  FILLER_16_394
timestamp 1586364061
transform 1 0 37352 0 -1 11424
box -38 -48 314 592
use scs8hd_decap_3  PHY_33
timestamp 1586364061
transform -1 0 38824 0 -1 11424
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_158
timestamp 1586364061
transform 1 0 37628 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_8  FILLER_16_398
timestamp 1586364061
transform 1 0 37720 0 -1 11424
box -38 -48 774 592
use scs8hd_fill_1  FILLER_16_406
timestamp 1586364061
transform 1 0 38456 0 -1 11424
box -38 -48 130 592
use scs8hd_mux2_2  mux_bottom_ipin_1.mux_l2_in_2_
timestamp 1586364061
transform 1 0 1932 0 1 11424
box -38 -48 866 592
use scs8hd_decap_3  PHY_34
timestamp 1586364061
transform 1 0 1104 0 1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.mux_l2_in_2__A0
timestamp 1586364061
transform 1 0 1748 0 1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_17_3
timestamp 1586364061
transform 1 0 1380 0 1 11424
box -38 -48 406 592
use scs8hd_fill_2  FILLER_17_18
timestamp 1586364061
transform 1 0 2760 0 1 11424
box -38 -48 222 592
use scs8hd_mux2_2  mux_bottom_ipin_0.mux_l4_in_0_
timestamp 1586364061
transform 1 0 3496 0 1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.mux_l1_in_2__A0
timestamp 1586364061
transform 1 0 4508 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__46__A
timestamp 1586364061
transform 1 0 2944 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l4_in_0__S
timestamp 1586364061
transform 1 0 3312 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_22
timestamp 1586364061
transform 1 0 3128 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_35
timestamp 1586364061
transform 1 0 4324 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_39
timestamp 1586364061
transform 1 0 4692 0 1 11424
box -38 -48 222 592
use scs8hd_mux2_2  mux_bottom_ipin_1.mux_l1_in_2_
timestamp 1586364061
transform 1 0 5060 0 1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.mux_l1_in_2__A1
timestamp 1586364061
transform 1 0 4876 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__39__A
timestamp 1586364061
transform 1 0 6440 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l3_in_1__S
timestamp 1586364061
transform 1 0 6072 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_52
timestamp 1586364061
transform 1 0 5888 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_56
timestamp 1586364061
transform 1 0 6256 0 1 11424
box -38 -48 222 592
use scs8hd_buf_2  _40_
timestamp 1586364061
transform 1 0 6808 0 1 11424
box -38 -48 406 592
use scs8hd_mux2_2  mux_bottom_ipin_0.mux_l2_in_0_
timestamp 1586364061
transform 1 0 8096 0 1 11424
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_159
timestamp 1586364061
transform 1 0 6716 0 1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 7912 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__40__A
timestamp 1586364061
transform 1 0 7360 0 1 11424
box -38 -48 222 592
use scs8hd_fill_1  FILLER_17_60
timestamp 1586364061
transform 1 0 6624 0 1 11424
box -38 -48 130 592
use scs8hd_fill_2  FILLER_17_66
timestamp 1586364061
transform 1 0 7176 0 1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_17_70
timestamp 1586364061
transform 1 0 7544 0 1 11424
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 9108 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 9476 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_85
timestamp 1586364061
transform 1 0 8924 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_89
timestamp 1586364061
transform 1 0 9292 0 1 11424
box -38 -48 222 592
use scs8hd_decap_8  FILLER_17_93
timestamp 1586364061
transform 1 0 9660 0 1 11424
box -38 -48 774 592
use scs8hd_buf_4  mux_bottom_ipin_5.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 11040 0 1 11424
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_5.mux_l4_in_0__S
timestamp 1586364061
transform 1 0 11776 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 10672 0 1 11424
box -38 -48 222 592
use scs8hd_decap_3  FILLER_17_101
timestamp 1586364061
transform 1 0 10396 0 1 11424
box -38 -48 314 592
use scs8hd_fill_2  FILLER_17_106
timestamp 1586364061
transform 1 0 10856 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_114
timestamp 1586364061
transform 1 0 11592 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_118
timestamp 1586364061
transform 1 0 11960 0 1 11424
box -38 -48 222 592
use scs8hd_mux2_2  mux_bottom_ipin_6.mux_l1_in_0_
timestamp 1586364061
transform 1 0 12880 0 1 11424
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_160
timestamp 1586364061
transform 1 0 12328 0 1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_6.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 12696 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_6.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 12144 0 1 11424
box -38 -48 222 592
use scs8hd_decap_3  FILLER_17_123
timestamp 1586364061
transform 1 0 12420 0 1 11424
box -38 -48 314 592
use scs8hd_decap_12  FILLER_17_137
timestamp 1586364061
transform 1 0 13708 0 1 11424
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_7.mux_l2_in_2__S
timestamp 1586364061
transform 1 0 15272 0 1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_17_149
timestamp 1586364061
transform 1 0 14812 0 1 11424
box -38 -48 406 592
use scs8hd_fill_1  FILLER_17_153
timestamp 1586364061
transform 1 0 15180 0 1 11424
box -38 -48 130 592
use scs8hd_decap_4  FILLER_17_156
timestamp 1586364061
transform 1 0 15456 0 1 11424
box -38 -48 406 592
use scs8hd_mux2_2  mux_bottom_ipin_7.mux_l2_in_3_
timestamp 1586364061
transform 1 0 16376 0 1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_7.mux_l2_in_3__A1
timestamp 1586364061
transform 1 0 16192 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_7.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 17388 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_7.mux_l4_in_0__A0
timestamp 1586364061
transform 1 0 15824 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_162
timestamp 1586364061
transform 1 0 16008 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_175
timestamp 1586364061
transform 1 0 17204 0 1 11424
box -38 -48 222 592
use scs8hd_conb_1  _16_
timestamp 1586364061
transform 1 0 18032 0 1 11424
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_161
timestamp 1586364061
transform 1 0 17940 0 1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_7.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 19228 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_7.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 17756 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_7.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 18492 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_179
timestamp 1586364061
transform 1 0 17572 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_187
timestamp 1586364061
transform 1 0 18308 0 1 11424
box -38 -48 222 592
use scs8hd_decap_6  FILLER_17_191
timestamp 1586364061
transform 1 0 18676 0 1 11424
box -38 -48 590 592
use scs8hd_dfxbp_1  mem_bottom_ipin_7.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 19412 0 1 11424
box -38 -48 1786 592
use scs8hd_fill_2  FILLER_17_218
timestamp 1586364061
transform 1 0 21160 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_8.mux_l2_in_3__A1
timestamp 1586364061
transform 1 0 21344 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_8.mux_l2_in_3__A0
timestamp 1586364061
transform 1 0 21712 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_8.mux_l2_in_3__S
timestamp 1586364061
transform 1 0 22080 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_9.mux_l3_in_1__A1
timestamp 1586364061
transform 1 0 23000 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_9.mux_l4_in_0__A1
timestamp 1586364061
transform 1 0 22632 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_222
timestamp 1586364061
transform 1 0 21528 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_226
timestamp 1586364061
transform 1 0 21896 0 1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_17_230
timestamp 1586364061
transform 1 0 22264 0 1 11424
box -38 -48 406 592
use scs8hd_fill_2  FILLER_17_236
timestamp 1586364061
transform 1 0 22816 0 1 11424
box -38 -48 222 592
use scs8hd_mux2_2  mux_bottom_ipin_9.mux_l3_in_1_
timestamp 1586364061
transform 1 0 23920 0 1 11424
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_162
timestamp 1586364061
transform 1 0 23552 0 1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_9.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 23368 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_240
timestamp 1586364061
transform 1 0 23184 0 1 11424
box -38 -48 222 592
use scs8hd_decap_3  FILLER_17_245
timestamp 1586364061
transform 1 0 23644 0 1 11424
box -38 -48 314 592
use scs8hd_fill_2  FILLER_17_257
timestamp 1586364061
transform 1 0 24748 0 1 11424
box -38 -48 222 592
use scs8hd_mux2_2  mux_bottom_ipin_9.mux_l2_in_2_
timestamp 1586364061
transform 1 0 25484 0 1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_9.mux_l2_in_2__A0
timestamp 1586364061
transform 1 0 25300 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_9.mux_l2_in_3__A1
timestamp 1586364061
transform 1 0 24932 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_9.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 26496 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_261
timestamp 1586364061
transform 1 0 25116 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_274
timestamp 1586364061
transform 1 0 26312 0 1 11424
box -38 -48 222 592
use scs8hd_mux2_2  mux_bottom_ipin_9.mux_l1_in_0_
timestamp 1586364061
transform 1 0 27048 0 1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_9.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 26864 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_278
timestamp 1586364061
transform 1 0 26680 0 1 11424
box -38 -48 222 592
use scs8hd_decap_12  FILLER_17_291
timestamp 1586364061
transform 1 0 27876 0 1 11424
box -38 -48 1142 592
use scs8hd_buf_2  _60_
timestamp 1586364061
transform 1 0 29348 0 1 11424
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_163
timestamp 1586364061
transform 1 0 29164 0 1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__60__A
timestamp 1586364061
transform 1 0 29900 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_14.mux_l4_in_0__S
timestamp 1586364061
transform 1 0 30268 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_303
timestamp 1586364061
transform 1 0 28980 0 1 11424
box -38 -48 222 592
use scs8hd_fill_1  FILLER_17_306
timestamp 1586364061
transform 1 0 29256 0 1 11424
box -38 -48 130 592
use scs8hd_fill_2  FILLER_17_311
timestamp 1586364061
transform 1 0 29716 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_315
timestamp 1586364061
transform 1 0 30084 0 1 11424
box -38 -48 222 592
use scs8hd_buf_2  _62_
timestamp 1586364061
transform 1 0 32108 0 1 11424
box -38 -48 406 592
use scs8hd_mux2_2  mux_bottom_ipin_14.mux_l4_in_0_
timestamp 1586364061
transform 1 0 30452 0 1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__59__A
timestamp 1586364061
transform 1 0 31464 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__62__A
timestamp 1586364061
transform 1 0 31924 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_328
timestamp 1586364061
transform 1 0 31280 0 1 11424
box -38 -48 222 592
use scs8hd_decap_3  FILLER_17_332
timestamp 1586364061
transform 1 0 31648 0 1 11424
box -38 -48 314 592
use scs8hd_mux2_2  mux_bottom_ipin_15.mux_l2_in_3_
timestamp 1586364061
transform 1 0 33212 0 1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__58__A
timestamp 1586364061
transform 1 0 32660 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_15.mux_l2_in_3__A1
timestamp 1586364061
transform 1 0 33028 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_341
timestamp 1586364061
transform 1 0 32476 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_345
timestamp 1586364061
transform 1 0 32844 0 1 11424
box -38 -48 222 592
use scs8hd_mux2_2  mux_bottom_ipin_15.mux_l2_in_1_
timestamp 1586364061
transform 1 0 34868 0 1 11424
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_164
timestamp 1586364061
transform 1 0 34776 0 1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_15.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 34592 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_15.scs8hd_dfxbp_1_3__CLK
timestamp 1586364061
transform 1 0 34224 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_358
timestamp 1586364061
transform 1 0 34040 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_362
timestamp 1586364061
transform 1 0 34408 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_376
timestamp 1586364061
transform 1 0 35696 0 1 11424
box -38 -48 222 592
use scs8hd_conb_1  _26_
timestamp 1586364061
transform 1 0 37536 0 1 11424
box -38 -48 314 592
use scs8hd_buf_2  _68_
timestamp 1586364061
transform 1 0 36432 0 1 11424
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__68__A
timestamp 1586364061
transform 1 0 36984 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_15.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 35880 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_15.scs8hd_dfxbp_1_3__D
timestamp 1586364061
transform 1 0 36248 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_380
timestamp 1586364061
transform 1 0 36064 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_388
timestamp 1586364061
transform 1 0 36800 0 1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_17_392
timestamp 1586364061
transform 1 0 37168 0 1 11424
box -38 -48 406 592
use scs8hd_decap_3  PHY_35
timestamp 1586364061
transform -1 0 38824 0 1 11424
box -38 -48 314 592
use scs8hd_decap_8  FILLER_17_399
timestamp 1586364061
transform 1 0 37812 0 1 11424
box -38 -48 774 592
use scs8hd_buf_2  _46_
timestamp 1586364061
transform 1 0 2668 0 -1 12512
box -38 -48 406 592
use scs8hd_buf_4  mux_bottom_ipin_0.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 1380 0 -1 12512
box -38 -48 590 592
use scs8hd_decap_3  PHY_36
timestamp 1586364061
transform 1 0 1104 0 -1 12512
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.mux_l2_in_2__S
timestamp 1586364061
transform 1 0 2116 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 2484 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_9
timestamp 1586364061
transform 1 0 1932 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_13
timestamp 1586364061
transform 1 0 2300 0 -1 12512
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_165
timestamp 1586364061
transform 1 0 3956 0 -1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 4232 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l3_in_1__A1
timestamp 1586364061
transform 1 0 4692 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l4_in_0__A0
timestamp 1586364061
transform 1 0 3496 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_18_21
timestamp 1586364061
transform 1 0 3036 0 -1 12512
box -38 -48 406 592
use scs8hd_fill_1  FILLER_18_25
timestamp 1586364061
transform 1 0 3404 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_3  FILLER_18_28
timestamp 1586364061
transform 1 0 3680 0 -1 12512
box -38 -48 314 592
use scs8hd_fill_2  FILLER_18_32
timestamp 1586364061
transform 1 0 4048 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_3  FILLER_18_36
timestamp 1586364061
transform 1 0 4416 0 -1 12512
box -38 -48 314 592
use scs8hd_buf_2  _39_
timestamp 1586364061
transform 1 0 6440 0 -1 12512
box -38 -48 406 592
use scs8hd_mux2_2  mux_bottom_ipin_0.mux_l3_in_1_
timestamp 1586364061
transform 1 0 4876 0 -1 12512
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.mux_l1_in_2__S
timestamp 1586364061
transform 1 0 5888 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_50
timestamp 1586364061
transform 1 0 5704 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_18_54
timestamp 1586364061
transform 1 0 6072 0 -1 12512
box -38 -48 406 592
use scs8hd_mux2_2  mux_bottom_ipin_0.mux_l2_in_1_
timestamp 1586364061
transform 1 0 7912 0 -1 12512
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 7728 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_8  FILLER_18_62
timestamp 1586364061
transform 1 0 6808 0 -1 12512
box -38 -48 774 592
use scs8hd_fill_2  FILLER_18_70
timestamp 1586364061
transform 1 0 7544 0 -1 12512
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_166
timestamp 1586364061
transform 1 0 9568 0 -1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 8924 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_83
timestamp 1586364061
transform 1 0 8740 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_18_87
timestamp 1586364061
transform 1 0 9108 0 -1 12512
box -38 -48 406 592
use scs8hd_fill_1  FILLER_18_91
timestamp 1586364061
transform 1 0 9476 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_12  FILLER_18_93
timestamp 1586364061
transform 1 0 9660 0 -1 12512
box -38 -48 1142 592
use scs8hd_mux2_2  mux_bottom_ipin_5.mux_l4_in_0_
timestamp 1586364061
transform 1 0 11408 0 -1 12512
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_5.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 11040 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_3  FILLER_18_105
timestamp 1586364061
transform 1 0 10764 0 -1 12512
box -38 -48 314 592
use scs8hd_fill_2  FILLER_18_110
timestamp 1586364061
transform 1 0 11224 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_6.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 12880 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_6  FILLER_18_121
timestamp 1586364061
transform 1 0 12236 0 -1 12512
box -38 -48 590 592
use scs8hd_fill_1  FILLER_18_127
timestamp 1586364061
transform 1 0 12788 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_12  FILLER_18_130
timestamp 1586364061
transform 1 0 13064 0 -1 12512
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_167
timestamp 1586364061
transform 1 0 15180 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_8  FILLER_18_142
timestamp 1586364061
transform 1 0 14168 0 -1 12512
box -38 -48 774 592
use scs8hd_decap_3  FILLER_18_150
timestamp 1586364061
transform 1 0 14904 0 -1 12512
box -38 -48 314 592
use scs8hd_decap_12  FILLER_18_154
timestamp 1586364061
transform 1 0 15272 0 -1 12512
box -38 -48 1142 592
use scs8hd_mux2_2  mux_bottom_ipin_7.mux_l3_in_0_
timestamp 1586364061
transform 1 0 17204 0 -1 12512
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_7.mux_l2_in_3__S
timestamp 1586364061
transform 1 0 16376 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_7.mux_l4_in_0__A1
timestamp 1586364061
transform 1 0 16836 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_3  FILLER_18_168
timestamp 1586364061
transform 1 0 16560 0 -1 12512
box -38 -48 314 592
use scs8hd_fill_2  FILLER_18_173
timestamp 1586364061
transform 1 0 17020 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_12  FILLER_18_184
timestamp 1586364061
transform 1 0 18032 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_18_196
timestamp 1586364061
transform 1 0 19136 0 -1 12512
box -38 -48 314 592
use scs8hd_mux2_2  mux_bottom_ipin_8.mux_l2_in_3_
timestamp 1586364061
transform 1 0 20884 0 -1 12512
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_168
timestamp 1586364061
transform 1 0 20792 0 -1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_7.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 19412 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_12  FILLER_18_201
timestamp 1586364061
transform 1 0 19596 0 -1 12512
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_18_213
timestamp 1586364061
transform 1 0 20700 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_12  FILLER_18_224
timestamp 1586364061
transform 1 0 21712 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_18_236
timestamp 1586364061
transform 1 0 22816 0 -1 12512
box -38 -48 774 592
use scs8hd_mux2_2  mux_bottom_ipin_9.mux_l2_in_3_
timestamp 1586364061
transform 1 0 24380 0 -1 12512
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_9.mux_l3_in_1__S
timestamp 1586364061
transform 1 0 23920 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_9.mux_l3_in_1__A0
timestamp 1586364061
transform 1 0 23552 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_246
timestamp 1586364061
transform 1 0 23736 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_3  FILLER_18_250
timestamp 1586364061
transform 1 0 24104 0 -1 12512
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_169
timestamp 1586364061
transform 1 0 26404 0 -1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_9.mux_l2_in_2__A1
timestamp 1586364061
transform 1 0 25484 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_3  FILLER_18_262
timestamp 1586364061
transform 1 0 25208 0 -1 12512
box -38 -48 314 592
use scs8hd_decap_8  FILLER_18_267
timestamp 1586364061
transform 1 0 25668 0 -1 12512
box -38 -48 774 592
use scs8hd_decap_6  FILLER_18_276
timestamp 1586364061
transform 1 0 26496 0 -1 12512
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_9.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 27048 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_12  FILLER_18_284
timestamp 1586364061
transform 1 0 27232 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_296
timestamp 1586364061
transform 1 0 28336 0 -1 12512
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_14.mux_l4_in_0__A0
timestamp 1586364061
transform 1 0 30084 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_6  FILLER_18_308
timestamp 1586364061
transform 1 0 29440 0 -1 12512
box -38 -48 590 592
use scs8hd_fill_1  FILLER_18_314
timestamp 1586364061
transform 1 0 29992 0 -1 12512
box -38 -48 130 592
use scs8hd_fill_2  FILLER_18_317
timestamp 1586364061
transform 1 0 30268 0 -1 12512
box -38 -48 222 592
use scs8hd_buf_2  _58_
timestamp 1586364061
transform 1 0 32108 0 -1 12512
box -38 -48 406 592
use scs8hd_buf_2  _59_
timestamp 1586364061
transform 1 0 30912 0 -1 12512
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_170
timestamp 1586364061
transform 1 0 32016 0 -1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_14.mux_l4_in_0__A1
timestamp 1586364061
transform 1 0 30452 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_3  FILLER_18_321
timestamp 1586364061
transform 1 0 30636 0 -1 12512
box -38 -48 314 592
use scs8hd_decap_8  FILLER_18_328
timestamp 1586364061
transform 1 0 31280 0 -1 12512
box -38 -48 774 592
use scs8hd_mux2_2  mux_bottom_ipin_15.mux_l3_in_1_
timestamp 1586364061
transform 1 0 33212 0 -1 12512
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_15.mux_l2_in_3__A0
timestamp 1586364061
transform 1 0 33028 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_15.mux_l3_in_1__S
timestamp 1586364061
transform 1 0 32660 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_341
timestamp 1586364061
transform 1 0 32476 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_345
timestamp 1586364061
transform 1 0 32844 0 -1 12512
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_bottom_ipin_15.scs8hd_dfxbp_1_3_
timestamp 1586364061
transform 1 0 34776 0 -1 12512
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_15.mux_l3_in_1__A1
timestamp 1586364061
transform 1 0 34224 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_15.mux_l3_in_1__A0
timestamp 1586364061
transform 1 0 34592 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_358
timestamp 1586364061
transform 1 0 34040 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_362
timestamp 1586364061
transform 1 0 34408 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_12  FILLER_18_385
timestamp 1586364061
transform 1 0 36524 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_3  PHY_37
timestamp 1586364061
transform -1 0 38824 0 -1 12512
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_171
timestamp 1586364061
transform 1 0 37628 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_8  FILLER_18_398
timestamp 1586364061
transform 1 0 37720 0 -1 12512
box -38 -48 774 592
use scs8hd_fill_1  FILLER_18_406
timestamp 1586364061
transform 1 0 38456 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_8  FILLER_20_7
timestamp 1586364061
transform 1 0 1748 0 -1 13600
box -38 -48 774 592
use scs8hd_fill_1  FILLER_19_7
timestamp 1586364061
transform 1 0 1748 0 1 12512
box -38 -48 130 592
use scs8hd_fill_2  FILLER_19_3
timestamp 1586364061
transform 1 0 1380 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__47__A
timestamp 1586364061
transform 1 0 1564 0 1 12512
box -38 -48 222 592
use scs8hd_decap_3  PHY_40
timestamp 1586364061
transform 1 0 1104 0 -1 13600
box -38 -48 314 592
use scs8hd_decap_3  PHY_38
timestamp 1586364061
transform 1 0 1104 0 1 12512
box -38 -48 314 592
use scs8hd_buf_4  mux_bottom_ipin_1.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 1840 0 1 12512
box -38 -48 590 592
use scs8hd_buf_2  _47_
timestamp 1586364061
transform 1 0 1380 0 -1 13600
box -38 -48 406 592
use scs8hd_fill_2  FILLER_20_15
timestamp 1586364061
transform 1 0 2484 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_14
timestamp 1586364061
transform 1 0 2392 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 2576 0 1 12512
box -38 -48 222 592
use scs8hd_buf_4  mux_bottom_ipin_2.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 2668 0 -1 13600
box -38 -48 590 592
use scs8hd_decap_4  FILLER_19_18
timestamp 1586364061
transform 1 0 2760 0 1 12512
box -38 -48 406 592
use scs8hd_decap_4  FILLER_20_27
timestamp 1586364061
transform 1 0 3588 0 -1 13600
box -38 -48 406 592
use scs8hd_fill_2  FILLER_20_23
timestamp 1586364061
transform 1 0 3220 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_29
timestamp 1586364061
transform 1 0 3772 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_25
timestamp 1586364061
transform 1 0 3404 0 1 12512
box -38 -48 222 592
use scs8hd_fill_1  FILLER_19_22
timestamp 1586364061
transform 1 0 3128 0 1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 3404 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 3220 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__41__A
timestamp 1586364061
transform 1 0 3588 0 1 12512
box -38 -48 222 592
use scs8hd_decap_8  FILLER_20_36
timestamp 1586364061
transform 1 0 4416 0 -1 13600
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 3956 0 1 12512
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_178
timestamp 1586364061
transform 1 0 3956 0 -1 13600
box -38 -48 130 592
use scs8hd_mux2_2  mux_bottom_ipin_1.mux_l2_in_1_
timestamp 1586364061
transform 1 0 4140 0 1 12512
box -38 -48 866 592
use scs8hd_buf_2  _41_
timestamp 1586364061
transform 1 0 4048 0 -1 13600
box -38 -48 406 592
use scs8hd_conb_1  _19_
timestamp 1586364061
transform 1 0 5704 0 1 12512
box -38 -48 314 592
use scs8hd_buf_2  _38_
timestamp 1586364061
transform 1 0 5152 0 -1 13600
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__38__A
timestamp 1586364061
transform 1 0 5152 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l3_in_1__A0
timestamp 1586364061
transform 1 0 5520 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_3.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 6532 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_42
timestamp 1586364061
transform 1 0 4968 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_46
timestamp 1586364061
transform 1 0 5336 0 1 12512
box -38 -48 222 592
use scs8hd_decap_6  FILLER_19_53
timestamp 1586364061
transform 1 0 5980 0 1 12512
box -38 -48 590 592
use scs8hd_decap_12  FILLER_20_48
timestamp 1586364061
transform 1 0 5520 0 -1 13600
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_20_60
timestamp 1586364061
transform 1 0 6624 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_68
timestamp 1586364061
transform 1 0 7360 0 1 12512
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_179
timestamp 1586364061
transform 1 0 6808 0 -1 13600
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_172
timestamp 1586364061
transform 1 0 6716 0 1 12512
box -38 -48 130 592
use scs8hd_buf_4  mux_bottom_ipin_3.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 6808 0 1 12512
box -38 -48 590 592
use scs8hd_buf_2  _35_
timestamp 1586364061
transform 1 0 6900 0 -1 13600
box -38 -48 406 592
use scs8hd_decap_4  FILLER_19_72
timestamp 1586364061
transform 1 0 7728 0 1 12512
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__35__A
timestamp 1586364061
transform 1 0 7544 0 1 12512
box -38 -48 222 592
use scs8hd_buf_2  _32_
timestamp 1586364061
transform 1 0 8096 0 1 12512
box -38 -48 406 592
use scs8hd_decap_12  FILLER_20_79
timestamp 1586364061
transform 1 0 8372 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_67
timestamp 1586364061
transform 1 0 7268 0 -1 13600
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_180
timestamp 1586364061
transform 1 0 9660 0 -1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__32__A
timestamp 1586364061
transform 1 0 8648 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_80
timestamp 1586364061
transform 1 0 8464 0 1 12512
box -38 -48 222 592
use scs8hd_decap_12  FILLER_19_84
timestamp 1586364061
transform 1 0 8832 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_19_96
timestamp 1586364061
transform 1 0 9936 0 1 12512
box -38 -48 406 592
use scs8hd_fill_2  FILLER_20_91
timestamp 1586364061
transform 1 0 9476 0 -1 13600
box -38 -48 222 592
use scs8hd_decap_12  FILLER_20_94
timestamp 1586364061
transform 1 0 9752 0 -1 13600
box -38 -48 1142 592
use scs8hd_buf_4  mux_bottom_ipin_4.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 10304 0 1 12512
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_4.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 11040 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_106
timestamp 1586364061
transform 1 0 10856 0 1 12512
box -38 -48 222 592
use scs8hd_decap_12  FILLER_19_110
timestamp 1586364061
transform 1 0 11224 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_106
timestamp 1586364061
transform 1 0 10856 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_20_118
timestamp 1586364061
transform 1 0 11960 0 -1 13600
box -38 -48 590 592
use scs8hd_buf_4  mux_bottom_ipin_6.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 12972 0 1 12512
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_173
timestamp 1586364061
transform 1 0 12328 0 1 12512
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_181
timestamp 1586364061
transform 1 0 12512 0 -1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_6.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 13708 0 1 12512
box -38 -48 222 592
use scs8hd_decap_6  FILLER_19_123
timestamp 1586364061
transform 1 0 12420 0 1 12512
box -38 -48 590 592
use scs8hd_fill_2  FILLER_19_135
timestamp 1586364061
transform 1 0 13524 0 1 12512
box -38 -48 222 592
use scs8hd_decap_12  FILLER_20_125
timestamp 1586364061
transform 1 0 12604 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_137
timestamp 1586364061
transform 1 0 13708 0 -1 13600
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_182
timestamp 1586364061
transform 1 0 15364 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_12  FILLER_19_139
timestamp 1586364061
transform 1 0 13892 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_151
timestamp 1586364061
transform 1 0 14996 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_20_149
timestamp 1586364061
transform 1 0 14812 0 -1 13600
box -38 -48 590 592
use scs8hd_decap_12  FILLER_20_156
timestamp 1586364061
transform 1 0 15456 0 -1 13600
box -38 -48 1142 592
use scs8hd_buf_4  mux_bottom_ipin_7.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 16192 0 1 12512
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_7.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 16928 0 1 12512
box -38 -48 222 592
use scs8hd_fill_1  FILLER_19_163
timestamp 1586364061
transform 1 0 16100 0 1 12512
box -38 -48 130 592
use scs8hd_fill_2  FILLER_19_170
timestamp 1586364061
transform 1 0 16744 0 1 12512
box -38 -48 222 592
use scs8hd_decap_8  FILLER_19_174
timestamp 1586364061
transform 1 0 17112 0 1 12512
box -38 -48 774 592
use scs8hd_decap_12  FILLER_20_168
timestamp 1586364061
transform 1 0 16560 0 -1 13600
box -38 -48 1142 592
use scs8hd_buf_4  mux_bottom_ipin_8.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 18768 0 1 12512
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_174
timestamp 1586364061
transform 1 0 17940 0 1 12512
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_183
timestamp 1586364061
transform 1 0 18216 0 -1 13600
box -38 -48 130 592
use scs8hd_fill_1  FILLER_19_182
timestamp 1586364061
transform 1 0 17848 0 1 12512
box -38 -48 130 592
use scs8hd_decap_8  FILLER_19_184
timestamp 1586364061
transform 1 0 18032 0 1 12512
box -38 -48 774 592
use scs8hd_fill_2  FILLER_19_198
timestamp 1586364061
transform 1 0 19320 0 1 12512
box -38 -48 222 592
use scs8hd_decap_6  FILLER_20_180
timestamp 1586364061
transform 1 0 17664 0 -1 13600
box -38 -48 590 592
use scs8hd_decap_12  FILLER_20_187
timestamp 1586364061
transform 1 0 18308 0 -1 13600
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_184
timestamp 1586364061
transform 1 0 21068 0 -1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_8.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 19504 0 1 12512
box -38 -48 222 592
use scs8hd_decap_12  FILLER_19_202
timestamp 1586364061
transform 1 0 19688 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_19_214
timestamp 1586364061
transform 1 0 20792 0 1 12512
box -38 -48 774 592
use scs8hd_decap_12  FILLER_20_199
timestamp 1586364061
transform 1 0 19412 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_20_211
timestamp 1586364061
transform 1 0 20516 0 -1 13600
box -38 -48 590 592
use scs8hd_decap_12  FILLER_20_218
timestamp 1586364061
transform 1 0 21160 0 -1 13600
box -38 -48 1142 592
use scs8hd_buf_4  mux_bottom_ipin_9.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 21804 0 1 12512
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_9.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 22540 0 1 12512
box -38 -48 222 592
use scs8hd_decap_3  FILLER_19_222
timestamp 1586364061
transform 1 0 21528 0 1 12512
box -38 -48 314 592
use scs8hd_fill_2  FILLER_19_231
timestamp 1586364061
transform 1 0 22356 0 1 12512
box -38 -48 222 592
use scs8hd_decap_6  FILLER_19_235
timestamp 1586364061
transform 1 0 22724 0 1 12512
box -38 -48 590 592
use scs8hd_decap_12  FILLER_20_230
timestamp 1586364061
transform 1 0 22264 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_20_242
timestamp 1586364061
transform 1 0 23368 0 -1 13600
box -38 -48 590 592
use scs8hd_decap_3  FILLER_19_245
timestamp 1586364061
transform 1 0 23644 0 1 12512
box -38 -48 314 592
use scs8hd_fill_1  FILLER_19_241
timestamp 1586364061
transform 1 0 23276 0 1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_11.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 23368 0 1 12512
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_175
timestamp 1586364061
transform 1 0 23552 0 1 12512
box -38 -48 130 592
use scs8hd_fill_2  FILLER_20_255
timestamp 1586364061
transform 1 0 24564 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_250
timestamp 1586364061
transform 1 0 24104 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_9.mux_l1_in_2__S
timestamp 1586364061
transform 1 0 24748 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_9.mux_l1_in_2__A0
timestamp 1586364061
transform 1 0 23920 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_9.mux_l1_in_2__A1
timestamp 1586364061
transform 1 0 24288 0 1 12512
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_185
timestamp 1586364061
transform 1 0 23920 0 -1 13600
box -38 -48 130 592
use scs8hd_mux2_2  mux_bottom_ipin_9.mux_l1_in_2_
timestamp 1586364061
transform 1 0 24472 0 1 12512
box -38 -48 866 592
use scs8hd_buf_4  mux_bottom_ipin_11.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 24012 0 -1 13600
box -38 -48 590 592
use scs8hd_decap_12  FILLER_19_263
timestamp 1586364061
transform 1 0 25300 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_19_275
timestamp 1586364061
transform 1 0 26404 0 1 12512
box -38 -48 774 592
use scs8hd_decap_12  FILLER_20_259
timestamp 1586364061
transform 1 0 24932 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_20_271
timestamp 1586364061
transform 1 0 26036 0 -1 13600
box -38 -48 774 592
use scs8hd_buf_4  mux_bottom_ipin_12.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 27324 0 1 12512
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_186
timestamp 1586364061
transform 1 0 26772 0 -1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_12.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 28060 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_283
timestamp 1586364061
transform 1 0 27140 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_291
timestamp 1586364061
transform 1 0 27876 0 1 12512
box -38 -48 222 592
use scs8hd_decap_8  FILLER_19_295
timestamp 1586364061
transform 1 0 28244 0 1 12512
box -38 -48 774 592
use scs8hd_decap_12  FILLER_20_280
timestamp 1586364061
transform 1 0 26864 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_292
timestamp 1586364061
transform 1 0 27968 0 -1 13600
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_176
timestamp 1586364061
transform 1 0 29164 0 1 12512
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_187
timestamp 1586364061
transform 1 0 29624 0 -1 13600
box -38 -48 130 592
use scs8hd_fill_2  FILLER_19_303
timestamp 1586364061
transform 1 0 28980 0 1 12512
box -38 -48 222 592
use scs8hd_decap_12  FILLER_19_306
timestamp 1586364061
transform 1 0 29256 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_20_304
timestamp 1586364061
transform 1 0 29072 0 -1 13600
box -38 -48 590 592
use scs8hd_decap_12  FILLER_20_311
timestamp 1586364061
transform 1 0 29716 0 -1 13600
box -38 -48 1142 592
use scs8hd_buf_2  _55_
timestamp 1586364061
transform 1 0 32108 0 1 12512
box -38 -48 406 592
use scs8hd_buf_4  mux_bottom_ipin_13.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 30820 0 1 12512
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_13.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 31556 0 1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_19_318
timestamp 1586364061
transform 1 0 30360 0 1 12512
box -38 -48 406 592
use scs8hd_fill_1  FILLER_19_322
timestamp 1586364061
transform 1 0 30728 0 1 12512
box -38 -48 130 592
use scs8hd_fill_2  FILLER_19_329
timestamp 1586364061
transform 1 0 31372 0 1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_19_333
timestamp 1586364061
transform 1 0 31740 0 1 12512
box -38 -48 406 592
use scs8hd_decap_12  FILLER_20_323
timestamp 1586364061
transform 1 0 30820 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_20_335
timestamp 1586364061
transform 1 0 31924 0 -1 13600
box -38 -48 590 592
use scs8hd_decap_6  FILLER_20_342
timestamp 1586364061
transform 1 0 32568 0 -1 13600
box -38 -48 590 592
use scs8hd_fill_2  FILLER_19_345
timestamp 1586364061
transform 1 0 32844 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_341
timestamp 1586364061
transform 1 0 32476 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__55__A
timestamp 1586364061
transform 1 0 32660 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_15.mux_l4_in_0__S
timestamp 1586364061
transform 1 0 33028 0 1 12512
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_188
timestamp 1586364061
transform 1 0 32476 0 -1 13600
box -38 -48 130 592
use scs8hd_fill_2  FILLER_20_356
timestamp 1586364061
transform 1 0 33856 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_352
timestamp 1586364061
transform 1 0 33488 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__54__A
timestamp 1586364061
transform 1 0 33672 0 -1 13600
box -38 -48 222 592
use scs8hd_mux2_2  mux_bottom_ipin_15.mux_l4_in_0_
timestamp 1586364061
transform 1 0 33212 0 1 12512
box -38 -48 866 592
use scs8hd_buf_2  _54_
timestamp 1586364061
transform 1 0 33120 0 -1 13600
box -38 -48 406 592
use scs8hd_fill_2  FILLER_19_362
timestamp 1586364061
transform 1 0 34408 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_358
timestamp 1586364061
transform 1 0 34040 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_15.mux_l4_in_0__A1
timestamp 1586364061
transform 1 0 34040 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__52__A
timestamp 1586364061
transform 1 0 34224 0 1 12512
box -38 -48 222 592
use scs8hd_buf_2  _52_
timestamp 1586364061
transform 1 0 34224 0 -1 13600
box -38 -48 406 592
use scs8hd_decap_3  FILLER_20_369
timestamp 1586364061
transform 1 0 35052 0 -1 13600
box -38 -48 314 592
use scs8hd_decap_3  FILLER_20_364
timestamp 1586364061
transform 1 0 34592 0 -1 13600
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_15.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 34868 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_15.mux_l4_in_0__A0
timestamp 1586364061
transform 1 0 34592 0 1 12512
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_177
timestamp 1586364061
transform 1 0 34776 0 1 12512
box -38 -48 130 592
use scs8hd_buf_4  mux_bottom_ipin_15.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 34868 0 1 12512
box -38 -48 590 592
use scs8hd_fill_2  FILLER_19_373
timestamp 1586364061
transform 1 0 35420 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__65__A
timestamp 1586364061
transform 1 0 35604 0 1 12512
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_189
timestamp 1586364061
transform 1 0 35328 0 -1 13600
box -38 -48 130 592
use scs8hd_buf_2  _65_
timestamp 1586364061
transform 1 0 35420 0 -1 13600
box -38 -48 406 592
use scs8hd_decap_8  FILLER_20_377
timestamp 1586364061
transform 1 0 35788 0 -1 13600
box -38 -48 774 592
use scs8hd_fill_2  FILLER_19_385
timestamp 1586364061
transform 1 0 36524 0 1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_19_377
timestamp 1586364061
transform 1 0 35788 0 1 12512
box -38 -48 406 592
use scs8hd_buf_2  _63_
timestamp 1586364061
transform 1 0 36524 0 -1 13600
box -38 -48 406 592
use scs8hd_buf_2  _53_
timestamp 1586364061
transform 1 0 36156 0 1 12512
box -38 -48 406 592
use scs8hd_fill_2  FILLER_19_389
timestamp 1586364061
transform 1 0 36892 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__63__A
timestamp 1586364061
transform 1 0 37076 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__53__A
timestamp 1586364061
transform 1 0 36708 0 1 12512
box -38 -48 222 592
use scs8hd_buf_2  _61_
timestamp 1586364061
transform 1 0 37260 0 1 12512
box -38 -48 406 592
use scs8hd_decap_12  FILLER_20_389
timestamp 1586364061
transform 1 0 36892 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_3  PHY_39
timestamp 1586364061
transform -1 0 38824 0 1 12512
box -38 -48 314 592
use scs8hd_decap_3  PHY_41
timestamp 1586364061
transform -1 0 38824 0 -1 13600
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_190
timestamp 1586364061
transform 1 0 38180 0 -1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__61__A
timestamp 1586364061
transform 1 0 37812 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_397
timestamp 1586364061
transform 1 0 37628 0 1 12512
box -38 -48 222 592
use scs8hd_decap_6  FILLER_19_401
timestamp 1586364061
transform 1 0 37996 0 1 12512
box -38 -48 590 592
use scs8hd_fill_2  FILLER_20_401
timestamp 1586364061
transform 1 0 37996 0 -1 13600
box -38 -48 222 592
use scs8hd_decap_3  FILLER_20_404
timestamp 1586364061
transform 1 0 38272 0 -1 13600
box -38 -48 314 592
<< labels >>
rlabel metal3 s 39520 15784 40000 15904 6 ccff_head
port 0 nsew default input
rlabel metal2 s 38750 15520 38806 16000 6 ccff_tail
port 1 nsew default tristate
rlabel metal3 s 0 144 480 264 6 chanx_left_in[0]
port 2 nsew default input
rlabel metal3 s 0 4088 480 4208 6 chanx_left_in[10]
port 3 nsew default input
rlabel metal3 s 0 4496 480 4616 6 chanx_left_in[11]
port 4 nsew default input
rlabel metal3 s 0 4904 480 5024 6 chanx_left_in[12]
port 5 nsew default input
rlabel metal3 s 0 5312 480 5432 6 chanx_left_in[13]
port 6 nsew default input
rlabel metal3 s 0 5720 480 5840 6 chanx_left_in[14]
port 7 nsew default input
rlabel metal3 s 0 6128 480 6248 6 chanx_left_in[15]
port 8 nsew default input
rlabel metal3 s 0 6536 480 6656 6 chanx_left_in[16]
port 9 nsew default input
rlabel metal3 s 0 6944 480 7064 6 chanx_left_in[17]
port 10 nsew default input
rlabel metal3 s 0 7352 480 7472 6 chanx_left_in[18]
port 11 nsew default input
rlabel metal3 s 0 7760 480 7880 6 chanx_left_in[19]
port 12 nsew default input
rlabel metal3 s 0 416 480 536 6 chanx_left_in[1]
port 13 nsew default input
rlabel metal3 s 0 824 480 944 6 chanx_left_in[2]
port 14 nsew default input
rlabel metal3 s 0 1232 480 1352 6 chanx_left_in[3]
port 15 nsew default input
rlabel metal3 s 0 1640 480 1760 6 chanx_left_in[4]
port 16 nsew default input
rlabel metal3 s 0 2048 480 2168 6 chanx_left_in[5]
port 17 nsew default input
rlabel metal3 s 0 2456 480 2576 6 chanx_left_in[6]
port 18 nsew default input
rlabel metal3 s 0 2864 480 2984 6 chanx_left_in[7]
port 19 nsew default input
rlabel metal3 s 0 3272 480 3392 6 chanx_left_in[8]
port 20 nsew default input
rlabel metal3 s 0 3680 480 3800 6 chanx_left_in[9]
port 21 nsew default input
rlabel metal3 s 0 8168 480 8288 6 chanx_left_out[0]
port 22 nsew default tristate
rlabel metal3 s 0 12112 480 12232 6 chanx_left_out[10]
port 23 nsew default tristate
rlabel metal3 s 0 12520 480 12640 6 chanx_left_out[11]
port 24 nsew default tristate
rlabel metal3 s 0 12928 480 13048 6 chanx_left_out[12]
port 25 nsew default tristate
rlabel metal3 s 0 13336 480 13456 6 chanx_left_out[13]
port 26 nsew default tristate
rlabel metal3 s 0 13744 480 13864 6 chanx_left_out[14]
port 27 nsew default tristate
rlabel metal3 s 0 14152 480 14272 6 chanx_left_out[15]
port 28 nsew default tristate
rlabel metal3 s 0 14560 480 14680 6 chanx_left_out[16]
port 29 nsew default tristate
rlabel metal3 s 0 14968 480 15088 6 chanx_left_out[17]
port 30 nsew default tristate
rlabel metal3 s 0 15376 480 15496 6 chanx_left_out[18]
port 31 nsew default tristate
rlabel metal3 s 0 15784 480 15904 6 chanx_left_out[19]
port 32 nsew default tristate
rlabel metal3 s 0 8440 480 8560 6 chanx_left_out[1]
port 33 nsew default tristate
rlabel metal3 s 0 8848 480 8968 6 chanx_left_out[2]
port 34 nsew default tristate
rlabel metal3 s 0 9256 480 9376 6 chanx_left_out[3]
port 35 nsew default tristate
rlabel metal3 s 0 9664 480 9784 6 chanx_left_out[4]
port 36 nsew default tristate
rlabel metal3 s 0 10072 480 10192 6 chanx_left_out[5]
port 37 nsew default tristate
rlabel metal3 s 0 10480 480 10600 6 chanx_left_out[6]
port 38 nsew default tristate
rlabel metal3 s 0 10888 480 11008 6 chanx_left_out[7]
port 39 nsew default tristate
rlabel metal3 s 0 11296 480 11416 6 chanx_left_out[8]
port 40 nsew default tristate
rlabel metal3 s 0 11704 480 11824 6 chanx_left_out[9]
port 41 nsew default tristate
rlabel metal3 s 39520 144 40000 264 6 chanx_right_in[0]
port 42 nsew default input
rlabel metal3 s 39520 3952 40000 4072 6 chanx_right_in[10]
port 43 nsew default input
rlabel metal3 s 39520 4360 40000 4480 6 chanx_right_in[11]
port 44 nsew default input
rlabel metal3 s 39520 4768 40000 4888 6 chanx_right_in[12]
port 45 nsew default input
rlabel metal3 s 39520 5176 40000 5296 6 chanx_right_in[13]
port 46 nsew default input
rlabel metal3 s 39520 5584 40000 5704 6 chanx_right_in[14]
port 47 nsew default input
rlabel metal3 s 39520 5992 40000 6112 6 chanx_right_in[15]
port 48 nsew default input
rlabel metal3 s 39520 6400 40000 6520 6 chanx_right_in[16]
port 49 nsew default input
rlabel metal3 s 39520 6672 40000 6792 6 chanx_right_in[17]
port 50 nsew default input
rlabel metal3 s 39520 7080 40000 7200 6 chanx_right_in[18]
port 51 nsew default input
rlabel metal3 s 39520 7488 40000 7608 6 chanx_right_in[19]
port 52 nsew default input
rlabel metal3 s 39520 416 40000 536 6 chanx_right_in[1]
port 53 nsew default input
rlabel metal3 s 39520 824 40000 944 6 chanx_right_in[2]
port 54 nsew default input
rlabel metal3 s 39520 1232 40000 1352 6 chanx_right_in[3]
port 55 nsew default input
rlabel metal3 s 39520 1640 40000 1760 6 chanx_right_in[4]
port 56 nsew default input
rlabel metal3 s 39520 2048 40000 2168 6 chanx_right_in[5]
port 57 nsew default input
rlabel metal3 s 39520 2456 40000 2576 6 chanx_right_in[6]
port 58 nsew default input
rlabel metal3 s 39520 2864 40000 2984 6 chanx_right_in[7]
port 59 nsew default input
rlabel metal3 s 39520 3272 40000 3392 6 chanx_right_in[8]
port 60 nsew default input
rlabel metal3 s 39520 3544 40000 3664 6 chanx_right_in[9]
port 61 nsew default input
rlabel metal3 s 39520 7896 40000 8016 6 chanx_right_out[0]
port 62 nsew default tristate
rlabel metal3 s 39520 11840 40000 11960 6 chanx_right_out[10]
port 63 nsew default tristate
rlabel metal3 s 39520 12248 40000 12368 6 chanx_right_out[11]
port 64 nsew default tristate
rlabel metal3 s 39520 12656 40000 12776 6 chanx_right_out[12]
port 65 nsew default tristate
rlabel metal3 s 39520 12928 40000 13048 6 chanx_right_out[13]
port 66 nsew default tristate
rlabel metal3 s 39520 13336 40000 13456 6 chanx_right_out[14]
port 67 nsew default tristate
rlabel metal3 s 39520 13744 40000 13864 6 chanx_right_out[15]
port 68 nsew default tristate
rlabel metal3 s 39520 14152 40000 14272 6 chanx_right_out[16]
port 69 nsew default tristate
rlabel metal3 s 39520 14560 40000 14680 6 chanx_right_out[17]
port 70 nsew default tristate
rlabel metal3 s 39520 14968 40000 15088 6 chanx_right_out[18]
port 71 nsew default tristate
rlabel metal3 s 39520 15376 40000 15496 6 chanx_right_out[19]
port 72 nsew default tristate
rlabel metal3 s 39520 8304 40000 8424 6 chanx_right_out[1]
port 73 nsew default tristate
rlabel metal3 s 39520 8712 40000 8832 6 chanx_right_out[2]
port 74 nsew default tristate
rlabel metal3 s 39520 9120 40000 9240 6 chanx_right_out[3]
port 75 nsew default tristate
rlabel metal3 s 39520 9528 40000 9648 6 chanx_right_out[4]
port 76 nsew default tristate
rlabel metal3 s 39520 9800 40000 9920 6 chanx_right_out[5]
port 77 nsew default tristate
rlabel metal3 s 39520 10208 40000 10328 6 chanx_right_out[6]
port 78 nsew default tristate
rlabel metal3 s 39520 10616 40000 10736 6 chanx_right_out[7]
port 79 nsew default tristate
rlabel metal3 s 39520 11024 40000 11144 6 chanx_right_out[8]
port 80 nsew default tristate
rlabel metal3 s 39520 11432 40000 11552 6 chanx_right_out[9]
port 81 nsew default tristate
rlabel metal2 s 19982 0 20038 480 6 prog_clk
port 82 nsew default input
rlabel metal2 s 1122 15520 1178 16000 6 top_grid_pin_16_
port 83 nsew default tristate
rlabel metal2 s 3422 15520 3478 16000 6 top_grid_pin_17_
port 84 nsew default tristate
rlabel metal2 s 5814 15520 5870 16000 6 top_grid_pin_18_
port 85 nsew default tristate
rlabel metal2 s 8114 15520 8170 16000 6 top_grid_pin_19_
port 86 nsew default tristate
rlabel metal2 s 10506 15520 10562 16000 6 top_grid_pin_20_
port 87 nsew default tristate
rlabel metal2 s 12806 15520 12862 16000 6 top_grid_pin_21_
port 88 nsew default tristate
rlabel metal2 s 15198 15520 15254 16000 6 top_grid_pin_22_
port 89 nsew default tristate
rlabel metal2 s 17590 15520 17646 16000 6 top_grid_pin_23_
port 90 nsew default tristate
rlabel metal2 s 19890 15520 19946 16000 6 top_grid_pin_24_
port 91 nsew default tristate
rlabel metal2 s 22282 15520 22338 16000 6 top_grid_pin_25_
port 92 nsew default tristate
rlabel metal2 s 24582 15520 24638 16000 6 top_grid_pin_26_
port 93 nsew default tristate
rlabel metal2 s 26974 15520 27030 16000 6 top_grid_pin_27_
port 94 nsew default tristate
rlabel metal2 s 29366 15520 29422 16000 6 top_grid_pin_28_
port 95 nsew default tristate
rlabel metal2 s 31666 15520 31722 16000 6 top_grid_pin_29_
port 96 nsew default tristate
rlabel metal2 s 34058 15520 34114 16000 6 top_grid_pin_30_
port 97 nsew default tristate
rlabel metal2 s 36358 15520 36414 16000 6 top_grid_pin_31_
port 98 nsew default tristate
rlabel metal4 s 7611 2128 7931 13648 6 vpwr
port 99 nsew default input
rlabel metal4 s 14277 2128 14597 13648 6 vgnd
port 100 nsew default input
<< properties >>
string FIXED_BBOX 0 0 40000 16000
<< end >>
