magic
tech EFS8A
magscale 1 2
timestamp 1602539824
<< locali >>
rect 220455 2839 220489 2907
rect 220455 2805 220461 2839
<< viali >>
rect 178233 7497 178267 7531
rect 92765 7293 92799 7327
rect 93317 7293 93351 7327
rect 178049 7293 178083 7327
rect 229385 7293 229419 7327
rect 229937 7293 229971 7327
rect 92949 7157 92983 7191
rect 178693 7157 178727 7191
rect 229569 7157 229603 7191
rect 170781 6953 170815 6987
rect 170597 6817 170631 6851
rect 88257 6749 88291 6783
rect 88441 6749 88475 6783
rect 225337 6749 225371 6783
rect 225521 6749 225555 6783
rect 88625 6613 88659 6647
rect 215677 6613 215711 6647
rect 225705 6613 225739 6647
rect 88257 6409 88291 6443
rect 225337 6409 225371 6443
rect 215953 6341 215987 6375
rect 215493 6273 215527 6307
rect 215585 6273 215619 6307
rect 215769 6273 215803 6307
rect 88717 6069 88751 6103
rect 170689 6069 170723 6103
rect 225889 6069 225923 6103
rect 215401 5729 215435 5763
rect 217333 5729 217367 5763
rect 215125 5661 215159 5695
rect 217517 5661 217551 5695
rect 216781 5525 216815 5559
rect 217701 5525 217735 5559
rect 215953 5321 215987 5355
rect 217885 5321 217919 5355
rect 221473 5321 221507 5355
rect 223957 5321 223991 5355
rect 209237 5253 209271 5287
rect 213193 5253 213227 5287
rect 216689 5253 216723 5287
rect 224417 5253 224451 5287
rect 216781 5185 216815 5219
rect 224049 5185 224083 5219
rect 93133 5117 93167 5151
rect 208869 5117 208903 5151
rect 209053 5117 209087 5151
rect 212273 5117 212307 5151
rect 214297 5117 214331 5151
rect 215033 5117 215067 5151
rect 217057 5117 217091 5151
rect 217517 5117 217551 5151
rect 220553 5117 220587 5151
rect 224233 5117 224267 5151
rect 212181 5049 212215 5083
rect 212635 5049 212669 5083
rect 214941 5049 214975 5083
rect 215354 5049 215388 5083
rect 216965 5049 216999 5083
rect 217149 5049 217183 5083
rect 220874 5049 220908 5083
rect 93317 4981 93351 5015
rect 93777 4981 93811 5015
rect 208593 4981 208627 5015
rect 216321 4981 216355 5015
rect 218161 4981 218195 5015
rect 220369 4981 220403 5015
rect 208961 4777 208995 4811
rect 214849 4777 214883 4811
rect 216229 4777 216263 4811
rect 220553 4777 220587 4811
rect 224141 4777 224175 4811
rect 215630 4709 215664 4743
rect 218339 4709 218373 4743
rect 213837 4641 213871 4675
rect 214481 4641 214515 4675
rect 215309 4573 215343 4607
rect 217977 4573 218011 4607
rect 212365 4437 212399 4471
rect 212825 4437 212859 4471
rect 215217 4437 215251 4471
rect 216873 4437 216907 4471
rect 218897 4437 218931 4471
rect 214297 4233 214331 4267
rect 215125 4233 215159 4267
rect 218069 4233 218103 4267
rect 212365 4029 212399 4063
rect 213101 4029 213135 4063
rect 215769 4029 215803 4063
rect 216045 4029 216079 4063
rect 216413 4029 216447 4063
rect 216965 4029 216999 4063
rect 212825 3961 212859 3995
rect 213193 3961 213227 3995
rect 213561 3961 213595 3995
rect 215401 3961 215435 3995
rect 217057 3961 217091 3995
rect 218345 3961 218379 3995
rect 212641 3893 212675 3927
rect 213009 3893 213043 3927
rect 213837 3893 213871 3927
rect 214757 3893 214791 3927
rect 217425 3893 217459 3927
rect 213377 3689 213411 3723
rect 216597 3689 216631 3723
rect 216965 3689 216999 3723
rect 220645 3689 220679 3723
rect 212549 3621 212583 3655
rect 215033 3621 215067 3655
rect 215585 3621 215619 3655
rect 215953 3621 215987 3655
rect 216321 3621 216355 3655
rect 220087 3621 220121 3655
rect 213285 3553 213319 3587
rect 213745 3553 213779 3587
rect 214113 3553 214147 3587
rect 214481 3553 214515 3587
rect 215769 3553 215803 3587
rect 215861 3553 215895 3587
rect 217517 3553 217551 3587
rect 219725 3485 219759 3519
rect 212917 3417 212951 3451
rect 215493 3417 215527 3451
rect 217793 3349 217827 3383
rect 211997 3145 212031 3179
rect 212273 3145 212307 3179
rect 214021 3145 214055 3179
rect 214665 3145 214699 3179
rect 215585 3145 215619 3179
rect 217517 3145 217551 3179
rect 213377 3077 213411 3111
rect 215217 3077 215251 3111
rect 211629 3009 211663 3043
rect 212457 3009 212491 3043
rect 214481 2941 214515 2975
rect 216045 2941 216079 2975
rect 216229 2941 216263 2975
rect 216597 2941 216631 2975
rect 216965 2941 216999 2975
rect 217241 2941 217275 2975
rect 220093 2941 220127 2975
rect 212778 2873 212812 2907
rect 217885 2873 217919 2907
rect 213653 2805 213687 2839
rect 218253 2805 218287 2839
rect 219541 2805 219575 2839
rect 219909 2805 219943 2839
rect 220461 2805 220495 2839
rect 221013 2805 221047 2839
rect 211629 2601 211663 2635
rect 212089 2601 212123 2635
rect 213009 2601 213043 2635
rect 213745 2601 213779 2635
rect 214573 2601 214607 2635
rect 214849 2601 214883 2635
rect 217333 2601 217367 2635
rect 217793 2601 217827 2635
rect 219725 2601 219759 2635
rect 220093 2601 220127 2635
rect 220553 2601 220587 2635
rect 221933 2601 221967 2635
rect 213653 2533 213687 2567
rect 213837 2533 213871 2567
rect 214205 2533 214239 2567
rect 216689 2533 216723 2567
rect 212273 2465 212307 2499
rect 213285 2465 213319 2499
rect 213469 2465 213503 2499
rect 215493 2465 215527 2499
rect 215677 2465 215711 2499
rect 216229 2465 216263 2499
rect 216413 2465 216447 2499
rect 216965 2465 216999 2499
rect 221473 2465 221507 2499
rect 228189 2465 228223 2499
rect 228741 2465 228775 2499
rect 309425 2465 309459 2499
rect 350825 2465 350859 2499
rect 351377 2465 351411 2499
rect 211353 2397 211387 2431
rect 221289 2397 221323 2431
rect 308597 2397 308631 2431
rect 309241 2397 309275 2431
rect 309057 2329 309091 2363
rect 309885 2329 309919 2363
rect 212457 2261 212491 2295
rect 221197 2261 221231 2295
rect 228373 2261 228407 2295
rect 351009 2261 351043 2295
<< metal1 >>
rect 106 8168 112 8220
rect 164 8208 170 8220
rect 178218 8208 178224 8220
rect 164 8180 178224 8208
rect 164 8168 170 8180
rect 178218 8168 178224 8180
rect 178276 8168 178282 8220
rect 1104 7642 422832 7664
rect 1104 7590 71648 7642
rect 71700 7590 71712 7642
rect 71764 7590 71776 7642
rect 71828 7590 71840 7642
rect 71892 7590 212982 7642
rect 213034 7590 213046 7642
rect 213098 7590 213110 7642
rect 213162 7590 213174 7642
rect 213226 7590 354315 7642
rect 354367 7590 354379 7642
rect 354431 7590 354443 7642
rect 354495 7590 354507 7642
rect 354559 7590 422832 7642
rect 1104 7568 422832 7590
rect 178218 7528 178224 7540
rect 178179 7500 178224 7528
rect 178218 7488 178224 7500
rect 178276 7488 178282 7540
rect 88610 7284 88616 7336
rect 88668 7324 88674 7336
rect 92753 7327 92811 7333
rect 92753 7324 92765 7327
rect 88668 7296 92765 7324
rect 88668 7284 88674 7296
rect 92753 7293 92765 7296
rect 92799 7324 92811 7327
rect 93305 7327 93363 7333
rect 93305 7324 93317 7327
rect 92799 7296 93317 7324
rect 92799 7293 92811 7296
rect 92753 7287 92811 7293
rect 93305 7293 93317 7296
rect 93351 7293 93363 7327
rect 93305 7287 93363 7293
rect 178037 7327 178095 7333
rect 178037 7293 178049 7327
rect 178083 7324 178095 7327
rect 178083 7296 178724 7324
rect 178083 7293 178095 7296
rect 178037 7287 178095 7293
rect 106090 7256 106096 7268
rect 93136 7228 106096 7256
rect 92937 7191 92995 7197
rect 92937 7157 92949 7191
rect 92983 7188 92995 7191
rect 93136 7188 93164 7228
rect 106090 7216 106096 7228
rect 106148 7216 106154 7268
rect 178696 7197 178724 7296
rect 225690 7284 225696 7336
rect 225748 7324 225754 7336
rect 229373 7327 229431 7333
rect 229373 7324 229385 7327
rect 225748 7296 229385 7324
rect 225748 7284 225754 7296
rect 229373 7293 229385 7296
rect 229419 7324 229431 7327
rect 229925 7327 229983 7333
rect 229925 7324 229937 7327
rect 229419 7296 229937 7324
rect 229419 7293 229431 7296
rect 229373 7287 229431 7293
rect 229925 7293 229937 7296
rect 229971 7293 229983 7327
rect 229925 7287 229983 7293
rect 92983 7160 93164 7188
rect 178681 7191 178739 7197
rect 92983 7157 92995 7160
rect 92937 7151 92995 7157
rect 178681 7157 178693 7191
rect 178727 7188 178739 7191
rect 190638 7188 190644 7200
rect 178727 7160 190644 7188
rect 178727 7157 178739 7160
rect 178681 7151 178739 7157
rect 190638 7148 190644 7160
rect 190696 7148 190702 7200
rect 229554 7188 229560 7200
rect 229515 7160 229560 7188
rect 229554 7148 229560 7160
rect 229612 7148 229618 7200
rect 1104 7098 422832 7120
rect 1104 7046 142315 7098
rect 142367 7046 142379 7098
rect 142431 7046 142443 7098
rect 142495 7046 142507 7098
rect 142559 7046 283648 7098
rect 283700 7046 283712 7098
rect 283764 7046 283776 7098
rect 283828 7046 283840 7098
rect 283892 7046 422832 7098
rect 1104 7024 422832 7046
rect 170769 6987 170827 6993
rect 170769 6953 170781 6987
rect 170815 6984 170827 6987
rect 176286 6984 176292 6996
rect 170815 6956 176292 6984
rect 170815 6953 170827 6956
rect 170769 6947 170827 6953
rect 176286 6944 176292 6956
rect 176344 6944 176350 6996
rect 170585 6851 170643 6857
rect 170585 6817 170597 6851
rect 170631 6848 170643 6851
rect 170674 6848 170680 6860
rect 170631 6820 170680 6848
rect 170631 6817 170643 6820
rect 170585 6811 170643 6817
rect 170674 6808 170680 6820
rect 170732 6808 170738 6860
rect 74994 6740 75000 6792
rect 75052 6780 75058 6792
rect 88242 6780 88248 6792
rect 75052 6752 88248 6780
rect 75052 6740 75058 6752
rect 88242 6740 88248 6752
rect 88300 6740 88306 6792
rect 88429 6783 88487 6789
rect 88429 6749 88441 6783
rect 88475 6780 88487 6783
rect 88702 6780 88708 6792
rect 88475 6752 88708 6780
rect 88475 6749 88487 6752
rect 88429 6743 88487 6749
rect 88702 6740 88708 6752
rect 88760 6740 88766 6792
rect 225322 6780 225328 6792
rect 225283 6752 225328 6780
rect 225322 6740 225328 6752
rect 225380 6740 225386 6792
rect 225506 6780 225512 6792
rect 225467 6752 225512 6780
rect 225506 6740 225512 6752
rect 225564 6740 225570 6792
rect 88610 6644 88616 6656
rect 88571 6616 88616 6644
rect 88610 6604 88616 6616
rect 88668 6604 88674 6656
rect 215662 6644 215668 6656
rect 215623 6616 215668 6644
rect 215662 6604 215668 6616
rect 215720 6604 215726 6656
rect 225690 6644 225696 6656
rect 225651 6616 225696 6644
rect 225690 6604 225696 6616
rect 225748 6604 225754 6656
rect 1104 6554 422832 6576
rect 1104 6502 71648 6554
rect 71700 6502 71712 6554
rect 71764 6502 71776 6554
rect 71828 6502 71840 6554
rect 71892 6502 212982 6554
rect 213034 6502 213046 6554
rect 213098 6502 213110 6554
rect 213162 6502 213174 6554
rect 213226 6502 354315 6554
rect 354367 6502 354379 6554
rect 354431 6502 354443 6554
rect 354495 6502 354507 6554
rect 354559 6502 422832 6554
rect 1104 6480 422832 6502
rect 88242 6440 88248 6452
rect 88203 6412 88248 6440
rect 88242 6400 88248 6412
rect 88300 6400 88306 6452
rect 225322 6440 225328 6452
rect 225283 6412 225328 6440
rect 225322 6400 225328 6412
rect 225380 6400 225386 6452
rect 215938 6372 215944 6384
rect 215899 6344 215944 6372
rect 215938 6332 215944 6344
rect 215996 6332 216002 6384
rect 215481 6307 215539 6313
rect 215481 6273 215493 6307
rect 215527 6304 215539 6307
rect 215570 6304 215576 6316
rect 215527 6276 215576 6304
rect 215527 6273 215539 6276
rect 215481 6267 215539 6273
rect 215570 6264 215576 6276
rect 215628 6264 215634 6316
rect 215662 6264 215668 6316
rect 215720 6304 215726 6316
rect 215757 6307 215815 6313
rect 215757 6304 215769 6307
rect 215720 6276 215769 6304
rect 215720 6264 215726 6276
rect 215757 6273 215769 6276
rect 215803 6273 215815 6307
rect 215757 6267 215815 6273
rect 88702 6100 88708 6112
rect 88663 6072 88708 6100
rect 88702 6060 88708 6072
rect 88760 6060 88766 6112
rect 170674 6100 170680 6112
rect 170635 6072 170680 6100
rect 170674 6060 170680 6072
rect 170732 6060 170738 6112
rect 221458 6060 221464 6112
rect 221516 6100 221522 6112
rect 225506 6100 225512 6112
rect 221516 6072 225512 6100
rect 221516 6060 221522 6072
rect 225506 6060 225512 6072
rect 225564 6100 225570 6112
rect 225877 6103 225935 6109
rect 225877 6100 225889 6103
rect 225564 6072 225889 6100
rect 225564 6060 225570 6072
rect 225877 6069 225889 6072
rect 225923 6069 225935 6103
rect 225877 6063 225935 6069
rect 1104 6010 422832 6032
rect 1104 5958 142315 6010
rect 142367 5958 142379 6010
rect 142431 5958 142443 6010
rect 142495 5958 142507 6010
rect 142559 5958 283648 6010
rect 283700 5958 283712 6010
rect 283764 5958 283776 6010
rect 283828 5958 283840 6010
rect 283892 5958 422832 6010
rect 1104 5936 422832 5958
rect 215386 5760 215392 5772
rect 215347 5732 215392 5760
rect 215386 5720 215392 5732
rect 215444 5720 215450 5772
rect 217321 5763 217379 5769
rect 217321 5729 217333 5763
rect 217367 5760 217379 5763
rect 217870 5760 217876 5772
rect 217367 5732 217876 5760
rect 217367 5729 217379 5732
rect 217321 5723 217379 5729
rect 217870 5720 217876 5732
rect 217928 5720 217934 5772
rect 215110 5692 215116 5704
rect 215071 5664 215116 5692
rect 215110 5652 215116 5664
rect 215168 5652 215174 5704
rect 217502 5692 217508 5704
rect 217463 5664 217508 5692
rect 217502 5652 217508 5664
rect 217560 5652 217566 5704
rect 216766 5556 216772 5568
rect 216727 5528 216772 5556
rect 216766 5516 216772 5528
rect 216824 5516 216830 5568
rect 217686 5556 217692 5568
rect 217647 5528 217692 5556
rect 217686 5516 217692 5528
rect 217744 5516 217750 5568
rect 223942 5516 223948 5568
rect 224000 5556 224006 5568
rect 423582 5556 423588 5568
rect 224000 5528 423588 5556
rect 224000 5516 224006 5528
rect 423582 5516 423588 5528
rect 423640 5516 423646 5568
rect 1104 5466 422832 5488
rect 1104 5414 71648 5466
rect 71700 5414 71712 5466
rect 71764 5414 71776 5466
rect 71828 5414 71840 5466
rect 71892 5414 212982 5466
rect 213034 5414 213046 5466
rect 213098 5414 213110 5466
rect 213162 5414 213174 5466
rect 213226 5414 354315 5466
rect 354367 5414 354379 5466
rect 354431 5414 354443 5466
rect 354495 5414 354507 5466
rect 354559 5414 422832 5466
rect 1104 5392 422832 5414
rect 215662 5312 215668 5364
rect 215720 5352 215726 5364
rect 215941 5355 215999 5361
rect 215941 5352 215953 5355
rect 215720 5324 215953 5352
rect 215720 5312 215726 5324
rect 215941 5321 215953 5324
rect 215987 5321 215999 5355
rect 217870 5352 217876 5364
rect 217831 5324 217876 5352
rect 215941 5315 215999 5321
rect 217870 5312 217876 5324
rect 217928 5312 217934 5364
rect 221458 5352 221464 5364
rect 221419 5324 221464 5352
rect 221458 5312 221464 5324
rect 221516 5312 221522 5364
rect 223942 5352 223948 5364
rect 223903 5324 223948 5352
rect 223942 5312 223948 5324
rect 224000 5312 224006 5364
rect 209222 5284 209228 5296
rect 209183 5256 209228 5284
rect 209222 5244 209228 5256
rect 209280 5244 209286 5296
rect 212810 5244 212816 5296
rect 212868 5284 212874 5296
rect 213181 5287 213239 5293
rect 213181 5284 213193 5287
rect 212868 5256 213193 5284
rect 212868 5244 212874 5256
rect 213181 5253 213193 5256
rect 213227 5253 213239 5287
rect 213181 5247 213239 5253
rect 214558 5244 214564 5296
rect 214616 5284 214622 5296
rect 216677 5287 216735 5293
rect 216677 5284 216689 5287
rect 214616 5256 216689 5284
rect 214616 5244 214622 5256
rect 216677 5253 216689 5256
rect 216723 5284 216735 5287
rect 216723 5256 217088 5284
rect 216723 5253 216735 5256
rect 216677 5247 216735 5253
rect 216766 5216 216772 5228
rect 216727 5188 216772 5216
rect 216766 5176 216772 5188
rect 216824 5176 216830 5228
rect 93121 5151 93179 5157
rect 93121 5117 93133 5151
rect 93167 5148 93179 5151
rect 208857 5151 208915 5157
rect 208857 5148 208869 5151
rect 93167 5120 93808 5148
rect 93167 5117 93179 5120
rect 93121 5111 93179 5117
rect 93780 5024 93808 5120
rect 208596 5120 208869 5148
rect 208596 5024 208624 5120
rect 208857 5117 208869 5120
rect 208903 5117 208915 5151
rect 209038 5148 209044 5160
rect 208999 5120 209044 5148
rect 208857 5111 208915 5117
rect 209038 5108 209044 5120
rect 209096 5108 209102 5160
rect 212261 5151 212319 5157
rect 212261 5117 212273 5151
rect 212307 5148 212319 5151
rect 212350 5148 212356 5160
rect 212307 5120 212356 5148
rect 212307 5117 212319 5120
rect 212261 5111 212319 5117
rect 212350 5108 212356 5120
rect 212408 5108 212414 5160
rect 214285 5151 214343 5157
rect 214285 5117 214297 5151
rect 214331 5148 214343 5151
rect 215021 5151 215079 5157
rect 215021 5148 215033 5151
rect 214331 5120 215033 5148
rect 214331 5117 214343 5120
rect 214285 5111 214343 5117
rect 215021 5117 215033 5120
rect 215067 5148 215079 5151
rect 216306 5148 216312 5160
rect 215067 5120 216312 5148
rect 215067 5117 215079 5120
rect 215021 5111 215079 5117
rect 216306 5108 216312 5120
rect 216364 5108 216370 5160
rect 217060 5157 217088 5256
rect 223960 5216 223988 5312
rect 224402 5284 224408 5296
rect 224363 5256 224408 5284
rect 224402 5244 224408 5256
rect 224460 5244 224466 5296
rect 224037 5219 224095 5225
rect 224037 5216 224049 5219
rect 223960 5188 224049 5216
rect 224037 5185 224049 5188
rect 224083 5185 224095 5219
rect 224037 5179 224095 5185
rect 217045 5151 217103 5157
rect 217045 5117 217057 5151
rect 217091 5117 217103 5151
rect 217045 5111 217103 5117
rect 217505 5151 217563 5157
rect 217505 5117 217517 5151
rect 217551 5148 217563 5151
rect 220538 5148 220544 5160
rect 217551 5120 220544 5148
rect 217551 5117 217563 5120
rect 217505 5111 217563 5117
rect 220538 5108 220544 5120
rect 220596 5108 220602 5160
rect 224218 5148 224224 5160
rect 224179 5120 224224 5148
rect 224218 5108 224224 5120
rect 224276 5108 224282 5160
rect 212166 5080 212172 5092
rect 212079 5052 212172 5080
rect 212166 5040 212172 5052
rect 212224 5080 212230 5092
rect 212623 5083 212681 5089
rect 212623 5080 212635 5083
rect 212224 5052 212635 5080
rect 212224 5040 212230 5052
rect 212623 5049 212635 5052
rect 212669 5080 212681 5083
rect 214926 5080 214932 5092
rect 212669 5052 214932 5080
rect 212669 5049 212681 5052
rect 212623 5043 212681 5049
rect 214926 5040 214932 5052
rect 214984 5080 214990 5092
rect 215342 5083 215400 5089
rect 215342 5080 215354 5083
rect 214984 5052 215354 5080
rect 214984 5040 214990 5052
rect 215342 5049 215354 5052
rect 215388 5049 215400 5083
rect 215342 5043 215400 5049
rect 216858 5040 216864 5092
rect 216916 5080 216922 5092
rect 216953 5083 217011 5089
rect 216953 5080 216965 5083
rect 216916 5052 216965 5080
rect 216916 5040 216922 5052
rect 216953 5049 216965 5052
rect 216999 5049 217011 5083
rect 217134 5080 217140 5092
rect 217095 5052 217140 5080
rect 216953 5043 217011 5049
rect 217134 5040 217140 5052
rect 217192 5040 217198 5092
rect 220862 5083 220920 5089
rect 220862 5049 220874 5083
rect 220908 5049 220920 5083
rect 220862 5043 220920 5049
rect 93302 5012 93308 5024
rect 93263 4984 93308 5012
rect 93302 4972 93308 4984
rect 93360 4972 93366 5024
rect 93762 5012 93768 5024
rect 93723 4984 93768 5012
rect 93762 4972 93768 4984
rect 93820 4972 93826 5024
rect 208578 5012 208584 5024
rect 208539 4984 208584 5012
rect 208578 4972 208584 4984
rect 208636 4972 208642 5024
rect 216309 5015 216367 5021
rect 216309 4981 216321 5015
rect 216355 5012 216367 5015
rect 216490 5012 216496 5024
rect 216355 4984 216496 5012
rect 216355 4981 216367 4984
rect 216309 4975 216367 4981
rect 216490 4972 216496 4984
rect 216548 4972 216554 5024
rect 218146 5012 218152 5024
rect 218107 4984 218152 5012
rect 218146 4972 218152 4984
rect 218204 4972 218210 5024
rect 220354 5012 220360 5024
rect 220315 4984 220360 5012
rect 220354 4972 220360 4984
rect 220412 5012 220418 5024
rect 220877 5012 220905 5043
rect 220412 4984 220905 5012
rect 220412 4972 220418 4984
rect 1104 4922 422832 4944
rect 1104 4870 142315 4922
rect 142367 4870 142379 4922
rect 142431 4870 142443 4922
rect 142495 4870 142507 4922
rect 142559 4870 283648 4922
rect 283700 4870 283712 4922
rect 283764 4870 283776 4922
rect 283828 4870 283840 4922
rect 283892 4870 422832 4922
rect 1104 4848 422832 4870
rect 208949 4811 209007 4817
rect 208949 4777 208961 4811
rect 208995 4808 209007 4811
rect 209038 4808 209044 4820
rect 208995 4780 209044 4808
rect 208995 4777 209007 4780
rect 208949 4771 209007 4777
rect 209038 4768 209044 4780
rect 209096 4768 209102 4820
rect 213730 4768 213736 4820
rect 213788 4808 213794 4820
rect 214837 4811 214895 4817
rect 214837 4808 214849 4811
rect 213788 4780 214849 4808
rect 213788 4768 213794 4780
rect 214837 4777 214849 4780
rect 214883 4808 214895 4811
rect 215110 4808 215116 4820
rect 214883 4780 215116 4808
rect 214883 4777 214895 4780
rect 214837 4771 214895 4777
rect 215110 4768 215116 4780
rect 215168 4768 215174 4820
rect 216217 4811 216275 4817
rect 216217 4777 216229 4811
rect 216263 4808 216275 4811
rect 220538 4808 220544 4820
rect 216263 4780 216812 4808
rect 220499 4780 220544 4808
rect 216263 4777 216275 4780
rect 216217 4771 216275 4777
rect 214926 4700 214932 4752
rect 214984 4740 214990 4752
rect 215618 4743 215676 4749
rect 215618 4740 215630 4743
rect 214984 4712 215630 4740
rect 214984 4700 214990 4712
rect 215618 4709 215630 4712
rect 215664 4709 215676 4743
rect 216784 4740 216812 4780
rect 220538 4768 220544 4780
rect 220596 4768 220602 4820
rect 224034 4768 224040 4820
rect 224092 4808 224098 4820
rect 224129 4811 224187 4817
rect 224129 4808 224141 4811
rect 224092 4780 224141 4808
rect 224092 4768 224098 4780
rect 224129 4777 224141 4780
rect 224175 4808 224187 4811
rect 224218 4808 224224 4820
rect 224175 4780 224224 4808
rect 224175 4777 224187 4780
rect 224129 4771 224187 4777
rect 224218 4768 224224 4780
rect 224276 4768 224282 4820
rect 217502 4740 217508 4752
rect 216784 4712 217508 4740
rect 215618 4703 215676 4709
rect 217502 4700 217508 4712
rect 217560 4740 217566 4752
rect 218146 4740 218152 4752
rect 217560 4712 218152 4740
rect 217560 4700 217566 4712
rect 218146 4700 218152 4712
rect 218204 4700 218210 4752
rect 218327 4743 218385 4749
rect 218327 4709 218339 4743
rect 218373 4740 218385 4743
rect 218422 4740 218428 4752
rect 218373 4712 218428 4740
rect 218373 4709 218385 4712
rect 218327 4703 218385 4709
rect 218422 4700 218428 4712
rect 218480 4740 218486 4752
rect 220354 4740 220360 4752
rect 218480 4712 220360 4740
rect 218480 4700 218486 4712
rect 220354 4700 220360 4712
rect 220412 4700 220418 4752
rect 213822 4672 213828 4684
rect 213783 4644 213828 4672
rect 213822 4632 213828 4644
rect 213880 4632 213886 4684
rect 214466 4672 214472 4684
rect 214379 4644 214472 4672
rect 214466 4632 214472 4644
rect 214524 4672 214530 4684
rect 216674 4672 216680 4684
rect 214524 4644 216680 4672
rect 214524 4632 214530 4644
rect 216674 4632 216680 4644
rect 216732 4632 216738 4684
rect 214282 4564 214288 4616
rect 214340 4604 214346 4616
rect 215297 4607 215355 4613
rect 215297 4604 215309 4607
rect 214340 4576 215309 4604
rect 214340 4564 214346 4576
rect 215297 4573 215309 4576
rect 215343 4573 215355 4607
rect 215297 4567 215355 4573
rect 217965 4607 218023 4613
rect 217965 4573 217977 4607
rect 218011 4604 218023 4607
rect 218330 4604 218336 4616
rect 218011 4576 218336 4604
rect 218011 4573 218023 4576
rect 217965 4567 218023 4573
rect 218330 4564 218336 4576
rect 218388 4564 218394 4616
rect 212350 4468 212356 4480
rect 212311 4440 212356 4468
rect 212350 4428 212356 4440
rect 212408 4428 212414 4480
rect 212810 4468 212816 4480
rect 212771 4440 212816 4468
rect 212810 4428 212816 4440
rect 212868 4428 212874 4480
rect 215205 4471 215263 4477
rect 215205 4437 215217 4471
rect 215251 4468 215263 4471
rect 215386 4468 215392 4480
rect 215251 4440 215392 4468
rect 215251 4437 215263 4440
rect 215205 4431 215263 4437
rect 215386 4428 215392 4440
rect 215444 4468 215450 4480
rect 216858 4468 216864 4480
rect 215444 4440 216864 4468
rect 215444 4428 215450 4440
rect 216858 4428 216864 4440
rect 216916 4428 216922 4480
rect 218885 4471 218943 4477
rect 218885 4437 218897 4471
rect 218931 4468 218943 4471
rect 220446 4468 220452 4480
rect 218931 4440 220452 4468
rect 218931 4437 218943 4440
rect 218885 4431 218943 4437
rect 220446 4428 220452 4440
rect 220504 4428 220510 4480
rect 1104 4378 422832 4400
rect 1104 4326 71648 4378
rect 71700 4326 71712 4378
rect 71764 4326 71776 4378
rect 71828 4326 71840 4378
rect 71892 4326 212982 4378
rect 213034 4326 213046 4378
rect 213098 4326 213110 4378
rect 213162 4326 213174 4378
rect 213226 4326 354315 4378
rect 354367 4326 354379 4378
rect 354431 4326 354443 4378
rect 354495 4326 354507 4378
rect 354559 4326 422832 4378
rect 1104 4304 422832 4326
rect 214282 4264 214288 4276
rect 214243 4236 214288 4264
rect 214282 4224 214288 4236
rect 214340 4224 214346 4276
rect 214926 4224 214932 4276
rect 214984 4264 214990 4276
rect 215113 4267 215171 4273
rect 215113 4264 215125 4267
rect 214984 4236 215125 4264
rect 214984 4224 214990 4236
rect 215113 4233 215125 4236
rect 215159 4264 215171 4267
rect 218057 4267 218115 4273
rect 218057 4264 218069 4267
rect 215159 4236 218069 4264
rect 215159 4233 215171 4236
rect 215113 4227 215171 4233
rect 218057 4233 218069 4236
rect 218103 4264 218115 4267
rect 218422 4264 218428 4276
rect 218103 4236 218428 4264
rect 218103 4233 218115 4236
rect 218057 4227 218115 4233
rect 218422 4224 218428 4236
rect 218480 4224 218486 4276
rect 215018 4088 215024 4140
rect 215076 4128 215082 4140
rect 215076 4100 215984 4128
rect 215076 4088 215082 4100
rect 212353 4063 212411 4069
rect 212353 4029 212365 4063
rect 212399 4060 212411 4063
rect 213089 4063 213147 4069
rect 213089 4060 213101 4063
rect 212399 4032 213101 4060
rect 212399 4029 212411 4032
rect 212353 4023 212411 4029
rect 213089 4029 213101 4032
rect 213135 4060 213147 4063
rect 214466 4060 214472 4072
rect 213135 4032 214472 4060
rect 213135 4029 213147 4032
rect 213089 4023 213147 4029
rect 214466 4020 214472 4032
rect 214524 4020 214530 4072
rect 215757 4063 215815 4069
rect 215757 4029 215769 4063
rect 215803 4029 215815 4063
rect 215956 4060 215984 4100
rect 216033 4063 216091 4069
rect 216033 4060 216045 4063
rect 215956 4032 216045 4060
rect 215757 4023 215815 4029
rect 216033 4029 216045 4032
rect 216079 4029 216091 4063
rect 216398 4060 216404 4072
rect 216359 4032 216404 4060
rect 216033 4023 216091 4029
rect 212810 3992 212816 4004
rect 212771 3964 212816 3992
rect 212810 3952 212816 3964
rect 212868 3952 212874 4004
rect 213178 3992 213184 4004
rect 213139 3964 213184 3992
rect 213178 3952 213184 3964
rect 213236 3952 213242 4004
rect 213546 3992 213552 4004
rect 213507 3964 213552 3992
rect 213546 3952 213552 3964
rect 213604 3952 213610 4004
rect 215386 3992 215392 4004
rect 213840 3964 215392 3992
rect 213840 3936 213868 3964
rect 215386 3952 215392 3964
rect 215444 3952 215450 4004
rect 212626 3924 212632 3936
rect 212587 3896 212632 3924
rect 212626 3884 212632 3896
rect 212684 3924 212690 3936
rect 212997 3927 213055 3933
rect 212997 3924 213009 3927
rect 212684 3896 213009 3924
rect 212684 3884 212690 3896
rect 212997 3893 213009 3896
rect 213043 3893 213055 3927
rect 212997 3887 213055 3893
rect 213270 3884 213276 3936
rect 213328 3924 213334 3936
rect 213822 3924 213828 3936
rect 213328 3896 213828 3924
rect 213328 3884 213334 3896
rect 213822 3884 213828 3896
rect 213880 3884 213886 3936
rect 214742 3924 214748 3936
rect 214703 3896 214748 3924
rect 214742 3884 214748 3896
rect 214800 3884 214806 3936
rect 215404 3924 215432 3952
rect 215772 3924 215800 4023
rect 216398 4020 216404 4032
rect 216456 4020 216462 4072
rect 216490 4020 216496 4072
rect 216548 4060 216554 4072
rect 216953 4063 217011 4069
rect 216953 4060 216965 4063
rect 216548 4032 216965 4060
rect 216548 4020 216554 4032
rect 216953 4029 216965 4032
rect 216999 4060 217011 4063
rect 217134 4060 217140 4072
rect 216999 4032 217140 4060
rect 216999 4029 217011 4032
rect 216953 4023 217011 4029
rect 217134 4020 217140 4032
rect 217192 4060 217198 4072
rect 217192 4032 217456 4060
rect 217192 4020 217198 4032
rect 217042 3992 217048 4004
rect 217003 3964 217048 3992
rect 217042 3952 217048 3964
rect 217100 3952 217106 4004
rect 217428 3933 217456 4032
rect 217594 3952 217600 4004
rect 217652 3992 217658 4004
rect 218330 3992 218336 4004
rect 217652 3964 218336 3992
rect 217652 3952 217658 3964
rect 218330 3952 218336 3964
rect 218388 3952 218394 4004
rect 215404 3896 215800 3924
rect 217413 3927 217471 3933
rect 217413 3893 217425 3927
rect 217459 3924 217471 3927
rect 217778 3924 217784 3936
rect 217459 3896 217784 3924
rect 217459 3893 217471 3896
rect 217413 3887 217471 3893
rect 217778 3884 217784 3896
rect 217836 3884 217842 3936
rect 1104 3834 422832 3856
rect 1104 3782 142315 3834
rect 142367 3782 142379 3834
rect 142431 3782 142443 3834
rect 142495 3782 142507 3834
rect 142559 3782 283648 3834
rect 283700 3782 283712 3834
rect 283764 3782 283776 3834
rect 283828 3782 283840 3834
rect 283892 3782 422832 3834
rect 1104 3760 422832 3782
rect 212350 3680 212356 3732
rect 212408 3720 212414 3732
rect 213365 3723 213423 3729
rect 213365 3720 213377 3723
rect 212408 3692 213377 3720
rect 212408 3680 212414 3692
rect 213365 3689 213377 3692
rect 213411 3689 213423 3723
rect 216398 3720 216404 3732
rect 213365 3683 213423 3689
rect 215588 3692 216404 3720
rect 212537 3655 212595 3661
rect 212537 3621 212549 3655
rect 212583 3652 212595 3655
rect 212810 3652 212816 3664
rect 212583 3624 212816 3652
rect 212583 3621 212595 3624
rect 212537 3615 212595 3621
rect 212810 3612 212816 3624
rect 212868 3652 212874 3664
rect 214742 3652 214748 3664
rect 212868 3624 214748 3652
rect 212868 3612 212874 3624
rect 213270 3584 213276 3596
rect 213231 3556 213276 3584
rect 213270 3544 213276 3556
rect 213328 3544 213334 3596
rect 213730 3584 213736 3596
rect 213643 3556 213736 3584
rect 213730 3544 213736 3556
rect 213788 3544 213794 3596
rect 214116 3593 214144 3624
rect 214742 3612 214748 3624
rect 214800 3652 214806 3664
rect 215588 3661 215616 3692
rect 216398 3680 216404 3692
rect 216456 3720 216462 3732
rect 216585 3723 216643 3729
rect 216585 3720 216597 3723
rect 216456 3692 216597 3720
rect 216456 3680 216462 3692
rect 216585 3689 216597 3692
rect 216631 3689 216643 3723
rect 216585 3683 216643 3689
rect 216674 3680 216680 3732
rect 216732 3720 216738 3732
rect 216953 3723 217011 3729
rect 216953 3720 216965 3723
rect 216732 3692 216965 3720
rect 216732 3680 216738 3692
rect 216953 3689 216965 3692
rect 216999 3689 217011 3723
rect 216953 3683 217011 3689
rect 220633 3723 220691 3729
rect 220633 3689 220645 3723
rect 220679 3720 220691 3723
rect 224034 3720 224040 3732
rect 220679 3692 224040 3720
rect 220679 3689 220691 3692
rect 220633 3683 220691 3689
rect 224034 3680 224040 3692
rect 224092 3680 224098 3732
rect 215021 3655 215079 3661
rect 215021 3652 215033 3655
rect 214800 3624 215033 3652
rect 214800 3612 214806 3624
rect 215021 3621 215033 3624
rect 215067 3652 215079 3655
rect 215573 3655 215631 3661
rect 215573 3652 215585 3655
rect 215067 3624 215585 3652
rect 215067 3621 215079 3624
rect 215021 3615 215079 3621
rect 215573 3621 215585 3624
rect 215619 3621 215631 3655
rect 215573 3615 215631 3621
rect 215941 3655 215999 3661
rect 215941 3621 215953 3655
rect 215987 3621 215999 3655
rect 216306 3652 216312 3664
rect 216267 3624 216312 3652
rect 215941 3615 215999 3621
rect 214101 3587 214159 3593
rect 214101 3553 214113 3587
rect 214147 3553 214159 3587
rect 214466 3584 214472 3596
rect 214427 3556 214472 3584
rect 214101 3547 214159 3553
rect 214466 3544 214472 3556
rect 214524 3584 214530 3596
rect 215754 3584 215760 3596
rect 214524 3556 215760 3584
rect 214524 3544 214530 3556
rect 215754 3544 215760 3556
rect 215812 3544 215818 3596
rect 215849 3587 215907 3593
rect 215849 3553 215861 3587
rect 215895 3553 215907 3587
rect 215849 3547 215907 3553
rect 215956 3584 215984 3615
rect 216306 3612 216312 3624
rect 216364 3612 216370 3664
rect 220075 3655 220133 3661
rect 220075 3621 220087 3655
rect 220121 3652 220133 3655
rect 220446 3652 220452 3664
rect 220121 3624 220452 3652
rect 220121 3621 220133 3624
rect 220075 3615 220133 3621
rect 220446 3612 220452 3624
rect 220504 3612 220510 3664
rect 216858 3584 216864 3596
rect 215956 3556 216864 3584
rect 211982 3476 211988 3528
rect 212040 3516 212046 3528
rect 213748 3516 213776 3544
rect 212040 3488 213776 3516
rect 212040 3476 212046 3488
rect 215386 3476 215392 3528
rect 215444 3516 215450 3528
rect 215864 3516 215892 3547
rect 215444 3488 215892 3516
rect 215444 3476 215450 3488
rect 212905 3451 212963 3457
rect 212905 3417 212917 3451
rect 212951 3448 212963 3451
rect 213178 3448 213184 3460
rect 212951 3420 213184 3448
rect 212951 3417 212963 3420
rect 212905 3411 212963 3417
rect 213178 3408 213184 3420
rect 213236 3448 213242 3460
rect 213638 3448 213644 3460
rect 213236 3420 213644 3448
rect 213236 3408 213242 3420
rect 213638 3408 213644 3420
rect 213696 3448 213702 3460
rect 215481 3451 215539 3457
rect 215481 3448 215493 3451
rect 213696 3420 215493 3448
rect 213696 3408 213702 3420
rect 215481 3417 215493 3420
rect 215527 3448 215539 3451
rect 215956 3448 215984 3556
rect 216858 3544 216864 3556
rect 216916 3544 216922 3596
rect 217502 3584 217508 3596
rect 217463 3556 217508 3584
rect 217502 3544 217508 3556
rect 217560 3544 217566 3596
rect 217042 3476 217048 3528
rect 217100 3516 217106 3528
rect 219710 3516 219716 3528
rect 217100 3488 219716 3516
rect 217100 3476 217106 3488
rect 219710 3476 219716 3488
rect 219768 3476 219774 3528
rect 217502 3448 217508 3460
rect 215527 3420 215984 3448
rect 216646 3420 217508 3448
rect 215527 3417 215539 3420
rect 215481 3411 215539 3417
rect 215754 3340 215760 3392
rect 215812 3380 215818 3392
rect 216646 3380 216674 3420
rect 217502 3408 217508 3420
rect 217560 3408 217566 3460
rect 217778 3380 217784 3392
rect 215812 3352 216674 3380
rect 217739 3352 217784 3380
rect 215812 3340 215818 3352
rect 217778 3340 217784 3352
rect 217836 3340 217842 3392
rect 1104 3290 422832 3312
rect 1104 3238 71648 3290
rect 71700 3238 71712 3290
rect 71764 3238 71776 3290
rect 71828 3238 71840 3290
rect 71892 3238 212982 3290
rect 213034 3238 213046 3290
rect 213098 3238 213110 3290
rect 213162 3238 213174 3290
rect 213226 3238 354315 3290
rect 354367 3238 354379 3290
rect 354431 3238 354443 3290
rect 354495 3238 354507 3290
rect 354559 3238 422832 3290
rect 1104 3216 422832 3238
rect 211982 3176 211988 3188
rect 211943 3148 211988 3176
rect 211982 3136 211988 3148
rect 212040 3136 212046 3188
rect 212166 3136 212172 3188
rect 212224 3176 212230 3188
rect 212261 3179 212319 3185
rect 212261 3176 212273 3179
rect 212224 3148 212273 3176
rect 212224 3136 212230 3148
rect 212261 3145 212273 3148
rect 212307 3145 212319 3179
rect 212261 3139 212319 3145
rect 212626 3136 212632 3188
rect 212684 3176 212690 3188
rect 214009 3179 214067 3185
rect 214009 3176 214021 3179
rect 212684 3148 214021 3176
rect 212684 3136 212690 3148
rect 214009 3145 214021 3148
rect 214055 3176 214067 3179
rect 214466 3176 214472 3188
rect 214055 3148 214472 3176
rect 214055 3145 214067 3148
rect 214009 3139 214067 3145
rect 214466 3136 214472 3148
rect 214524 3136 214530 3188
rect 214653 3179 214711 3185
rect 214653 3145 214665 3179
rect 214699 3176 214711 3179
rect 214742 3176 214748 3188
rect 214699 3148 214748 3176
rect 214699 3145 214711 3148
rect 214653 3139 214711 3145
rect 214742 3136 214748 3148
rect 214800 3136 214806 3188
rect 215386 3136 215392 3188
rect 215444 3176 215450 3188
rect 215573 3179 215631 3185
rect 215573 3176 215585 3179
rect 215444 3148 215585 3176
rect 215444 3136 215450 3148
rect 215573 3145 215585 3148
rect 215619 3145 215631 3179
rect 217502 3176 217508 3188
rect 217463 3148 217508 3176
rect 215573 3139 215631 3145
rect 217502 3136 217508 3148
rect 217560 3136 217566 3188
rect 208946 3068 208952 3120
rect 209004 3108 209010 3120
rect 213365 3111 213423 3117
rect 213365 3108 213377 3111
rect 209004 3080 213377 3108
rect 209004 3068 209010 3080
rect 213365 3077 213377 3080
rect 213411 3077 213423 3111
rect 214484 3108 214512 3136
rect 214834 3108 214840 3120
rect 214484 3080 214840 3108
rect 213365 3071 213423 3077
rect 214834 3068 214840 3080
rect 214892 3108 214898 3120
rect 215205 3111 215263 3117
rect 215205 3108 215217 3111
rect 214892 3080 215217 3108
rect 214892 3068 214898 3080
rect 215205 3077 215217 3080
rect 215251 3077 215263 3111
rect 215205 3071 215263 3077
rect 211617 3043 211675 3049
rect 211617 3009 211629 3043
rect 211663 3040 211675 3043
rect 212445 3043 212503 3049
rect 212445 3040 212457 3043
rect 211663 3012 212457 3040
rect 211663 3009 211675 3012
rect 211617 3003 211675 3009
rect 212445 3009 212457 3012
rect 212491 3040 212503 3043
rect 213546 3040 213552 3052
rect 212491 3012 213552 3040
rect 212491 3009 212503 3012
rect 212445 3003 212503 3009
rect 213546 3000 213552 3012
rect 213604 3000 213610 3052
rect 216674 3040 216680 3052
rect 216048 3012 216680 3040
rect 214469 2975 214527 2981
rect 214469 2941 214481 2975
rect 214515 2972 214527 2975
rect 214558 2972 214564 2984
rect 214515 2944 214564 2972
rect 214515 2941 214527 2944
rect 214469 2935 214527 2941
rect 214558 2932 214564 2944
rect 214616 2932 214622 2984
rect 216048 2981 216076 3012
rect 216674 3000 216680 3012
rect 216732 3000 216738 3052
rect 216033 2975 216091 2981
rect 216033 2941 216045 2975
rect 216079 2941 216091 2975
rect 216033 2935 216091 2941
rect 216122 2932 216128 2984
rect 216180 2972 216186 2984
rect 216217 2975 216275 2981
rect 216217 2972 216229 2975
rect 216180 2944 216229 2972
rect 216180 2932 216186 2944
rect 216217 2941 216229 2944
rect 216263 2941 216275 2975
rect 216217 2935 216275 2941
rect 216398 2932 216404 2984
rect 216456 2972 216462 2984
rect 216585 2975 216643 2981
rect 216585 2972 216597 2975
rect 216456 2944 216597 2972
rect 216456 2932 216462 2944
rect 216585 2941 216597 2944
rect 216631 2941 216643 2975
rect 216585 2935 216643 2941
rect 216953 2975 217011 2981
rect 216953 2941 216965 2975
rect 216999 2941 217011 2975
rect 216953 2935 217011 2941
rect 217229 2975 217287 2981
rect 217229 2941 217241 2975
rect 217275 2972 217287 2975
rect 220078 2972 220084 2984
rect 217275 2944 220084 2972
rect 217275 2941 217287 2944
rect 217229 2935 217287 2941
rect 212166 2864 212172 2916
rect 212224 2904 212230 2916
rect 212766 2907 212824 2913
rect 212766 2904 212778 2907
rect 212224 2876 212778 2904
rect 212224 2864 212230 2876
rect 212766 2873 212778 2876
rect 212812 2873 212824 2907
rect 212766 2867 212824 2873
rect 214098 2864 214104 2916
rect 214156 2904 214162 2916
rect 216968 2904 216996 2935
rect 220078 2932 220084 2944
rect 220136 2932 220142 2984
rect 217778 2904 217784 2916
rect 214156 2876 217784 2904
rect 214156 2864 214162 2876
rect 217778 2864 217784 2876
rect 217836 2904 217842 2916
rect 217873 2907 217931 2913
rect 217873 2904 217885 2907
rect 217836 2876 217885 2904
rect 217836 2864 217842 2876
rect 217873 2873 217885 2876
rect 217919 2873 217931 2907
rect 217873 2867 217931 2873
rect 213270 2796 213276 2848
rect 213328 2836 213334 2848
rect 213641 2839 213699 2845
rect 213641 2836 213653 2839
rect 213328 2808 213653 2836
rect 213328 2796 213334 2808
rect 213641 2805 213653 2808
rect 213687 2805 213699 2839
rect 218238 2836 218244 2848
rect 218199 2808 218244 2836
rect 213641 2799 213699 2805
rect 218238 2796 218244 2808
rect 218296 2796 218302 2848
rect 219529 2839 219587 2845
rect 219529 2805 219541 2839
rect 219575 2836 219587 2839
rect 219897 2839 219955 2845
rect 219897 2836 219909 2839
rect 219575 2808 219909 2836
rect 219575 2805 219587 2808
rect 219529 2799 219587 2805
rect 219897 2805 219909 2808
rect 219943 2836 219955 2839
rect 220446 2836 220452 2848
rect 219943 2808 220452 2836
rect 219943 2805 219955 2808
rect 219897 2799 219955 2805
rect 220446 2796 220452 2808
rect 220504 2796 220510 2848
rect 220998 2836 221004 2848
rect 220959 2808 221004 2836
rect 220998 2796 221004 2808
rect 221056 2796 221062 2848
rect 1104 2746 422832 2768
rect 1104 2694 142315 2746
rect 142367 2694 142379 2746
rect 142431 2694 142443 2746
rect 142495 2694 142507 2746
rect 142559 2694 283648 2746
rect 283700 2694 283712 2746
rect 283764 2694 283776 2746
rect 283828 2694 283840 2746
rect 283892 2694 422832 2746
rect 1104 2672 422832 2694
rect 209222 2592 209228 2644
rect 209280 2632 209286 2644
rect 211617 2635 211675 2641
rect 211617 2632 211629 2635
rect 209280 2604 211629 2632
rect 209280 2592 209286 2604
rect 211617 2601 211629 2604
rect 211663 2601 211675 2635
rect 211617 2595 211675 2601
rect 212077 2635 212135 2641
rect 212077 2601 212089 2635
rect 212123 2632 212135 2635
rect 212994 2632 213000 2644
rect 212123 2604 212534 2632
rect 212907 2604 213000 2632
rect 212123 2601 212135 2604
rect 212077 2595 212135 2601
rect 211632 2496 211660 2595
rect 212506 2564 212534 2604
rect 212994 2592 213000 2604
rect 213052 2632 213058 2644
rect 213733 2635 213791 2641
rect 213733 2632 213745 2635
rect 213052 2604 213745 2632
rect 213052 2592 213058 2604
rect 213733 2601 213745 2604
rect 213779 2632 213791 2635
rect 214558 2632 214564 2644
rect 213779 2604 214564 2632
rect 213779 2601 213791 2604
rect 213733 2595 213791 2601
rect 214558 2592 214564 2604
rect 214616 2592 214622 2644
rect 214834 2632 214840 2644
rect 214795 2604 214840 2632
rect 214834 2592 214840 2604
rect 214892 2592 214898 2644
rect 216766 2632 216772 2644
rect 215496 2604 216772 2632
rect 213638 2564 213644 2576
rect 212506 2536 213644 2564
rect 213638 2524 213644 2536
rect 213696 2524 213702 2576
rect 213825 2567 213883 2573
rect 213825 2533 213837 2567
rect 213871 2564 213883 2567
rect 214098 2564 214104 2576
rect 213871 2536 214104 2564
rect 213871 2533 213883 2536
rect 213825 2527 213883 2533
rect 212261 2499 212319 2505
rect 212261 2496 212273 2499
rect 211632 2468 212273 2496
rect 212261 2465 212273 2468
rect 212307 2465 212319 2499
rect 213270 2496 213276 2508
rect 213231 2468 213276 2496
rect 212261 2459 212319 2465
rect 213270 2456 213276 2468
rect 213328 2496 213334 2508
rect 213457 2499 213515 2505
rect 213457 2496 213469 2499
rect 213328 2468 213469 2496
rect 213328 2456 213334 2468
rect 213457 2465 213469 2468
rect 213503 2465 213515 2499
rect 213840 2496 213868 2527
rect 214098 2524 214104 2536
rect 214156 2524 214162 2576
rect 214193 2567 214251 2573
rect 214193 2533 214205 2567
rect 214239 2564 214251 2567
rect 214282 2564 214288 2576
rect 214239 2536 214288 2564
rect 214239 2533 214251 2536
rect 214193 2527 214251 2533
rect 214282 2524 214288 2536
rect 214340 2524 214346 2576
rect 215496 2505 215524 2604
rect 216766 2592 216772 2604
rect 216824 2632 216830 2644
rect 217321 2635 217379 2641
rect 217321 2632 217333 2635
rect 216824 2604 217333 2632
rect 216824 2592 216830 2604
rect 217321 2601 217333 2604
rect 217367 2601 217379 2635
rect 217321 2595 217379 2601
rect 217781 2635 217839 2641
rect 217781 2601 217793 2635
rect 217827 2632 217839 2635
rect 218238 2632 218244 2644
rect 217827 2604 218244 2632
rect 217827 2601 217839 2604
rect 217781 2595 217839 2601
rect 215754 2524 215760 2576
rect 215812 2564 215818 2576
rect 216677 2567 216735 2573
rect 215812 2536 216444 2564
rect 215812 2524 215818 2536
rect 213457 2459 213515 2465
rect 213656 2468 213868 2496
rect 215481 2499 215539 2505
rect 211341 2431 211399 2437
rect 211341 2397 211353 2431
rect 211387 2428 211399 2431
rect 213656 2428 213684 2468
rect 215481 2465 215493 2499
rect 215527 2465 215539 2499
rect 215481 2459 215539 2465
rect 215665 2499 215723 2505
rect 215665 2465 215677 2499
rect 215711 2496 215723 2499
rect 216122 2496 216128 2508
rect 215711 2468 216128 2496
rect 215711 2465 215723 2468
rect 215665 2459 215723 2465
rect 211387 2400 213684 2428
rect 211387 2397 211399 2400
rect 211341 2391 211399 2397
rect 213730 2388 213736 2440
rect 213788 2428 213794 2440
rect 215680 2428 215708 2459
rect 216122 2456 216128 2468
rect 216180 2456 216186 2508
rect 216217 2499 216275 2505
rect 216217 2465 216229 2499
rect 216263 2496 216275 2499
rect 216306 2496 216312 2508
rect 216263 2468 216312 2496
rect 216263 2465 216275 2468
rect 216217 2459 216275 2465
rect 216306 2456 216312 2468
rect 216364 2456 216370 2508
rect 216416 2505 216444 2536
rect 216677 2533 216689 2567
rect 216723 2564 216735 2567
rect 217594 2564 217600 2576
rect 216723 2536 217600 2564
rect 216723 2533 216735 2536
rect 216677 2527 216735 2533
rect 217594 2524 217600 2536
rect 217652 2524 217658 2576
rect 216401 2499 216459 2505
rect 216401 2465 216413 2499
rect 216447 2465 216459 2499
rect 216953 2499 217011 2505
rect 216953 2496 216965 2499
rect 216401 2459 216459 2465
rect 216646 2468 216965 2496
rect 213788 2400 215708 2428
rect 213788 2388 213794 2400
rect 216140 2360 216168 2456
rect 216324 2428 216352 2456
rect 216646 2428 216674 2468
rect 216953 2465 216965 2468
rect 216999 2465 217011 2499
rect 216953 2459 217011 2465
rect 216324 2400 216674 2428
rect 217796 2360 217824 2595
rect 218238 2592 218244 2604
rect 218296 2592 218302 2644
rect 219710 2632 219716 2644
rect 219671 2604 219716 2632
rect 219710 2592 219716 2604
rect 219768 2592 219774 2644
rect 220078 2632 220084 2644
rect 220039 2604 220084 2632
rect 220078 2592 220084 2604
rect 220136 2592 220142 2644
rect 220538 2632 220544 2644
rect 220499 2604 220544 2632
rect 220538 2592 220544 2604
rect 220596 2592 220602 2644
rect 221918 2632 221924 2644
rect 221879 2604 221924 2632
rect 221918 2592 221924 2604
rect 221976 2592 221982 2644
rect 220556 2496 220584 2592
rect 221461 2499 221519 2505
rect 221461 2496 221473 2499
rect 220556 2468 221473 2496
rect 221461 2465 221473 2468
rect 221507 2465 221519 2499
rect 221461 2459 221519 2465
rect 224402 2456 224408 2508
rect 224460 2496 224466 2508
rect 228177 2499 228235 2505
rect 228177 2496 228189 2499
rect 224460 2468 228189 2496
rect 224460 2456 224466 2468
rect 228177 2465 228189 2468
rect 228223 2496 228235 2499
rect 228729 2499 228787 2505
rect 228729 2496 228741 2499
rect 228223 2468 228741 2496
rect 228223 2465 228235 2468
rect 228177 2459 228235 2465
rect 228729 2465 228741 2468
rect 228775 2465 228787 2499
rect 309413 2499 309471 2505
rect 309413 2496 309425 2499
rect 228729 2459 228787 2465
rect 308600 2468 309425 2496
rect 308600 2440 308628 2468
rect 309413 2465 309425 2468
rect 309459 2465 309471 2499
rect 350810 2496 350816 2508
rect 350771 2468 350816 2496
rect 309413 2459 309471 2465
rect 350810 2456 350816 2468
rect 350868 2496 350874 2508
rect 351365 2499 351423 2505
rect 351365 2496 351377 2499
rect 350868 2468 351377 2496
rect 350868 2456 350874 2468
rect 351365 2465 351377 2468
rect 351411 2465 351423 2499
rect 351365 2459 351423 2465
rect 221277 2431 221335 2437
rect 221277 2397 221289 2431
rect 221323 2397 221335 2431
rect 308582 2428 308588 2440
rect 308543 2400 308588 2428
rect 221277 2391 221335 2397
rect 216140 2332 217824 2360
rect 212442 2292 212448 2304
rect 212403 2264 212448 2292
rect 212442 2252 212448 2264
rect 212500 2252 212506 2304
rect 221182 2292 221188 2304
rect 221143 2264 221188 2292
rect 221182 2252 221188 2264
rect 221240 2292 221246 2304
rect 221292 2292 221320 2391
rect 308582 2388 308588 2400
rect 308640 2388 308646 2440
rect 309229 2431 309287 2437
rect 309229 2397 309241 2431
rect 309275 2397 309287 2431
rect 309229 2391 309287 2397
rect 309045 2363 309103 2369
rect 309045 2329 309057 2363
rect 309091 2360 309103 2363
rect 309244 2360 309272 2391
rect 309870 2360 309876 2372
rect 309091 2332 309272 2360
rect 309831 2332 309876 2360
rect 309091 2329 309103 2332
rect 309045 2323 309103 2329
rect 228358 2292 228364 2304
rect 221240 2264 221320 2292
rect 228319 2264 228364 2292
rect 221240 2252 221246 2264
rect 228358 2252 228364 2264
rect 228416 2252 228422 2304
rect 309244 2292 309272 2332
rect 309870 2320 309876 2332
rect 309928 2320 309934 2372
rect 318058 2292 318064 2304
rect 309244 2264 318064 2292
rect 318058 2252 318064 2264
rect 318116 2252 318122 2304
rect 350994 2292 351000 2304
rect 350955 2264 351000 2292
rect 350994 2252 351000 2264
rect 351052 2252 351058 2304
rect 1104 2202 422832 2224
rect 1104 2150 71648 2202
rect 71700 2150 71712 2202
rect 71764 2150 71776 2202
rect 71828 2150 71840 2202
rect 71892 2150 212982 2202
rect 213034 2150 213046 2202
rect 213098 2150 213110 2202
rect 213162 2150 213174 2202
rect 213226 2150 354315 2202
rect 354367 2150 354379 2202
rect 354431 2150 354443 2202
rect 354495 2150 354507 2202
rect 354559 2150 422832 2202
rect 1104 2128 422832 2150
<< via1 >>
rect 112 8168 164 8220
rect 178224 8168 178276 8220
rect 71648 7590 71700 7642
rect 71712 7590 71764 7642
rect 71776 7590 71828 7642
rect 71840 7590 71892 7642
rect 212982 7590 213034 7642
rect 213046 7590 213098 7642
rect 213110 7590 213162 7642
rect 213174 7590 213226 7642
rect 354315 7590 354367 7642
rect 354379 7590 354431 7642
rect 354443 7590 354495 7642
rect 354507 7590 354559 7642
rect 178224 7531 178276 7540
rect 178224 7497 178233 7531
rect 178233 7497 178267 7531
rect 178267 7497 178276 7531
rect 178224 7488 178276 7497
rect 88616 7284 88668 7336
rect 106096 7216 106148 7268
rect 225696 7284 225748 7336
rect 190644 7148 190696 7200
rect 229560 7191 229612 7200
rect 229560 7157 229569 7191
rect 229569 7157 229603 7191
rect 229603 7157 229612 7191
rect 229560 7148 229612 7157
rect 142315 7046 142367 7098
rect 142379 7046 142431 7098
rect 142443 7046 142495 7098
rect 142507 7046 142559 7098
rect 283648 7046 283700 7098
rect 283712 7046 283764 7098
rect 283776 7046 283828 7098
rect 283840 7046 283892 7098
rect 176292 6944 176344 6996
rect 170680 6808 170732 6860
rect 75000 6740 75052 6792
rect 88248 6783 88300 6792
rect 88248 6749 88257 6783
rect 88257 6749 88291 6783
rect 88291 6749 88300 6783
rect 88248 6740 88300 6749
rect 88708 6740 88760 6792
rect 225328 6783 225380 6792
rect 225328 6749 225337 6783
rect 225337 6749 225371 6783
rect 225371 6749 225380 6783
rect 225328 6740 225380 6749
rect 225512 6783 225564 6792
rect 225512 6749 225521 6783
rect 225521 6749 225555 6783
rect 225555 6749 225564 6783
rect 225512 6740 225564 6749
rect 88616 6647 88668 6656
rect 88616 6613 88625 6647
rect 88625 6613 88659 6647
rect 88659 6613 88668 6647
rect 88616 6604 88668 6613
rect 215668 6647 215720 6656
rect 215668 6613 215677 6647
rect 215677 6613 215711 6647
rect 215711 6613 215720 6647
rect 215668 6604 215720 6613
rect 225696 6647 225748 6656
rect 225696 6613 225705 6647
rect 225705 6613 225739 6647
rect 225739 6613 225748 6647
rect 225696 6604 225748 6613
rect 71648 6502 71700 6554
rect 71712 6502 71764 6554
rect 71776 6502 71828 6554
rect 71840 6502 71892 6554
rect 212982 6502 213034 6554
rect 213046 6502 213098 6554
rect 213110 6502 213162 6554
rect 213174 6502 213226 6554
rect 354315 6502 354367 6554
rect 354379 6502 354431 6554
rect 354443 6502 354495 6554
rect 354507 6502 354559 6554
rect 88248 6443 88300 6452
rect 88248 6409 88257 6443
rect 88257 6409 88291 6443
rect 88291 6409 88300 6443
rect 88248 6400 88300 6409
rect 225328 6443 225380 6452
rect 225328 6409 225337 6443
rect 225337 6409 225371 6443
rect 225371 6409 225380 6443
rect 225328 6400 225380 6409
rect 215944 6375 215996 6384
rect 215944 6341 215953 6375
rect 215953 6341 215987 6375
rect 215987 6341 215996 6375
rect 215944 6332 215996 6341
rect 215576 6307 215628 6316
rect 215576 6273 215585 6307
rect 215585 6273 215619 6307
rect 215619 6273 215628 6307
rect 215576 6264 215628 6273
rect 215668 6264 215720 6316
rect 88708 6103 88760 6112
rect 88708 6069 88717 6103
rect 88717 6069 88751 6103
rect 88751 6069 88760 6103
rect 88708 6060 88760 6069
rect 170680 6103 170732 6112
rect 170680 6069 170689 6103
rect 170689 6069 170723 6103
rect 170723 6069 170732 6103
rect 170680 6060 170732 6069
rect 221464 6060 221516 6112
rect 225512 6060 225564 6112
rect 142315 5958 142367 6010
rect 142379 5958 142431 6010
rect 142443 5958 142495 6010
rect 142507 5958 142559 6010
rect 283648 5958 283700 6010
rect 283712 5958 283764 6010
rect 283776 5958 283828 6010
rect 283840 5958 283892 6010
rect 215392 5763 215444 5772
rect 215392 5729 215401 5763
rect 215401 5729 215435 5763
rect 215435 5729 215444 5763
rect 215392 5720 215444 5729
rect 217876 5720 217928 5772
rect 215116 5695 215168 5704
rect 215116 5661 215125 5695
rect 215125 5661 215159 5695
rect 215159 5661 215168 5695
rect 215116 5652 215168 5661
rect 217508 5695 217560 5704
rect 217508 5661 217517 5695
rect 217517 5661 217551 5695
rect 217551 5661 217560 5695
rect 217508 5652 217560 5661
rect 216772 5559 216824 5568
rect 216772 5525 216781 5559
rect 216781 5525 216815 5559
rect 216815 5525 216824 5559
rect 216772 5516 216824 5525
rect 217692 5559 217744 5568
rect 217692 5525 217701 5559
rect 217701 5525 217735 5559
rect 217735 5525 217744 5559
rect 217692 5516 217744 5525
rect 223948 5516 224000 5568
rect 423588 5516 423640 5568
rect 71648 5414 71700 5466
rect 71712 5414 71764 5466
rect 71776 5414 71828 5466
rect 71840 5414 71892 5466
rect 212982 5414 213034 5466
rect 213046 5414 213098 5466
rect 213110 5414 213162 5466
rect 213174 5414 213226 5466
rect 354315 5414 354367 5466
rect 354379 5414 354431 5466
rect 354443 5414 354495 5466
rect 354507 5414 354559 5466
rect 215668 5312 215720 5364
rect 217876 5355 217928 5364
rect 217876 5321 217885 5355
rect 217885 5321 217919 5355
rect 217919 5321 217928 5355
rect 217876 5312 217928 5321
rect 221464 5355 221516 5364
rect 221464 5321 221473 5355
rect 221473 5321 221507 5355
rect 221507 5321 221516 5355
rect 221464 5312 221516 5321
rect 223948 5355 224000 5364
rect 223948 5321 223957 5355
rect 223957 5321 223991 5355
rect 223991 5321 224000 5355
rect 223948 5312 224000 5321
rect 209228 5287 209280 5296
rect 209228 5253 209237 5287
rect 209237 5253 209271 5287
rect 209271 5253 209280 5287
rect 209228 5244 209280 5253
rect 212816 5244 212868 5296
rect 214564 5244 214616 5296
rect 216772 5219 216824 5228
rect 216772 5185 216781 5219
rect 216781 5185 216815 5219
rect 216815 5185 216824 5219
rect 216772 5176 216824 5185
rect 209044 5151 209096 5160
rect 209044 5117 209053 5151
rect 209053 5117 209087 5151
rect 209087 5117 209096 5151
rect 209044 5108 209096 5117
rect 212356 5108 212408 5160
rect 216312 5108 216364 5160
rect 224408 5287 224460 5296
rect 224408 5253 224417 5287
rect 224417 5253 224451 5287
rect 224451 5253 224460 5287
rect 224408 5244 224460 5253
rect 220544 5151 220596 5160
rect 220544 5117 220553 5151
rect 220553 5117 220587 5151
rect 220587 5117 220596 5151
rect 220544 5108 220596 5117
rect 224224 5151 224276 5160
rect 224224 5117 224233 5151
rect 224233 5117 224267 5151
rect 224267 5117 224276 5151
rect 224224 5108 224276 5117
rect 212172 5083 212224 5092
rect 212172 5049 212181 5083
rect 212181 5049 212215 5083
rect 212215 5049 212224 5083
rect 212172 5040 212224 5049
rect 214932 5083 214984 5092
rect 214932 5049 214941 5083
rect 214941 5049 214975 5083
rect 214975 5049 214984 5083
rect 214932 5040 214984 5049
rect 216864 5040 216916 5092
rect 217140 5083 217192 5092
rect 217140 5049 217149 5083
rect 217149 5049 217183 5083
rect 217183 5049 217192 5083
rect 217140 5040 217192 5049
rect 93308 5015 93360 5024
rect 93308 4981 93317 5015
rect 93317 4981 93351 5015
rect 93351 4981 93360 5015
rect 93308 4972 93360 4981
rect 93768 5015 93820 5024
rect 93768 4981 93777 5015
rect 93777 4981 93811 5015
rect 93811 4981 93820 5015
rect 93768 4972 93820 4981
rect 208584 5015 208636 5024
rect 208584 4981 208593 5015
rect 208593 4981 208627 5015
rect 208627 4981 208636 5015
rect 208584 4972 208636 4981
rect 216496 4972 216548 5024
rect 218152 5015 218204 5024
rect 218152 4981 218161 5015
rect 218161 4981 218195 5015
rect 218195 4981 218204 5015
rect 218152 4972 218204 4981
rect 220360 5015 220412 5024
rect 220360 4981 220369 5015
rect 220369 4981 220403 5015
rect 220403 4981 220412 5015
rect 220360 4972 220412 4981
rect 142315 4870 142367 4922
rect 142379 4870 142431 4922
rect 142443 4870 142495 4922
rect 142507 4870 142559 4922
rect 283648 4870 283700 4922
rect 283712 4870 283764 4922
rect 283776 4870 283828 4922
rect 283840 4870 283892 4922
rect 209044 4768 209096 4820
rect 213736 4768 213788 4820
rect 215116 4768 215168 4820
rect 220544 4811 220596 4820
rect 214932 4700 214984 4752
rect 220544 4777 220553 4811
rect 220553 4777 220587 4811
rect 220587 4777 220596 4811
rect 220544 4768 220596 4777
rect 224040 4768 224092 4820
rect 224224 4768 224276 4820
rect 217508 4700 217560 4752
rect 218152 4700 218204 4752
rect 218428 4700 218480 4752
rect 220360 4700 220412 4752
rect 213828 4675 213880 4684
rect 213828 4641 213837 4675
rect 213837 4641 213871 4675
rect 213871 4641 213880 4675
rect 213828 4632 213880 4641
rect 214472 4675 214524 4684
rect 214472 4641 214481 4675
rect 214481 4641 214515 4675
rect 214515 4641 214524 4675
rect 214472 4632 214524 4641
rect 216680 4632 216732 4684
rect 214288 4564 214340 4616
rect 218336 4564 218388 4616
rect 212356 4471 212408 4480
rect 212356 4437 212365 4471
rect 212365 4437 212399 4471
rect 212399 4437 212408 4471
rect 212356 4428 212408 4437
rect 212816 4471 212868 4480
rect 212816 4437 212825 4471
rect 212825 4437 212859 4471
rect 212859 4437 212868 4471
rect 212816 4428 212868 4437
rect 215392 4428 215444 4480
rect 216864 4471 216916 4480
rect 216864 4437 216873 4471
rect 216873 4437 216907 4471
rect 216907 4437 216916 4471
rect 216864 4428 216916 4437
rect 220452 4428 220504 4480
rect 71648 4326 71700 4378
rect 71712 4326 71764 4378
rect 71776 4326 71828 4378
rect 71840 4326 71892 4378
rect 212982 4326 213034 4378
rect 213046 4326 213098 4378
rect 213110 4326 213162 4378
rect 213174 4326 213226 4378
rect 354315 4326 354367 4378
rect 354379 4326 354431 4378
rect 354443 4326 354495 4378
rect 354507 4326 354559 4378
rect 214288 4267 214340 4276
rect 214288 4233 214297 4267
rect 214297 4233 214331 4267
rect 214331 4233 214340 4267
rect 214288 4224 214340 4233
rect 214932 4224 214984 4276
rect 218428 4224 218480 4276
rect 215024 4088 215076 4140
rect 214472 4020 214524 4072
rect 216404 4063 216456 4072
rect 212816 3995 212868 4004
rect 212816 3961 212825 3995
rect 212825 3961 212859 3995
rect 212859 3961 212868 3995
rect 212816 3952 212868 3961
rect 213184 3995 213236 4004
rect 213184 3961 213193 3995
rect 213193 3961 213227 3995
rect 213227 3961 213236 3995
rect 213184 3952 213236 3961
rect 213552 3995 213604 4004
rect 213552 3961 213561 3995
rect 213561 3961 213595 3995
rect 213595 3961 213604 3995
rect 213552 3952 213604 3961
rect 215392 3995 215444 4004
rect 215392 3961 215401 3995
rect 215401 3961 215435 3995
rect 215435 3961 215444 3995
rect 215392 3952 215444 3961
rect 212632 3927 212684 3936
rect 212632 3893 212641 3927
rect 212641 3893 212675 3927
rect 212675 3893 212684 3927
rect 212632 3884 212684 3893
rect 213276 3884 213328 3936
rect 213828 3927 213880 3936
rect 213828 3893 213837 3927
rect 213837 3893 213871 3927
rect 213871 3893 213880 3927
rect 213828 3884 213880 3893
rect 214748 3927 214800 3936
rect 214748 3893 214757 3927
rect 214757 3893 214791 3927
rect 214791 3893 214800 3927
rect 214748 3884 214800 3893
rect 216404 4029 216413 4063
rect 216413 4029 216447 4063
rect 216447 4029 216456 4063
rect 216404 4020 216456 4029
rect 216496 4020 216548 4072
rect 217140 4020 217192 4072
rect 217048 3995 217100 4004
rect 217048 3961 217057 3995
rect 217057 3961 217091 3995
rect 217091 3961 217100 3995
rect 217048 3952 217100 3961
rect 217600 3952 217652 4004
rect 218336 3995 218388 4004
rect 218336 3961 218345 3995
rect 218345 3961 218379 3995
rect 218379 3961 218388 3995
rect 218336 3952 218388 3961
rect 217784 3884 217836 3936
rect 142315 3782 142367 3834
rect 142379 3782 142431 3834
rect 142443 3782 142495 3834
rect 142507 3782 142559 3834
rect 283648 3782 283700 3834
rect 283712 3782 283764 3834
rect 283776 3782 283828 3834
rect 283840 3782 283892 3834
rect 212356 3680 212408 3732
rect 212816 3612 212868 3664
rect 213276 3587 213328 3596
rect 213276 3553 213285 3587
rect 213285 3553 213319 3587
rect 213319 3553 213328 3587
rect 213276 3544 213328 3553
rect 213736 3587 213788 3596
rect 213736 3553 213745 3587
rect 213745 3553 213779 3587
rect 213779 3553 213788 3587
rect 213736 3544 213788 3553
rect 214748 3612 214800 3664
rect 216404 3680 216456 3732
rect 216680 3680 216732 3732
rect 224040 3680 224092 3732
rect 216312 3655 216364 3664
rect 214472 3587 214524 3596
rect 214472 3553 214481 3587
rect 214481 3553 214515 3587
rect 214515 3553 214524 3587
rect 215760 3587 215812 3596
rect 214472 3544 214524 3553
rect 215760 3553 215769 3587
rect 215769 3553 215803 3587
rect 215803 3553 215812 3587
rect 215760 3544 215812 3553
rect 216312 3621 216321 3655
rect 216321 3621 216355 3655
rect 216355 3621 216364 3655
rect 216312 3612 216364 3621
rect 220452 3612 220504 3664
rect 211988 3476 212040 3528
rect 215392 3476 215444 3528
rect 213184 3408 213236 3460
rect 213644 3408 213696 3460
rect 216864 3544 216916 3596
rect 217508 3587 217560 3596
rect 217508 3553 217517 3587
rect 217517 3553 217551 3587
rect 217551 3553 217560 3587
rect 217508 3544 217560 3553
rect 217048 3476 217100 3528
rect 219716 3519 219768 3528
rect 219716 3485 219725 3519
rect 219725 3485 219759 3519
rect 219759 3485 219768 3519
rect 219716 3476 219768 3485
rect 215760 3340 215812 3392
rect 217508 3408 217560 3460
rect 217784 3383 217836 3392
rect 217784 3349 217793 3383
rect 217793 3349 217827 3383
rect 217827 3349 217836 3383
rect 217784 3340 217836 3349
rect 71648 3238 71700 3290
rect 71712 3238 71764 3290
rect 71776 3238 71828 3290
rect 71840 3238 71892 3290
rect 212982 3238 213034 3290
rect 213046 3238 213098 3290
rect 213110 3238 213162 3290
rect 213174 3238 213226 3290
rect 354315 3238 354367 3290
rect 354379 3238 354431 3290
rect 354443 3238 354495 3290
rect 354507 3238 354559 3290
rect 211988 3179 212040 3188
rect 211988 3145 211997 3179
rect 211997 3145 212031 3179
rect 212031 3145 212040 3179
rect 211988 3136 212040 3145
rect 212172 3136 212224 3188
rect 212632 3136 212684 3188
rect 214472 3136 214524 3188
rect 214748 3136 214800 3188
rect 215392 3136 215444 3188
rect 217508 3179 217560 3188
rect 217508 3145 217517 3179
rect 217517 3145 217551 3179
rect 217551 3145 217560 3179
rect 217508 3136 217560 3145
rect 208952 3068 209004 3120
rect 214840 3068 214892 3120
rect 213552 3000 213604 3052
rect 214564 2932 214616 2984
rect 216680 3000 216732 3052
rect 216128 2932 216180 2984
rect 216404 2932 216456 2984
rect 220084 2975 220136 2984
rect 212172 2864 212224 2916
rect 214104 2864 214156 2916
rect 220084 2941 220093 2975
rect 220093 2941 220127 2975
rect 220127 2941 220136 2975
rect 220084 2932 220136 2941
rect 217784 2864 217836 2916
rect 213276 2796 213328 2848
rect 218244 2839 218296 2848
rect 218244 2805 218253 2839
rect 218253 2805 218287 2839
rect 218287 2805 218296 2839
rect 218244 2796 218296 2805
rect 220452 2839 220504 2848
rect 220452 2805 220461 2839
rect 220461 2805 220495 2839
rect 220495 2805 220504 2839
rect 220452 2796 220504 2805
rect 221004 2839 221056 2848
rect 221004 2805 221013 2839
rect 221013 2805 221047 2839
rect 221047 2805 221056 2839
rect 221004 2796 221056 2805
rect 142315 2694 142367 2746
rect 142379 2694 142431 2746
rect 142443 2694 142495 2746
rect 142507 2694 142559 2746
rect 283648 2694 283700 2746
rect 283712 2694 283764 2746
rect 283776 2694 283828 2746
rect 283840 2694 283892 2746
rect 209228 2592 209280 2644
rect 213000 2635 213052 2644
rect 213000 2601 213009 2635
rect 213009 2601 213043 2635
rect 213043 2601 213052 2635
rect 213000 2592 213052 2601
rect 214564 2635 214616 2644
rect 214564 2601 214573 2635
rect 214573 2601 214607 2635
rect 214607 2601 214616 2635
rect 214564 2592 214616 2601
rect 214840 2635 214892 2644
rect 214840 2601 214849 2635
rect 214849 2601 214883 2635
rect 214883 2601 214892 2635
rect 214840 2592 214892 2601
rect 213644 2567 213696 2576
rect 213644 2533 213653 2567
rect 213653 2533 213687 2567
rect 213687 2533 213696 2567
rect 213644 2524 213696 2533
rect 213276 2499 213328 2508
rect 213276 2465 213285 2499
rect 213285 2465 213319 2499
rect 213319 2465 213328 2499
rect 213276 2456 213328 2465
rect 214104 2524 214156 2576
rect 214288 2524 214340 2576
rect 216772 2592 216824 2644
rect 215760 2524 215812 2576
rect 213736 2388 213788 2440
rect 216128 2456 216180 2508
rect 216312 2456 216364 2508
rect 217600 2524 217652 2576
rect 218244 2592 218296 2644
rect 219716 2635 219768 2644
rect 219716 2601 219725 2635
rect 219725 2601 219759 2635
rect 219759 2601 219768 2635
rect 219716 2592 219768 2601
rect 220084 2635 220136 2644
rect 220084 2601 220093 2635
rect 220093 2601 220127 2635
rect 220127 2601 220136 2635
rect 220084 2592 220136 2601
rect 220544 2635 220596 2644
rect 220544 2601 220553 2635
rect 220553 2601 220587 2635
rect 220587 2601 220596 2635
rect 220544 2592 220596 2601
rect 221924 2635 221976 2644
rect 221924 2601 221933 2635
rect 221933 2601 221967 2635
rect 221967 2601 221976 2635
rect 221924 2592 221976 2601
rect 224408 2456 224460 2508
rect 350816 2499 350868 2508
rect 350816 2465 350825 2499
rect 350825 2465 350859 2499
rect 350859 2465 350868 2499
rect 350816 2456 350868 2465
rect 308588 2431 308640 2440
rect 212448 2295 212500 2304
rect 212448 2261 212457 2295
rect 212457 2261 212491 2295
rect 212491 2261 212500 2295
rect 212448 2252 212500 2261
rect 221188 2295 221240 2304
rect 221188 2261 221197 2295
rect 221197 2261 221231 2295
rect 221231 2261 221240 2295
rect 308588 2397 308597 2431
rect 308597 2397 308631 2431
rect 308631 2397 308640 2431
rect 308588 2388 308640 2397
rect 309876 2363 309928 2372
rect 228364 2295 228416 2304
rect 221188 2252 221240 2261
rect 228364 2261 228373 2295
rect 228373 2261 228407 2295
rect 228407 2261 228416 2295
rect 228364 2252 228416 2261
rect 309876 2329 309885 2363
rect 309885 2329 309919 2363
rect 309919 2329 309928 2363
rect 309876 2320 309928 2329
rect 318064 2252 318116 2304
rect 351000 2295 351052 2304
rect 351000 2261 351009 2295
rect 351009 2261 351043 2295
rect 351043 2261 351052 2295
rect 351000 2252 351052 2261
rect 71648 2150 71700 2202
rect 71712 2150 71764 2202
rect 71776 2150 71828 2202
rect 71840 2150 71892 2202
rect 212982 2150 213034 2202
rect 213046 2150 213098 2202
rect 213110 2150 213162 2202
rect 213174 2150 213226 2202
rect 354315 2150 354367 2202
rect 354379 2150 354431 2202
rect 354443 2150 354495 2202
rect 354507 2150 354559 2202
<< metal2 >>
rect 35346 9602 35402 10000
rect 106002 9602 106058 10000
rect 176658 9602 176714 10000
rect 35346 9574 35664 9602
rect 35346 9520 35402 9574
rect 110 9344 166 9353
rect 110 9279 166 9288
rect 124 8226 152 9279
rect 112 8220 164 8226
rect 112 8162 164 8168
rect 18 8120 74 8129
rect 18 8055 74 8064
rect 32 4729 60 8055
rect 35636 6905 35664 9574
rect 106002 9574 106136 9602
rect 106002 9520 106058 9574
rect 71622 7644 71918 7664
rect 71678 7642 71702 7644
rect 71758 7642 71782 7644
rect 71838 7642 71862 7644
rect 71700 7590 71702 7642
rect 71764 7590 71776 7642
rect 71838 7590 71840 7642
rect 71678 7588 71702 7590
rect 71758 7588 71782 7590
rect 71838 7588 71862 7590
rect 71622 7568 71918 7588
rect 88616 7336 88668 7342
rect 88616 7278 88668 7284
rect 110 6896 166 6905
rect 110 6831 166 6840
rect 35622 6896 35678 6905
rect 35622 6831 35678 6840
rect 74998 6896 75054 6905
rect 74998 6831 75054 6840
rect 124 5273 152 6831
rect 75012 6798 75040 6831
rect 75000 6792 75052 6798
rect 75000 6734 75052 6740
rect 88248 6792 88300 6798
rect 88248 6734 88300 6740
rect 71622 6556 71918 6576
rect 71678 6554 71702 6556
rect 71758 6554 71782 6556
rect 71838 6554 71862 6556
rect 71700 6502 71702 6554
rect 71764 6502 71776 6554
rect 71838 6502 71840 6554
rect 71678 6500 71702 6502
rect 71758 6500 71782 6502
rect 71838 6500 71862 6502
rect 71622 6480 71918 6500
rect 88260 6458 88288 6734
rect 88628 6662 88656 7278
rect 106108 7274 106136 9574
rect 176304 9574 176714 9602
rect 106096 7268 106148 7274
rect 106096 7210 106148 7216
rect 142289 7100 142585 7120
rect 142345 7098 142369 7100
rect 142425 7098 142449 7100
rect 142505 7098 142529 7100
rect 142367 7046 142369 7098
rect 142431 7046 142443 7098
rect 142505 7046 142507 7098
rect 142345 7044 142369 7046
rect 142425 7044 142449 7046
rect 142505 7044 142529 7046
rect 142289 7024 142585 7044
rect 176304 7002 176332 9574
rect 176658 9520 176714 9574
rect 247314 9602 247370 10000
rect 317970 9602 318026 10000
rect 388626 9602 388682 10000
rect 247314 9574 247448 9602
rect 247314 9520 247370 9574
rect 178224 8220 178276 8226
rect 178224 8162 178276 8168
rect 178236 7546 178264 8162
rect 212956 7644 213252 7664
rect 213012 7642 213036 7644
rect 213092 7642 213116 7644
rect 213172 7642 213196 7644
rect 213034 7590 213036 7642
rect 213098 7590 213110 7642
rect 213172 7590 213174 7642
rect 213012 7588 213036 7590
rect 213092 7588 213116 7590
rect 213172 7588 213196 7590
rect 212956 7568 213252 7588
rect 178224 7540 178276 7546
rect 178224 7482 178276 7488
rect 225696 7336 225748 7342
rect 225696 7278 225748 7284
rect 190644 7200 190696 7206
rect 190644 7142 190696 7148
rect 176292 6996 176344 7002
rect 176292 6938 176344 6944
rect 170680 6860 170732 6866
rect 170680 6802 170732 6808
rect 88708 6792 88760 6798
rect 88708 6734 88760 6740
rect 88616 6656 88668 6662
rect 88616 6598 88668 6604
rect 88248 6452 88300 6458
rect 88248 6394 88300 6400
rect 71622 5468 71918 5488
rect 71678 5466 71702 5468
rect 71758 5466 71782 5468
rect 71838 5466 71862 5468
rect 71700 5414 71702 5466
rect 71764 5414 71776 5466
rect 71838 5414 71840 5466
rect 71678 5412 71702 5414
rect 71758 5412 71782 5414
rect 71838 5412 71862 5414
rect 71622 5392 71918 5412
rect 110 5264 166 5273
rect 110 5199 166 5208
rect 18 4720 74 4729
rect 18 4655 74 4664
rect 71622 4380 71918 4400
rect 71678 4378 71702 4380
rect 71758 4378 71782 4380
rect 71838 4378 71862 4380
rect 71700 4326 71702 4378
rect 71764 4326 71776 4378
rect 71838 4326 71840 4378
rect 71678 4324 71702 4326
rect 71758 4324 71782 4326
rect 71838 4324 71862 4326
rect 71622 4304 71918 4324
rect 88628 4185 88656 6598
rect 88720 6118 88748 6734
rect 170692 6118 170720 6802
rect 88708 6112 88760 6118
rect 88708 6054 88760 6060
rect 170680 6112 170732 6118
rect 170680 6054 170732 6060
rect 88720 5409 88748 6054
rect 142289 6012 142585 6032
rect 142345 6010 142369 6012
rect 142425 6010 142449 6012
rect 142505 6010 142529 6012
rect 142367 5958 142369 6010
rect 142431 5958 142443 6010
rect 142505 5958 142507 6010
rect 142345 5956 142369 5958
rect 142425 5956 142449 5958
rect 142505 5956 142529 5958
rect 142289 5936 142585 5956
rect 88706 5400 88762 5409
rect 88706 5335 88762 5344
rect 170692 5273 170720 6054
rect 170678 5264 170734 5273
rect 170678 5199 170734 5208
rect 190656 5137 190684 7142
rect 225326 6896 225382 6905
rect 225326 6831 225382 6840
rect 225340 6798 225368 6831
rect 225328 6792 225380 6798
rect 225328 6734 225380 6740
rect 225512 6792 225564 6798
rect 225512 6734 225564 6740
rect 215668 6656 215720 6662
rect 215668 6598 215720 6604
rect 212956 6556 213252 6576
rect 213012 6554 213036 6556
rect 213092 6554 213116 6556
rect 213172 6554 213196 6556
rect 213034 6502 213036 6554
rect 213098 6502 213110 6554
rect 213172 6502 213174 6554
rect 213012 6500 213036 6502
rect 213092 6500 213116 6502
rect 213172 6500 213196 6502
rect 212956 6480 213252 6500
rect 215680 6322 215708 6598
rect 225340 6458 225368 6734
rect 225328 6452 225380 6458
rect 225328 6394 225380 6400
rect 215944 6384 215996 6390
rect 215944 6326 215996 6332
rect 215576 6316 215628 6322
rect 215576 6258 215628 6264
rect 215668 6316 215720 6322
rect 215668 6258 215720 6264
rect 215588 6225 215616 6258
rect 215574 6216 215630 6225
rect 215574 6151 215630 6160
rect 215392 5772 215444 5778
rect 215392 5714 215444 5720
rect 215116 5704 215168 5710
rect 215116 5646 215168 5652
rect 212956 5468 213252 5488
rect 213012 5466 213036 5468
rect 213092 5466 213116 5468
rect 213172 5466 213196 5468
rect 213034 5414 213036 5466
rect 213098 5414 213110 5466
rect 213172 5414 213174 5466
rect 213012 5412 213036 5414
rect 213092 5412 213116 5414
rect 213172 5412 213196 5414
rect 212814 5400 212870 5409
rect 212956 5392 213252 5412
rect 212814 5335 212870 5344
rect 212828 5302 212856 5335
rect 209228 5296 209280 5302
rect 209228 5238 209280 5244
rect 212816 5296 212868 5302
rect 212816 5238 212868 5244
rect 214564 5296 214616 5302
rect 214564 5238 214616 5244
rect 209044 5160 209096 5166
rect 93306 5128 93362 5137
rect 93306 5063 93362 5072
rect 190642 5128 190698 5137
rect 209044 5102 209096 5108
rect 190642 5063 190698 5072
rect 93320 5030 93348 5063
rect 93308 5024 93360 5030
rect 93308 4966 93360 4972
rect 93768 5024 93820 5030
rect 93768 4966 93820 4972
rect 88614 4176 88670 4185
rect 88614 4111 88670 4120
rect 93780 4049 93808 4966
rect 142289 4924 142585 4944
rect 142345 4922 142369 4924
rect 142425 4922 142449 4924
rect 142505 4922 142529 4924
rect 142367 4870 142369 4922
rect 142431 4870 142443 4922
rect 142505 4870 142507 4922
rect 142345 4868 142369 4870
rect 142425 4868 142449 4870
rect 142505 4868 142529 4870
rect 142289 4848 142585 4868
rect 93766 4040 93822 4049
rect 93766 3975 93822 3984
rect 105634 4040 105690 4049
rect 105634 3975 105690 3984
rect 105648 3505 105676 3975
rect 142289 3836 142585 3856
rect 142345 3834 142369 3836
rect 142425 3834 142449 3836
rect 142505 3834 142529 3836
rect 142367 3782 142369 3834
rect 142431 3782 142443 3834
rect 142505 3782 142507 3834
rect 142345 3780 142369 3782
rect 142425 3780 142449 3782
rect 142505 3780 142529 3782
rect 142289 3760 142585 3780
rect 105634 3496 105690 3505
rect 105634 3431 105690 3440
rect 71622 3292 71918 3312
rect 71678 3290 71702 3292
rect 71758 3290 71782 3292
rect 71838 3290 71862 3292
rect 71700 3238 71702 3290
rect 71764 3238 71776 3290
rect 71838 3238 71840 3290
rect 71678 3236 71702 3238
rect 71758 3236 71782 3238
rect 71838 3236 71862 3238
rect 71622 3216 71918 3236
rect 63774 2952 63830 2961
rect 63774 2887 63830 2896
rect 21454 1456 21510 1465
rect 21454 1391 21510 1400
rect 21178 82 21234 480
rect 21468 82 21496 1391
rect 21178 54 21496 82
rect 63498 82 63554 480
rect 63788 82 63816 2887
rect 71622 2204 71918 2224
rect 71678 2202 71702 2204
rect 71758 2202 71782 2204
rect 71838 2202 71862 2204
rect 71700 2150 71702 2202
rect 71764 2150 71776 2202
rect 71838 2150 71840 2202
rect 71678 2148 71702 2150
rect 71758 2148 71782 2150
rect 71838 2148 71862 2150
rect 71622 2128 71918 2148
rect 63498 54 63816 82
rect 105648 82 105676 3431
rect 148598 3088 148654 3097
rect 148598 3023 148654 3032
rect 142289 2748 142585 2768
rect 142345 2746 142369 2748
rect 142425 2746 142449 2748
rect 142505 2746 142529 2748
rect 142367 2694 142369 2746
rect 142431 2694 142443 2746
rect 142505 2694 142507 2746
rect 142345 2692 142369 2694
rect 142425 2692 142449 2694
rect 142505 2692 142529 2694
rect 142289 2672 142585 2692
rect 105910 82 105966 480
rect 105648 54 105966 82
rect 21178 0 21234 54
rect 63498 0 63554 54
rect 105910 0 105966 54
rect 148322 82 148378 480
rect 148612 82 148640 3023
rect 148322 54 148640 82
rect 190656 82 190684 5063
rect 208584 5024 208636 5030
rect 208584 4966 208636 4972
rect 208596 4729 208624 4966
rect 209056 4826 209084 5102
rect 209044 4820 209096 4826
rect 209044 4762 209096 4768
rect 208582 4720 208638 4729
rect 208582 4655 208638 4664
rect 209056 4154 209084 4762
rect 208964 4126 209084 4154
rect 208964 3126 208992 4126
rect 208952 3120 209004 3126
rect 209240 3097 209268 5238
rect 212356 5160 212408 5166
rect 212356 5102 212408 5108
rect 212172 5092 212224 5098
rect 212172 5034 212224 5040
rect 211988 3528 212040 3534
rect 211988 3470 212040 3476
rect 212000 3194 212028 3470
rect 212184 3194 212212 5034
rect 212368 4486 212396 5102
rect 213736 4820 213788 4826
rect 213736 4762 213788 4768
rect 212356 4480 212408 4486
rect 212356 4422 212408 4428
rect 212816 4480 212868 4486
rect 212816 4422 212868 4428
rect 212368 3738 212396 4422
rect 212630 4040 212686 4049
rect 212828 4010 212856 4422
rect 212956 4380 213252 4400
rect 213012 4378 213036 4380
rect 213092 4378 213116 4380
rect 213172 4378 213196 4380
rect 213034 4326 213036 4378
rect 213098 4326 213110 4378
rect 213172 4326 213174 4378
rect 213012 4324 213036 4326
rect 213092 4324 213116 4326
rect 213172 4324 213196 4326
rect 212956 4304 213252 4324
rect 212630 3975 212686 3984
rect 212816 4004 212868 4010
rect 212644 3942 212672 3975
rect 212816 3946 212868 3952
rect 213184 4004 213236 4010
rect 213184 3946 213236 3952
rect 213552 4004 213604 4010
rect 213552 3946 213604 3952
rect 212632 3936 212684 3942
rect 212632 3878 212684 3884
rect 212356 3732 212408 3738
rect 212356 3674 212408 3680
rect 212644 3194 212672 3878
rect 212828 3670 212856 3946
rect 212816 3664 212868 3670
rect 212816 3606 212868 3612
rect 213196 3466 213224 3946
rect 213276 3936 213328 3942
rect 213276 3878 213328 3884
rect 213288 3602 213316 3878
rect 213276 3596 213328 3602
rect 213276 3538 213328 3544
rect 213184 3460 213236 3466
rect 213184 3402 213236 3408
rect 212956 3292 213252 3312
rect 213012 3290 213036 3292
rect 213092 3290 213116 3292
rect 213172 3290 213196 3292
rect 213034 3238 213036 3290
rect 213098 3238 213110 3290
rect 213172 3238 213174 3290
rect 213012 3236 213036 3238
rect 213092 3236 213116 3238
rect 213172 3236 213196 3238
rect 212956 3216 213252 3236
rect 211988 3188 212040 3194
rect 211988 3130 212040 3136
rect 212172 3188 212224 3194
rect 212172 3130 212224 3136
rect 212632 3188 212684 3194
rect 212632 3130 212684 3136
rect 208952 3062 209004 3068
rect 209226 3088 209282 3097
rect 209226 3023 209282 3032
rect 209240 2650 209268 3023
rect 212184 2922 212212 3130
rect 212172 2916 212224 2922
rect 212172 2858 212224 2864
rect 213288 2854 213316 3538
rect 213564 3058 213592 3946
rect 213748 3602 213776 4762
rect 213828 4684 213880 4690
rect 213828 4626 213880 4632
rect 214472 4684 214524 4690
rect 214472 4626 214524 4632
rect 213840 3942 213868 4626
rect 214288 4616 214340 4622
rect 214288 4558 214340 4564
rect 214300 4282 214328 4558
rect 214288 4276 214340 4282
rect 214288 4218 214340 4224
rect 213828 3936 213880 3942
rect 213828 3878 213880 3884
rect 213736 3596 213788 3602
rect 213736 3538 213788 3544
rect 213644 3460 213696 3466
rect 213644 3402 213696 3408
rect 213552 3052 213604 3058
rect 213552 2994 213604 3000
rect 213276 2848 213328 2854
rect 213276 2790 213328 2796
rect 209228 2644 209280 2650
rect 209228 2586 209280 2592
rect 213000 2644 213052 2650
rect 213000 2586 213052 2592
rect 213012 2553 213040 2586
rect 200946 2544 201002 2553
rect 200946 2479 201002 2488
rect 212998 2544 213054 2553
rect 213288 2514 213316 2790
rect 213656 2582 213684 3402
rect 213644 2576 213696 2582
rect 213644 2518 213696 2524
rect 212998 2479 213054 2488
rect 213276 2508 213328 2514
rect 200960 1465 200988 2479
rect 213276 2450 213328 2456
rect 213288 2417 213316 2450
rect 213748 2446 213776 3538
rect 214104 2916 214156 2922
rect 214104 2858 214156 2864
rect 214116 2582 214144 2858
rect 214300 2582 214328 4218
rect 214484 4078 214512 4626
rect 214472 4072 214524 4078
rect 214472 4014 214524 4020
rect 214472 3596 214524 3602
rect 214472 3538 214524 3544
rect 214484 3194 214512 3538
rect 214472 3188 214524 3194
rect 214472 3130 214524 3136
rect 214576 2990 214604 5238
rect 214932 5092 214984 5098
rect 214932 5034 214984 5040
rect 214944 4758 214972 5034
rect 215128 4826 215156 5646
rect 215116 4820 215168 4826
rect 215116 4762 215168 4768
rect 214932 4752 214984 4758
rect 214932 4694 214984 4700
rect 214944 4282 214972 4694
rect 214932 4276 214984 4282
rect 214932 4218 214984 4224
rect 215128 4154 215156 4762
rect 215404 4486 215432 5714
rect 215680 5370 215708 6258
rect 215668 5364 215720 5370
rect 215668 5306 215720 5312
rect 215956 5137 215984 6326
rect 225524 6118 225552 6734
rect 225708 6662 225736 7278
rect 229560 7200 229612 7206
rect 229560 7142 229612 7148
rect 229572 6769 229600 7142
rect 247420 6905 247448 9574
rect 317970 9574 318104 9602
rect 317970 9520 318026 9574
rect 283622 7100 283918 7120
rect 283678 7098 283702 7100
rect 283758 7098 283782 7100
rect 283838 7098 283862 7100
rect 283700 7046 283702 7098
rect 283764 7046 283776 7098
rect 283838 7046 283840 7098
rect 283678 7044 283702 7046
rect 283758 7044 283782 7046
rect 283838 7044 283862 7046
rect 283622 7024 283918 7044
rect 247406 6896 247462 6905
rect 247406 6831 247462 6840
rect 318076 6769 318104 9574
rect 388626 9574 388760 9602
rect 388626 9520 388682 9574
rect 354289 7644 354585 7664
rect 354345 7642 354369 7644
rect 354425 7642 354449 7644
rect 354505 7642 354529 7644
rect 354367 7590 354369 7642
rect 354431 7590 354443 7642
rect 354505 7590 354507 7642
rect 354345 7588 354369 7590
rect 354425 7588 354449 7590
rect 354505 7588 354529 7590
rect 354289 7568 354585 7588
rect 229558 6760 229614 6769
rect 229558 6695 229614 6704
rect 318062 6760 318118 6769
rect 318062 6695 318118 6704
rect 225696 6656 225748 6662
rect 225696 6598 225748 6604
rect 225708 6361 225736 6598
rect 354289 6556 354585 6576
rect 354345 6554 354369 6556
rect 354425 6554 354449 6556
rect 354505 6554 354529 6556
rect 354367 6502 354369 6554
rect 354431 6502 354443 6554
rect 354505 6502 354507 6554
rect 354345 6500 354369 6502
rect 354425 6500 354449 6502
rect 354505 6500 354529 6502
rect 354289 6480 354585 6500
rect 225694 6352 225750 6361
rect 225694 6287 225750 6296
rect 388732 6225 388760 9574
rect 423586 9208 423642 9217
rect 423416 9166 423586 9194
rect 388718 6216 388774 6225
rect 388718 6151 388774 6160
rect 221464 6112 221516 6118
rect 221464 6054 221516 6060
rect 225512 6112 225564 6118
rect 225512 6054 225564 6060
rect 217874 5808 217930 5817
rect 217874 5743 217876 5752
rect 217928 5743 217930 5752
rect 217876 5714 217928 5720
rect 217508 5704 217560 5710
rect 217508 5646 217560 5652
rect 216772 5568 216824 5574
rect 216772 5510 216824 5516
rect 216784 5234 216812 5510
rect 216772 5228 216824 5234
rect 216692 5188 216772 5216
rect 216312 5160 216364 5166
rect 215942 5128 215998 5137
rect 216312 5102 216364 5108
rect 215942 5063 215998 5072
rect 215392 4480 215444 4486
rect 215392 4422 215444 4428
rect 215036 4146 215156 4154
rect 215024 4140 215156 4146
rect 215076 4126 215156 4140
rect 215024 4082 215076 4088
rect 215392 4004 215444 4010
rect 215392 3946 215444 3952
rect 214748 3936 214800 3942
rect 214748 3878 214800 3884
rect 214760 3670 214788 3878
rect 214748 3664 214800 3670
rect 214748 3606 214800 3612
rect 214760 3194 214788 3606
rect 215404 3534 215432 3946
rect 216324 3670 216352 5102
rect 216496 5024 216548 5030
rect 216496 4966 216548 4972
rect 216508 4078 216536 4966
rect 216692 4690 216720 5188
rect 216772 5170 216824 5176
rect 216864 5092 216916 5098
rect 216864 5034 216916 5040
rect 217140 5092 217192 5098
rect 217140 5034 217192 5040
rect 216680 4684 216732 4690
rect 216680 4626 216732 4632
rect 216404 4072 216456 4078
rect 216404 4014 216456 4020
rect 216496 4072 216548 4078
rect 216496 4014 216548 4020
rect 216416 3738 216444 4014
rect 216692 3738 216720 4626
rect 216876 4486 216904 5034
rect 216864 4480 216916 4486
rect 216864 4422 216916 4428
rect 216404 3732 216456 3738
rect 216404 3674 216456 3680
rect 216680 3732 216732 3738
rect 216680 3674 216732 3680
rect 216312 3664 216364 3670
rect 216312 3606 216364 3612
rect 215760 3596 215812 3602
rect 215760 3538 215812 3544
rect 215392 3528 215444 3534
rect 215392 3470 215444 3476
rect 215404 3194 215432 3470
rect 215772 3398 215800 3538
rect 215760 3392 215812 3398
rect 215760 3334 215812 3340
rect 214748 3188 214800 3194
rect 214748 3130 214800 3136
rect 215392 3188 215444 3194
rect 215392 3130 215444 3136
rect 214840 3120 214892 3126
rect 214840 3062 214892 3068
rect 214564 2984 214616 2990
rect 214564 2926 214616 2932
rect 214576 2650 214604 2926
rect 214852 2650 214880 3062
rect 214564 2644 214616 2650
rect 214564 2586 214616 2592
rect 214840 2644 214892 2650
rect 214840 2586 214892 2592
rect 215772 2582 215800 3334
rect 216416 2990 216444 3674
rect 216692 3058 216720 3674
rect 216876 3602 216904 4422
rect 217152 4078 217180 5034
rect 217520 4758 217548 5646
rect 217692 5568 217744 5574
rect 217692 5510 217744 5516
rect 217508 4752 217560 4758
rect 217508 4694 217560 4700
rect 217140 4072 217192 4078
rect 217140 4014 217192 4020
rect 217048 4004 217100 4010
rect 217048 3946 217100 3952
rect 217600 4004 217652 4010
rect 217600 3946 217652 3952
rect 216864 3596 216916 3602
rect 216864 3538 216916 3544
rect 216680 3052 216732 3058
rect 216680 2994 216732 3000
rect 216128 2984 216180 2990
rect 216128 2926 216180 2932
rect 216404 2984 216456 2990
rect 216404 2926 216456 2932
rect 214104 2576 214156 2582
rect 214104 2518 214156 2524
rect 214288 2576 214340 2582
rect 214288 2518 214340 2524
rect 215760 2576 215812 2582
rect 215760 2518 215812 2524
rect 216140 2514 216168 2926
rect 216128 2508 216180 2514
rect 216128 2450 216180 2456
rect 216312 2508 216364 2514
rect 216416 2496 216444 2926
rect 216692 2632 216720 2994
rect 216772 2644 216824 2650
rect 216692 2604 216772 2632
rect 216772 2586 216824 2592
rect 216364 2468 216444 2496
rect 216312 2450 216364 2456
rect 213736 2440 213788 2446
rect 213274 2408 213330 2417
rect 213736 2382 213788 2388
rect 213274 2343 213330 2352
rect 212448 2304 212500 2310
rect 212448 2246 212500 2252
rect 200946 1456 201002 1465
rect 200946 1391 201002 1400
rect 212460 921 212488 2246
rect 212956 2204 213252 2224
rect 213012 2202 213036 2204
rect 213092 2202 213116 2204
rect 213172 2202 213196 2204
rect 213034 2150 213036 2202
rect 213098 2150 213110 2202
rect 213172 2150 213174 2202
rect 213012 2148 213036 2150
rect 213092 2148 213116 2150
rect 213172 2148 213196 2150
rect 212956 2128 213252 2148
rect 212446 912 212502 921
rect 212446 847 212502 856
rect 190734 82 190790 480
rect 216876 241 216904 3538
rect 217060 3534 217088 3946
rect 217508 3596 217560 3602
rect 217508 3538 217560 3544
rect 217048 3528 217100 3534
rect 217048 3470 217100 3476
rect 217520 3466 217548 3538
rect 217508 3460 217560 3466
rect 217508 3402 217560 3408
rect 217520 3194 217548 3402
rect 217508 3188 217560 3194
rect 217508 3130 217560 3136
rect 217612 2582 217640 3946
rect 217704 3505 217732 5510
rect 217888 5370 217916 5714
rect 221476 5370 221504 6054
rect 283622 6012 283918 6032
rect 283678 6010 283702 6012
rect 283758 6010 283782 6012
rect 283838 6010 283862 6012
rect 283700 5958 283702 6010
rect 283764 5958 283776 6010
rect 283838 5958 283840 6010
rect 283678 5956 283702 5958
rect 283758 5956 283782 5958
rect 283838 5956 283862 5958
rect 283622 5936 283918 5956
rect 423416 5817 423444 9166
rect 423586 9143 423642 9152
rect 423586 7576 423642 7585
rect 423586 7511 423642 7520
rect 423402 5808 423458 5817
rect 423402 5743 423458 5752
rect 423600 5574 423628 7511
rect 423678 5944 423734 5953
rect 423678 5879 423734 5888
rect 223948 5568 224000 5574
rect 223948 5510 224000 5516
rect 423588 5568 423640 5574
rect 423588 5510 423640 5516
rect 223960 5370 223988 5510
rect 354289 5468 354585 5488
rect 354345 5466 354369 5468
rect 354425 5466 354449 5468
rect 354505 5466 354529 5468
rect 354367 5414 354369 5466
rect 354431 5414 354443 5466
rect 354505 5414 354507 5466
rect 354345 5412 354369 5414
rect 354425 5412 354449 5414
rect 354505 5412 354529 5414
rect 354289 5392 354585 5412
rect 217876 5364 217928 5370
rect 217876 5306 217928 5312
rect 221464 5364 221516 5370
rect 221464 5306 221516 5312
rect 223948 5364 224000 5370
rect 223948 5306 224000 5312
rect 224408 5296 224460 5302
rect 221922 5264 221978 5273
rect 224408 5238 224460 5244
rect 221922 5199 221978 5208
rect 220544 5160 220596 5166
rect 220544 5102 220596 5108
rect 218152 5024 218204 5030
rect 218152 4966 218204 4972
rect 220360 5024 220412 5030
rect 220360 4966 220412 4972
rect 218164 4758 218192 4966
rect 220372 4758 220400 4966
rect 220556 4826 220584 5102
rect 220544 4820 220596 4826
rect 220544 4762 220596 4768
rect 218152 4752 218204 4758
rect 218152 4694 218204 4700
rect 218428 4752 218480 4758
rect 218428 4694 218480 4700
rect 220360 4752 220412 4758
rect 220360 4694 220412 4700
rect 218336 4616 218388 4622
rect 218336 4558 218388 4564
rect 218348 4010 218376 4558
rect 218440 4282 218468 4694
rect 218428 4276 218480 4282
rect 218428 4218 218480 4224
rect 218336 4004 218388 4010
rect 218336 3946 218388 3952
rect 217784 3936 217836 3942
rect 217784 3878 217836 3884
rect 217690 3496 217746 3505
rect 217690 3431 217746 3440
rect 217796 3398 217824 3878
rect 220372 3652 220400 4694
rect 220452 4480 220504 4486
rect 220504 4440 220584 4468
rect 220452 4422 220504 4428
rect 220452 3664 220504 3670
rect 220372 3624 220452 3652
rect 220452 3606 220504 3612
rect 219716 3528 219768 3534
rect 219716 3470 219768 3476
rect 217784 3392 217836 3398
rect 217784 3334 217836 3340
rect 217796 2922 217824 3334
rect 217784 2916 217836 2922
rect 217784 2858 217836 2864
rect 218244 2848 218296 2854
rect 218244 2790 218296 2796
rect 218256 2650 218284 2790
rect 219728 2650 219756 3470
rect 220084 2984 220136 2990
rect 220084 2926 220136 2932
rect 220096 2650 220124 2926
rect 220464 2854 220492 3606
rect 220452 2848 220504 2854
rect 220452 2790 220504 2796
rect 218244 2644 218296 2650
rect 218244 2586 218296 2592
rect 219716 2644 219768 2650
rect 219716 2586 219768 2592
rect 220084 2644 220136 2650
rect 220084 2586 220136 2592
rect 217600 2576 217652 2582
rect 217600 2518 217652 2524
rect 220464 1465 220492 2790
rect 220556 2650 220584 4440
rect 221936 4185 221964 5199
rect 224224 5160 224276 5166
rect 224224 5102 224276 5108
rect 224236 4826 224264 5102
rect 224040 4820 224092 4826
rect 224040 4762 224092 4768
rect 224224 4820 224276 4826
rect 224224 4762 224276 4768
rect 221922 4176 221978 4185
rect 221922 4111 221978 4120
rect 221004 2848 221056 2854
rect 221004 2790 221056 2796
rect 220544 2644 220596 2650
rect 220544 2586 220596 2592
rect 221016 2553 221044 2790
rect 221936 2650 221964 4111
rect 224052 3738 224080 4762
rect 224040 3732 224092 3738
rect 224040 3674 224092 3680
rect 224420 2961 224448 5238
rect 283622 4924 283918 4944
rect 283678 4922 283702 4924
rect 283758 4922 283782 4924
rect 283838 4922 283862 4924
rect 283700 4870 283702 4922
rect 283764 4870 283776 4922
rect 283838 4870 283840 4922
rect 283678 4868 283702 4870
rect 283758 4868 283782 4870
rect 283838 4868 283862 4870
rect 283622 4848 283918 4868
rect 354289 4380 354585 4400
rect 354345 4378 354369 4380
rect 354425 4378 354449 4380
rect 354505 4378 354529 4380
rect 354367 4326 354369 4378
rect 354431 4326 354443 4378
rect 354505 4326 354507 4378
rect 354345 4324 354369 4326
rect 354425 4324 354449 4326
rect 354505 4324 354529 4326
rect 354289 4304 354585 4324
rect 283622 3836 283918 3856
rect 283678 3834 283702 3836
rect 283758 3834 283782 3836
rect 283838 3834 283862 3836
rect 283700 3782 283702 3834
rect 283764 3782 283776 3834
rect 283838 3782 283840 3834
rect 283678 3780 283702 3782
rect 283758 3780 283782 3782
rect 283838 3780 283862 3782
rect 283622 3760 283918 3780
rect 354289 3292 354585 3312
rect 354345 3290 354369 3292
rect 354425 3290 354449 3292
rect 354505 3290 354529 3292
rect 354367 3238 354369 3290
rect 354431 3238 354443 3290
rect 354505 3238 354507 3290
rect 354345 3236 354369 3238
rect 354425 3236 354449 3238
rect 354505 3236 354529 3238
rect 354289 3216 354585 3236
rect 224406 2952 224462 2961
rect 224406 2887 224462 2896
rect 221924 2644 221976 2650
rect 221924 2586 221976 2592
rect 221002 2544 221058 2553
rect 224420 2514 224448 2887
rect 423692 2825 423720 5879
rect 423678 2816 423734 2825
rect 283622 2748 283918 2768
rect 423678 2751 423734 2760
rect 283678 2746 283702 2748
rect 283758 2746 283782 2748
rect 283838 2746 283862 2748
rect 283700 2694 283702 2746
rect 283764 2694 283776 2746
rect 283838 2694 283840 2746
rect 283678 2692 283702 2694
rect 283758 2692 283782 2694
rect 283838 2692 283862 2694
rect 283622 2672 283918 2692
rect 308586 2544 308642 2553
rect 221002 2479 221058 2488
rect 224408 2508 224460 2514
rect 423586 2544 423642 2553
rect 308586 2479 308642 2488
rect 350816 2508 350868 2514
rect 224408 2450 224460 2456
rect 308600 2446 308628 2479
rect 423586 2479 423642 2488
rect 350816 2450 350868 2456
rect 308588 2440 308640 2446
rect 350828 2417 350856 2450
rect 309966 2408 310022 2417
rect 308588 2382 308640 2388
rect 309888 2378 309966 2394
rect 309876 2372 309966 2378
rect 309928 2366 309966 2372
rect 309966 2343 310022 2352
rect 350814 2408 350870 2417
rect 350814 2343 350870 2352
rect 309876 2314 309928 2320
rect 221188 2304 221240 2310
rect 221188 2246 221240 2252
rect 228364 2304 228416 2310
rect 228364 2246 228416 2252
rect 318064 2304 318116 2310
rect 318064 2246 318116 2252
rect 351000 2304 351052 2310
rect 351000 2246 351052 2252
rect 220450 1456 220506 1465
rect 220450 1391 220506 1400
rect 216862 232 216918 241
rect 216862 167 216918 176
rect 221200 105 221228 2246
rect 228376 1193 228404 2246
rect 228362 1184 228418 1193
rect 228362 1119 228418 1128
rect 275282 1184 275338 1193
rect 275282 1119 275338 1128
rect 190656 54 190790 82
rect 148322 0 148378 54
rect 190734 0 190790 54
rect 221186 96 221242 105
rect 221186 31 221242 40
rect 233146 96 233202 480
rect 275296 82 275324 1119
rect 275558 82 275614 480
rect 275296 54 275614 82
rect 233146 0 233202 40
rect 275558 0 275614 54
rect 317970 82 318026 480
rect 318076 82 318104 2246
rect 351012 1193 351040 2246
rect 354289 2204 354585 2224
rect 354345 2202 354369 2204
rect 354425 2202 354449 2204
rect 354505 2202 354529 2204
rect 354367 2150 354369 2202
rect 354431 2150 354443 2202
rect 354505 2150 354507 2202
rect 354345 2148 354369 2150
rect 354425 2148 354449 2150
rect 354505 2148 354529 2150
rect 354289 2128 354585 2148
rect 423600 1465 423628 2479
rect 423586 1456 423642 1465
rect 423586 1391 423642 1400
rect 350998 1184 351054 1193
rect 350998 1119 351054 1128
rect 360106 1184 360162 1193
rect 360106 1119 360162 1128
rect 317970 54 318104 82
rect 360120 82 360148 1119
rect 402886 912 402942 921
rect 402886 847 402942 856
rect 360382 82 360438 480
rect 360120 54 360438 82
rect 317970 0 318026 54
rect 360382 0 360438 54
rect 402794 82 402850 480
rect 402900 82 402928 847
rect 402794 54 402928 82
rect 402794 0 402850 54
<< via2 >>
rect 110 9288 166 9344
rect 18 8064 74 8120
rect 71622 7642 71678 7644
rect 71702 7642 71758 7644
rect 71782 7642 71838 7644
rect 71862 7642 71918 7644
rect 71622 7590 71648 7642
rect 71648 7590 71678 7642
rect 71702 7590 71712 7642
rect 71712 7590 71758 7642
rect 71782 7590 71828 7642
rect 71828 7590 71838 7642
rect 71862 7590 71892 7642
rect 71892 7590 71918 7642
rect 71622 7588 71678 7590
rect 71702 7588 71758 7590
rect 71782 7588 71838 7590
rect 71862 7588 71918 7590
rect 110 6840 166 6896
rect 35622 6840 35678 6896
rect 74998 6840 75054 6896
rect 71622 6554 71678 6556
rect 71702 6554 71758 6556
rect 71782 6554 71838 6556
rect 71862 6554 71918 6556
rect 71622 6502 71648 6554
rect 71648 6502 71678 6554
rect 71702 6502 71712 6554
rect 71712 6502 71758 6554
rect 71782 6502 71828 6554
rect 71828 6502 71838 6554
rect 71862 6502 71892 6554
rect 71892 6502 71918 6554
rect 71622 6500 71678 6502
rect 71702 6500 71758 6502
rect 71782 6500 71838 6502
rect 71862 6500 71918 6502
rect 142289 7098 142345 7100
rect 142369 7098 142425 7100
rect 142449 7098 142505 7100
rect 142529 7098 142585 7100
rect 142289 7046 142315 7098
rect 142315 7046 142345 7098
rect 142369 7046 142379 7098
rect 142379 7046 142425 7098
rect 142449 7046 142495 7098
rect 142495 7046 142505 7098
rect 142529 7046 142559 7098
rect 142559 7046 142585 7098
rect 142289 7044 142345 7046
rect 142369 7044 142425 7046
rect 142449 7044 142505 7046
rect 142529 7044 142585 7046
rect 212956 7642 213012 7644
rect 213036 7642 213092 7644
rect 213116 7642 213172 7644
rect 213196 7642 213252 7644
rect 212956 7590 212982 7642
rect 212982 7590 213012 7642
rect 213036 7590 213046 7642
rect 213046 7590 213092 7642
rect 213116 7590 213162 7642
rect 213162 7590 213172 7642
rect 213196 7590 213226 7642
rect 213226 7590 213252 7642
rect 212956 7588 213012 7590
rect 213036 7588 213092 7590
rect 213116 7588 213172 7590
rect 213196 7588 213252 7590
rect 71622 5466 71678 5468
rect 71702 5466 71758 5468
rect 71782 5466 71838 5468
rect 71862 5466 71918 5468
rect 71622 5414 71648 5466
rect 71648 5414 71678 5466
rect 71702 5414 71712 5466
rect 71712 5414 71758 5466
rect 71782 5414 71828 5466
rect 71828 5414 71838 5466
rect 71862 5414 71892 5466
rect 71892 5414 71918 5466
rect 71622 5412 71678 5414
rect 71702 5412 71758 5414
rect 71782 5412 71838 5414
rect 71862 5412 71918 5414
rect 110 5208 166 5264
rect 18 4664 74 4720
rect 71622 4378 71678 4380
rect 71702 4378 71758 4380
rect 71782 4378 71838 4380
rect 71862 4378 71918 4380
rect 71622 4326 71648 4378
rect 71648 4326 71678 4378
rect 71702 4326 71712 4378
rect 71712 4326 71758 4378
rect 71782 4326 71828 4378
rect 71828 4326 71838 4378
rect 71862 4326 71892 4378
rect 71892 4326 71918 4378
rect 71622 4324 71678 4326
rect 71702 4324 71758 4326
rect 71782 4324 71838 4326
rect 71862 4324 71918 4326
rect 142289 6010 142345 6012
rect 142369 6010 142425 6012
rect 142449 6010 142505 6012
rect 142529 6010 142585 6012
rect 142289 5958 142315 6010
rect 142315 5958 142345 6010
rect 142369 5958 142379 6010
rect 142379 5958 142425 6010
rect 142449 5958 142495 6010
rect 142495 5958 142505 6010
rect 142529 5958 142559 6010
rect 142559 5958 142585 6010
rect 142289 5956 142345 5958
rect 142369 5956 142425 5958
rect 142449 5956 142505 5958
rect 142529 5956 142585 5958
rect 88706 5344 88762 5400
rect 170678 5208 170734 5264
rect 225326 6840 225382 6896
rect 212956 6554 213012 6556
rect 213036 6554 213092 6556
rect 213116 6554 213172 6556
rect 213196 6554 213252 6556
rect 212956 6502 212982 6554
rect 212982 6502 213012 6554
rect 213036 6502 213046 6554
rect 213046 6502 213092 6554
rect 213116 6502 213162 6554
rect 213162 6502 213172 6554
rect 213196 6502 213226 6554
rect 213226 6502 213252 6554
rect 212956 6500 213012 6502
rect 213036 6500 213092 6502
rect 213116 6500 213172 6502
rect 213196 6500 213252 6502
rect 215574 6160 215630 6216
rect 212956 5466 213012 5468
rect 213036 5466 213092 5468
rect 213116 5466 213172 5468
rect 213196 5466 213252 5468
rect 212956 5414 212982 5466
rect 212982 5414 213012 5466
rect 213036 5414 213046 5466
rect 213046 5414 213092 5466
rect 213116 5414 213162 5466
rect 213162 5414 213172 5466
rect 213196 5414 213226 5466
rect 213226 5414 213252 5466
rect 212956 5412 213012 5414
rect 213036 5412 213092 5414
rect 213116 5412 213172 5414
rect 213196 5412 213252 5414
rect 212814 5344 212870 5400
rect 93306 5072 93362 5128
rect 190642 5072 190698 5128
rect 88614 4120 88670 4176
rect 142289 4922 142345 4924
rect 142369 4922 142425 4924
rect 142449 4922 142505 4924
rect 142529 4922 142585 4924
rect 142289 4870 142315 4922
rect 142315 4870 142345 4922
rect 142369 4870 142379 4922
rect 142379 4870 142425 4922
rect 142449 4870 142495 4922
rect 142495 4870 142505 4922
rect 142529 4870 142559 4922
rect 142559 4870 142585 4922
rect 142289 4868 142345 4870
rect 142369 4868 142425 4870
rect 142449 4868 142505 4870
rect 142529 4868 142585 4870
rect 93766 3984 93822 4040
rect 105634 3984 105690 4040
rect 142289 3834 142345 3836
rect 142369 3834 142425 3836
rect 142449 3834 142505 3836
rect 142529 3834 142585 3836
rect 142289 3782 142315 3834
rect 142315 3782 142345 3834
rect 142369 3782 142379 3834
rect 142379 3782 142425 3834
rect 142449 3782 142495 3834
rect 142495 3782 142505 3834
rect 142529 3782 142559 3834
rect 142559 3782 142585 3834
rect 142289 3780 142345 3782
rect 142369 3780 142425 3782
rect 142449 3780 142505 3782
rect 142529 3780 142585 3782
rect 105634 3440 105690 3496
rect 71622 3290 71678 3292
rect 71702 3290 71758 3292
rect 71782 3290 71838 3292
rect 71862 3290 71918 3292
rect 71622 3238 71648 3290
rect 71648 3238 71678 3290
rect 71702 3238 71712 3290
rect 71712 3238 71758 3290
rect 71782 3238 71828 3290
rect 71828 3238 71838 3290
rect 71862 3238 71892 3290
rect 71892 3238 71918 3290
rect 71622 3236 71678 3238
rect 71702 3236 71758 3238
rect 71782 3236 71838 3238
rect 71862 3236 71918 3238
rect 63774 2896 63830 2952
rect 21454 1400 21510 1456
rect 71622 2202 71678 2204
rect 71702 2202 71758 2204
rect 71782 2202 71838 2204
rect 71862 2202 71918 2204
rect 71622 2150 71648 2202
rect 71648 2150 71678 2202
rect 71702 2150 71712 2202
rect 71712 2150 71758 2202
rect 71782 2150 71828 2202
rect 71828 2150 71838 2202
rect 71862 2150 71892 2202
rect 71892 2150 71918 2202
rect 71622 2148 71678 2150
rect 71702 2148 71758 2150
rect 71782 2148 71838 2150
rect 71862 2148 71918 2150
rect 148598 3032 148654 3088
rect 142289 2746 142345 2748
rect 142369 2746 142425 2748
rect 142449 2746 142505 2748
rect 142529 2746 142585 2748
rect 142289 2694 142315 2746
rect 142315 2694 142345 2746
rect 142369 2694 142379 2746
rect 142379 2694 142425 2746
rect 142449 2694 142495 2746
rect 142495 2694 142505 2746
rect 142529 2694 142559 2746
rect 142559 2694 142585 2746
rect 142289 2692 142345 2694
rect 142369 2692 142425 2694
rect 142449 2692 142505 2694
rect 142529 2692 142585 2694
rect 208582 4664 208638 4720
rect 212630 3984 212686 4040
rect 212956 4378 213012 4380
rect 213036 4378 213092 4380
rect 213116 4378 213172 4380
rect 213196 4378 213252 4380
rect 212956 4326 212982 4378
rect 212982 4326 213012 4378
rect 213036 4326 213046 4378
rect 213046 4326 213092 4378
rect 213116 4326 213162 4378
rect 213162 4326 213172 4378
rect 213196 4326 213226 4378
rect 213226 4326 213252 4378
rect 212956 4324 213012 4326
rect 213036 4324 213092 4326
rect 213116 4324 213172 4326
rect 213196 4324 213252 4326
rect 212956 3290 213012 3292
rect 213036 3290 213092 3292
rect 213116 3290 213172 3292
rect 213196 3290 213252 3292
rect 212956 3238 212982 3290
rect 212982 3238 213012 3290
rect 213036 3238 213046 3290
rect 213046 3238 213092 3290
rect 213116 3238 213162 3290
rect 213162 3238 213172 3290
rect 213196 3238 213226 3290
rect 213226 3238 213252 3290
rect 212956 3236 213012 3238
rect 213036 3236 213092 3238
rect 213116 3236 213172 3238
rect 213196 3236 213252 3238
rect 209226 3032 209282 3088
rect 200946 2488 201002 2544
rect 212998 2488 213054 2544
rect 283622 7098 283678 7100
rect 283702 7098 283758 7100
rect 283782 7098 283838 7100
rect 283862 7098 283918 7100
rect 283622 7046 283648 7098
rect 283648 7046 283678 7098
rect 283702 7046 283712 7098
rect 283712 7046 283758 7098
rect 283782 7046 283828 7098
rect 283828 7046 283838 7098
rect 283862 7046 283892 7098
rect 283892 7046 283918 7098
rect 283622 7044 283678 7046
rect 283702 7044 283758 7046
rect 283782 7044 283838 7046
rect 283862 7044 283918 7046
rect 247406 6840 247462 6896
rect 354289 7642 354345 7644
rect 354369 7642 354425 7644
rect 354449 7642 354505 7644
rect 354529 7642 354585 7644
rect 354289 7590 354315 7642
rect 354315 7590 354345 7642
rect 354369 7590 354379 7642
rect 354379 7590 354425 7642
rect 354449 7590 354495 7642
rect 354495 7590 354505 7642
rect 354529 7590 354559 7642
rect 354559 7590 354585 7642
rect 354289 7588 354345 7590
rect 354369 7588 354425 7590
rect 354449 7588 354505 7590
rect 354529 7588 354585 7590
rect 229558 6704 229614 6760
rect 318062 6704 318118 6760
rect 354289 6554 354345 6556
rect 354369 6554 354425 6556
rect 354449 6554 354505 6556
rect 354529 6554 354585 6556
rect 354289 6502 354315 6554
rect 354315 6502 354345 6554
rect 354369 6502 354379 6554
rect 354379 6502 354425 6554
rect 354449 6502 354495 6554
rect 354495 6502 354505 6554
rect 354529 6502 354559 6554
rect 354559 6502 354585 6554
rect 354289 6500 354345 6502
rect 354369 6500 354425 6502
rect 354449 6500 354505 6502
rect 354529 6500 354585 6502
rect 225694 6296 225750 6352
rect 388718 6160 388774 6216
rect 217874 5772 217930 5808
rect 217874 5752 217876 5772
rect 217876 5752 217928 5772
rect 217928 5752 217930 5772
rect 215942 5072 215998 5128
rect 213274 2352 213330 2408
rect 200946 1400 201002 1456
rect 212956 2202 213012 2204
rect 213036 2202 213092 2204
rect 213116 2202 213172 2204
rect 213196 2202 213252 2204
rect 212956 2150 212982 2202
rect 212982 2150 213012 2202
rect 213036 2150 213046 2202
rect 213046 2150 213092 2202
rect 213116 2150 213162 2202
rect 213162 2150 213172 2202
rect 213196 2150 213226 2202
rect 213226 2150 213252 2202
rect 212956 2148 213012 2150
rect 213036 2148 213092 2150
rect 213116 2148 213172 2150
rect 213196 2148 213252 2150
rect 212446 856 212502 912
rect 283622 6010 283678 6012
rect 283702 6010 283758 6012
rect 283782 6010 283838 6012
rect 283862 6010 283918 6012
rect 283622 5958 283648 6010
rect 283648 5958 283678 6010
rect 283702 5958 283712 6010
rect 283712 5958 283758 6010
rect 283782 5958 283828 6010
rect 283828 5958 283838 6010
rect 283862 5958 283892 6010
rect 283892 5958 283918 6010
rect 283622 5956 283678 5958
rect 283702 5956 283758 5958
rect 283782 5956 283838 5958
rect 283862 5956 283918 5958
rect 423586 9152 423642 9208
rect 423586 7520 423642 7576
rect 423402 5752 423458 5808
rect 423678 5888 423734 5944
rect 354289 5466 354345 5468
rect 354369 5466 354425 5468
rect 354449 5466 354505 5468
rect 354529 5466 354585 5468
rect 354289 5414 354315 5466
rect 354315 5414 354345 5466
rect 354369 5414 354379 5466
rect 354379 5414 354425 5466
rect 354449 5414 354495 5466
rect 354495 5414 354505 5466
rect 354529 5414 354559 5466
rect 354559 5414 354585 5466
rect 354289 5412 354345 5414
rect 354369 5412 354425 5414
rect 354449 5412 354505 5414
rect 354529 5412 354585 5414
rect 221922 5208 221978 5264
rect 217690 3440 217746 3496
rect 221922 4120 221978 4176
rect 283622 4922 283678 4924
rect 283702 4922 283758 4924
rect 283782 4922 283838 4924
rect 283862 4922 283918 4924
rect 283622 4870 283648 4922
rect 283648 4870 283678 4922
rect 283702 4870 283712 4922
rect 283712 4870 283758 4922
rect 283782 4870 283828 4922
rect 283828 4870 283838 4922
rect 283862 4870 283892 4922
rect 283892 4870 283918 4922
rect 283622 4868 283678 4870
rect 283702 4868 283758 4870
rect 283782 4868 283838 4870
rect 283862 4868 283918 4870
rect 354289 4378 354345 4380
rect 354369 4378 354425 4380
rect 354449 4378 354505 4380
rect 354529 4378 354585 4380
rect 354289 4326 354315 4378
rect 354315 4326 354345 4378
rect 354369 4326 354379 4378
rect 354379 4326 354425 4378
rect 354449 4326 354495 4378
rect 354495 4326 354505 4378
rect 354529 4326 354559 4378
rect 354559 4326 354585 4378
rect 354289 4324 354345 4326
rect 354369 4324 354425 4326
rect 354449 4324 354505 4326
rect 354529 4324 354585 4326
rect 283622 3834 283678 3836
rect 283702 3834 283758 3836
rect 283782 3834 283838 3836
rect 283862 3834 283918 3836
rect 283622 3782 283648 3834
rect 283648 3782 283678 3834
rect 283702 3782 283712 3834
rect 283712 3782 283758 3834
rect 283782 3782 283828 3834
rect 283828 3782 283838 3834
rect 283862 3782 283892 3834
rect 283892 3782 283918 3834
rect 283622 3780 283678 3782
rect 283702 3780 283758 3782
rect 283782 3780 283838 3782
rect 283862 3780 283918 3782
rect 354289 3290 354345 3292
rect 354369 3290 354425 3292
rect 354449 3290 354505 3292
rect 354529 3290 354585 3292
rect 354289 3238 354315 3290
rect 354315 3238 354345 3290
rect 354369 3238 354379 3290
rect 354379 3238 354425 3290
rect 354449 3238 354495 3290
rect 354495 3238 354505 3290
rect 354529 3238 354559 3290
rect 354559 3238 354585 3290
rect 354289 3236 354345 3238
rect 354369 3236 354425 3238
rect 354449 3236 354505 3238
rect 354529 3236 354585 3238
rect 224406 2896 224462 2952
rect 221002 2488 221058 2544
rect 423678 2760 423734 2816
rect 283622 2746 283678 2748
rect 283702 2746 283758 2748
rect 283782 2746 283838 2748
rect 283862 2746 283918 2748
rect 283622 2694 283648 2746
rect 283648 2694 283678 2746
rect 283702 2694 283712 2746
rect 283712 2694 283758 2746
rect 283782 2694 283828 2746
rect 283828 2694 283838 2746
rect 283862 2694 283892 2746
rect 283892 2694 283918 2746
rect 283622 2692 283678 2694
rect 283702 2692 283758 2694
rect 283782 2692 283838 2694
rect 283862 2692 283918 2694
rect 308586 2488 308642 2544
rect 423586 2488 423642 2544
rect 309966 2352 310022 2408
rect 350814 2352 350870 2408
rect 220450 1400 220506 1456
rect 216862 176 216918 232
rect 228362 1128 228418 1184
rect 275282 1128 275338 1184
rect 221186 40 221242 96
rect 233146 40 233202 96
rect 354289 2202 354345 2204
rect 354369 2202 354425 2204
rect 354449 2202 354505 2204
rect 354529 2202 354585 2204
rect 354289 2150 354315 2202
rect 354315 2150 354345 2202
rect 354369 2150 354379 2202
rect 354379 2150 354425 2202
rect 354449 2150 354495 2202
rect 354495 2150 354505 2202
rect 354529 2150 354559 2202
rect 354559 2150 354585 2202
rect 354289 2148 354345 2150
rect 354369 2148 354425 2150
rect 354449 2148 354505 2150
rect 354529 2148 354585 2150
rect 423586 1400 423642 1456
rect 350998 1128 351054 1184
rect 360106 1128 360162 1184
rect 402886 856 402942 912
<< metal3 >>
rect 0 9344 480 9376
rect 0 9288 110 9344
rect 166 9288 480 9344
rect 0 9256 480 9288
rect 423520 9208 424000 9240
rect 423520 9152 423586 9208
rect 423642 9152 424000 9208
rect 423520 9120 424000 9152
rect 0 8120 480 8152
rect 0 8064 18 8120
rect 74 8064 480 8120
rect 0 8032 480 8064
rect 71610 7648 71930 7649
rect 71610 7584 71618 7648
rect 71682 7584 71698 7648
rect 71762 7584 71778 7648
rect 71842 7584 71858 7648
rect 71922 7584 71930 7648
rect 71610 7583 71930 7584
rect 212944 7648 213264 7649
rect 212944 7584 212952 7648
rect 213016 7584 213032 7648
rect 213096 7584 213112 7648
rect 213176 7584 213192 7648
rect 213256 7584 213264 7648
rect 212944 7583 213264 7584
rect 354277 7648 354597 7649
rect 354277 7584 354285 7648
rect 354349 7584 354365 7648
rect 354429 7584 354445 7648
rect 354509 7584 354525 7648
rect 354589 7584 354597 7648
rect 354277 7583 354597 7584
rect 423520 7576 424000 7608
rect 423520 7520 423586 7576
rect 423642 7520 424000 7576
rect 423520 7488 424000 7520
rect 142277 7104 142597 7105
rect 142277 7040 142285 7104
rect 142349 7040 142365 7104
rect 142429 7040 142445 7104
rect 142509 7040 142525 7104
rect 142589 7040 142597 7104
rect 142277 7039 142597 7040
rect 283610 7104 283930 7105
rect 283610 7040 283618 7104
rect 283682 7040 283698 7104
rect 283762 7040 283778 7104
rect 283842 7040 283858 7104
rect 283922 7040 283930 7104
rect 283610 7039 283930 7040
rect 0 6896 480 6928
rect 0 6840 110 6896
rect 166 6840 480 6896
rect 0 6808 480 6840
rect 35617 6898 35683 6901
rect 74993 6898 75059 6901
rect 35617 6896 75059 6898
rect 35617 6840 35622 6896
rect 35678 6840 74998 6896
rect 75054 6840 75059 6896
rect 35617 6838 75059 6840
rect 35617 6835 35683 6838
rect 74993 6835 75059 6838
rect 225321 6898 225387 6901
rect 247401 6898 247467 6901
rect 225321 6896 247467 6898
rect 225321 6840 225326 6896
rect 225382 6840 247406 6896
rect 247462 6840 247467 6896
rect 225321 6838 247467 6840
rect 225321 6835 225387 6838
rect 247401 6835 247467 6838
rect 229553 6762 229619 6765
rect 318057 6762 318123 6765
rect 229553 6760 318123 6762
rect 229553 6704 229558 6760
rect 229614 6704 318062 6760
rect 318118 6704 318123 6760
rect 229553 6702 318123 6704
rect 229553 6699 229619 6702
rect 318057 6699 318123 6702
rect 71610 6560 71930 6561
rect 71610 6496 71618 6560
rect 71682 6496 71698 6560
rect 71762 6496 71778 6560
rect 71842 6496 71858 6560
rect 71922 6496 71930 6560
rect 71610 6495 71930 6496
rect 212944 6560 213264 6561
rect 212944 6496 212952 6560
rect 213016 6496 213032 6560
rect 213096 6496 213112 6560
rect 213176 6496 213192 6560
rect 213256 6496 213264 6560
rect 212944 6495 213264 6496
rect 354277 6560 354597 6561
rect 354277 6496 354285 6560
rect 354349 6496 354365 6560
rect 354429 6496 354445 6560
rect 354509 6496 354525 6560
rect 354589 6496 354597 6560
rect 354277 6495 354597 6496
rect 225689 6354 225755 6357
rect 62 6352 225755 6354
rect 62 6296 225694 6352
rect 225750 6296 225755 6352
rect 62 6294 225755 6296
rect 62 5704 122 6294
rect 225689 6291 225755 6294
rect 215569 6218 215635 6221
rect 388713 6218 388779 6221
rect 215569 6216 388779 6218
rect 215569 6160 215574 6216
rect 215630 6160 388718 6216
rect 388774 6160 388779 6216
rect 215569 6158 388779 6160
rect 215569 6155 215635 6158
rect 388713 6155 388779 6158
rect 142277 6016 142597 6017
rect 142277 5952 142285 6016
rect 142349 5952 142365 6016
rect 142429 5952 142445 6016
rect 142509 5952 142525 6016
rect 142589 5952 142597 6016
rect 142277 5951 142597 5952
rect 283610 6016 283930 6017
rect 283610 5952 283618 6016
rect 283682 5952 283698 6016
rect 283762 5952 283778 6016
rect 283842 5952 283858 6016
rect 283922 5952 283930 6016
rect 283610 5951 283930 5952
rect 423520 5944 424000 5976
rect 423520 5888 423678 5944
rect 423734 5888 424000 5944
rect 423520 5856 424000 5888
rect 217869 5810 217935 5813
rect 423397 5810 423463 5813
rect 217869 5808 423463 5810
rect 217869 5752 217874 5808
rect 217930 5752 423402 5808
rect 423458 5752 423463 5808
rect 217869 5750 423463 5752
rect 217869 5747 217935 5750
rect 423397 5747 423463 5750
rect 0 5584 480 5704
rect 71610 5472 71930 5473
rect 71610 5408 71618 5472
rect 71682 5408 71698 5472
rect 71762 5408 71778 5472
rect 71842 5408 71858 5472
rect 71922 5408 71930 5472
rect 71610 5407 71930 5408
rect 212944 5472 213264 5473
rect 212944 5408 212952 5472
rect 213016 5408 213032 5472
rect 213096 5408 213112 5472
rect 213176 5408 213192 5472
rect 213256 5408 213264 5472
rect 212944 5407 213264 5408
rect 354277 5472 354597 5473
rect 354277 5408 354285 5472
rect 354349 5408 354365 5472
rect 354429 5408 354445 5472
rect 354509 5408 354525 5472
rect 354589 5408 354597 5472
rect 354277 5407 354597 5408
rect 88701 5402 88767 5405
rect 212809 5402 212875 5405
rect 88701 5400 212875 5402
rect 88701 5344 88706 5400
rect 88762 5344 212814 5400
rect 212870 5344 212875 5400
rect 88701 5342 212875 5344
rect 88701 5339 88767 5342
rect 212809 5339 212875 5342
rect 105 5266 171 5269
rect 170673 5266 170739 5269
rect 221917 5266 221983 5269
rect 105 5264 81450 5266
rect 105 5208 110 5264
rect 166 5208 81450 5264
rect 105 5206 81450 5208
rect 105 5203 171 5206
rect 81390 5130 81450 5206
rect 170673 5264 221983 5266
rect 170673 5208 170678 5264
rect 170734 5208 221922 5264
rect 221978 5208 221983 5264
rect 170673 5206 221983 5208
rect 170673 5203 170739 5206
rect 221917 5203 221983 5206
rect 93301 5130 93367 5133
rect 81390 5128 93367 5130
rect 81390 5072 93306 5128
rect 93362 5072 93367 5128
rect 81390 5070 93367 5072
rect 93301 5067 93367 5070
rect 190637 5130 190703 5133
rect 215937 5130 216003 5133
rect 190637 5128 216003 5130
rect 190637 5072 190642 5128
rect 190698 5072 215942 5128
rect 215998 5072 216003 5128
rect 190637 5070 216003 5072
rect 190637 5067 190703 5070
rect 215937 5067 216003 5070
rect 142277 4928 142597 4929
rect 142277 4864 142285 4928
rect 142349 4864 142365 4928
rect 142429 4864 142445 4928
rect 142509 4864 142525 4928
rect 142589 4864 142597 4928
rect 142277 4863 142597 4864
rect 283610 4928 283930 4929
rect 283610 4864 283618 4928
rect 283682 4864 283698 4928
rect 283762 4864 283778 4928
rect 283842 4864 283858 4928
rect 283922 4864 283930 4928
rect 283610 4863 283930 4864
rect 13 4722 79 4725
rect 208577 4722 208643 4725
rect 13 4720 208643 4722
rect 13 4664 18 4720
rect 74 4664 208582 4720
rect 208638 4664 208643 4720
rect 13 4662 208643 4664
rect 13 4659 79 4662
rect 208577 4659 208643 4662
rect 423622 4450 423628 4452
rect 415350 4390 423628 4450
rect 71610 4384 71930 4385
rect 0 4316 480 4344
rect 71610 4320 71618 4384
rect 71682 4320 71698 4384
rect 71762 4320 71778 4384
rect 71842 4320 71858 4384
rect 71922 4320 71930 4384
rect 71610 4319 71930 4320
rect 212944 4384 213264 4385
rect 212944 4320 212952 4384
rect 213016 4320 213032 4384
rect 213096 4320 213112 4384
rect 213176 4320 213192 4384
rect 213256 4320 213264 4384
rect 212944 4319 213264 4320
rect 354277 4384 354597 4385
rect 354277 4320 354285 4384
rect 354349 4320 354365 4384
rect 354429 4320 354445 4384
rect 354509 4320 354525 4384
rect 354589 4320 354597 4384
rect 354277 4319 354597 4320
rect 0 4252 60 4316
rect 124 4252 480 4316
rect 415350 4314 415410 4390
rect 423622 4388 423628 4390
rect 423692 4388 423698 4452
rect 0 4224 480 4252
rect 409830 4254 415410 4314
rect 88609 4178 88675 4181
rect 9630 4176 88675 4178
rect 9630 4120 88614 4176
rect 88670 4120 88675 4176
rect 9630 4118 88675 4120
rect 54 3980 60 4044
rect 124 4042 130 4044
rect 9630 4042 9690 4118
rect 88609 4115 88675 4118
rect 221917 4178 221983 4181
rect 409830 4178 409890 4254
rect 423520 4180 424000 4208
rect 423520 4178 423628 4180
rect 221917 4176 409890 4178
rect 221917 4120 221922 4176
rect 221978 4120 409890 4176
rect 221917 4118 409890 4120
rect 423500 4118 423628 4178
rect 221917 4115 221983 4118
rect 423520 4116 423628 4118
rect 423692 4116 424000 4180
rect 423520 4088 424000 4116
rect 124 3982 9690 4042
rect 93761 4042 93827 4045
rect 105629 4042 105695 4045
rect 212625 4042 212691 4045
rect 93761 4040 105695 4042
rect 93761 3984 93766 4040
rect 93822 3984 105634 4040
rect 105690 3984 105695 4040
rect 93761 3982 105695 3984
rect 124 3980 130 3982
rect 93761 3979 93827 3982
rect 105629 3979 105695 3982
rect 197310 4040 212691 4042
rect 197310 3984 212630 4040
rect 212686 3984 212691 4040
rect 197310 3982 212691 3984
rect 142277 3840 142597 3841
rect 142277 3776 142285 3840
rect 142349 3776 142365 3840
rect 142429 3776 142445 3840
rect 142509 3776 142525 3840
rect 142589 3776 142597 3840
rect 142277 3775 142597 3776
rect 197310 3634 197370 3982
rect 212625 3979 212691 3982
rect 283610 3840 283930 3841
rect 283610 3776 283618 3840
rect 283682 3776 283698 3840
rect 283762 3776 283778 3840
rect 283842 3776 283858 3840
rect 283922 3776 283930 3840
rect 283610 3775 283930 3776
rect 62 3574 197370 3634
rect 62 3120 122 3574
rect 105629 3498 105695 3501
rect 217685 3498 217751 3501
rect 105629 3496 217751 3498
rect 105629 3440 105634 3496
rect 105690 3440 217690 3496
rect 217746 3440 217751 3496
rect 105629 3438 217751 3440
rect 105629 3435 105695 3438
rect 217685 3435 217751 3438
rect 71610 3296 71930 3297
rect 71610 3232 71618 3296
rect 71682 3232 71698 3296
rect 71762 3232 71778 3296
rect 71842 3232 71858 3296
rect 71922 3232 71930 3296
rect 71610 3231 71930 3232
rect 212944 3296 213264 3297
rect 212944 3232 212952 3296
rect 213016 3232 213032 3296
rect 213096 3232 213112 3296
rect 213176 3232 213192 3296
rect 213256 3232 213264 3296
rect 212944 3231 213264 3232
rect 354277 3296 354597 3297
rect 354277 3232 354285 3296
rect 354349 3232 354365 3296
rect 354429 3232 354445 3296
rect 354509 3232 354525 3296
rect 354589 3232 354597 3296
rect 354277 3231 354597 3232
rect 0 3000 480 3120
rect 148593 3090 148659 3093
rect 209221 3090 209287 3093
rect 148593 3088 209287 3090
rect 148593 3032 148598 3088
rect 148654 3032 209226 3088
rect 209282 3032 209287 3088
rect 148593 3030 209287 3032
rect 148593 3027 148659 3030
rect 209221 3027 209287 3030
rect 63769 2954 63835 2957
rect 224401 2954 224467 2957
rect 63769 2952 224467 2954
rect 63769 2896 63774 2952
rect 63830 2896 224406 2952
rect 224462 2896 224467 2952
rect 63769 2894 224467 2896
rect 63769 2891 63835 2894
rect 224401 2891 224467 2894
rect 423673 2818 423739 2821
rect 415350 2816 423739 2818
rect 415350 2760 423678 2816
rect 423734 2760 423739 2816
rect 415350 2758 423739 2760
rect 142277 2752 142597 2753
rect 142277 2688 142285 2752
rect 142349 2688 142365 2752
rect 142429 2688 142445 2752
rect 142509 2688 142525 2752
rect 142589 2688 142597 2752
rect 142277 2687 142597 2688
rect 283610 2752 283930 2753
rect 283610 2688 283618 2752
rect 283682 2688 283698 2752
rect 283762 2688 283778 2752
rect 283842 2688 283858 2752
rect 283922 2688 283930 2752
rect 283610 2687 283930 2688
rect 415350 2682 415410 2758
rect 423673 2755 423739 2758
rect 409830 2622 415410 2682
rect 200941 2546 201007 2549
rect 212993 2546 213059 2549
rect 200941 2544 213059 2546
rect 200941 2488 200946 2544
rect 201002 2488 212998 2544
rect 213054 2488 213059 2544
rect 200941 2486 213059 2488
rect 200941 2483 201007 2486
rect 212993 2483 213059 2486
rect 220997 2546 221063 2549
rect 308581 2546 308647 2549
rect 409830 2546 409890 2622
rect 220997 2544 308647 2546
rect 220997 2488 221002 2544
rect 221058 2488 308586 2544
rect 308642 2488 308647 2544
rect 220997 2486 308647 2488
rect 220997 2483 221063 2486
rect 308581 2483 308647 2486
rect 351870 2486 409890 2546
rect 423520 2544 424000 2576
rect 423520 2488 423586 2544
rect 423642 2488 424000 2544
rect 213269 2410 213335 2413
rect 197310 2408 213335 2410
rect 197310 2352 213274 2408
rect 213330 2352 213335 2408
rect 197310 2350 213335 2352
rect 71610 2208 71930 2209
rect 71610 2144 71618 2208
rect 71682 2144 71698 2208
rect 71762 2144 71778 2208
rect 71842 2144 71858 2208
rect 71922 2144 71930 2208
rect 71610 2143 71930 2144
rect 54 2076 60 2140
rect 124 2138 130 2140
rect 124 2078 9690 2138
rect 124 2076 130 2078
rect 9630 2002 9690 2078
rect 197310 2002 197370 2350
rect 213269 2347 213335 2350
rect 309961 2410 310027 2413
rect 350809 2410 350875 2413
rect 351870 2410 351930 2486
rect 423520 2456 424000 2488
rect 309961 2408 351930 2410
rect 309961 2352 309966 2408
rect 310022 2352 350814 2408
rect 350870 2352 351930 2408
rect 309961 2350 351930 2352
rect 309961 2347 310027 2350
rect 350809 2347 350875 2350
rect 212944 2208 213264 2209
rect 212944 2144 212952 2208
rect 213016 2144 213032 2208
rect 213096 2144 213112 2208
rect 213176 2144 213192 2208
rect 213256 2144 213264 2208
rect 212944 2143 213264 2144
rect 354277 2208 354597 2209
rect 354277 2144 354285 2208
rect 354349 2144 354365 2208
rect 354429 2144 354445 2208
rect 354509 2144 354525 2208
rect 354589 2144 354597 2208
rect 354277 2143 354597 2144
rect 9630 1942 197370 2002
rect 0 1868 480 1896
rect 0 1804 60 1868
rect 124 1804 480 1868
rect 0 1776 480 1804
rect 21449 1458 21515 1461
rect 200941 1458 201007 1461
rect 21449 1456 201007 1458
rect 21449 1400 21454 1456
rect 21510 1400 200946 1456
rect 201002 1400 201007 1456
rect 21449 1398 201007 1400
rect 21449 1395 21515 1398
rect 200941 1395 201007 1398
rect 220445 1458 220511 1461
rect 423581 1458 423647 1461
rect 220445 1456 423647 1458
rect 220445 1400 220450 1456
rect 220506 1400 423586 1456
rect 423642 1400 423647 1456
rect 220445 1398 423647 1400
rect 220445 1395 220511 1398
rect 423581 1395 423647 1398
rect 228357 1186 228423 1189
rect 275277 1186 275343 1189
rect 228357 1184 275343 1186
rect 228357 1128 228362 1184
rect 228418 1128 275282 1184
rect 275338 1128 275343 1184
rect 228357 1126 275343 1128
rect 228357 1123 228423 1126
rect 275277 1123 275343 1126
rect 350993 1186 351059 1189
rect 360101 1186 360167 1189
rect 350993 1184 360167 1186
rect 350993 1128 350998 1184
rect 351054 1128 360106 1184
rect 360162 1128 360167 1184
rect 350993 1126 360167 1128
rect 350993 1123 351059 1126
rect 360101 1123 360167 1126
rect 212441 914 212507 917
rect 402881 914 402947 917
rect 212441 912 402947 914
rect 212441 856 212446 912
rect 212502 856 402886 912
rect 402942 856 402947 912
rect 212441 854 402947 856
rect 212441 851 212507 854
rect 402881 851 402947 854
rect 423520 824 424000 944
rect 0 552 480 672
rect 216857 234 216923 237
rect 423630 234 423690 824
rect 216857 232 423690 234
rect 216857 176 216862 232
rect 216918 176 423690 232
rect 216857 174 423690 176
rect 216857 171 216923 174
rect 221181 98 221247 101
rect 233141 98 233207 101
rect 221181 96 233207 98
rect 221181 40 221186 96
rect 221242 40 233146 96
rect 233202 40 233207 96
rect 221181 38 233207 40
rect 221181 35 221247 38
rect 233141 35 233207 38
<< via3 >>
rect 71618 7644 71682 7648
rect 71618 7588 71622 7644
rect 71622 7588 71678 7644
rect 71678 7588 71682 7644
rect 71618 7584 71682 7588
rect 71698 7644 71762 7648
rect 71698 7588 71702 7644
rect 71702 7588 71758 7644
rect 71758 7588 71762 7644
rect 71698 7584 71762 7588
rect 71778 7644 71842 7648
rect 71778 7588 71782 7644
rect 71782 7588 71838 7644
rect 71838 7588 71842 7644
rect 71778 7584 71842 7588
rect 71858 7644 71922 7648
rect 71858 7588 71862 7644
rect 71862 7588 71918 7644
rect 71918 7588 71922 7644
rect 71858 7584 71922 7588
rect 212952 7644 213016 7648
rect 212952 7588 212956 7644
rect 212956 7588 213012 7644
rect 213012 7588 213016 7644
rect 212952 7584 213016 7588
rect 213032 7644 213096 7648
rect 213032 7588 213036 7644
rect 213036 7588 213092 7644
rect 213092 7588 213096 7644
rect 213032 7584 213096 7588
rect 213112 7644 213176 7648
rect 213112 7588 213116 7644
rect 213116 7588 213172 7644
rect 213172 7588 213176 7644
rect 213112 7584 213176 7588
rect 213192 7644 213256 7648
rect 213192 7588 213196 7644
rect 213196 7588 213252 7644
rect 213252 7588 213256 7644
rect 213192 7584 213256 7588
rect 354285 7644 354349 7648
rect 354285 7588 354289 7644
rect 354289 7588 354345 7644
rect 354345 7588 354349 7644
rect 354285 7584 354349 7588
rect 354365 7644 354429 7648
rect 354365 7588 354369 7644
rect 354369 7588 354425 7644
rect 354425 7588 354429 7644
rect 354365 7584 354429 7588
rect 354445 7644 354509 7648
rect 354445 7588 354449 7644
rect 354449 7588 354505 7644
rect 354505 7588 354509 7644
rect 354445 7584 354509 7588
rect 354525 7644 354589 7648
rect 354525 7588 354529 7644
rect 354529 7588 354585 7644
rect 354585 7588 354589 7644
rect 354525 7584 354589 7588
rect 142285 7100 142349 7104
rect 142285 7044 142289 7100
rect 142289 7044 142345 7100
rect 142345 7044 142349 7100
rect 142285 7040 142349 7044
rect 142365 7100 142429 7104
rect 142365 7044 142369 7100
rect 142369 7044 142425 7100
rect 142425 7044 142429 7100
rect 142365 7040 142429 7044
rect 142445 7100 142509 7104
rect 142445 7044 142449 7100
rect 142449 7044 142505 7100
rect 142505 7044 142509 7100
rect 142445 7040 142509 7044
rect 142525 7100 142589 7104
rect 142525 7044 142529 7100
rect 142529 7044 142585 7100
rect 142585 7044 142589 7100
rect 142525 7040 142589 7044
rect 283618 7100 283682 7104
rect 283618 7044 283622 7100
rect 283622 7044 283678 7100
rect 283678 7044 283682 7100
rect 283618 7040 283682 7044
rect 283698 7100 283762 7104
rect 283698 7044 283702 7100
rect 283702 7044 283758 7100
rect 283758 7044 283762 7100
rect 283698 7040 283762 7044
rect 283778 7100 283842 7104
rect 283778 7044 283782 7100
rect 283782 7044 283838 7100
rect 283838 7044 283842 7100
rect 283778 7040 283842 7044
rect 283858 7100 283922 7104
rect 283858 7044 283862 7100
rect 283862 7044 283918 7100
rect 283918 7044 283922 7100
rect 283858 7040 283922 7044
rect 71618 6556 71682 6560
rect 71618 6500 71622 6556
rect 71622 6500 71678 6556
rect 71678 6500 71682 6556
rect 71618 6496 71682 6500
rect 71698 6556 71762 6560
rect 71698 6500 71702 6556
rect 71702 6500 71758 6556
rect 71758 6500 71762 6556
rect 71698 6496 71762 6500
rect 71778 6556 71842 6560
rect 71778 6500 71782 6556
rect 71782 6500 71838 6556
rect 71838 6500 71842 6556
rect 71778 6496 71842 6500
rect 71858 6556 71922 6560
rect 71858 6500 71862 6556
rect 71862 6500 71918 6556
rect 71918 6500 71922 6556
rect 71858 6496 71922 6500
rect 212952 6556 213016 6560
rect 212952 6500 212956 6556
rect 212956 6500 213012 6556
rect 213012 6500 213016 6556
rect 212952 6496 213016 6500
rect 213032 6556 213096 6560
rect 213032 6500 213036 6556
rect 213036 6500 213092 6556
rect 213092 6500 213096 6556
rect 213032 6496 213096 6500
rect 213112 6556 213176 6560
rect 213112 6500 213116 6556
rect 213116 6500 213172 6556
rect 213172 6500 213176 6556
rect 213112 6496 213176 6500
rect 213192 6556 213256 6560
rect 213192 6500 213196 6556
rect 213196 6500 213252 6556
rect 213252 6500 213256 6556
rect 213192 6496 213256 6500
rect 354285 6556 354349 6560
rect 354285 6500 354289 6556
rect 354289 6500 354345 6556
rect 354345 6500 354349 6556
rect 354285 6496 354349 6500
rect 354365 6556 354429 6560
rect 354365 6500 354369 6556
rect 354369 6500 354425 6556
rect 354425 6500 354429 6556
rect 354365 6496 354429 6500
rect 354445 6556 354509 6560
rect 354445 6500 354449 6556
rect 354449 6500 354505 6556
rect 354505 6500 354509 6556
rect 354445 6496 354509 6500
rect 354525 6556 354589 6560
rect 354525 6500 354529 6556
rect 354529 6500 354585 6556
rect 354585 6500 354589 6556
rect 354525 6496 354589 6500
rect 142285 6012 142349 6016
rect 142285 5956 142289 6012
rect 142289 5956 142345 6012
rect 142345 5956 142349 6012
rect 142285 5952 142349 5956
rect 142365 6012 142429 6016
rect 142365 5956 142369 6012
rect 142369 5956 142425 6012
rect 142425 5956 142429 6012
rect 142365 5952 142429 5956
rect 142445 6012 142509 6016
rect 142445 5956 142449 6012
rect 142449 5956 142505 6012
rect 142505 5956 142509 6012
rect 142445 5952 142509 5956
rect 142525 6012 142589 6016
rect 142525 5956 142529 6012
rect 142529 5956 142585 6012
rect 142585 5956 142589 6012
rect 142525 5952 142589 5956
rect 283618 6012 283682 6016
rect 283618 5956 283622 6012
rect 283622 5956 283678 6012
rect 283678 5956 283682 6012
rect 283618 5952 283682 5956
rect 283698 6012 283762 6016
rect 283698 5956 283702 6012
rect 283702 5956 283758 6012
rect 283758 5956 283762 6012
rect 283698 5952 283762 5956
rect 283778 6012 283842 6016
rect 283778 5956 283782 6012
rect 283782 5956 283838 6012
rect 283838 5956 283842 6012
rect 283778 5952 283842 5956
rect 283858 6012 283922 6016
rect 283858 5956 283862 6012
rect 283862 5956 283918 6012
rect 283918 5956 283922 6012
rect 283858 5952 283922 5956
rect 71618 5468 71682 5472
rect 71618 5412 71622 5468
rect 71622 5412 71678 5468
rect 71678 5412 71682 5468
rect 71618 5408 71682 5412
rect 71698 5468 71762 5472
rect 71698 5412 71702 5468
rect 71702 5412 71758 5468
rect 71758 5412 71762 5468
rect 71698 5408 71762 5412
rect 71778 5468 71842 5472
rect 71778 5412 71782 5468
rect 71782 5412 71838 5468
rect 71838 5412 71842 5468
rect 71778 5408 71842 5412
rect 71858 5468 71922 5472
rect 71858 5412 71862 5468
rect 71862 5412 71918 5468
rect 71918 5412 71922 5468
rect 71858 5408 71922 5412
rect 212952 5468 213016 5472
rect 212952 5412 212956 5468
rect 212956 5412 213012 5468
rect 213012 5412 213016 5468
rect 212952 5408 213016 5412
rect 213032 5468 213096 5472
rect 213032 5412 213036 5468
rect 213036 5412 213092 5468
rect 213092 5412 213096 5468
rect 213032 5408 213096 5412
rect 213112 5468 213176 5472
rect 213112 5412 213116 5468
rect 213116 5412 213172 5468
rect 213172 5412 213176 5468
rect 213112 5408 213176 5412
rect 213192 5468 213256 5472
rect 213192 5412 213196 5468
rect 213196 5412 213252 5468
rect 213252 5412 213256 5468
rect 213192 5408 213256 5412
rect 354285 5468 354349 5472
rect 354285 5412 354289 5468
rect 354289 5412 354345 5468
rect 354345 5412 354349 5468
rect 354285 5408 354349 5412
rect 354365 5468 354429 5472
rect 354365 5412 354369 5468
rect 354369 5412 354425 5468
rect 354425 5412 354429 5468
rect 354365 5408 354429 5412
rect 354445 5468 354509 5472
rect 354445 5412 354449 5468
rect 354449 5412 354505 5468
rect 354505 5412 354509 5468
rect 354445 5408 354509 5412
rect 354525 5468 354589 5472
rect 354525 5412 354529 5468
rect 354529 5412 354585 5468
rect 354585 5412 354589 5468
rect 354525 5408 354589 5412
rect 142285 4924 142349 4928
rect 142285 4868 142289 4924
rect 142289 4868 142345 4924
rect 142345 4868 142349 4924
rect 142285 4864 142349 4868
rect 142365 4924 142429 4928
rect 142365 4868 142369 4924
rect 142369 4868 142425 4924
rect 142425 4868 142429 4924
rect 142365 4864 142429 4868
rect 142445 4924 142509 4928
rect 142445 4868 142449 4924
rect 142449 4868 142505 4924
rect 142505 4868 142509 4924
rect 142445 4864 142509 4868
rect 142525 4924 142589 4928
rect 142525 4868 142529 4924
rect 142529 4868 142585 4924
rect 142585 4868 142589 4924
rect 142525 4864 142589 4868
rect 283618 4924 283682 4928
rect 283618 4868 283622 4924
rect 283622 4868 283678 4924
rect 283678 4868 283682 4924
rect 283618 4864 283682 4868
rect 283698 4924 283762 4928
rect 283698 4868 283702 4924
rect 283702 4868 283758 4924
rect 283758 4868 283762 4924
rect 283698 4864 283762 4868
rect 283778 4924 283842 4928
rect 283778 4868 283782 4924
rect 283782 4868 283838 4924
rect 283838 4868 283842 4924
rect 283778 4864 283842 4868
rect 283858 4924 283922 4928
rect 283858 4868 283862 4924
rect 283862 4868 283918 4924
rect 283918 4868 283922 4924
rect 283858 4864 283922 4868
rect 71618 4380 71682 4384
rect 71618 4324 71622 4380
rect 71622 4324 71678 4380
rect 71678 4324 71682 4380
rect 71618 4320 71682 4324
rect 71698 4380 71762 4384
rect 71698 4324 71702 4380
rect 71702 4324 71758 4380
rect 71758 4324 71762 4380
rect 71698 4320 71762 4324
rect 71778 4380 71842 4384
rect 71778 4324 71782 4380
rect 71782 4324 71838 4380
rect 71838 4324 71842 4380
rect 71778 4320 71842 4324
rect 71858 4380 71922 4384
rect 71858 4324 71862 4380
rect 71862 4324 71918 4380
rect 71918 4324 71922 4380
rect 71858 4320 71922 4324
rect 212952 4380 213016 4384
rect 212952 4324 212956 4380
rect 212956 4324 213012 4380
rect 213012 4324 213016 4380
rect 212952 4320 213016 4324
rect 213032 4380 213096 4384
rect 213032 4324 213036 4380
rect 213036 4324 213092 4380
rect 213092 4324 213096 4380
rect 213032 4320 213096 4324
rect 213112 4380 213176 4384
rect 213112 4324 213116 4380
rect 213116 4324 213172 4380
rect 213172 4324 213176 4380
rect 213112 4320 213176 4324
rect 213192 4380 213256 4384
rect 213192 4324 213196 4380
rect 213196 4324 213252 4380
rect 213252 4324 213256 4380
rect 213192 4320 213256 4324
rect 354285 4380 354349 4384
rect 354285 4324 354289 4380
rect 354289 4324 354345 4380
rect 354345 4324 354349 4380
rect 354285 4320 354349 4324
rect 354365 4380 354429 4384
rect 354365 4324 354369 4380
rect 354369 4324 354425 4380
rect 354425 4324 354429 4380
rect 354365 4320 354429 4324
rect 354445 4380 354509 4384
rect 354445 4324 354449 4380
rect 354449 4324 354505 4380
rect 354505 4324 354509 4380
rect 354445 4320 354509 4324
rect 354525 4380 354589 4384
rect 354525 4324 354529 4380
rect 354529 4324 354585 4380
rect 354585 4324 354589 4380
rect 354525 4320 354589 4324
rect 60 4252 124 4316
rect 423628 4388 423692 4452
rect 60 3980 124 4044
rect 423628 4116 423692 4180
rect 142285 3836 142349 3840
rect 142285 3780 142289 3836
rect 142289 3780 142345 3836
rect 142345 3780 142349 3836
rect 142285 3776 142349 3780
rect 142365 3836 142429 3840
rect 142365 3780 142369 3836
rect 142369 3780 142425 3836
rect 142425 3780 142429 3836
rect 142365 3776 142429 3780
rect 142445 3836 142509 3840
rect 142445 3780 142449 3836
rect 142449 3780 142505 3836
rect 142505 3780 142509 3836
rect 142445 3776 142509 3780
rect 142525 3836 142589 3840
rect 142525 3780 142529 3836
rect 142529 3780 142585 3836
rect 142585 3780 142589 3836
rect 142525 3776 142589 3780
rect 283618 3836 283682 3840
rect 283618 3780 283622 3836
rect 283622 3780 283678 3836
rect 283678 3780 283682 3836
rect 283618 3776 283682 3780
rect 283698 3836 283762 3840
rect 283698 3780 283702 3836
rect 283702 3780 283758 3836
rect 283758 3780 283762 3836
rect 283698 3776 283762 3780
rect 283778 3836 283842 3840
rect 283778 3780 283782 3836
rect 283782 3780 283838 3836
rect 283838 3780 283842 3836
rect 283778 3776 283842 3780
rect 283858 3836 283922 3840
rect 283858 3780 283862 3836
rect 283862 3780 283918 3836
rect 283918 3780 283922 3836
rect 283858 3776 283922 3780
rect 71618 3292 71682 3296
rect 71618 3236 71622 3292
rect 71622 3236 71678 3292
rect 71678 3236 71682 3292
rect 71618 3232 71682 3236
rect 71698 3292 71762 3296
rect 71698 3236 71702 3292
rect 71702 3236 71758 3292
rect 71758 3236 71762 3292
rect 71698 3232 71762 3236
rect 71778 3292 71842 3296
rect 71778 3236 71782 3292
rect 71782 3236 71838 3292
rect 71838 3236 71842 3292
rect 71778 3232 71842 3236
rect 71858 3292 71922 3296
rect 71858 3236 71862 3292
rect 71862 3236 71918 3292
rect 71918 3236 71922 3292
rect 71858 3232 71922 3236
rect 212952 3292 213016 3296
rect 212952 3236 212956 3292
rect 212956 3236 213012 3292
rect 213012 3236 213016 3292
rect 212952 3232 213016 3236
rect 213032 3292 213096 3296
rect 213032 3236 213036 3292
rect 213036 3236 213092 3292
rect 213092 3236 213096 3292
rect 213032 3232 213096 3236
rect 213112 3292 213176 3296
rect 213112 3236 213116 3292
rect 213116 3236 213172 3292
rect 213172 3236 213176 3292
rect 213112 3232 213176 3236
rect 213192 3292 213256 3296
rect 213192 3236 213196 3292
rect 213196 3236 213252 3292
rect 213252 3236 213256 3292
rect 213192 3232 213256 3236
rect 354285 3292 354349 3296
rect 354285 3236 354289 3292
rect 354289 3236 354345 3292
rect 354345 3236 354349 3292
rect 354285 3232 354349 3236
rect 354365 3292 354429 3296
rect 354365 3236 354369 3292
rect 354369 3236 354425 3292
rect 354425 3236 354429 3292
rect 354365 3232 354429 3236
rect 354445 3292 354509 3296
rect 354445 3236 354449 3292
rect 354449 3236 354505 3292
rect 354505 3236 354509 3292
rect 354445 3232 354509 3236
rect 354525 3292 354589 3296
rect 354525 3236 354529 3292
rect 354529 3236 354585 3292
rect 354585 3236 354589 3292
rect 354525 3232 354589 3236
rect 142285 2748 142349 2752
rect 142285 2692 142289 2748
rect 142289 2692 142345 2748
rect 142345 2692 142349 2748
rect 142285 2688 142349 2692
rect 142365 2748 142429 2752
rect 142365 2692 142369 2748
rect 142369 2692 142425 2748
rect 142425 2692 142429 2748
rect 142365 2688 142429 2692
rect 142445 2748 142509 2752
rect 142445 2692 142449 2748
rect 142449 2692 142505 2748
rect 142505 2692 142509 2748
rect 142445 2688 142509 2692
rect 142525 2748 142589 2752
rect 142525 2692 142529 2748
rect 142529 2692 142585 2748
rect 142585 2692 142589 2748
rect 142525 2688 142589 2692
rect 283618 2748 283682 2752
rect 283618 2692 283622 2748
rect 283622 2692 283678 2748
rect 283678 2692 283682 2748
rect 283618 2688 283682 2692
rect 283698 2748 283762 2752
rect 283698 2692 283702 2748
rect 283702 2692 283758 2748
rect 283758 2692 283762 2748
rect 283698 2688 283762 2692
rect 283778 2748 283842 2752
rect 283778 2692 283782 2748
rect 283782 2692 283838 2748
rect 283838 2692 283842 2748
rect 283778 2688 283842 2692
rect 283858 2748 283922 2752
rect 283858 2692 283862 2748
rect 283862 2692 283918 2748
rect 283918 2692 283922 2748
rect 283858 2688 283922 2692
rect 71618 2204 71682 2208
rect 71618 2148 71622 2204
rect 71622 2148 71678 2204
rect 71678 2148 71682 2204
rect 71618 2144 71682 2148
rect 71698 2204 71762 2208
rect 71698 2148 71702 2204
rect 71702 2148 71758 2204
rect 71758 2148 71762 2204
rect 71698 2144 71762 2148
rect 71778 2204 71842 2208
rect 71778 2148 71782 2204
rect 71782 2148 71838 2204
rect 71838 2148 71842 2204
rect 71778 2144 71842 2148
rect 71858 2204 71922 2208
rect 71858 2148 71862 2204
rect 71862 2148 71918 2204
rect 71918 2148 71922 2204
rect 71858 2144 71922 2148
rect 60 2076 124 2140
rect 212952 2204 213016 2208
rect 212952 2148 212956 2204
rect 212956 2148 213012 2204
rect 213012 2148 213016 2204
rect 212952 2144 213016 2148
rect 213032 2204 213096 2208
rect 213032 2148 213036 2204
rect 213036 2148 213092 2204
rect 213092 2148 213096 2204
rect 213032 2144 213096 2148
rect 213112 2204 213176 2208
rect 213112 2148 213116 2204
rect 213116 2148 213172 2204
rect 213172 2148 213176 2204
rect 213112 2144 213176 2148
rect 213192 2204 213256 2208
rect 213192 2148 213196 2204
rect 213196 2148 213252 2204
rect 213252 2148 213256 2204
rect 213192 2144 213256 2148
rect 354285 2204 354349 2208
rect 354285 2148 354289 2204
rect 354289 2148 354345 2204
rect 354345 2148 354349 2204
rect 354285 2144 354349 2148
rect 354365 2204 354429 2208
rect 354365 2148 354369 2204
rect 354369 2148 354425 2204
rect 354425 2148 354429 2204
rect 354365 2144 354429 2148
rect 354445 2204 354509 2208
rect 354445 2148 354449 2204
rect 354449 2148 354505 2204
rect 354505 2148 354509 2204
rect 354445 2144 354509 2148
rect 354525 2204 354589 2208
rect 354525 2148 354529 2204
rect 354529 2148 354585 2204
rect 354585 2148 354589 2204
rect 354525 2144 354589 2148
rect 60 1804 124 1868
<< metal4 >>
rect 71610 7648 71931 7664
rect 71610 7584 71618 7648
rect 71682 7584 71698 7648
rect 71762 7584 71778 7648
rect 71842 7584 71858 7648
rect 71922 7584 71931 7648
rect 71610 6560 71931 7584
rect 71610 6496 71618 6560
rect 71682 6496 71698 6560
rect 71762 6496 71778 6560
rect 71842 6496 71858 6560
rect 71922 6496 71931 6560
rect 71610 5472 71931 6496
rect 71610 5408 71618 5472
rect 71682 5408 71698 5472
rect 71762 5408 71778 5472
rect 71842 5408 71858 5472
rect 71922 5408 71931 5472
rect 71610 4384 71931 5408
rect 71610 4320 71618 4384
rect 71682 4320 71698 4384
rect 71762 4320 71778 4384
rect 71842 4320 71858 4384
rect 71922 4320 71931 4384
rect 59 4316 125 4317
rect 59 4252 60 4316
rect 124 4252 125 4316
rect 59 4251 125 4252
rect 62 4045 122 4251
rect 59 4044 125 4045
rect 59 3980 60 4044
rect 124 3980 125 4044
rect 59 3979 125 3980
rect 71610 3296 71931 4320
rect 71610 3232 71618 3296
rect 71682 3232 71698 3296
rect 71762 3232 71778 3296
rect 71842 3232 71858 3296
rect 71922 3232 71931 3296
rect 71610 2208 71931 3232
rect 71610 2144 71618 2208
rect 71682 2144 71698 2208
rect 71762 2144 71778 2208
rect 71842 2144 71858 2208
rect 71922 2144 71931 2208
rect 59 2140 125 2141
rect 59 2076 60 2140
rect 124 2076 125 2140
rect 71610 2128 71931 2144
rect 142277 7104 142597 7664
rect 142277 7040 142285 7104
rect 142349 7040 142365 7104
rect 142429 7040 142445 7104
rect 142509 7040 142525 7104
rect 142589 7040 142597 7104
rect 142277 6016 142597 7040
rect 142277 5952 142285 6016
rect 142349 5952 142365 6016
rect 142429 5952 142445 6016
rect 142509 5952 142525 6016
rect 142589 5952 142597 6016
rect 142277 4928 142597 5952
rect 142277 4864 142285 4928
rect 142349 4864 142365 4928
rect 142429 4864 142445 4928
rect 142509 4864 142525 4928
rect 142589 4864 142597 4928
rect 142277 3840 142597 4864
rect 142277 3776 142285 3840
rect 142349 3776 142365 3840
rect 142429 3776 142445 3840
rect 142509 3776 142525 3840
rect 142589 3776 142597 3840
rect 142277 2752 142597 3776
rect 142277 2688 142285 2752
rect 142349 2688 142365 2752
rect 142429 2688 142445 2752
rect 142509 2688 142525 2752
rect 142589 2688 142597 2752
rect 142277 2128 142597 2688
rect 212944 7648 213264 7664
rect 212944 7584 212952 7648
rect 213016 7584 213032 7648
rect 213096 7584 213112 7648
rect 213176 7584 213192 7648
rect 213256 7584 213264 7648
rect 212944 6560 213264 7584
rect 212944 6496 212952 6560
rect 213016 6496 213032 6560
rect 213096 6496 213112 6560
rect 213176 6496 213192 6560
rect 213256 6496 213264 6560
rect 212944 5472 213264 6496
rect 212944 5408 212952 5472
rect 213016 5408 213032 5472
rect 213096 5408 213112 5472
rect 213176 5408 213192 5472
rect 213256 5408 213264 5472
rect 212944 4384 213264 5408
rect 212944 4320 212952 4384
rect 213016 4320 213032 4384
rect 213096 4320 213112 4384
rect 213176 4320 213192 4384
rect 213256 4320 213264 4384
rect 212944 3296 213264 4320
rect 212944 3232 212952 3296
rect 213016 3232 213032 3296
rect 213096 3232 213112 3296
rect 213176 3232 213192 3296
rect 213256 3232 213264 3296
rect 212944 2208 213264 3232
rect 212944 2144 212952 2208
rect 213016 2144 213032 2208
rect 213096 2144 213112 2208
rect 213176 2144 213192 2208
rect 213256 2144 213264 2208
rect 212944 2128 213264 2144
rect 283610 7104 283930 7664
rect 283610 7040 283618 7104
rect 283682 7040 283698 7104
rect 283762 7040 283778 7104
rect 283842 7040 283858 7104
rect 283922 7040 283930 7104
rect 283610 6016 283930 7040
rect 283610 5952 283618 6016
rect 283682 5952 283698 6016
rect 283762 5952 283778 6016
rect 283842 5952 283858 6016
rect 283922 5952 283930 6016
rect 283610 4928 283930 5952
rect 283610 4864 283618 4928
rect 283682 4864 283698 4928
rect 283762 4864 283778 4928
rect 283842 4864 283858 4928
rect 283922 4864 283930 4928
rect 283610 3840 283930 4864
rect 283610 3776 283618 3840
rect 283682 3776 283698 3840
rect 283762 3776 283778 3840
rect 283842 3776 283858 3840
rect 283922 3776 283930 3840
rect 283610 2752 283930 3776
rect 283610 2688 283618 2752
rect 283682 2688 283698 2752
rect 283762 2688 283778 2752
rect 283842 2688 283858 2752
rect 283922 2688 283930 2752
rect 283610 2128 283930 2688
rect 354277 7648 354597 7664
rect 354277 7584 354285 7648
rect 354349 7584 354365 7648
rect 354429 7584 354445 7648
rect 354509 7584 354525 7648
rect 354589 7584 354597 7648
rect 354277 6560 354597 7584
rect 354277 6496 354285 6560
rect 354349 6496 354365 6560
rect 354429 6496 354445 6560
rect 354509 6496 354525 6560
rect 354589 6496 354597 6560
rect 354277 5472 354597 6496
rect 354277 5408 354285 5472
rect 354349 5408 354365 5472
rect 354429 5408 354445 5472
rect 354509 5408 354525 5472
rect 354589 5408 354597 5472
rect 354277 4384 354597 5408
rect 423627 4452 423693 4453
rect 423627 4388 423628 4452
rect 423692 4388 423693 4452
rect 423627 4387 423693 4388
rect 354277 4320 354285 4384
rect 354349 4320 354365 4384
rect 354429 4320 354445 4384
rect 354509 4320 354525 4384
rect 354589 4320 354597 4384
rect 354277 3296 354597 4320
rect 423630 4181 423690 4387
rect 423627 4180 423693 4181
rect 423627 4116 423628 4180
rect 423692 4116 423693 4180
rect 423627 4115 423693 4116
rect 354277 3232 354285 3296
rect 354349 3232 354365 3296
rect 354429 3232 354445 3296
rect 354509 3232 354525 3296
rect 354589 3232 354597 3296
rect 354277 2208 354597 3232
rect 354277 2144 354285 2208
rect 354349 2144 354365 2208
rect 354429 2144 354445 2208
rect 354509 2144 354525 2208
rect 354589 2144 354597 2208
rect 354277 2128 354597 2144
rect 59 2075 125 2076
rect 62 1869 122 2075
rect 59 1868 125 1869
rect 59 1804 60 1868
rect 124 1804 125 1868
rect 59 1803 125 1804
use scs8hd_decap_3  PHY_0 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1104 0 -1 2720
box -38 -48 314 592
use scs8hd_decap_3  PHY_2
timestamp 1586364061
transform 1 0 1104 0 1 2720
box -38 -48 314 592
use scs8hd_decap_12  FILLER_0_3 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1380 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_15
timestamp 1586364061
transform 1 0 2484 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_3
timestamp 1586364061
transform 1 0 1380 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_15
timestamp 1586364061
transform 1 0 2484 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_20 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 3956 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_4  FILLER_0_27 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 3588 0 -1 2720
box -38 -48 406 592
use scs8hd_decap_12  FILLER_0_32
timestamp 1586364061
transform 1 0 4048 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_27
timestamp 1586364061
transform 1 0 3588 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_44
timestamp 1586364061
transform 1 0 5152 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_39
timestamp 1586364061
transform 1 0 4692 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_1_51 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 5796 0 1 2720
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_21
timestamp 1586364061
transform 1 0 6808 0 -1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_167
timestamp 1586364061
transform 1 0 6716 0 1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_56 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 6256 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_0_63
timestamp 1586364061
transform 1 0 6900 0 -1 2720
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_1_59 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 6532 0 1 2720
box -38 -48 222 592
use scs8hd_decap_12  FILLER_1_62
timestamp 1586364061
transform 1 0 6808 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_75
timestamp 1586364061
transform 1 0 8004 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_0_87
timestamp 1586364061
transform 1 0 9108 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_1_74
timestamp 1586364061
transform 1 0 7912 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_86
timestamp 1586364061
transform 1 0 9016 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_22
timestamp 1586364061
transform 1 0 9660 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_12  FILLER_0_94
timestamp 1586364061
transform 1 0 9752 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_106
timestamp 1586364061
transform 1 0 10856 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_98
timestamp 1586364061
transform 1 0 10120 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_23
timestamp 1586364061
transform 1 0 12512 0 -1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_168
timestamp 1586364061
transform 1 0 12328 0 1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_118
timestamp 1586364061
transform 1 0 11960 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_1_110
timestamp 1586364061
transform 1 0 11224 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_123
timestamp 1586364061
transform 1 0 12420 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_125
timestamp 1586364061
transform 1 0 12604 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_137
timestamp 1586364061
transform 1 0 13708 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_135
timestamp 1586364061
transform 1 0 13524 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_24
timestamp 1586364061
transform 1 0 15364 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_149
timestamp 1586364061
transform 1 0 14812 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_0_156
timestamp 1586364061
transform 1 0 15456 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_147
timestamp 1586364061
transform 1 0 14628 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_159
timestamp 1586364061
transform 1 0 15732 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_168
timestamp 1586364061
transform 1 0 16560 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_171
timestamp 1586364061
transform 1 0 16836 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_25
timestamp 1586364061
transform 1 0 18216 0 -1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_169
timestamp 1586364061
transform 1 0 17940 0 1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_180
timestamp 1586364061
transform 1 0 17664 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_0_187
timestamp 1586364061
transform 1 0 18308 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_184
timestamp 1586364061
transform 1 0 18032 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_196
timestamp 1586364061
transform 1 0 19136 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_199
timestamp 1586364061
transform 1 0 19412 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_0_211
timestamp 1586364061
transform 1 0 20516 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_1_208
timestamp 1586364061
transform 1 0 20240 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_26
timestamp 1586364061
transform 1 0 21068 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_12  FILLER_0_218
timestamp 1586364061
transform 1 0 21160 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_230
timestamp 1586364061
transform 1 0 22264 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_220
timestamp 1586364061
transform 1 0 21344 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_27
timestamp 1586364061
transform 1 0 23920 0 -1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_170
timestamp 1586364061
transform 1 0 23552 0 1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_242
timestamp 1586364061
transform 1 0 23368 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_0_249
timestamp 1586364061
transform 1 0 24012 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_232
timestamp 1586364061
transform 1 0 22448 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_245
timestamp 1586364061
transform 1 0 23644 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_261
timestamp 1586364061
transform 1 0 25116 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_257
timestamp 1586364061
transform 1 0 24748 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_28
timestamp 1586364061
transform 1 0 26772 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_273
timestamp 1586364061
transform 1 0 26220 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_0_280
timestamp 1586364061
transform 1 0 26864 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_269
timestamp 1586364061
transform 1 0 25852 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_281
timestamp 1586364061
transform 1 0 26956 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_292
timestamp 1586364061
transform 1 0 27968 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_293
timestamp 1586364061
transform 1 0 28060 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_29
timestamp 1586364061
transform 1 0 29624 0 -1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_171
timestamp 1586364061
transform 1 0 29164 0 1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_304
timestamp 1586364061
transform 1 0 29072 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_0_311
timestamp 1586364061
transform 1 0 29716 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_306
timestamp 1586364061
transform 1 0 29256 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_318
timestamp 1586364061
transform 1 0 30360 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_323
timestamp 1586364061
transform 1 0 30820 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_0_335
timestamp 1586364061
transform 1 0 31924 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_1_330
timestamp 1586364061
transform 1 0 31464 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_30
timestamp 1586364061
transform 1 0 32476 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_12  FILLER_0_342
timestamp 1586364061
transform 1 0 32568 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_354
timestamp 1586364061
transform 1 0 33672 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_342
timestamp 1586364061
transform 1 0 32568 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_354
timestamp 1586364061
transform 1 0 33672 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_31
timestamp 1586364061
transform 1 0 35328 0 -1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_172
timestamp 1586364061
transform 1 0 34776 0 1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_366
timestamp 1586364061
transform 1 0 34776 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_0_373
timestamp 1586364061
transform 1 0 35420 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_367
timestamp 1586364061
transform 1 0 34868 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_385
timestamp 1586364061
transform 1 0 36524 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_379
timestamp 1586364061
transform 1 0 35972 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_391
timestamp 1586364061
transform 1 0 37076 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_32
timestamp 1586364061
transform 1 0 38180 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_397
timestamp 1586364061
transform 1 0 37628 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_0_404
timestamp 1586364061
transform 1 0 38272 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_403
timestamp 1586364061
transform 1 0 38180 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_173
timestamp 1586364061
transform 1 0 40388 0 1 2720
box -38 -48 130 592
use scs8hd_decap_12  FILLER_0_416
timestamp 1586364061
transform 1 0 39376 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_0_428
timestamp 1586364061
transform 1 0 40480 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_1_415
timestamp 1586364061
transform 1 0 39284 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_428
timestamp 1586364061
transform 1 0 40480 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_33
timestamp 1586364061
transform 1 0 41032 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_12  FILLER_0_435
timestamp 1586364061
transform 1 0 41124 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_440
timestamp 1586364061
transform 1 0 41584 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_447
timestamp 1586364061
transform 1 0 42228 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_0_459
timestamp 1586364061
transform 1 0 43332 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_1_452
timestamp 1586364061
transform 1 0 42688 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_34
timestamp 1586364061
transform 1 0 43884 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_12  FILLER_0_466
timestamp 1586364061
transform 1 0 43976 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_478
timestamp 1586364061
transform 1 0 45080 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_464
timestamp 1586364061
transform 1 0 43792 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_476
timestamp 1586364061
transform 1 0 44896 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_35
timestamp 1586364061
transform 1 0 46736 0 -1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_174
timestamp 1586364061
transform 1 0 46000 0 1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_490
timestamp 1586364061
transform 1 0 46184 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_0_497
timestamp 1586364061
transform 1 0 46828 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_489
timestamp 1586364061
transform 1 0 46092 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_509
timestamp 1586364061
transform 1 0 47932 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_501
timestamp 1586364061
transform 1 0 47196 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_513
timestamp 1586364061
transform 1 0 48300 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_36
timestamp 1586364061
transform 1 0 49588 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_521
timestamp 1586364061
transform 1 0 49036 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_0_528
timestamp 1586364061
transform 1 0 49680 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_525
timestamp 1586364061
transform 1 0 49404 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_175
timestamp 1586364061
transform 1 0 51612 0 1 2720
box -38 -48 130 592
use scs8hd_decap_12  FILLER_0_540
timestamp 1586364061
transform 1 0 50784 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_0_552
timestamp 1586364061
transform 1 0 51888 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_1_537
timestamp 1586364061
transform 1 0 50508 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_550
timestamp 1586364061
transform 1 0 51704 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_37
timestamp 1586364061
transform 1 0 52440 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_12  FILLER_0_559
timestamp 1586364061
transform 1 0 52532 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_562
timestamp 1586364061
transform 1 0 52808 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_571
timestamp 1586364061
transform 1 0 53636 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_0_583
timestamp 1586364061
transform 1 0 54740 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_1_574
timestamp 1586364061
transform 1 0 53912 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_586
timestamp 1586364061
transform 1 0 55016 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_38
timestamp 1586364061
transform 1 0 55292 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_12  FILLER_0_590
timestamp 1586364061
transform 1 0 55384 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_602
timestamp 1586364061
transform 1 0 56488 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_598
timestamp 1586364061
transform 1 0 56120 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_39
timestamp 1586364061
transform 1 0 58144 0 -1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_176
timestamp 1586364061
transform 1 0 57224 0 1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_614
timestamp 1586364061
transform 1 0 57592 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_0_621
timestamp 1586364061
transform 1 0 58236 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_611
timestamp 1586364061
transform 1 0 57316 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_623
timestamp 1586364061
transform 1 0 58420 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_633
timestamp 1586364061
transform 1 0 59340 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_635
timestamp 1586364061
transform 1 0 59524 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_40
timestamp 1586364061
transform 1 0 60996 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_645
timestamp 1586364061
transform 1 0 60444 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_0_652
timestamp 1586364061
transform 1 0 61088 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_647
timestamp 1586364061
transform 1 0 60628 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_659
timestamp 1586364061
transform 1 0 61732 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_177
timestamp 1586364061
transform 1 0 62836 0 1 2720
box -38 -48 130 592
use scs8hd_decap_12  FILLER_0_664
timestamp 1586364061
transform 1 0 62192 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_0_676
timestamp 1586364061
transform 1 0 63296 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_1_672
timestamp 1586364061
transform 1 0 62928 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_41
timestamp 1586364061
transform 1 0 63848 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_12  FILLER_0_683
timestamp 1586364061
transform 1 0 63940 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_695
timestamp 1586364061
transform 1 0 65044 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_684
timestamp 1586364061
transform 1 0 64032 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_42
timestamp 1586364061
transform 1 0 66700 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_707
timestamp 1586364061
transform 1 0 66148 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_1_696
timestamp 1586364061
transform 1 0 65136 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_708
timestamp 1586364061
transform 1 0 66240 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_714
timestamp 1586364061
transform 1 0 66792 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_726
timestamp 1586364061
transform 1 0 67896 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_720
timestamp 1586364061
transform 1 0 67344 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_43
timestamp 1586364061
transform 1 0 69552 0 -1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_178
timestamp 1586364061
transform 1 0 68448 0 1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_738
timestamp 1586364061
transform 1 0 69000 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_0_745
timestamp 1586364061
transform 1 0 69644 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_733
timestamp 1586364061
transform 1 0 68540 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_745
timestamp 1586364061
transform 1 0 69644 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_757
timestamp 1586364061
transform 1 0 70748 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_757
timestamp 1586364061
transform 1 0 70748 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_44
timestamp 1586364061
transform 1 0 72404 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_769
timestamp 1586364061
transform 1 0 71852 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_0_776
timestamp 1586364061
transform 1 0 72496 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_769
timestamp 1586364061
transform 1 0 71852 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_781
timestamp 1586364061
transform 1 0 72956 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_179
timestamp 1586364061
transform 1 0 74060 0 1 2720
box -38 -48 130 592
use scs8hd_decap_12  FILLER_0_788
timestamp 1586364061
transform 1 0 73600 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_0_800
timestamp 1586364061
transform 1 0 74704 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_1_794
timestamp 1586364061
transform 1 0 74152 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_45
timestamp 1586364061
transform 1 0 75256 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_12  FILLER_0_807
timestamp 1586364061
transform 1 0 75348 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_819
timestamp 1586364061
transform 1 0 76452 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_806
timestamp 1586364061
transform 1 0 75256 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_818
timestamp 1586364061
transform 1 0 76360 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_46
timestamp 1586364061
transform 1 0 78108 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_831
timestamp 1586364061
transform 1 0 77556 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_0_838
timestamp 1586364061
transform 1 0 78200 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_830
timestamp 1586364061
transform 1 0 77464 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_180
timestamp 1586364061
transform 1 0 79672 0 1 2720
box -38 -48 130 592
use scs8hd_decap_12  FILLER_0_850
timestamp 1586364061
transform 1 0 79304 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_842
timestamp 1586364061
transform 1 0 78568 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_855
timestamp 1586364061
transform 1 0 79764 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_47
timestamp 1586364061
transform 1 0 80960 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_862
timestamp 1586364061
transform 1 0 80408 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_0_869
timestamp 1586364061
transform 1 0 81052 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_867
timestamp 1586364061
transform 1 0 80868 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_881
timestamp 1586364061
transform 1 0 82156 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_879
timestamp 1586364061
transform 1 0 81972 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_891
timestamp 1586364061
transform 1 0 83076 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_48
timestamp 1586364061
transform 1 0 83812 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_893
timestamp 1586364061
transform 1 0 83260 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_0_900
timestamp 1586364061
transform 1 0 83904 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_903
timestamp 1586364061
transform 1 0 84180 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_181
timestamp 1586364061
transform 1 0 85284 0 1 2720
box -38 -48 130 592
use scs8hd_decap_12  FILLER_0_912
timestamp 1586364061
transform 1 0 85008 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_0_924
timestamp 1586364061
transform 1 0 86112 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_1_916
timestamp 1586364061
transform 1 0 85376 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_49
timestamp 1586364061
transform 1 0 86664 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_12  FILLER_0_931
timestamp 1586364061
transform 1 0 86756 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_943
timestamp 1586364061
transform 1 0 87860 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_928
timestamp 1586364061
transform 1 0 86480 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_940
timestamp 1586364061
transform 1 0 87584 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_50
timestamp 1586364061
transform 1 0 89516 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_955
timestamp 1586364061
transform 1 0 88964 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_0_962
timestamp 1586364061
transform 1 0 89608 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_952
timestamp 1586364061
transform 1 0 88688 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_182
timestamp 1586364061
transform 1 0 90896 0 1 2720
box -38 -48 130 592
use scs8hd_decap_12  FILLER_0_974
timestamp 1586364061
transform 1 0 90712 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_964
timestamp 1586364061
transform 1 0 89792 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_977
timestamp 1586364061
transform 1 0 90988 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_51
timestamp 1586364061
transform 1 0 92368 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_986
timestamp 1586364061
transform 1 0 91816 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_0_993
timestamp 1586364061
transform 1 0 92460 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_989
timestamp 1586364061
transform 1 0 92092 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_1005
timestamp 1586364061
transform 1 0 93564 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_1001
timestamp 1586364061
transform 1 0 93196 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_1013
timestamp 1586364061
transform 1 0 94300 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_52
timestamp 1586364061
transform 1 0 95220 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_1017
timestamp 1586364061
transform 1 0 94668 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_0_1024
timestamp 1586364061
transform 1 0 95312 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_1025
timestamp 1586364061
transform 1 0 95404 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_183
timestamp 1586364061
transform 1 0 96508 0 1 2720
box -38 -48 130 592
use scs8hd_decap_12  FILLER_0_1036
timestamp 1586364061
transform 1 0 96416 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_0_1048
timestamp 1586364061
transform 1 0 97520 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_1_1038
timestamp 1586364061
transform 1 0 96600 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_1050
timestamp 1586364061
transform 1 0 97704 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_53
timestamp 1586364061
transform 1 0 98072 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_12  FILLER_0_1055
timestamp 1586364061
transform 1 0 98164 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_1067
timestamp 1586364061
transform 1 0 99268 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_1062
timestamp 1586364061
transform 1 0 98808 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_54
timestamp 1586364061
transform 1 0 100924 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_1079
timestamp 1586364061
transform 1 0 100372 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_0_1086
timestamp 1586364061
transform 1 0 101016 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_1074
timestamp 1586364061
transform 1 0 99912 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_1086
timestamp 1586364061
transform 1 0 101016 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_184
timestamp 1586364061
transform 1 0 102120 0 1 2720
box -38 -48 130 592
use scs8hd_decap_12  FILLER_0_1098
timestamp 1586364061
transform 1 0 102120 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_1099
timestamp 1586364061
transform 1 0 102212 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_55
timestamp 1586364061
transform 1 0 103776 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_1110
timestamp 1586364061
transform 1 0 103224 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_0_1117
timestamp 1586364061
transform 1 0 103868 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_1111
timestamp 1586364061
transform 1 0 103316 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_1123
timestamp 1586364061
transform 1 0 104420 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_1129
timestamp 1586364061
transform 1 0 104972 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_0_1141
timestamp 1586364061
transform 1 0 106076 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_1_1135
timestamp 1586364061
transform 1 0 105524 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_56
timestamp 1586364061
transform 1 0 106628 0 -1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_185
timestamp 1586364061
transform 1 0 107732 0 1 2720
box -38 -48 130 592
use scs8hd_decap_12  FILLER_0_1148
timestamp 1586364061
transform 1 0 106720 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_1147
timestamp 1586364061
transform 1 0 106628 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_1160
timestamp 1586364061
transform 1 0 107824 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_0_1172
timestamp 1586364061
transform 1 0 108928 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_1_1160
timestamp 1586364061
transform 1 0 107824 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_1172
timestamp 1586364061
transform 1 0 108928 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_57
timestamp 1586364061
transform 1 0 109480 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_12  FILLER_0_1179
timestamp 1586364061
transform 1 0 109572 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_1191
timestamp 1586364061
transform 1 0 110676 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_1184
timestamp 1586364061
transform 1 0 110032 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_58
timestamp 1586364061
transform 1 0 112332 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_1203
timestamp 1586364061
transform 1 0 111780 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_0_1210
timestamp 1586364061
transform 1 0 112424 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_1196
timestamp 1586364061
transform 1 0 111136 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_1208
timestamp 1586364061
transform 1 0 112240 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_186
timestamp 1586364061
transform 1 0 113344 0 1 2720
box -38 -48 130 592
use scs8hd_decap_12  FILLER_0_1222
timestamp 1586364061
transform 1 0 113528 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_1221
timestamp 1586364061
transform 1 0 113436 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_59
timestamp 1586364061
transform 1 0 115184 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_1234
timestamp 1586364061
transform 1 0 114632 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_0_1241
timestamp 1586364061
transform 1 0 115276 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_1233
timestamp 1586364061
transform 1 0 114540 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_1245
timestamp 1586364061
transform 1 0 115644 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_1253
timestamp 1586364061
transform 1 0 116380 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_0_1265
timestamp 1586364061
transform 1 0 117484 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_1_1257
timestamp 1586364061
transform 1 0 116748 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_60
timestamp 1586364061
transform 1 0 118036 0 -1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_187
timestamp 1586364061
transform 1 0 118956 0 1 2720
box -38 -48 130 592
use scs8hd_decap_12  FILLER_0_1272
timestamp 1586364061
transform 1 0 118128 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_1284
timestamp 1586364061
transform 1 0 119232 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_1269
timestamp 1586364061
transform 1 0 117852 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_1282
timestamp 1586364061
transform 1 0 119048 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_61
timestamp 1586364061
transform 1 0 120888 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_1296
timestamp 1586364061
transform 1 0 120336 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_1_1294
timestamp 1586364061
transform 1 0 120152 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_1303
timestamp 1586364061
transform 1 0 120980 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_1315
timestamp 1586364061
transform 1 0 122084 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_1306
timestamp 1586364061
transform 1 0 121256 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_1318
timestamp 1586364061
transform 1 0 122360 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_62
timestamp 1586364061
transform 1 0 123740 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_1327
timestamp 1586364061
transform 1 0 123188 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_0_1334
timestamp 1586364061
transform 1 0 123832 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_1330
timestamp 1586364061
transform 1 0 123464 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_188
timestamp 1586364061
transform 1 0 124568 0 1 2720
box -38 -48 130 592
use scs8hd_decap_12  FILLER_0_1346
timestamp 1586364061
transform 1 0 124936 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_1343
timestamp 1586364061
transform 1 0 124660 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_1355
timestamp 1586364061
transform 1 0 125764 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_63
timestamp 1586364061
transform 1 0 126592 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_1358
timestamp 1586364061
transform 1 0 126040 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_0_1365
timestamp 1586364061
transform 1 0 126684 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_1367
timestamp 1586364061
transform 1 0 126868 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_1377
timestamp 1586364061
transform 1 0 127788 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_0_1389
timestamp 1586364061
transform 1 0 128892 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_1_1379
timestamp 1586364061
transform 1 0 127972 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_1391
timestamp 1586364061
transform 1 0 129076 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_64
timestamp 1586364061
transform 1 0 129444 0 -1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_189
timestamp 1586364061
transform 1 0 130180 0 1 2720
box -38 -48 130 592
use scs8hd_decap_12  FILLER_0_1396
timestamp 1586364061
transform 1 0 129536 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_1408
timestamp 1586364061
transform 1 0 130640 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_1404
timestamp 1586364061
transform 1 0 130272 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_65
timestamp 1586364061
transform 1 0 132296 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_1420
timestamp 1586364061
transform 1 0 131744 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_1_1416
timestamp 1586364061
transform 1 0 131376 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_1427
timestamp 1586364061
transform 1 0 132388 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_1439
timestamp 1586364061
transform 1 0 133492 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_1428
timestamp 1586364061
transform 1 0 132480 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_1440
timestamp 1586364061
transform 1 0 133584 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_66
timestamp 1586364061
transform 1 0 135148 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_1451
timestamp 1586364061
transform 1 0 134596 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_0_1458
timestamp 1586364061
transform 1 0 135240 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_1452
timestamp 1586364061
transform 1 0 134688 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_190
timestamp 1586364061
transform 1 0 135792 0 1 2720
box -38 -48 130 592
use scs8hd_decap_12  FILLER_0_1470
timestamp 1586364061
transform 1 0 136344 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_1465
timestamp 1586364061
transform 1 0 135884 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_1477
timestamp 1586364061
transform 1 0 136988 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_67
timestamp 1586364061
transform 1 0 138000 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_1482
timestamp 1586364061
transform 1 0 137448 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_0_1489
timestamp 1586364061
transform 1 0 138092 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_1489
timestamp 1586364061
transform 1 0 138092 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_1501
timestamp 1586364061
transform 1 0 139196 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_0_1513
timestamp 1586364061
transform 1 0 140300 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_1_1501
timestamp 1586364061
transform 1 0 139196 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_1513
timestamp 1586364061
transform 1 0 140300 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_68
timestamp 1586364061
transform 1 0 140852 0 -1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_191
timestamp 1586364061
transform 1 0 141404 0 1 2720
box -38 -48 130 592
use scs8hd_decap_12  FILLER_0_1520
timestamp 1586364061
transform 1 0 140944 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_1532
timestamp 1586364061
transform 1 0 142048 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_1526
timestamp 1586364061
transform 1 0 141496 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_69
timestamp 1586364061
transform 1 0 143704 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_1544
timestamp 1586364061
transform 1 0 143152 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_0_1551
timestamp 1586364061
transform 1 0 143796 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_1538
timestamp 1586364061
transform 1 0 142600 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_1550
timestamp 1586364061
transform 1 0 143704 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_1563
timestamp 1586364061
transform 1 0 144900 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_1562
timestamp 1586364061
transform 1 0 144808 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_70
timestamp 1586364061
transform 1 0 146556 0 -1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_192
timestamp 1586364061
transform 1 0 147016 0 1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_1575
timestamp 1586364061
transform 1 0 146004 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_0_1582
timestamp 1586364061
transform 1 0 146648 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_1574
timestamp 1586364061
transform 1 0 145912 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_1587
timestamp 1586364061
transform 1 0 147108 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_1594
timestamp 1586364061
transform 1 0 147752 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_1599
timestamp 1586364061
transform 1 0 148212 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_71
timestamp 1586364061
transform 1 0 149408 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_1606
timestamp 1586364061
transform 1 0 148856 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_0_1613
timestamp 1586364061
transform 1 0 149500 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_1611
timestamp 1586364061
transform 1 0 149316 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_1623
timestamp 1586364061
transform 1 0 150420 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_1625
timestamp 1586364061
transform 1 0 150604 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_0_1637
timestamp 1586364061
transform 1 0 151708 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_1_1635
timestamp 1586364061
transform 1 0 151524 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_72
timestamp 1586364061
transform 1 0 152260 0 -1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_193
timestamp 1586364061
transform 1 0 152628 0 1 2720
box -38 -48 130 592
use scs8hd_decap_12  FILLER_0_1644
timestamp 1586364061
transform 1 0 152352 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_1656
timestamp 1586364061
transform 1 0 153456 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_1648
timestamp 1586364061
transform 1 0 152720 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_73
timestamp 1586364061
transform 1 0 155112 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_1668
timestamp 1586364061
transform 1 0 154560 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_0_1675
timestamp 1586364061
transform 1 0 155204 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_1660
timestamp 1586364061
transform 1 0 153824 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_1672
timestamp 1586364061
transform 1 0 154928 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_1687
timestamp 1586364061
transform 1 0 156308 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_1684
timestamp 1586364061
transform 1 0 156032 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_74
timestamp 1586364061
transform 1 0 157964 0 -1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_194
timestamp 1586364061
transform 1 0 158240 0 1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_1699
timestamp 1586364061
transform 1 0 157412 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_0_1706
timestamp 1586364061
transform 1 0 158056 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_1696
timestamp 1586364061
transform 1 0 157136 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_1709
timestamp 1586364061
transform 1 0 158332 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_1718
timestamp 1586364061
transform 1 0 159160 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_0_1730
timestamp 1586364061
transform 1 0 160264 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_1_1721
timestamp 1586364061
transform 1 0 159436 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_75
timestamp 1586364061
transform 1 0 160816 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_12  FILLER_0_1737
timestamp 1586364061
transform 1 0 160908 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_1733
timestamp 1586364061
transform 1 0 160540 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_1745
timestamp 1586364061
transform 1 0 161644 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_1749
timestamp 1586364061
transform 1 0 162012 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_0_1761
timestamp 1586364061
transform 1 0 163116 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_1_1757
timestamp 1586364061
transform 1 0 162748 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_76
timestamp 1586364061
transform 1 0 163668 0 -1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_195
timestamp 1586364061
transform 1 0 163852 0 1 2720
box -38 -48 130 592
use scs8hd_decap_12  FILLER_0_1768
timestamp 1586364061
transform 1 0 163760 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_1780
timestamp 1586364061
transform 1 0 164864 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_1770
timestamp 1586364061
transform 1 0 163944 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_1782
timestamp 1586364061
transform 1 0 165048 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_77
timestamp 1586364061
transform 1 0 166520 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_1792
timestamp 1586364061
transform 1 0 165968 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_0_1799
timestamp 1586364061
transform 1 0 166612 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_1794
timestamp 1586364061
transform 1 0 166152 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_1811
timestamp 1586364061
transform 1 0 167716 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_1806
timestamp 1586364061
transform 1 0 167256 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_1818
timestamp 1586364061
transform 1 0 168360 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_78
timestamp 1586364061
transform 1 0 169372 0 -1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_196
timestamp 1586364061
transform 1 0 169464 0 1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_1823
timestamp 1586364061
transform 1 0 168820 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_0_1830
timestamp 1586364061
transform 1 0 169464 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_1831
timestamp 1586364061
transform 1 0 169556 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_1842
timestamp 1586364061
transform 1 0 170568 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_0_1854
timestamp 1586364061
transform 1 0 171672 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_1_1843
timestamp 1586364061
transform 1 0 170660 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_1855
timestamp 1586364061
transform 1 0 171764 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_79
timestamp 1586364061
transform 1 0 172224 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_12  FILLER_0_1861
timestamp 1586364061
transform 1 0 172316 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_1867
timestamp 1586364061
transform 1 0 172868 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_1873
timestamp 1586364061
transform 1 0 173420 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_0_1885
timestamp 1586364061
transform 1 0 174524 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_1_1879
timestamp 1586364061
transform 1 0 173972 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_80
timestamp 1586364061
transform 1 0 175076 0 -1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_197
timestamp 1586364061
transform 1 0 175076 0 1 2720
box -38 -48 130 592
use scs8hd_decap_12  FILLER_0_1892
timestamp 1586364061
transform 1 0 175168 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_1904
timestamp 1586364061
transform 1 0 176272 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_1892
timestamp 1586364061
transform 1 0 175168 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_1904
timestamp 1586364061
transform 1 0 176272 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_81
timestamp 1586364061
transform 1 0 177928 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_1916
timestamp 1586364061
transform 1 0 177376 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_0_1923
timestamp 1586364061
transform 1 0 178020 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_1916
timestamp 1586364061
transform 1 0 177376 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_1935
timestamp 1586364061
transform 1 0 179124 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_1928
timestamp 1586364061
transform 1 0 178480 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_1940
timestamp 1586364061
transform 1 0 179584 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_82
timestamp 1586364061
transform 1 0 180780 0 -1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_198
timestamp 1586364061
transform 1 0 180688 0 1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_1947
timestamp 1586364061
transform 1 0 180228 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_0_1954
timestamp 1586364061
transform 1 0 180872 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_1953
timestamp 1586364061
transform 1 0 180780 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_1966
timestamp 1586364061
transform 1 0 181976 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_0_1978
timestamp 1586364061
transform 1 0 183080 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_1_1965
timestamp 1586364061
transform 1 0 181884 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_1977
timestamp 1586364061
transform 1 0 182988 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_83
timestamp 1586364061
transform 1 0 183632 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_12  FILLER_0_1985
timestamp 1586364061
transform 1 0 183724 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_1997
timestamp 1586364061
transform 1 0 184828 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_1989
timestamp 1586364061
transform 1 0 184092 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_84
timestamp 1586364061
transform 1 0 186484 0 -1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_199
timestamp 1586364061
transform 1 0 186300 0 1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_2009
timestamp 1586364061
transform 1 0 185932 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_1_2001
timestamp 1586364061
transform 1 0 185196 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_2014
timestamp 1586364061
transform 1 0 186392 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_2016
timestamp 1586364061
transform 1 0 186576 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_2028
timestamp 1586364061
transform 1 0 187680 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_2026
timestamp 1586364061
transform 1 0 187496 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_85
timestamp 1586364061
transform 1 0 189336 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_2040
timestamp 1586364061
transform 1 0 188784 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_0_2047
timestamp 1586364061
transform 1 0 189428 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_2038
timestamp 1586364061
transform 1 0 188600 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_2050
timestamp 1586364061
transform 1 0 189704 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_2059
timestamp 1586364061
transform 1 0 190532 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_2062
timestamp 1586364061
transform 1 0 190808 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_86
timestamp 1586364061
transform 1 0 192188 0 -1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_200
timestamp 1586364061
transform 1 0 191912 0 1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_2071
timestamp 1586364061
transform 1 0 191636 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_0_2078
timestamp 1586364061
transform 1 0 192280 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_2075
timestamp 1586364061
transform 1 0 192004 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_2090
timestamp 1586364061
transform 1 0 193384 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_0_2102
timestamp 1586364061
transform 1 0 194488 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_1_2087
timestamp 1586364061
transform 1 0 193108 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_2099
timestamp 1586364061
transform 1 0 194212 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_87
timestamp 1586364061
transform 1 0 195040 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_12  FILLER_0_2109
timestamp 1586364061
transform 1 0 195132 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_2121
timestamp 1586364061
transform 1 0 196236 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_2111
timestamp 1586364061
transform 1 0 195316 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_88
timestamp 1586364061
transform 1 0 197892 0 -1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_201
timestamp 1586364061
transform 1 0 197524 0 1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_2133
timestamp 1586364061
transform 1 0 197340 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_0_2140
timestamp 1586364061
transform 1 0 197984 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_2123
timestamp 1586364061
transform 1 0 196420 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_2136
timestamp 1586364061
transform 1 0 197616 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_2152
timestamp 1586364061
transform 1 0 199088 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_2148
timestamp 1586364061
transform 1 0 198720 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_89
timestamp 1586364061
transform 1 0 200744 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_2164
timestamp 1586364061
transform 1 0 200192 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_0_2171
timestamp 1586364061
transform 1 0 200836 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_2160
timestamp 1586364061
transform 1 0 199824 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_2172
timestamp 1586364061
transform 1 0 200928 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_2183
timestamp 1586364061
transform 1 0 201940 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_2184
timestamp 1586364061
transform 1 0 202032 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_90
timestamp 1586364061
transform 1 0 203596 0 -1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_202
timestamp 1586364061
transform 1 0 203136 0 1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_2195
timestamp 1586364061
transform 1 0 203044 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_0_2202
timestamp 1586364061
transform 1 0 203688 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_2197
timestamp 1586364061
transform 1 0 203228 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_2209
timestamp 1586364061
transform 1 0 204332 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_2214
timestamp 1586364061
transform 1 0 204792 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_0_2226
timestamp 1586364061
transform 1 0 205896 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_1_2221
timestamp 1586364061
transform 1 0 205436 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_91
timestamp 1586364061
transform 1 0 206448 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_12  FILLER_0_2233
timestamp 1586364061
transform 1 0 206540 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_2245
timestamp 1586364061
transform 1 0 207644 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_2233
timestamp 1586364061
transform 1 0 206540 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_2245
timestamp 1586364061
transform 1 0 207644 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_92
timestamp 1586364061
transform 1 0 209300 0 -1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_203
timestamp 1586364061
transform 1 0 208748 0 1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_2257
timestamp 1586364061
transform 1 0 208748 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_0_2264
timestamp 1586364061
transform 1 0 209392 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_2258
timestamp 1586364061
transform 1 0 208840 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_0_2276
timestamp 1586364061
transform 1 0 210496 0 -1 2720
box -38 -48 774 592
use scs8hd_decap_12  FILLER_1_2270
timestamp 1586364061
transform 1 0 209944 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_1_2282
timestamp 1586364061
transform 1 0 211048 0 1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_1_2289
timestamp 1586364061
transform 1 0 211692 0 1 2720
box -38 -48 222 592
use scs8hd_fill_1  FILLER_1_2286 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 211416 0 1 2720
box -38 -48 130 592
use scs8hd_fill_2  FILLER_0_2290
timestamp 1586364061
transform 1 0 211784 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_2286
timestamp 1586364061
transform 1 0 211416 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.LATCH_0_.latch_SLEEPB tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 211508 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__15__B
timestamp 1586364061
transform 1 0 211876 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__09__D
timestamp 1586364061
transform 1 0 211232 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__17__A
timestamp 1586364061
transform 1 0 211600 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__09__B
timestamp 1586364061
transform 1 0 211968 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_2293
timestamp 1586364061
transform 1 0 212060 0 1 2720
box -38 -48 222 592
use scs8hd_decap_3  FILLER_0_2299
timestamp 1586364061
transform 1 0 212612 0 -1 2720
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 212244 0 1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_93
timestamp 1586364061
transform 1 0 212152 0 -1 2720
box -38 -48 130 592
use scs8hd_buf_2  _17_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 212244 0 -1 2720
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.LATCH_0_.latch tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 212428 0 1 2720
box -38 -48 1050 592
use scs8hd_fill_2  FILLER_1_2308
timestamp 1586364061
transform 1 0 213440 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_2304
timestamp 1586364061
transform 1 0 213072 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__09__C
timestamp 1586364061
transform 1 0 212888 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__09__A
timestamp 1586364061
transform 1 0 213256 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_2316
timestamp 1586364061
transform 1 0 214176 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_2312
timestamp 1586364061
transform 1 0 213808 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_2317
timestamp 1586364061
transform 1 0 214268 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__15__D
timestamp 1586364061
transform 1 0 213992 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__15__A
timestamp 1586364061
transform 1 0 213624 0 1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_204
timestamp 1586364061
transform 1 0 214360 0 1 2720
box -38 -48 130 592
use scs8hd_and4_4  _09_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 213440 0 -1 2720
box -38 -48 866 592
use scs8hd_fill_1  FILLER_1_2326
timestamp 1586364061
transform 1 0 215096 0 1 2720
box -38 -48 130 592
use scs8hd_decap_4  FILLER_1_2322
timestamp 1586364061
transform 1 0 214728 0 1 2720
box -38 -48 406 592
use scs8hd_fill_1  FILLER_0_2326
timestamp 1586364061
transform 1 0 215096 0 -1 2720
box -38 -48 130 592
use scs8hd_fill_2  FILLER_0_2321
timestamp 1586364061
transform 1 0 214636 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__04__A
timestamp 1586364061
transform 1 0 214452 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__05__B
timestamp 1586364061
transform 1 0 215188 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__14__D
timestamp 1586364061
transform 1 0 214820 0 -1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_94
timestamp 1586364061
transform 1 0 215004 0 -1 2720
box -38 -48 130 592
use scs8hd_buf_1  _04_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 214452 0 1 2720
box -38 -48 314 592
use scs8hd_fill_2  FILLER_1_2329
timestamp 1586364061
transform 1 0 215372 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__05__C
timestamp 1586364061
transform 1 0 215556 0 1 2720
box -38 -48 222 592
use scs8hd_nor4_4  _14_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 215188 0 -1 2720
box -38 -48 1602 592
use scs8hd_nor4_4  _12_
timestamp 1586364061
transform 1 0 215740 0 1 2720
box -38 -48 1602 592
use scs8hd_diode_2  ANTENNA__08__A
timestamp 1586364061
transform 1 0 217488 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__14__C
timestamp 1586364061
transform 1 0 216936 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__14__A
timestamp 1586364061
transform 1 0 217304 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__14__B
timestamp 1586364061
transform 1 0 217672 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_2344
timestamp 1586364061
transform 1 0 216752 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_2348
timestamp 1586364061
transform 1 0 217120 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_2352
timestamp 1586364061
transform 1 0 217488 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_2350
timestamp 1586364061
transform 1 0 217304 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_2354
timestamp 1586364061
transform 1 0 217672 0 1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_95
timestamp 1586364061
transform 1 0 217856 0 -1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__12__D
timestamp 1586364061
transform 1 0 217856 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__12__B
timestamp 1586364061
transform 1 0 218224 0 1 2720
box -38 -48 222 592
use scs8hd_decap_12  FILLER_0_2357
timestamp 1586364061
transform 1 0 217948 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_0_2369
timestamp 1586364061
transform 1 0 219052 0 -1 2720
box -38 -48 590 592
use scs8hd_fill_2  FILLER_1_2358
timestamp 1586364061
transform 1 0 218040 0 1 2720
box -38 -48 222 592
use scs8hd_decap_8  FILLER_1_2362
timestamp 1586364061
transform 1 0 218408 0 1 2720
box -38 -48 774 592
use scs8hd_decap_3  FILLER_1_2370
timestamp 1586364061
transform 1 0 219144 0 1 2720
box -38 -48 314 592
use scs8hd_fill_2  FILLER_1_2375
timestamp 1586364061
transform 1 0 219604 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_2378
timestamp 1586364061
transform 1 0 219880 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_1  FILLER_0_2375
timestamp 1586364061
transform 1 0 219604 0 -1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 220064 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 219696 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 219420 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 219788 0 1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_205
timestamp 1586364061
transform 1 0 219972 0 1 2720
box -38 -48 130 592
use scs8hd_decap_3  FILLER_0_2388
timestamp 1586364061
transform 1 0 220800 0 -1 2720
box -38 -48 314 592
use scs8hd_decap_3  FILLER_0_2382
timestamp 1586364061
transform 1 0 220248 0 -1 2720
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer_TEB
timestamp 1586364061
transform 1 0 220524 0 -1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_96
timestamp 1586364061
transform 1 0 220708 0 -1 2720
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.LATCH_0_.latch
timestamp 1586364061
transform 1 0 220064 0 1 2720
box -38 -48 1050 592
use scs8hd_ebufn_1  logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 221260 0 -1 2720
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA_logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer_A
timestamp 1586364061
transform 1 0 221076 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_12  FILLER_0_2401
timestamp 1586364061
transform 1 0 221996 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_2391
timestamp 1586364061
transform 1 0 221076 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_2403
timestamp 1586364061
transform 1 0 222180 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_97
timestamp 1586364061
transform 1 0 223560 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_4  FILLER_0_2413
timestamp 1586364061
transform 1 0 223100 0 -1 2720
box -38 -48 406 592
use scs8hd_fill_1  FILLER_0_2417
timestamp 1586364061
transform 1 0 223468 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_12  FILLER_0_2419
timestamp 1586364061
transform 1 0 223652 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_2415
timestamp 1586364061
transform 1 0 223284 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_206
timestamp 1586364061
transform 1 0 225584 0 1 2720
box -38 -48 130 592
use scs8hd_decap_12  FILLER_0_2431
timestamp 1586364061
transform 1 0 224756 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_0_2443
timestamp 1586364061
transform 1 0 225860 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_1_2427
timestamp 1586364061
transform 1 0 224388 0 1 2720
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_1_2439
timestamp 1586364061
transform 1 0 225492 0 1 2720
box -38 -48 130 592
use scs8hd_decap_12  FILLER_1_2441
timestamp 1586364061
transform 1 0 225676 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_98
timestamp 1586364061
transform 1 0 226412 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_12  FILLER_0_2450
timestamp 1586364061
transform 1 0 226504 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_2453
timestamp 1586364061
transform 1 0 226780 0 1 2720
box -38 -48 1142 592
use scs8hd_buf_2  _21_
timestamp 1586364061
transform 1 0 228160 0 -1 2720
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__21__A
timestamp 1586364061
transform 1 0 228712 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_6  FILLER_0_2462
timestamp 1586364061
transform 1 0 227608 0 -1 2720
box -38 -48 590 592
use scs8hd_fill_2  FILLER_0_2472
timestamp 1586364061
transform 1 0 228528 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_0_2476
timestamp 1586364061
transform 1 0 228896 0 -1 2720
box -38 -48 406 592
use scs8hd_decap_12  FILLER_1_2465
timestamp 1586364061
transform 1 0 227884 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_2477
timestamp 1586364061
transform 1 0 228988 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_99
timestamp 1586364061
transform 1 0 229264 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_12  FILLER_0_2481
timestamp 1586364061
transform 1 0 229356 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_2493
timestamp 1586364061
transform 1 0 230460 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_2489
timestamp 1586364061
transform 1 0 230092 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_100
timestamp 1586364061
transform 1 0 232116 0 -1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_207
timestamp 1586364061
transform 1 0 231196 0 1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_2505
timestamp 1586364061
transform 1 0 231564 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_0_2512
timestamp 1586364061
transform 1 0 232208 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_2502
timestamp 1586364061
transform 1 0 231288 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_2514
timestamp 1586364061
transform 1 0 232392 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_2524
timestamp 1586364061
transform 1 0 233312 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_2526
timestamp 1586364061
transform 1 0 233496 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_101
timestamp 1586364061
transform 1 0 234968 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_2536
timestamp 1586364061
transform 1 0 234416 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_0_2543
timestamp 1586364061
transform 1 0 235060 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_2538
timestamp 1586364061
transform 1 0 234600 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_2550
timestamp 1586364061
transform 1 0 235704 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_208
timestamp 1586364061
transform 1 0 236808 0 1 2720
box -38 -48 130 592
use scs8hd_decap_12  FILLER_0_2555
timestamp 1586364061
transform 1 0 236164 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_0_2567
timestamp 1586364061
transform 1 0 237268 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_1_2563
timestamp 1586364061
transform 1 0 236900 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_102
timestamp 1586364061
transform 1 0 237820 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_12  FILLER_0_2574
timestamp 1586364061
transform 1 0 237912 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_2586
timestamp 1586364061
transform 1 0 239016 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_2575
timestamp 1586364061
transform 1 0 238004 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_103
timestamp 1586364061
transform 1 0 240672 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_2598
timestamp 1586364061
transform 1 0 240120 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_1_2587
timestamp 1586364061
transform 1 0 239108 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_2599
timestamp 1586364061
transform 1 0 240212 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_2605
timestamp 1586364061
transform 1 0 240764 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_2617
timestamp 1586364061
transform 1 0 241868 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_2611
timestamp 1586364061
transform 1 0 241316 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_104
timestamp 1586364061
transform 1 0 243524 0 -1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_209
timestamp 1586364061
transform 1 0 242420 0 1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_2629
timestamp 1586364061
transform 1 0 242972 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_0_2636
timestamp 1586364061
transform 1 0 243616 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_2624
timestamp 1586364061
transform 1 0 242512 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_2636
timestamp 1586364061
transform 1 0 243616 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_2648
timestamp 1586364061
transform 1 0 244720 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_2648
timestamp 1586364061
transform 1 0 244720 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_105
timestamp 1586364061
transform 1 0 246376 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_2660
timestamp 1586364061
transform 1 0 245824 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_0_2667
timestamp 1586364061
transform 1 0 246468 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_2660
timestamp 1586364061
transform 1 0 245824 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_2672
timestamp 1586364061
transform 1 0 246928 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_210
timestamp 1586364061
transform 1 0 248032 0 1 2720
box -38 -48 130 592
use scs8hd_decap_12  FILLER_0_2679
timestamp 1586364061
transform 1 0 247572 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_0_2691
timestamp 1586364061
transform 1 0 248676 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_1_2685
timestamp 1586364061
transform 1 0 248124 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_106
timestamp 1586364061
transform 1 0 249228 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_12  FILLER_0_2698
timestamp 1586364061
transform 1 0 249320 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_2710
timestamp 1586364061
transform 1 0 250424 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_2697
timestamp 1586364061
transform 1 0 249228 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_2709
timestamp 1586364061
transform 1 0 250332 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_107
timestamp 1586364061
transform 1 0 252080 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_2722
timestamp 1586364061
transform 1 0 251528 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_0_2729
timestamp 1586364061
transform 1 0 252172 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_2721
timestamp 1586364061
transform 1 0 251436 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_211
timestamp 1586364061
transform 1 0 253644 0 1 2720
box -38 -48 130 592
use scs8hd_decap_12  FILLER_0_2741
timestamp 1586364061
transform 1 0 253276 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_2733
timestamp 1586364061
transform 1 0 252540 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_2746
timestamp 1586364061
transform 1 0 253736 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_108
timestamp 1586364061
transform 1 0 254932 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_2753
timestamp 1586364061
transform 1 0 254380 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_0_2760
timestamp 1586364061
transform 1 0 255024 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_2758
timestamp 1586364061
transform 1 0 254840 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_2772
timestamp 1586364061
transform 1 0 256128 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_2770
timestamp 1586364061
transform 1 0 255944 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_2782
timestamp 1586364061
transform 1 0 257048 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_109
timestamp 1586364061
transform 1 0 257784 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_2784
timestamp 1586364061
transform 1 0 257232 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_0_2791
timestamp 1586364061
transform 1 0 257876 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_2794
timestamp 1586364061
transform 1 0 258152 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_212
timestamp 1586364061
transform 1 0 259256 0 1 2720
box -38 -48 130 592
use scs8hd_decap_12  FILLER_0_2803
timestamp 1586364061
transform 1 0 258980 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_0_2815
timestamp 1586364061
transform 1 0 260084 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_1_2807
timestamp 1586364061
transform 1 0 259348 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_110
timestamp 1586364061
transform 1 0 260636 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_12  FILLER_0_2822
timestamp 1586364061
transform 1 0 260728 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_2834
timestamp 1586364061
transform 1 0 261832 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_2819
timestamp 1586364061
transform 1 0 260452 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_2831
timestamp 1586364061
transform 1 0 261556 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_111
timestamp 1586364061
transform 1 0 263488 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_2846
timestamp 1586364061
transform 1 0 262936 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_0_2853
timestamp 1586364061
transform 1 0 263580 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_2843
timestamp 1586364061
transform 1 0 262660 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_213
timestamp 1586364061
transform 1 0 264868 0 1 2720
box -38 -48 130 592
use scs8hd_decap_12  FILLER_0_2865
timestamp 1586364061
transform 1 0 264684 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_2855
timestamp 1586364061
transform 1 0 263764 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_2868
timestamp 1586364061
transform 1 0 264960 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_112
timestamp 1586364061
transform 1 0 266340 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_2877
timestamp 1586364061
transform 1 0 265788 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_0_2884
timestamp 1586364061
transform 1 0 266432 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_2880
timestamp 1586364061
transform 1 0 266064 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_2896
timestamp 1586364061
transform 1 0 267536 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_2892
timestamp 1586364061
transform 1 0 267168 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_2904
timestamp 1586364061
transform 1 0 268272 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_113
timestamp 1586364061
transform 1 0 269192 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_2908
timestamp 1586364061
transform 1 0 268640 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_0_2915
timestamp 1586364061
transform 1 0 269284 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_2916
timestamp 1586364061
transform 1 0 269376 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_214
timestamp 1586364061
transform 1 0 270480 0 1 2720
box -38 -48 130 592
use scs8hd_decap_12  FILLER_0_2927
timestamp 1586364061
transform 1 0 270388 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_0_2939
timestamp 1586364061
transform 1 0 271492 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_1_2929
timestamp 1586364061
transform 1 0 270572 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_2941
timestamp 1586364061
transform 1 0 271676 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_114
timestamp 1586364061
transform 1 0 272044 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_12  FILLER_0_2946
timestamp 1586364061
transform 1 0 272136 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_2958
timestamp 1586364061
transform 1 0 273240 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_2953
timestamp 1586364061
transform 1 0 272780 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_115
timestamp 1586364061
transform 1 0 274896 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_2970
timestamp 1586364061
transform 1 0 274344 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_0_2977
timestamp 1586364061
transform 1 0 274988 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_2965
timestamp 1586364061
transform 1 0 273884 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_2977
timestamp 1586364061
transform 1 0 274988 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_215
timestamp 1586364061
transform 1 0 276092 0 1 2720
box -38 -48 130 592
use scs8hd_decap_12  FILLER_0_2989
timestamp 1586364061
transform 1 0 276092 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_2990
timestamp 1586364061
transform 1 0 276184 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_116
timestamp 1586364061
transform 1 0 277748 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_3001
timestamp 1586364061
transform 1 0 277196 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_0_3008
timestamp 1586364061
transform 1 0 277840 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_3002
timestamp 1586364061
transform 1 0 277288 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_3014
timestamp 1586364061
transform 1 0 278392 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_3020
timestamp 1586364061
transform 1 0 278944 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_0_3032
timestamp 1586364061
transform 1 0 280048 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_1_3026
timestamp 1586364061
transform 1 0 279496 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_117
timestamp 1586364061
transform 1 0 280600 0 -1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_216
timestamp 1586364061
transform 1 0 281704 0 1 2720
box -38 -48 130 592
use scs8hd_decap_12  FILLER_0_3039
timestamp 1586364061
transform 1 0 280692 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_3038
timestamp 1586364061
transform 1 0 280600 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_3051
timestamp 1586364061
transform 1 0 281796 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_0_3063
timestamp 1586364061
transform 1 0 282900 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_1_3051
timestamp 1586364061
transform 1 0 281796 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_3063
timestamp 1586364061
transform 1 0 282900 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_118
timestamp 1586364061
transform 1 0 283452 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_12  FILLER_0_3070
timestamp 1586364061
transform 1 0 283544 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_3082
timestamp 1586364061
transform 1 0 284648 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_3075
timestamp 1586364061
transform 1 0 284004 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_119
timestamp 1586364061
transform 1 0 286304 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_3094
timestamp 1586364061
transform 1 0 285752 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_0_3101
timestamp 1586364061
transform 1 0 286396 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_3087
timestamp 1586364061
transform 1 0 285108 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_3099
timestamp 1586364061
transform 1 0 286212 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_217
timestamp 1586364061
transform 1 0 287316 0 1 2720
box -38 -48 130 592
use scs8hd_decap_12  FILLER_0_3113
timestamp 1586364061
transform 1 0 287500 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_3112
timestamp 1586364061
transform 1 0 287408 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_120
timestamp 1586364061
transform 1 0 289156 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_3125
timestamp 1586364061
transform 1 0 288604 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_0_3132
timestamp 1586364061
transform 1 0 289248 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_3124
timestamp 1586364061
transform 1 0 288512 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_3136
timestamp 1586364061
transform 1 0 289616 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_3144
timestamp 1586364061
transform 1 0 290352 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_0_3156
timestamp 1586364061
transform 1 0 291456 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_1_3148
timestamp 1586364061
transform 1 0 290720 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_121
timestamp 1586364061
transform 1 0 292008 0 -1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_218
timestamp 1586364061
transform 1 0 292928 0 1 2720
box -38 -48 130 592
use scs8hd_decap_12  FILLER_0_3163
timestamp 1586364061
transform 1 0 292100 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_3160
timestamp 1586364061
transform 1 0 291824 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_3173
timestamp 1586364061
transform 1 0 293020 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_3175
timestamp 1586364061
transform 1 0 293204 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_0_3187
timestamp 1586364061
transform 1 0 294308 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_1_3185
timestamp 1586364061
transform 1 0 294124 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_122
timestamp 1586364061
transform 1 0 294860 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_12  FILLER_0_3194
timestamp 1586364061
transform 1 0 294952 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_3206
timestamp 1586364061
transform 1 0 296056 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_3197
timestamp 1586364061
transform 1 0 295228 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_3209
timestamp 1586364061
transform 1 0 296332 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_123
timestamp 1586364061
transform 1 0 297712 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_3218
timestamp 1586364061
transform 1 0 297160 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_0_3225
timestamp 1586364061
transform 1 0 297804 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_3221
timestamp 1586364061
transform 1 0 297436 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_219
timestamp 1586364061
transform 1 0 298540 0 1 2720
box -38 -48 130 592
use scs8hd_decap_12  FILLER_0_3237
timestamp 1586364061
transform 1 0 298908 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_3234
timestamp 1586364061
transform 1 0 298632 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_3246
timestamp 1586364061
transform 1 0 299736 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_124
timestamp 1586364061
transform 1 0 300564 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_3249
timestamp 1586364061
transform 1 0 300012 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_0_3256
timestamp 1586364061
transform 1 0 300656 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_3258
timestamp 1586364061
transform 1 0 300840 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_3268
timestamp 1586364061
transform 1 0 301760 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_0_3280
timestamp 1586364061
transform 1 0 302864 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_1_3270
timestamp 1586364061
transform 1 0 301944 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_125
timestamp 1586364061
transform 1 0 303416 0 -1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_220
timestamp 1586364061
transform 1 0 304152 0 1 2720
box -38 -48 130 592
use scs8hd_decap_12  FILLER_0_3287
timestamp 1586364061
transform 1 0 303508 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_3299
timestamp 1586364061
transform 1 0 304612 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_3282
timestamp 1586364061
transform 1 0 303048 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_3295
timestamp 1586364061
transform 1 0 304244 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_126
timestamp 1586364061
transform 1 0 306268 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_3311
timestamp 1586364061
transform 1 0 305716 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_1_3307
timestamp 1586364061
transform 1 0 305348 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_3318
timestamp 1586364061
transform 1 0 306360 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_3330
timestamp 1586364061
transform 1 0 307464 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_3319
timestamp 1586364061
transform 1 0 306452 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_3331
timestamp 1586364061
transform 1 0 307556 0 1 2720
box -38 -48 1142 592
use scs8hd_ebufn_1  logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer
timestamp 1586364061
transform 1 0 309212 0 -1 2720
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_127
timestamp 1586364061
transform 1 0 309120 0 -1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer_A
timestamp 1586364061
transform 1 0 308936 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer_TEB
timestamp 1586364061
transform 1 0 308568 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_3344
timestamp 1586364061
transform 1 0 308752 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_12  FILLER_1_3343
timestamp 1586364061
transform 1 0 308660 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_221
timestamp 1586364061
transform 1 0 309764 0 1 2720
box -38 -48 130 592
use scs8hd_decap_12  FILLER_0_3357
timestamp 1586364061
transform 1 0 309948 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_0_3369
timestamp 1586364061
transform 1 0 311052 0 -1 2720
box -38 -48 774 592
use scs8hd_decap_12  FILLER_1_3356
timestamp 1586364061
transform 1 0 309856 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_3368
timestamp 1586364061
transform 1 0 310960 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_128
timestamp 1586364061
transform 1 0 311972 0 -1 2720
box -38 -48 130 592
use scs8hd_fill_2  FILLER_0_3377
timestamp 1586364061
transform 1 0 311788 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_12  FILLER_0_3380
timestamp 1586364061
transform 1 0 312064 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_3380
timestamp 1586364061
transform 1 0 312064 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_3392
timestamp 1586364061
transform 1 0 313168 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_0_3404
timestamp 1586364061
transform 1 0 314272 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_1_3392
timestamp 1586364061
transform 1 0 313168 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_3404
timestamp 1586364061
transform 1 0 314272 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_129
timestamp 1586364061
transform 1 0 314824 0 -1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_222
timestamp 1586364061
transform 1 0 315376 0 1 2720
box -38 -48 130 592
use scs8hd_decap_12  FILLER_0_3411
timestamp 1586364061
transform 1 0 314916 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_3423
timestamp 1586364061
transform 1 0 316020 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_3417
timestamp 1586364061
transform 1 0 315468 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_130
timestamp 1586364061
transform 1 0 317676 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_3435
timestamp 1586364061
transform 1 0 317124 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_0_3442
timestamp 1586364061
transform 1 0 317768 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_3429
timestamp 1586364061
transform 1 0 316572 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_3441
timestamp 1586364061
transform 1 0 317676 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_3454
timestamp 1586364061
transform 1 0 318872 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_3453
timestamp 1586364061
transform 1 0 318780 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_131
timestamp 1586364061
transform 1 0 320528 0 -1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_223
timestamp 1586364061
transform 1 0 320988 0 1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_3466
timestamp 1586364061
transform 1 0 319976 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_0_3473
timestamp 1586364061
transform 1 0 320620 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_3465
timestamp 1586364061
transform 1 0 319884 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_3478
timestamp 1586364061
transform 1 0 321080 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_3485
timestamp 1586364061
transform 1 0 321724 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_3490
timestamp 1586364061
transform 1 0 322184 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_132
timestamp 1586364061
transform 1 0 323380 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_3497
timestamp 1586364061
transform 1 0 322828 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_0_3504
timestamp 1586364061
transform 1 0 323472 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_3502
timestamp 1586364061
transform 1 0 323288 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_3516
timestamp 1586364061
transform 1 0 324576 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_0_3528
timestamp 1586364061
transform 1 0 325680 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_1_3514
timestamp 1586364061
transform 1 0 324392 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_3526
timestamp 1586364061
transform 1 0 325496 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_133
timestamp 1586364061
transform 1 0 326232 0 -1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_224
timestamp 1586364061
transform 1 0 326600 0 1 2720
box -38 -48 130 592
use scs8hd_decap_12  FILLER_0_3535
timestamp 1586364061
transform 1 0 326324 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_3547
timestamp 1586364061
transform 1 0 327428 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_3539
timestamp 1586364061
transform 1 0 326692 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_134
timestamp 1586364061
transform 1 0 329084 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_3559
timestamp 1586364061
transform 1 0 328532 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_0_3566
timestamp 1586364061
transform 1 0 329176 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_3551
timestamp 1586364061
transform 1 0 327796 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_3563
timestamp 1586364061
transform 1 0 328900 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_3578
timestamp 1586364061
transform 1 0 330280 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_3575
timestamp 1586364061
transform 1 0 330004 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_135
timestamp 1586364061
transform 1 0 331936 0 -1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_225
timestamp 1586364061
transform 1 0 332212 0 1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_3590
timestamp 1586364061
transform 1 0 331384 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_0_3597
timestamp 1586364061
transform 1 0 332028 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_3587
timestamp 1586364061
transform 1 0 331108 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_3600
timestamp 1586364061
transform 1 0 332304 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_3609
timestamp 1586364061
transform 1 0 333132 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_3612
timestamp 1586364061
transform 1 0 333408 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_136
timestamp 1586364061
transform 1 0 334788 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_3621
timestamp 1586364061
transform 1 0 334236 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_0_3628
timestamp 1586364061
transform 1 0 334880 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_3624
timestamp 1586364061
transform 1 0 334512 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_3636
timestamp 1586364061
transform 1 0 335616 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_3640
timestamp 1586364061
transform 1 0 335984 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_0_3652
timestamp 1586364061
transform 1 0 337088 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_1_3648
timestamp 1586364061
transform 1 0 336720 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_137
timestamp 1586364061
transform 1 0 337640 0 -1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_226
timestamp 1586364061
transform 1 0 337824 0 1 2720
box -38 -48 130 592
use scs8hd_decap_12  FILLER_0_3659
timestamp 1586364061
transform 1 0 337732 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_3671
timestamp 1586364061
transform 1 0 338836 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_3661
timestamp 1586364061
transform 1 0 337916 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_3673
timestamp 1586364061
transform 1 0 339020 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_138
timestamp 1586364061
transform 1 0 340492 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_3683
timestamp 1586364061
transform 1 0 339940 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_0_3690
timestamp 1586364061
transform 1 0 340584 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_3685
timestamp 1586364061
transform 1 0 340124 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_3702
timestamp 1586364061
transform 1 0 341688 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_3697
timestamp 1586364061
transform 1 0 341228 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_3709
timestamp 1586364061
transform 1 0 342332 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_139
timestamp 1586364061
transform 1 0 343344 0 -1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_227
timestamp 1586364061
transform 1 0 343436 0 1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_3714
timestamp 1586364061
transform 1 0 342792 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_0_3721
timestamp 1586364061
transform 1 0 343436 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_3722
timestamp 1586364061
transform 1 0 343528 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_3733
timestamp 1586364061
transform 1 0 344540 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_0_3745
timestamp 1586364061
transform 1 0 345644 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_1_3734
timestamp 1586364061
transform 1 0 344632 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_140
timestamp 1586364061
transform 1 0 346196 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_12  FILLER_0_3752
timestamp 1586364061
transform 1 0 346288 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_3746
timestamp 1586364061
transform 1 0 345736 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_3758
timestamp 1586364061
transform 1 0 346840 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_3764
timestamp 1586364061
transform 1 0 347392 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_0_3776
timestamp 1586364061
transform 1 0 348496 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_1_3770
timestamp 1586364061
transform 1 0 347944 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_141
timestamp 1586364061
transform 1 0 349048 0 -1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_228
timestamp 1586364061
transform 1 0 349048 0 1 2720
box -38 -48 130 592
use scs8hd_decap_12  FILLER_0_3783
timestamp 1586364061
transform 1 0 349140 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_0_3795
timestamp 1586364061
transform 1 0 350244 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_1_3783
timestamp 1586364061
transform 1 0 349140 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_3795
timestamp 1586364061
transform 1 0 350244 0 1 2720
box -38 -48 1142 592
use scs8hd_buf_2  _22_
timestamp 1586364061
transform 1 0 350796 0 -1 2720
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_142
timestamp 1586364061
transform 1 0 351900 0 -1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__22__A
timestamp 1586364061
transform 1 0 351348 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_3805
timestamp 1586364061
transform 1 0 351164 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_0_3809
timestamp 1586364061
transform 1 0 351532 0 -1 2720
box -38 -48 406 592
use scs8hd_decap_12  FILLER_0_3814
timestamp 1586364061
transform 1 0 351992 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_3807
timestamp 1586364061
transform 1 0 351348 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_3826
timestamp 1586364061
transform 1 0 353096 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_3819
timestamp 1586364061
transform 1 0 352452 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_3831
timestamp 1586364061
transform 1 0 353556 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_143
timestamp 1586364061
transform 1 0 354752 0 -1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_229
timestamp 1586364061
transform 1 0 354660 0 1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_3838
timestamp 1586364061
transform 1 0 354200 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_0_3845
timestamp 1586364061
transform 1 0 354844 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_3844
timestamp 1586364061
transform 1 0 354752 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_3857
timestamp 1586364061
transform 1 0 355948 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_0_3869
timestamp 1586364061
transform 1 0 357052 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_1_3856
timestamp 1586364061
transform 1 0 355856 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_3868
timestamp 1586364061
transform 1 0 356960 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_144
timestamp 1586364061
transform 1 0 357604 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_12  FILLER_0_3876
timestamp 1586364061
transform 1 0 357696 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_3888
timestamp 1586364061
transform 1 0 358800 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_3880
timestamp 1586364061
transform 1 0 358064 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_145
timestamp 1586364061
transform 1 0 360456 0 -1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_230
timestamp 1586364061
transform 1 0 360272 0 1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_3900
timestamp 1586364061
transform 1 0 359904 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_1_3892
timestamp 1586364061
transform 1 0 359168 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_3905
timestamp 1586364061
transform 1 0 360364 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_3907
timestamp 1586364061
transform 1 0 360548 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_3919
timestamp 1586364061
transform 1 0 361652 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_3917
timestamp 1586364061
transform 1 0 361468 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_146
timestamp 1586364061
transform 1 0 363308 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_3931
timestamp 1586364061
transform 1 0 362756 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_0_3938
timestamp 1586364061
transform 1 0 363400 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_3929
timestamp 1586364061
transform 1 0 362572 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_3941
timestamp 1586364061
transform 1 0 363676 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_3950
timestamp 1586364061
transform 1 0 364504 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_3953
timestamp 1586364061
transform 1 0 364780 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_147
timestamp 1586364061
transform 1 0 366160 0 -1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_231
timestamp 1586364061
transform 1 0 365884 0 1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_3962
timestamp 1586364061
transform 1 0 365608 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_0_3969
timestamp 1586364061
transform 1 0 366252 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_3966
timestamp 1586364061
transform 1 0 365976 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_3981
timestamp 1586364061
transform 1 0 367356 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_0_3993
timestamp 1586364061
transform 1 0 368460 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_1_3978
timestamp 1586364061
transform 1 0 367080 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_3990
timestamp 1586364061
transform 1 0 368184 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_148
timestamp 1586364061
transform 1 0 369012 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_12  FILLER_0_4000
timestamp 1586364061
transform 1 0 369104 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_4012
timestamp 1586364061
transform 1 0 370208 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_4002
timestamp 1586364061
transform 1 0 369288 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_149
timestamp 1586364061
transform 1 0 371864 0 -1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_232
timestamp 1586364061
transform 1 0 371496 0 1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_4024
timestamp 1586364061
transform 1 0 371312 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_0_4031
timestamp 1586364061
transform 1 0 371956 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_4014
timestamp 1586364061
transform 1 0 370392 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_4027
timestamp 1586364061
transform 1 0 371588 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_4043
timestamp 1586364061
transform 1 0 373060 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_4039
timestamp 1586364061
transform 1 0 372692 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_150
timestamp 1586364061
transform 1 0 374716 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_4055
timestamp 1586364061
transform 1 0 374164 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_0_4062
timestamp 1586364061
transform 1 0 374808 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_4051
timestamp 1586364061
transform 1 0 373796 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_4063
timestamp 1586364061
transform 1 0 374900 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_4074
timestamp 1586364061
transform 1 0 375912 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_4075
timestamp 1586364061
transform 1 0 376004 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_151
timestamp 1586364061
transform 1 0 377568 0 -1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_233
timestamp 1586364061
transform 1 0 377108 0 1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_4086
timestamp 1586364061
transform 1 0 377016 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_0_4093
timestamp 1586364061
transform 1 0 377660 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_4088
timestamp 1586364061
transform 1 0 377200 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_4100
timestamp 1586364061
transform 1 0 378304 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_4105
timestamp 1586364061
transform 1 0 378764 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_0_4117
timestamp 1586364061
transform 1 0 379868 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_1_4112
timestamp 1586364061
transform 1 0 379408 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_152
timestamp 1586364061
transform 1 0 380420 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_12  FILLER_0_4124
timestamp 1586364061
transform 1 0 380512 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_4136
timestamp 1586364061
transform 1 0 381616 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_4124
timestamp 1586364061
transform 1 0 380512 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_4136
timestamp 1586364061
transform 1 0 381616 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_153
timestamp 1586364061
transform 1 0 383272 0 -1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_234
timestamp 1586364061
transform 1 0 382720 0 1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_4148
timestamp 1586364061
transform 1 0 382720 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_0_4155
timestamp 1586364061
transform 1 0 383364 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_4149
timestamp 1586364061
transform 1 0 382812 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_4167
timestamp 1586364061
transform 1 0 384468 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_4161
timestamp 1586364061
transform 1 0 383916 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_4173
timestamp 1586364061
transform 1 0 385020 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_154
timestamp 1586364061
transform 1 0 386124 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_4179
timestamp 1586364061
transform 1 0 385572 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_0_4186
timestamp 1586364061
transform 1 0 386216 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_4185
timestamp 1586364061
transform 1 0 386124 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_235
timestamp 1586364061
transform 1 0 388332 0 1 2720
box -38 -48 130 592
use scs8hd_decap_12  FILLER_0_4198
timestamp 1586364061
transform 1 0 387320 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_4197
timestamp 1586364061
transform 1 0 387228 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_155
timestamp 1586364061
transform 1 0 388976 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_4210
timestamp 1586364061
transform 1 0 388424 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_0_4217
timestamp 1586364061
transform 1 0 389068 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_4210
timestamp 1586364061
transform 1 0 388424 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_4222
timestamp 1586364061
transform 1 0 389528 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_4229
timestamp 1586364061
transform 1 0 390172 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_0_4241
timestamp 1586364061
transform 1 0 391276 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_1_4234
timestamp 1586364061
transform 1 0 390632 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_156
timestamp 1586364061
transform 1 0 391828 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_12  FILLER_0_4248
timestamp 1586364061
transform 1 0 391920 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_4260
timestamp 1586364061
transform 1 0 393024 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_4246
timestamp 1586364061
transform 1 0 391736 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_4258
timestamp 1586364061
transform 1 0 392840 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_157
timestamp 1586364061
transform 1 0 394680 0 -1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_236
timestamp 1586364061
transform 1 0 393944 0 1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_4272
timestamp 1586364061
transform 1 0 394128 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_0_4279
timestamp 1586364061
transform 1 0 394772 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_4271
timestamp 1586364061
transform 1 0 394036 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_4291
timestamp 1586364061
transform 1 0 395876 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_4283
timestamp 1586364061
transform 1 0 395140 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_4295
timestamp 1586364061
transform 1 0 396244 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_158
timestamp 1586364061
transform 1 0 397532 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_4303
timestamp 1586364061
transform 1 0 396980 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_0_4310
timestamp 1586364061
transform 1 0 397624 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_4307
timestamp 1586364061
transform 1 0 397348 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_237
timestamp 1586364061
transform 1 0 399556 0 1 2720
box -38 -48 130 592
use scs8hd_decap_12  FILLER_0_4322
timestamp 1586364061
transform 1 0 398728 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_0_4334
timestamp 1586364061
transform 1 0 399832 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_1_4319
timestamp 1586364061
transform 1 0 398452 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_4332
timestamp 1586364061
transform 1 0 399648 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_159
timestamp 1586364061
transform 1 0 400384 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_12  FILLER_0_4341
timestamp 1586364061
transform 1 0 400476 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_4344
timestamp 1586364061
transform 1 0 400752 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_4353
timestamp 1586364061
transform 1 0 401580 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_0_4365
timestamp 1586364061
transform 1 0 402684 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_1_4356
timestamp 1586364061
transform 1 0 401856 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_4368
timestamp 1586364061
transform 1 0 402960 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_160
timestamp 1586364061
transform 1 0 403236 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_12  FILLER_0_4372
timestamp 1586364061
transform 1 0 403328 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_4384
timestamp 1586364061
transform 1 0 404432 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_4380
timestamp 1586364061
transform 1 0 404064 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_161
timestamp 1586364061
transform 1 0 406088 0 -1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_238
timestamp 1586364061
transform 1 0 405168 0 1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_4396
timestamp 1586364061
transform 1 0 405536 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_0_4403
timestamp 1586364061
transform 1 0 406180 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_4393
timestamp 1586364061
transform 1 0 405260 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_4405
timestamp 1586364061
transform 1 0 406364 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_4415
timestamp 1586364061
transform 1 0 407284 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_4417
timestamp 1586364061
transform 1 0 407468 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_162
timestamp 1586364061
transform 1 0 408940 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_4427
timestamp 1586364061
transform 1 0 408388 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_0_4434
timestamp 1586364061
transform 1 0 409032 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_4429
timestamp 1586364061
transform 1 0 408572 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_4441
timestamp 1586364061
transform 1 0 409676 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_239
timestamp 1586364061
transform 1 0 410780 0 1 2720
box -38 -48 130 592
use scs8hd_decap_12  FILLER_0_4446
timestamp 1586364061
transform 1 0 410136 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_0_4458
timestamp 1586364061
transform 1 0 411240 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_1_4454
timestamp 1586364061
transform 1 0 410872 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_163
timestamp 1586364061
transform 1 0 411792 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_12  FILLER_0_4465
timestamp 1586364061
transform 1 0 411884 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_4477
timestamp 1586364061
transform 1 0 412988 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_4466
timestamp 1586364061
transform 1 0 411976 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_0_4489
timestamp 1586364061
transform 1 0 414092 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_1_4478
timestamp 1586364061
transform 1 0 413080 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_4490
timestamp 1586364061
transform 1 0 414184 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_164
timestamp 1586364061
transform 1 0 414644 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_12  FILLER_0_4496
timestamp 1586364061
transform 1 0 414736 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_4508
timestamp 1586364061
transform 1 0 415840 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_4502
timestamp 1586364061
transform 1 0 415288 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_165
timestamp 1586364061
transform 1 0 417496 0 -1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_240
timestamp 1586364061
transform 1 0 416392 0 1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_4520
timestamp 1586364061
transform 1 0 416944 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_0_4527
timestamp 1586364061
transform 1 0 417588 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_4515
timestamp 1586364061
transform 1 0 416484 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_4527
timestamp 1586364061
transform 1 0 417588 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_4539
timestamp 1586364061
transform 1 0 418692 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_4539
timestamp 1586364061
transform 1 0 418692 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_166
timestamp 1586364061
transform 1 0 420348 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_4551
timestamp 1586364061
transform 1 0 419796 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_0_4558
timestamp 1586364061
transform 1 0 420440 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_4551
timestamp 1586364061
transform 1 0 419796 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_4563
timestamp 1586364061
transform 1 0 420900 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_3  PHY_1
timestamp 1586364061
transform -1 0 422832 0 -1 2720
box -38 -48 314 592
use scs8hd_decap_3  PHY_3
timestamp 1586364061
transform -1 0 422832 0 1 2720
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_241
timestamp 1586364061
transform 1 0 422004 0 1 2720
box -38 -48 130 592
use scs8hd_decap_8  FILLER_0_4570
timestamp 1586364061
transform 1 0 421544 0 -1 2720
box -38 -48 774 592
use scs8hd_decap_3  FILLER_0_4578
timestamp 1586364061
transform 1 0 422280 0 -1 2720
box -38 -48 314 592
use scs8hd_decap_4  FILLER_1_4576
timestamp 1586364061
transform 1 0 422096 0 1 2720
box -38 -48 406 592
use scs8hd_fill_1  FILLER_1_4580
timestamp 1586364061
transform 1 0 422464 0 1 2720
box -38 -48 130 592
use scs8hd_decap_3  PHY_4
timestamp 1586364061
transform 1 0 1104 0 -1 3808
box -38 -48 314 592
use scs8hd_decap_12  FILLER_2_3
timestamp 1586364061
transform 1 0 1380 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_15
timestamp 1586364061
transform 1 0 2484 0 -1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_242
timestamp 1586364061
transform 1 0 3956 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_4  FILLER_2_27
timestamp 1586364061
transform 1 0 3588 0 -1 3808
box -38 -48 406 592
use scs8hd_decap_12  FILLER_2_32
timestamp 1586364061
transform 1 0 4048 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_44
timestamp 1586364061
transform 1 0 5152 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_56
timestamp 1586364061
transform 1 0 6256 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_68
timestamp 1586364061
transform 1 0 7360 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_80
timestamp 1586364061
transform 1 0 8464 0 -1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_243
timestamp 1586364061
transform 1 0 9568 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_2_93
timestamp 1586364061
transform 1 0 9660 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_105
timestamp 1586364061
transform 1 0 10764 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_117
timestamp 1586364061
transform 1 0 11868 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_129
timestamp 1586364061
transform 1 0 12972 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_141
timestamp 1586364061
transform 1 0 14076 0 -1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_244
timestamp 1586364061
transform 1 0 15180 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_2_154
timestamp 1586364061
transform 1 0 15272 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_166
timestamp 1586364061
transform 1 0 16376 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_178
timestamp 1586364061
transform 1 0 17480 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_190
timestamp 1586364061
transform 1 0 18584 0 -1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_245
timestamp 1586364061
transform 1 0 20792 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_2_202
timestamp 1586364061
transform 1 0 19688 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_215
timestamp 1586364061
transform 1 0 20884 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_227
timestamp 1586364061
transform 1 0 21988 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_239
timestamp 1586364061
transform 1 0 23092 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_251
timestamp 1586364061
transform 1 0 24196 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_263
timestamp 1586364061
transform 1 0 25300 0 -1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_246
timestamp 1586364061
transform 1 0 26404 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_2_276
timestamp 1586364061
transform 1 0 26496 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_288
timestamp 1586364061
transform 1 0 27600 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_300
timestamp 1586364061
transform 1 0 28704 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_312
timestamp 1586364061
transform 1 0 29808 0 -1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_247
timestamp 1586364061
transform 1 0 32016 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_2_324
timestamp 1586364061
transform 1 0 30912 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_337
timestamp 1586364061
transform 1 0 32108 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_349
timestamp 1586364061
transform 1 0 33212 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_361
timestamp 1586364061
transform 1 0 34316 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_373
timestamp 1586364061
transform 1 0 35420 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_385
timestamp 1586364061
transform 1 0 36524 0 -1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_248
timestamp 1586364061
transform 1 0 37628 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_2_398
timestamp 1586364061
transform 1 0 37720 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_410
timestamp 1586364061
transform 1 0 38824 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_422
timestamp 1586364061
transform 1 0 39928 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_434
timestamp 1586364061
transform 1 0 41032 0 -1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_249
timestamp 1586364061
transform 1 0 43240 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_2_446
timestamp 1586364061
transform 1 0 42136 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_459
timestamp 1586364061
transform 1 0 43332 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_471
timestamp 1586364061
transform 1 0 44436 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_483
timestamp 1586364061
transform 1 0 45540 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_495
timestamp 1586364061
transform 1 0 46644 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_507
timestamp 1586364061
transform 1 0 47748 0 -1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_250
timestamp 1586364061
transform 1 0 48852 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_2_520
timestamp 1586364061
transform 1 0 48944 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_532
timestamp 1586364061
transform 1 0 50048 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_544
timestamp 1586364061
transform 1 0 51152 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_556
timestamp 1586364061
transform 1 0 52256 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_568
timestamp 1586364061
transform 1 0 53360 0 -1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_251
timestamp 1586364061
transform 1 0 54464 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_2_581
timestamp 1586364061
transform 1 0 54556 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_593
timestamp 1586364061
transform 1 0 55660 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_605
timestamp 1586364061
transform 1 0 56764 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_617
timestamp 1586364061
transform 1 0 57868 0 -1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_252
timestamp 1586364061
transform 1 0 60076 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_2_629
timestamp 1586364061
transform 1 0 58972 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_642
timestamp 1586364061
transform 1 0 60168 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_654
timestamp 1586364061
transform 1 0 61272 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_666
timestamp 1586364061
transform 1 0 62376 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_678
timestamp 1586364061
transform 1 0 63480 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_690
timestamp 1586364061
transform 1 0 64584 0 -1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_253
timestamp 1586364061
transform 1 0 65688 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_2_703
timestamp 1586364061
transform 1 0 65780 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_715
timestamp 1586364061
transform 1 0 66884 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_727
timestamp 1586364061
transform 1 0 67988 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_739
timestamp 1586364061
transform 1 0 69092 0 -1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_254
timestamp 1586364061
transform 1 0 71300 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_2_751
timestamp 1586364061
transform 1 0 70196 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_764
timestamp 1586364061
transform 1 0 71392 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_776
timestamp 1586364061
transform 1 0 72496 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_788
timestamp 1586364061
transform 1 0 73600 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_800
timestamp 1586364061
transform 1 0 74704 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_812
timestamp 1586364061
transform 1 0 75808 0 -1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_255
timestamp 1586364061
transform 1 0 76912 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_2_825
timestamp 1586364061
transform 1 0 77004 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_837
timestamp 1586364061
transform 1 0 78108 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_849
timestamp 1586364061
transform 1 0 79212 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_861
timestamp 1586364061
transform 1 0 80316 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_873
timestamp 1586364061
transform 1 0 81420 0 -1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_256
timestamp 1586364061
transform 1 0 82524 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_2_886
timestamp 1586364061
transform 1 0 82616 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_898
timestamp 1586364061
transform 1 0 83720 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_910
timestamp 1586364061
transform 1 0 84824 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_922
timestamp 1586364061
transform 1 0 85928 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_934
timestamp 1586364061
transform 1 0 87032 0 -1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_257
timestamp 1586364061
transform 1 0 88136 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_2_947
timestamp 1586364061
transform 1 0 88228 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_959
timestamp 1586364061
transform 1 0 89332 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_971
timestamp 1586364061
transform 1 0 90436 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_983
timestamp 1586364061
transform 1 0 91540 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_995
timestamp 1586364061
transform 1 0 92644 0 -1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_258
timestamp 1586364061
transform 1 0 93748 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_2_1008
timestamp 1586364061
transform 1 0 93840 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_1020
timestamp 1586364061
transform 1 0 94944 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_1032
timestamp 1586364061
transform 1 0 96048 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_1044
timestamp 1586364061
transform 1 0 97152 0 -1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_259
timestamp 1586364061
transform 1 0 99360 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_2_1056
timestamp 1586364061
transform 1 0 98256 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_1069
timestamp 1586364061
transform 1 0 99452 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_1081
timestamp 1586364061
transform 1 0 100556 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_1093
timestamp 1586364061
transform 1 0 101660 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_1105
timestamp 1586364061
transform 1 0 102764 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_1117
timestamp 1586364061
transform 1 0 103868 0 -1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_260
timestamp 1586364061
transform 1 0 104972 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_2_1130
timestamp 1586364061
transform 1 0 105064 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_1142
timestamp 1586364061
transform 1 0 106168 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_1154
timestamp 1586364061
transform 1 0 107272 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_1166
timestamp 1586364061
transform 1 0 108376 0 -1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_261
timestamp 1586364061
transform 1 0 110584 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_2_1178
timestamp 1586364061
transform 1 0 109480 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_1191
timestamp 1586364061
transform 1 0 110676 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_1203
timestamp 1586364061
transform 1 0 111780 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_1215
timestamp 1586364061
transform 1 0 112884 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_1227
timestamp 1586364061
transform 1 0 113988 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_1239
timestamp 1586364061
transform 1 0 115092 0 -1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_262
timestamp 1586364061
transform 1 0 116196 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_2_1252
timestamp 1586364061
transform 1 0 116288 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_1264
timestamp 1586364061
transform 1 0 117392 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_1276
timestamp 1586364061
transform 1 0 118496 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_1288
timestamp 1586364061
transform 1 0 119600 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_1300
timestamp 1586364061
transform 1 0 120704 0 -1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_263
timestamp 1586364061
transform 1 0 121808 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_2_1313
timestamp 1586364061
transform 1 0 121900 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_1325
timestamp 1586364061
transform 1 0 123004 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_1337
timestamp 1586364061
transform 1 0 124108 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_1349
timestamp 1586364061
transform 1 0 125212 0 -1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_264
timestamp 1586364061
transform 1 0 127420 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_2_1361
timestamp 1586364061
transform 1 0 126316 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_1374
timestamp 1586364061
transform 1 0 127512 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_1386
timestamp 1586364061
transform 1 0 128616 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_1398
timestamp 1586364061
transform 1 0 129720 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_1410
timestamp 1586364061
transform 1 0 130824 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_1422
timestamp 1586364061
transform 1 0 131928 0 -1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_265
timestamp 1586364061
transform 1 0 133032 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_2_1435
timestamp 1586364061
transform 1 0 133124 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_1447
timestamp 1586364061
transform 1 0 134228 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_1459
timestamp 1586364061
transform 1 0 135332 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_1471
timestamp 1586364061
transform 1 0 136436 0 -1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_266
timestamp 1586364061
transform 1 0 138644 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_2_1483
timestamp 1586364061
transform 1 0 137540 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_1496
timestamp 1586364061
transform 1 0 138736 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_1508
timestamp 1586364061
transform 1 0 139840 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_1520
timestamp 1586364061
transform 1 0 140944 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_1532
timestamp 1586364061
transform 1 0 142048 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_1544
timestamp 1586364061
transform 1 0 143152 0 -1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_267
timestamp 1586364061
transform 1 0 144256 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_2_1557
timestamp 1586364061
transform 1 0 144348 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_1569
timestamp 1586364061
transform 1 0 145452 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_1581
timestamp 1586364061
transform 1 0 146556 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_1593
timestamp 1586364061
transform 1 0 147660 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_1605
timestamp 1586364061
transform 1 0 148764 0 -1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_268
timestamp 1586364061
transform 1 0 149868 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_2_1618
timestamp 1586364061
transform 1 0 149960 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_1630
timestamp 1586364061
transform 1 0 151064 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_1642
timestamp 1586364061
transform 1 0 152168 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_1654
timestamp 1586364061
transform 1 0 153272 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_1666
timestamp 1586364061
transform 1 0 154376 0 -1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_269
timestamp 1586364061
transform 1 0 155480 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_2_1679
timestamp 1586364061
transform 1 0 155572 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_1691
timestamp 1586364061
transform 1 0 156676 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_1703
timestamp 1586364061
transform 1 0 157780 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_1715
timestamp 1586364061
transform 1 0 158884 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_1727
timestamp 1586364061
transform 1 0 159988 0 -1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_270
timestamp 1586364061
transform 1 0 161092 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_2_1740
timestamp 1586364061
transform 1 0 161184 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_1752
timestamp 1586364061
transform 1 0 162288 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_1764
timestamp 1586364061
transform 1 0 163392 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_1776
timestamp 1586364061
transform 1 0 164496 0 -1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_271
timestamp 1586364061
transform 1 0 166704 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_2_1788
timestamp 1586364061
transform 1 0 165600 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_1801
timestamp 1586364061
transform 1 0 166796 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_1813
timestamp 1586364061
transform 1 0 167900 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_1825
timestamp 1586364061
transform 1 0 169004 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_1837
timestamp 1586364061
transform 1 0 170108 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_1849
timestamp 1586364061
transform 1 0 171212 0 -1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_272
timestamp 1586364061
transform 1 0 172316 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_2_1862
timestamp 1586364061
transform 1 0 172408 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_1874
timestamp 1586364061
transform 1 0 173512 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_1886
timestamp 1586364061
transform 1 0 174616 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_1898
timestamp 1586364061
transform 1 0 175720 0 -1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_273
timestamp 1586364061
transform 1 0 177928 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_2_1910
timestamp 1586364061
transform 1 0 176824 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_1923
timestamp 1586364061
transform 1 0 178020 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_1935
timestamp 1586364061
transform 1 0 179124 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_1947
timestamp 1586364061
transform 1 0 180228 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_1959
timestamp 1586364061
transform 1 0 181332 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_1971
timestamp 1586364061
transform 1 0 182436 0 -1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_274
timestamp 1586364061
transform 1 0 183540 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_2_1984
timestamp 1586364061
transform 1 0 183632 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_1996
timestamp 1586364061
transform 1 0 184736 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_2008
timestamp 1586364061
transform 1 0 185840 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_2020
timestamp 1586364061
transform 1 0 186944 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_2032
timestamp 1586364061
transform 1 0 188048 0 -1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_275
timestamp 1586364061
transform 1 0 189152 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_2_2045
timestamp 1586364061
transform 1 0 189244 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_2057
timestamp 1586364061
transform 1 0 190348 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_2069
timestamp 1586364061
transform 1 0 191452 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_2081
timestamp 1586364061
transform 1 0 192556 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_2093
timestamp 1586364061
transform 1 0 193660 0 -1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_276
timestamp 1586364061
transform 1 0 194764 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_2_2106
timestamp 1586364061
transform 1 0 194856 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_2118
timestamp 1586364061
transform 1 0 195960 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_2130
timestamp 1586364061
transform 1 0 197064 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_2142
timestamp 1586364061
transform 1 0 198168 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_2154
timestamp 1586364061
transform 1 0 199272 0 -1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_277
timestamp 1586364061
transform 1 0 200376 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_2_2167
timestamp 1586364061
transform 1 0 200468 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_2179
timestamp 1586364061
transform 1 0 201572 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_2191
timestamp 1586364061
transform 1 0 202676 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_2203
timestamp 1586364061
transform 1 0 203780 0 -1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_278
timestamp 1586364061
transform 1 0 205988 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_2_2215
timestamp 1586364061
transform 1 0 204884 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_2228
timestamp 1586364061
transform 1 0 206080 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_2240
timestamp 1586364061
transform 1 0 207184 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_2252
timestamp 1586364061
transform 1 0 208288 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_2264
timestamp 1586364061
transform 1 0 209392 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_2276
timestamp 1586364061
transform 1 0 210496 0 -1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_279
timestamp 1586364061
transform 1 0 211600 0 -1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__15__C
timestamp 1586364061
transform 1 0 212428 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_8  FILLER_2_2289
timestamp 1586364061
transform 1 0 211692 0 -1 3808
box -38 -48 774 592
use scs8hd_fill_2  FILLER_2_2299
timestamp 1586364061
transform 1 0 212612 0 -1 3808
box -38 -48 222 592
use scs8hd_nor4_4  _15_
timestamp 1586364061
transform 1 0 213256 0 -1 3808
box -38 -48 1602 592
use scs8hd_diode_2  ANTENNA__07__D
timestamp 1586364061
transform 1 0 212796 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_3  FILLER_2_2303
timestamp 1586364061
transform 1 0 212980 0 -1 3808
box -38 -48 314 592
use scs8hd_and4_4  _05_
timestamp 1586364061
transform 1 0 215556 0 -1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__05__D
timestamp 1586364061
transform 1 0 215372 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__05__A
timestamp 1586364061
transform 1 0 215004 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_2323
timestamp 1586364061
transform 1 0 214820 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_2327
timestamp 1586364061
transform 1 0 215188 0 -1 3808
box -38 -48 222 592
use scs8hd_inv_8  _08_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 217304 0 -1 3808
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_280
timestamp 1586364061
transform 1 0 217212 0 -1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__12__C
timestamp 1586364061
transform 1 0 216568 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__12__A
timestamp 1586364061
transform 1 0 216936 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_2340
timestamp 1586364061
transform 1 0 216384 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_2344
timestamp 1586364061
transform 1 0 216752 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_1  FILLER_2_2348
timestamp 1586364061
transform 1 0 217120 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_2_2359
timestamp 1586364061
transform 1 0 218132 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_2_2371
timestamp 1586364061
transform 1 0 219236 0 -1 3808
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.LATCH_0_.latch
timestamp 1586364061
transform 1 0 219696 0 -1 3808
box -38 -48 1050 592
use scs8hd_fill_1  FILLER_2_2375
timestamp 1586364061
transform 1 0 219604 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_2_2387
timestamp 1586364061
transform 1 0 220708 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_2_2399
timestamp 1586364061
transform 1 0 221812 0 -1 3808
box -38 -48 774 592
use scs8hd_decap_3  FILLER_2_2407
timestamp 1586364061
transform 1 0 222548 0 -1 3808
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_281
timestamp 1586364061
transform 1 0 222824 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_2_2411
timestamp 1586364061
transform 1 0 222916 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_2423
timestamp 1586364061
transform 1 0 224020 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_2435
timestamp 1586364061
transform 1 0 225124 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_2447
timestamp 1586364061
transform 1 0 226228 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_2459
timestamp 1586364061
transform 1 0 227332 0 -1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_282
timestamp 1586364061
transform 1 0 228436 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_2_2472
timestamp 1586364061
transform 1 0 228528 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_2484
timestamp 1586364061
transform 1 0 229632 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_2496
timestamp 1586364061
transform 1 0 230736 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_2508
timestamp 1586364061
transform 1 0 231840 0 -1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_283
timestamp 1586364061
transform 1 0 234048 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_2_2520
timestamp 1586364061
transform 1 0 232944 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_2533
timestamp 1586364061
transform 1 0 234140 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_2545
timestamp 1586364061
transform 1 0 235244 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_2557
timestamp 1586364061
transform 1 0 236348 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_2569
timestamp 1586364061
transform 1 0 237452 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_2581
timestamp 1586364061
transform 1 0 238556 0 -1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_284
timestamp 1586364061
transform 1 0 239660 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_2_2594
timestamp 1586364061
transform 1 0 239752 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_2606
timestamp 1586364061
transform 1 0 240856 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_2618
timestamp 1586364061
transform 1 0 241960 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_2630
timestamp 1586364061
transform 1 0 243064 0 -1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_285
timestamp 1586364061
transform 1 0 245272 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_2_2642
timestamp 1586364061
transform 1 0 244168 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_2655
timestamp 1586364061
transform 1 0 245364 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_2667
timestamp 1586364061
transform 1 0 246468 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_2679
timestamp 1586364061
transform 1 0 247572 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_2691
timestamp 1586364061
transform 1 0 248676 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_2703
timestamp 1586364061
transform 1 0 249780 0 -1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_286
timestamp 1586364061
transform 1 0 250884 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_2_2716
timestamp 1586364061
transform 1 0 250976 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_2728
timestamp 1586364061
transform 1 0 252080 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_2740
timestamp 1586364061
transform 1 0 253184 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_2752
timestamp 1586364061
transform 1 0 254288 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_2764
timestamp 1586364061
transform 1 0 255392 0 -1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_287
timestamp 1586364061
transform 1 0 256496 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_2_2777
timestamp 1586364061
transform 1 0 256588 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_2789
timestamp 1586364061
transform 1 0 257692 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_2801
timestamp 1586364061
transform 1 0 258796 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_2813
timestamp 1586364061
transform 1 0 259900 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_2825
timestamp 1586364061
transform 1 0 261004 0 -1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_288
timestamp 1586364061
transform 1 0 262108 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_2_2838
timestamp 1586364061
transform 1 0 262200 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_2850
timestamp 1586364061
transform 1 0 263304 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_2862
timestamp 1586364061
transform 1 0 264408 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_2874
timestamp 1586364061
transform 1 0 265512 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_2886
timestamp 1586364061
transform 1 0 266616 0 -1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_289
timestamp 1586364061
transform 1 0 267720 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_2_2899
timestamp 1586364061
transform 1 0 267812 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_2911
timestamp 1586364061
transform 1 0 268916 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_2923
timestamp 1586364061
transform 1 0 270020 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_2935
timestamp 1586364061
transform 1 0 271124 0 -1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_290
timestamp 1586364061
transform 1 0 273332 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_2_2947
timestamp 1586364061
transform 1 0 272228 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_2960
timestamp 1586364061
transform 1 0 273424 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_2972
timestamp 1586364061
transform 1 0 274528 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_2984
timestamp 1586364061
transform 1 0 275632 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_2996
timestamp 1586364061
transform 1 0 276736 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_3008
timestamp 1586364061
transform 1 0 277840 0 -1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_291
timestamp 1586364061
transform 1 0 278944 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_2_3021
timestamp 1586364061
transform 1 0 279036 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_3033
timestamp 1586364061
transform 1 0 280140 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_3045
timestamp 1586364061
transform 1 0 281244 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_3057
timestamp 1586364061
transform 1 0 282348 0 -1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_292
timestamp 1586364061
transform 1 0 284556 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_2_3069
timestamp 1586364061
transform 1 0 283452 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_3082
timestamp 1586364061
transform 1 0 284648 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_3094
timestamp 1586364061
transform 1 0 285752 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_3106
timestamp 1586364061
transform 1 0 286856 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_3118
timestamp 1586364061
transform 1 0 287960 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_3130
timestamp 1586364061
transform 1 0 289064 0 -1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_293
timestamp 1586364061
transform 1 0 290168 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_2_3143
timestamp 1586364061
transform 1 0 290260 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_3155
timestamp 1586364061
transform 1 0 291364 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_3167
timestamp 1586364061
transform 1 0 292468 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_3179
timestamp 1586364061
transform 1 0 293572 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_3191
timestamp 1586364061
transform 1 0 294676 0 -1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_294
timestamp 1586364061
transform 1 0 295780 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_2_3204
timestamp 1586364061
transform 1 0 295872 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_3216
timestamp 1586364061
transform 1 0 296976 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_3228
timestamp 1586364061
transform 1 0 298080 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_3240
timestamp 1586364061
transform 1 0 299184 0 -1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_295
timestamp 1586364061
transform 1 0 301392 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_2_3252
timestamp 1586364061
transform 1 0 300288 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_3265
timestamp 1586364061
transform 1 0 301484 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_3277
timestamp 1586364061
transform 1 0 302588 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_3289
timestamp 1586364061
transform 1 0 303692 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_3301
timestamp 1586364061
transform 1 0 304796 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_3313
timestamp 1586364061
transform 1 0 305900 0 -1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_296
timestamp 1586364061
transform 1 0 307004 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_2_3326
timestamp 1586364061
transform 1 0 307096 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_3338
timestamp 1586364061
transform 1 0 308200 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_3350
timestamp 1586364061
transform 1 0 309304 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_3362
timestamp 1586364061
transform 1 0 310408 0 -1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_297
timestamp 1586364061
transform 1 0 312616 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_2_3374
timestamp 1586364061
transform 1 0 311512 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_3387
timestamp 1586364061
transform 1 0 312708 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_3399
timestamp 1586364061
transform 1 0 313812 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_3411
timestamp 1586364061
transform 1 0 314916 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_3423
timestamp 1586364061
transform 1 0 316020 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_3435
timestamp 1586364061
transform 1 0 317124 0 -1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_298
timestamp 1586364061
transform 1 0 318228 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_2_3448
timestamp 1586364061
transform 1 0 318320 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_3460
timestamp 1586364061
transform 1 0 319424 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_3472
timestamp 1586364061
transform 1 0 320528 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_3484
timestamp 1586364061
transform 1 0 321632 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_3496
timestamp 1586364061
transform 1 0 322736 0 -1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_299
timestamp 1586364061
transform 1 0 323840 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_2_3509
timestamp 1586364061
transform 1 0 323932 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_3521
timestamp 1586364061
transform 1 0 325036 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_3533
timestamp 1586364061
transform 1 0 326140 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_3545
timestamp 1586364061
transform 1 0 327244 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_3557
timestamp 1586364061
transform 1 0 328348 0 -1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_300
timestamp 1586364061
transform 1 0 329452 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_2_3570
timestamp 1586364061
transform 1 0 329544 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_3582
timestamp 1586364061
transform 1 0 330648 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_3594
timestamp 1586364061
transform 1 0 331752 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_3606
timestamp 1586364061
transform 1 0 332856 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_3618
timestamp 1586364061
transform 1 0 333960 0 -1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_301
timestamp 1586364061
transform 1 0 335064 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_2_3631
timestamp 1586364061
transform 1 0 335156 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_3643
timestamp 1586364061
transform 1 0 336260 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_3655
timestamp 1586364061
transform 1 0 337364 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_3667
timestamp 1586364061
transform 1 0 338468 0 -1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_302
timestamp 1586364061
transform 1 0 340676 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_2_3679
timestamp 1586364061
transform 1 0 339572 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_3692
timestamp 1586364061
transform 1 0 340768 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_3704
timestamp 1586364061
transform 1 0 341872 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_3716
timestamp 1586364061
transform 1 0 342976 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_3728
timestamp 1586364061
transform 1 0 344080 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_3740
timestamp 1586364061
transform 1 0 345184 0 -1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_303
timestamp 1586364061
transform 1 0 346288 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_2_3753
timestamp 1586364061
transform 1 0 346380 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_3765
timestamp 1586364061
transform 1 0 347484 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_3777
timestamp 1586364061
transform 1 0 348588 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_3789
timestamp 1586364061
transform 1 0 349692 0 -1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_304
timestamp 1586364061
transform 1 0 351900 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_2_3801
timestamp 1586364061
transform 1 0 350796 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_3814
timestamp 1586364061
transform 1 0 351992 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_3826
timestamp 1586364061
transform 1 0 353096 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_3838
timestamp 1586364061
transform 1 0 354200 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_3850
timestamp 1586364061
transform 1 0 355304 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_3862
timestamp 1586364061
transform 1 0 356408 0 -1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_305
timestamp 1586364061
transform 1 0 357512 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_2_3875
timestamp 1586364061
transform 1 0 357604 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_3887
timestamp 1586364061
transform 1 0 358708 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_3899
timestamp 1586364061
transform 1 0 359812 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_3911
timestamp 1586364061
transform 1 0 360916 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_3923
timestamp 1586364061
transform 1 0 362020 0 -1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_306
timestamp 1586364061
transform 1 0 363124 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_2_3936
timestamp 1586364061
transform 1 0 363216 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_3948
timestamp 1586364061
transform 1 0 364320 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_3960
timestamp 1586364061
transform 1 0 365424 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_3972
timestamp 1586364061
transform 1 0 366528 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_3984
timestamp 1586364061
transform 1 0 367632 0 -1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_307
timestamp 1586364061
transform 1 0 368736 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_2_3997
timestamp 1586364061
transform 1 0 368828 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_4009
timestamp 1586364061
transform 1 0 369932 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_4021
timestamp 1586364061
transform 1 0 371036 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_4033
timestamp 1586364061
transform 1 0 372140 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_4045
timestamp 1586364061
transform 1 0 373244 0 -1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_308
timestamp 1586364061
transform 1 0 374348 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_2_4058
timestamp 1586364061
transform 1 0 374440 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_4070
timestamp 1586364061
transform 1 0 375544 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_4082
timestamp 1586364061
transform 1 0 376648 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_4094
timestamp 1586364061
transform 1 0 377752 0 -1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_309
timestamp 1586364061
transform 1 0 379960 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_2_4106
timestamp 1586364061
transform 1 0 378856 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_4119
timestamp 1586364061
transform 1 0 380052 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_4131
timestamp 1586364061
transform 1 0 381156 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_4143
timestamp 1586364061
transform 1 0 382260 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_4155
timestamp 1586364061
transform 1 0 383364 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_4167
timestamp 1586364061
transform 1 0 384468 0 -1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_310
timestamp 1586364061
transform 1 0 385572 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_2_4180
timestamp 1586364061
transform 1 0 385664 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_4192
timestamp 1586364061
transform 1 0 386768 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_4204
timestamp 1586364061
transform 1 0 387872 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_4216
timestamp 1586364061
transform 1 0 388976 0 -1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_311
timestamp 1586364061
transform 1 0 391184 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_2_4228
timestamp 1586364061
transform 1 0 390080 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_4241
timestamp 1586364061
transform 1 0 391276 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_4253
timestamp 1586364061
transform 1 0 392380 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_4265
timestamp 1586364061
transform 1 0 393484 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_4277
timestamp 1586364061
transform 1 0 394588 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_4289
timestamp 1586364061
transform 1 0 395692 0 -1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_312
timestamp 1586364061
transform 1 0 396796 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_2_4302
timestamp 1586364061
transform 1 0 396888 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_4314
timestamp 1586364061
transform 1 0 397992 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_4326
timestamp 1586364061
transform 1 0 399096 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_4338
timestamp 1586364061
transform 1 0 400200 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_4350
timestamp 1586364061
transform 1 0 401304 0 -1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_313
timestamp 1586364061
transform 1 0 402408 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_2_4363
timestamp 1586364061
transform 1 0 402500 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_4375
timestamp 1586364061
transform 1 0 403604 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_4387
timestamp 1586364061
transform 1 0 404708 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_4399
timestamp 1586364061
transform 1 0 405812 0 -1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_314
timestamp 1586364061
transform 1 0 408020 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_2_4411
timestamp 1586364061
transform 1 0 406916 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_4424
timestamp 1586364061
transform 1 0 408112 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_4436
timestamp 1586364061
transform 1 0 409216 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_4448
timestamp 1586364061
transform 1 0 410320 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_4460
timestamp 1586364061
transform 1 0 411424 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_4472
timestamp 1586364061
transform 1 0 412528 0 -1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_315
timestamp 1586364061
transform 1 0 413632 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_2_4485
timestamp 1586364061
transform 1 0 413724 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_4497
timestamp 1586364061
transform 1 0 414828 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_4509
timestamp 1586364061
transform 1 0 415932 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_4521
timestamp 1586364061
transform 1 0 417036 0 -1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_316
timestamp 1586364061
transform 1 0 419244 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_2_4533
timestamp 1586364061
transform 1 0 418140 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_4546
timestamp 1586364061
transform 1 0 419336 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_4558
timestamp 1586364061
transform 1 0 420440 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_3  PHY_5
timestamp 1586364061
transform -1 0 422832 0 -1 3808
box -38 -48 314 592
use scs8hd_decap_8  FILLER_2_4570
timestamp 1586364061
transform 1 0 421544 0 -1 3808
box -38 -48 774 592
use scs8hd_decap_3  FILLER_2_4578
timestamp 1586364061
transform 1 0 422280 0 -1 3808
box -38 -48 314 592
use scs8hd_decap_3  PHY_6
timestamp 1586364061
transform 1 0 1104 0 1 3808
box -38 -48 314 592
use scs8hd_decap_12  FILLER_3_3
timestamp 1586364061
transform 1 0 1380 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_15
timestamp 1586364061
transform 1 0 2484 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_27
timestamp 1586364061
transform 1 0 3588 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_39
timestamp 1586364061
transform 1 0 4692 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_3_51
timestamp 1586364061
transform 1 0 5796 0 1 3808
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_317
timestamp 1586364061
transform 1 0 6716 0 1 3808
box -38 -48 130 592
use scs8hd_fill_2  FILLER_3_59
timestamp 1586364061
transform 1 0 6532 0 1 3808
box -38 -48 222 592
use scs8hd_decap_12  FILLER_3_62
timestamp 1586364061
transform 1 0 6808 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_74
timestamp 1586364061
transform 1 0 7912 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_86
timestamp 1586364061
transform 1 0 9016 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_98
timestamp 1586364061
transform 1 0 10120 0 1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_318
timestamp 1586364061
transform 1 0 12328 0 1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_3_110
timestamp 1586364061
transform 1 0 11224 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_123
timestamp 1586364061
transform 1 0 12420 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_135
timestamp 1586364061
transform 1 0 13524 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_147
timestamp 1586364061
transform 1 0 14628 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_159
timestamp 1586364061
transform 1 0 15732 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_171
timestamp 1586364061
transform 1 0 16836 0 1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_319
timestamp 1586364061
transform 1 0 17940 0 1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_3_184
timestamp 1586364061
transform 1 0 18032 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_196
timestamp 1586364061
transform 1 0 19136 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_208
timestamp 1586364061
transform 1 0 20240 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_220
timestamp 1586364061
transform 1 0 21344 0 1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_320
timestamp 1586364061
transform 1 0 23552 0 1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_3_232
timestamp 1586364061
transform 1 0 22448 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_245
timestamp 1586364061
transform 1 0 23644 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_257
timestamp 1586364061
transform 1 0 24748 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_269
timestamp 1586364061
transform 1 0 25852 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_281
timestamp 1586364061
transform 1 0 26956 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_293
timestamp 1586364061
transform 1 0 28060 0 1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_321
timestamp 1586364061
transform 1 0 29164 0 1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_3_306
timestamp 1586364061
transform 1 0 29256 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_318
timestamp 1586364061
transform 1 0 30360 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_330
timestamp 1586364061
transform 1 0 31464 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_342
timestamp 1586364061
transform 1 0 32568 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_354
timestamp 1586364061
transform 1 0 33672 0 1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_322
timestamp 1586364061
transform 1 0 34776 0 1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_3_367
timestamp 1586364061
transform 1 0 34868 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_379
timestamp 1586364061
transform 1 0 35972 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_391
timestamp 1586364061
transform 1 0 37076 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_403
timestamp 1586364061
transform 1 0 38180 0 1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_323
timestamp 1586364061
transform 1 0 40388 0 1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_3_415
timestamp 1586364061
transform 1 0 39284 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_428
timestamp 1586364061
transform 1 0 40480 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_440
timestamp 1586364061
transform 1 0 41584 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_452
timestamp 1586364061
transform 1 0 42688 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_464
timestamp 1586364061
transform 1 0 43792 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_476
timestamp 1586364061
transform 1 0 44896 0 1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_324
timestamp 1586364061
transform 1 0 46000 0 1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_3_489
timestamp 1586364061
transform 1 0 46092 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_501
timestamp 1586364061
transform 1 0 47196 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_513
timestamp 1586364061
transform 1 0 48300 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_525
timestamp 1586364061
transform 1 0 49404 0 1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_325
timestamp 1586364061
transform 1 0 51612 0 1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_3_537
timestamp 1586364061
transform 1 0 50508 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_550
timestamp 1586364061
transform 1 0 51704 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_562
timestamp 1586364061
transform 1 0 52808 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_574
timestamp 1586364061
transform 1 0 53912 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_586
timestamp 1586364061
transform 1 0 55016 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_598
timestamp 1586364061
transform 1 0 56120 0 1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_326
timestamp 1586364061
transform 1 0 57224 0 1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_3_611
timestamp 1586364061
transform 1 0 57316 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_623
timestamp 1586364061
transform 1 0 58420 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_635
timestamp 1586364061
transform 1 0 59524 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_647
timestamp 1586364061
transform 1 0 60628 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_659
timestamp 1586364061
transform 1 0 61732 0 1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_327
timestamp 1586364061
transform 1 0 62836 0 1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_3_672
timestamp 1586364061
transform 1 0 62928 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_684
timestamp 1586364061
transform 1 0 64032 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_696
timestamp 1586364061
transform 1 0 65136 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_708
timestamp 1586364061
transform 1 0 66240 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_720
timestamp 1586364061
transform 1 0 67344 0 1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_328
timestamp 1586364061
transform 1 0 68448 0 1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_3_733
timestamp 1586364061
transform 1 0 68540 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_745
timestamp 1586364061
transform 1 0 69644 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_757
timestamp 1586364061
transform 1 0 70748 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_769
timestamp 1586364061
transform 1 0 71852 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_781
timestamp 1586364061
transform 1 0 72956 0 1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_329
timestamp 1586364061
transform 1 0 74060 0 1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_3_794
timestamp 1586364061
transform 1 0 74152 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_806
timestamp 1586364061
transform 1 0 75256 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_818
timestamp 1586364061
transform 1 0 76360 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_830
timestamp 1586364061
transform 1 0 77464 0 1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_330
timestamp 1586364061
transform 1 0 79672 0 1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_3_842
timestamp 1586364061
transform 1 0 78568 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_855
timestamp 1586364061
transform 1 0 79764 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_867
timestamp 1586364061
transform 1 0 80868 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_879
timestamp 1586364061
transform 1 0 81972 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_891
timestamp 1586364061
transform 1 0 83076 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_903
timestamp 1586364061
transform 1 0 84180 0 1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_331
timestamp 1586364061
transform 1 0 85284 0 1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_3_916
timestamp 1586364061
transform 1 0 85376 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_928
timestamp 1586364061
transform 1 0 86480 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_940
timestamp 1586364061
transform 1 0 87584 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_952
timestamp 1586364061
transform 1 0 88688 0 1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_332
timestamp 1586364061
transform 1 0 90896 0 1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_3_964
timestamp 1586364061
transform 1 0 89792 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_977
timestamp 1586364061
transform 1 0 90988 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_989
timestamp 1586364061
transform 1 0 92092 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_1001
timestamp 1586364061
transform 1 0 93196 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_1013
timestamp 1586364061
transform 1 0 94300 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_1025
timestamp 1586364061
transform 1 0 95404 0 1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_333
timestamp 1586364061
transform 1 0 96508 0 1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_3_1038
timestamp 1586364061
transform 1 0 96600 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_1050
timestamp 1586364061
transform 1 0 97704 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_1062
timestamp 1586364061
transform 1 0 98808 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_1074
timestamp 1586364061
transform 1 0 99912 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_1086
timestamp 1586364061
transform 1 0 101016 0 1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_334
timestamp 1586364061
transform 1 0 102120 0 1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_3_1099
timestamp 1586364061
transform 1 0 102212 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_1111
timestamp 1586364061
transform 1 0 103316 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_1123
timestamp 1586364061
transform 1 0 104420 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_1135
timestamp 1586364061
transform 1 0 105524 0 1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_335
timestamp 1586364061
transform 1 0 107732 0 1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_3_1147
timestamp 1586364061
transform 1 0 106628 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_1160
timestamp 1586364061
transform 1 0 107824 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_1172
timestamp 1586364061
transform 1 0 108928 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_1184
timestamp 1586364061
transform 1 0 110032 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_1196
timestamp 1586364061
transform 1 0 111136 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_1208
timestamp 1586364061
transform 1 0 112240 0 1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_336
timestamp 1586364061
transform 1 0 113344 0 1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_3_1221
timestamp 1586364061
transform 1 0 113436 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_1233
timestamp 1586364061
transform 1 0 114540 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_1245
timestamp 1586364061
transform 1 0 115644 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_1257
timestamp 1586364061
transform 1 0 116748 0 1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_337
timestamp 1586364061
transform 1 0 118956 0 1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_3_1269
timestamp 1586364061
transform 1 0 117852 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_1282
timestamp 1586364061
transform 1 0 119048 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_1294
timestamp 1586364061
transform 1 0 120152 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_1306
timestamp 1586364061
transform 1 0 121256 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_1318
timestamp 1586364061
transform 1 0 122360 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_1330
timestamp 1586364061
transform 1 0 123464 0 1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_338
timestamp 1586364061
transform 1 0 124568 0 1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_3_1343
timestamp 1586364061
transform 1 0 124660 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_1355
timestamp 1586364061
transform 1 0 125764 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_1367
timestamp 1586364061
transform 1 0 126868 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_1379
timestamp 1586364061
transform 1 0 127972 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_1391
timestamp 1586364061
transform 1 0 129076 0 1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_339
timestamp 1586364061
transform 1 0 130180 0 1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_3_1404
timestamp 1586364061
transform 1 0 130272 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_1416
timestamp 1586364061
transform 1 0 131376 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_1428
timestamp 1586364061
transform 1 0 132480 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_1440
timestamp 1586364061
transform 1 0 133584 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_1452
timestamp 1586364061
transform 1 0 134688 0 1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_340
timestamp 1586364061
transform 1 0 135792 0 1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_3_1465
timestamp 1586364061
transform 1 0 135884 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_1477
timestamp 1586364061
transform 1 0 136988 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_1489
timestamp 1586364061
transform 1 0 138092 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_1501
timestamp 1586364061
transform 1 0 139196 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_1513
timestamp 1586364061
transform 1 0 140300 0 1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_341
timestamp 1586364061
transform 1 0 141404 0 1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_3_1526
timestamp 1586364061
transform 1 0 141496 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_1538
timestamp 1586364061
transform 1 0 142600 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_1550
timestamp 1586364061
transform 1 0 143704 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_1562
timestamp 1586364061
transform 1 0 144808 0 1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_342
timestamp 1586364061
transform 1 0 147016 0 1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_3_1574
timestamp 1586364061
transform 1 0 145912 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_1587
timestamp 1586364061
transform 1 0 147108 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_1599
timestamp 1586364061
transform 1 0 148212 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_1611
timestamp 1586364061
transform 1 0 149316 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_1623
timestamp 1586364061
transform 1 0 150420 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_1635
timestamp 1586364061
transform 1 0 151524 0 1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_343
timestamp 1586364061
transform 1 0 152628 0 1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_3_1648
timestamp 1586364061
transform 1 0 152720 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_1660
timestamp 1586364061
transform 1 0 153824 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_1672
timestamp 1586364061
transform 1 0 154928 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_1684
timestamp 1586364061
transform 1 0 156032 0 1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_344
timestamp 1586364061
transform 1 0 158240 0 1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_3_1696
timestamp 1586364061
transform 1 0 157136 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_1709
timestamp 1586364061
transform 1 0 158332 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_1721
timestamp 1586364061
transform 1 0 159436 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_1733
timestamp 1586364061
transform 1 0 160540 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_1745
timestamp 1586364061
transform 1 0 161644 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_1757
timestamp 1586364061
transform 1 0 162748 0 1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_345
timestamp 1586364061
transform 1 0 163852 0 1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_3_1770
timestamp 1586364061
transform 1 0 163944 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_1782
timestamp 1586364061
transform 1 0 165048 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_1794
timestamp 1586364061
transform 1 0 166152 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_1806
timestamp 1586364061
transform 1 0 167256 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_1818
timestamp 1586364061
transform 1 0 168360 0 1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_346
timestamp 1586364061
transform 1 0 169464 0 1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_3_1831
timestamp 1586364061
transform 1 0 169556 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_1843
timestamp 1586364061
transform 1 0 170660 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_1855
timestamp 1586364061
transform 1 0 171764 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_1867
timestamp 1586364061
transform 1 0 172868 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_1879
timestamp 1586364061
transform 1 0 173972 0 1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_347
timestamp 1586364061
transform 1 0 175076 0 1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_3_1892
timestamp 1586364061
transform 1 0 175168 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_1904
timestamp 1586364061
transform 1 0 176272 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_1916
timestamp 1586364061
transform 1 0 177376 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_1928
timestamp 1586364061
transform 1 0 178480 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_1940
timestamp 1586364061
transform 1 0 179584 0 1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_348
timestamp 1586364061
transform 1 0 180688 0 1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_3_1953
timestamp 1586364061
transform 1 0 180780 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_1965
timestamp 1586364061
transform 1 0 181884 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_1977
timestamp 1586364061
transform 1 0 182988 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_1989
timestamp 1586364061
transform 1 0 184092 0 1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_349
timestamp 1586364061
transform 1 0 186300 0 1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_3_2001
timestamp 1586364061
transform 1 0 185196 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_2014
timestamp 1586364061
transform 1 0 186392 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_2026
timestamp 1586364061
transform 1 0 187496 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_2038
timestamp 1586364061
transform 1 0 188600 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_2050
timestamp 1586364061
transform 1 0 189704 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_2062
timestamp 1586364061
transform 1 0 190808 0 1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_350
timestamp 1586364061
transform 1 0 191912 0 1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_3_2075
timestamp 1586364061
transform 1 0 192004 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_2087
timestamp 1586364061
transform 1 0 193108 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_2099
timestamp 1586364061
transform 1 0 194212 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_2111
timestamp 1586364061
transform 1 0 195316 0 1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_351
timestamp 1586364061
transform 1 0 197524 0 1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_3_2123
timestamp 1586364061
transform 1 0 196420 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_2136
timestamp 1586364061
transform 1 0 197616 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_2148
timestamp 1586364061
transform 1 0 198720 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_2160
timestamp 1586364061
transform 1 0 199824 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_2172
timestamp 1586364061
transform 1 0 200928 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_2184
timestamp 1586364061
transform 1 0 202032 0 1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_352
timestamp 1586364061
transform 1 0 203136 0 1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_3_2197
timestamp 1586364061
transform 1 0 203228 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_2209
timestamp 1586364061
transform 1 0 204332 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_2221
timestamp 1586364061
transform 1 0 205436 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_2233
timestamp 1586364061
transform 1 0 206540 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_2245
timestamp 1586364061
transform 1 0 207644 0 1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_353
timestamp 1586364061
transform 1 0 208748 0 1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_3_2258
timestamp 1586364061
transform 1 0 208840 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_2270
timestamp 1586364061
transform 1 0 209944 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_2282
timestamp 1586364061
transform 1 0 211048 0 1 3808
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA__07__B
timestamp 1586364061
transform 1 0 212612 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__07__C
timestamp 1586364061
transform 1 0 212244 0 1 3808
box -38 -48 222 592
use scs8hd_fill_1  FILLER_3_2294
timestamp 1586364061
transform 1 0 212152 0 1 3808
box -38 -48 130 592
use scs8hd_fill_2  FILLER_3_2297
timestamp 1586364061
transform 1 0 212428 0 1 3808
box -38 -48 222 592
use scs8hd_and4_4  _07_
timestamp 1586364061
transform 1 0 212796 0 1 3808
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_354
timestamp 1586364061
transform 1 0 214360 0 1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__06__A
timestamp 1586364061
transform 1 0 213808 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 214176 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_2310
timestamp 1586364061
transform 1 0 213624 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_2314
timestamp 1586364061
transform 1 0 213992 0 1 3808
box -38 -48 222 592
use scs8hd_nor4_4  _13_
timestamp 1586364061
transform 1 0 215556 0 1 3808
box -38 -48 1602 592
use scs8hd_diode_2  ANTENNA__13__A
timestamp 1586364061
transform 1 0 215372 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 215004 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__13__C
timestamp 1586364061
transform 1 0 214636 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_2319
timestamp 1586364061
transform 1 0 214452 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_2323
timestamp 1586364061
transform 1 0 214820 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_2327
timestamp 1586364061
transform 1 0 215188 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__13__D
timestamp 1586364061
transform 1 0 217304 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_2348
timestamp 1586364061
transform 1 0 217120 0 1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_3_2352
timestamp 1586364061
transform 1 0 217488 0 1 3808
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 217948 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 218316 0 1 3808
box -38 -48 222 592
use scs8hd_fill_1  FILLER_3_2356
timestamp 1586364061
transform 1 0 217856 0 1 3808
box -38 -48 130 592
use scs8hd_fill_2  FILLER_3_2359
timestamp 1586364061
transform 1 0 218132 0 1 3808
box -38 -48 222 592
use scs8hd_decap_12  FILLER_3_2363
timestamp 1586364061
transform 1 0 218500 0 1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_355
timestamp 1586364061
transform 1 0 219972 0 1 3808
box -38 -48 130 592
use scs8hd_decap_4  FILLER_3_2375
timestamp 1586364061
transform 1 0 219604 0 1 3808
box -38 -48 406 592
use scs8hd_decap_12  FILLER_3_2380
timestamp 1586364061
transform 1 0 220064 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_2392
timestamp 1586364061
transform 1 0 221168 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_2404
timestamp 1586364061
transform 1 0 222272 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_2416
timestamp 1586364061
transform 1 0 223376 0 1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_356
timestamp 1586364061
transform 1 0 225584 0 1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_3_2428
timestamp 1586364061
transform 1 0 224480 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_2441
timestamp 1586364061
transform 1 0 225676 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_2453
timestamp 1586364061
transform 1 0 226780 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_2465
timestamp 1586364061
transform 1 0 227884 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_2477
timestamp 1586364061
transform 1 0 228988 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_2489
timestamp 1586364061
transform 1 0 230092 0 1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_357
timestamp 1586364061
transform 1 0 231196 0 1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_3_2502
timestamp 1586364061
transform 1 0 231288 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_2514
timestamp 1586364061
transform 1 0 232392 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_2526
timestamp 1586364061
transform 1 0 233496 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_2538
timestamp 1586364061
transform 1 0 234600 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_2550
timestamp 1586364061
transform 1 0 235704 0 1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_358
timestamp 1586364061
transform 1 0 236808 0 1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_3_2563
timestamp 1586364061
transform 1 0 236900 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_2575
timestamp 1586364061
transform 1 0 238004 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_2587
timestamp 1586364061
transform 1 0 239108 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_2599
timestamp 1586364061
transform 1 0 240212 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_2611
timestamp 1586364061
transform 1 0 241316 0 1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_359
timestamp 1586364061
transform 1 0 242420 0 1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_3_2624
timestamp 1586364061
transform 1 0 242512 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_2636
timestamp 1586364061
transform 1 0 243616 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_2648
timestamp 1586364061
transform 1 0 244720 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_2660
timestamp 1586364061
transform 1 0 245824 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_2672
timestamp 1586364061
transform 1 0 246928 0 1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_360
timestamp 1586364061
transform 1 0 248032 0 1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_3_2685
timestamp 1586364061
transform 1 0 248124 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_2697
timestamp 1586364061
transform 1 0 249228 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_2709
timestamp 1586364061
transform 1 0 250332 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_2721
timestamp 1586364061
transform 1 0 251436 0 1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_361
timestamp 1586364061
transform 1 0 253644 0 1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_3_2733
timestamp 1586364061
transform 1 0 252540 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_2746
timestamp 1586364061
transform 1 0 253736 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_2758
timestamp 1586364061
transform 1 0 254840 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_2770
timestamp 1586364061
transform 1 0 255944 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_2782
timestamp 1586364061
transform 1 0 257048 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_2794
timestamp 1586364061
transform 1 0 258152 0 1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_362
timestamp 1586364061
transform 1 0 259256 0 1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_3_2807
timestamp 1586364061
transform 1 0 259348 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_2819
timestamp 1586364061
transform 1 0 260452 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_2831
timestamp 1586364061
transform 1 0 261556 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_2843
timestamp 1586364061
transform 1 0 262660 0 1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_363
timestamp 1586364061
transform 1 0 264868 0 1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_3_2855
timestamp 1586364061
transform 1 0 263764 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_2868
timestamp 1586364061
transform 1 0 264960 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_2880
timestamp 1586364061
transform 1 0 266064 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_2892
timestamp 1586364061
transform 1 0 267168 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_2904
timestamp 1586364061
transform 1 0 268272 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_2916
timestamp 1586364061
transform 1 0 269376 0 1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_364
timestamp 1586364061
transform 1 0 270480 0 1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_3_2929
timestamp 1586364061
transform 1 0 270572 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_2941
timestamp 1586364061
transform 1 0 271676 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_2953
timestamp 1586364061
transform 1 0 272780 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_2965
timestamp 1586364061
transform 1 0 273884 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_2977
timestamp 1586364061
transform 1 0 274988 0 1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_365
timestamp 1586364061
transform 1 0 276092 0 1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_3_2990
timestamp 1586364061
transform 1 0 276184 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_3002
timestamp 1586364061
transform 1 0 277288 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_3014
timestamp 1586364061
transform 1 0 278392 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_3026
timestamp 1586364061
transform 1 0 279496 0 1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_366
timestamp 1586364061
transform 1 0 281704 0 1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_3_3038
timestamp 1586364061
transform 1 0 280600 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_3051
timestamp 1586364061
transform 1 0 281796 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_3063
timestamp 1586364061
transform 1 0 282900 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_3075
timestamp 1586364061
transform 1 0 284004 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_3087
timestamp 1586364061
transform 1 0 285108 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_3099
timestamp 1586364061
transform 1 0 286212 0 1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_367
timestamp 1586364061
transform 1 0 287316 0 1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_3_3112
timestamp 1586364061
transform 1 0 287408 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_3124
timestamp 1586364061
transform 1 0 288512 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_3136
timestamp 1586364061
transform 1 0 289616 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_3148
timestamp 1586364061
transform 1 0 290720 0 1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_368
timestamp 1586364061
transform 1 0 292928 0 1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_3_3160
timestamp 1586364061
transform 1 0 291824 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_3173
timestamp 1586364061
transform 1 0 293020 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_3185
timestamp 1586364061
transform 1 0 294124 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_3197
timestamp 1586364061
transform 1 0 295228 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_3209
timestamp 1586364061
transform 1 0 296332 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_3221
timestamp 1586364061
transform 1 0 297436 0 1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_369
timestamp 1586364061
transform 1 0 298540 0 1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_3_3234
timestamp 1586364061
transform 1 0 298632 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_3246
timestamp 1586364061
transform 1 0 299736 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_3258
timestamp 1586364061
transform 1 0 300840 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_3270
timestamp 1586364061
transform 1 0 301944 0 1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_370
timestamp 1586364061
transform 1 0 304152 0 1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_3_3282
timestamp 1586364061
transform 1 0 303048 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_3295
timestamp 1586364061
transform 1 0 304244 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_3307
timestamp 1586364061
transform 1 0 305348 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_3319
timestamp 1586364061
transform 1 0 306452 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_3331
timestamp 1586364061
transform 1 0 307556 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_3343
timestamp 1586364061
transform 1 0 308660 0 1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_371
timestamp 1586364061
transform 1 0 309764 0 1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_3_3356
timestamp 1586364061
transform 1 0 309856 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_3368
timestamp 1586364061
transform 1 0 310960 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_3380
timestamp 1586364061
transform 1 0 312064 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_3392
timestamp 1586364061
transform 1 0 313168 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_3404
timestamp 1586364061
transform 1 0 314272 0 1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_372
timestamp 1586364061
transform 1 0 315376 0 1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_3_3417
timestamp 1586364061
transform 1 0 315468 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_3429
timestamp 1586364061
transform 1 0 316572 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_3441
timestamp 1586364061
transform 1 0 317676 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_3453
timestamp 1586364061
transform 1 0 318780 0 1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_373
timestamp 1586364061
transform 1 0 320988 0 1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_3_3465
timestamp 1586364061
transform 1 0 319884 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_3478
timestamp 1586364061
transform 1 0 321080 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_3490
timestamp 1586364061
transform 1 0 322184 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_3502
timestamp 1586364061
transform 1 0 323288 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_3514
timestamp 1586364061
transform 1 0 324392 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_3526
timestamp 1586364061
transform 1 0 325496 0 1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_374
timestamp 1586364061
transform 1 0 326600 0 1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_3_3539
timestamp 1586364061
transform 1 0 326692 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_3551
timestamp 1586364061
transform 1 0 327796 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_3563
timestamp 1586364061
transform 1 0 328900 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_3575
timestamp 1586364061
transform 1 0 330004 0 1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_375
timestamp 1586364061
transform 1 0 332212 0 1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_3_3587
timestamp 1586364061
transform 1 0 331108 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_3600
timestamp 1586364061
transform 1 0 332304 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_3612
timestamp 1586364061
transform 1 0 333408 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_3624
timestamp 1586364061
transform 1 0 334512 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_3636
timestamp 1586364061
transform 1 0 335616 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_3648
timestamp 1586364061
transform 1 0 336720 0 1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_376
timestamp 1586364061
transform 1 0 337824 0 1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_3_3661
timestamp 1586364061
transform 1 0 337916 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_3673
timestamp 1586364061
transform 1 0 339020 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_3685
timestamp 1586364061
transform 1 0 340124 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_3697
timestamp 1586364061
transform 1 0 341228 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_3709
timestamp 1586364061
transform 1 0 342332 0 1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_377
timestamp 1586364061
transform 1 0 343436 0 1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_3_3722
timestamp 1586364061
transform 1 0 343528 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_3734
timestamp 1586364061
transform 1 0 344632 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_3746
timestamp 1586364061
transform 1 0 345736 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_3758
timestamp 1586364061
transform 1 0 346840 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_3770
timestamp 1586364061
transform 1 0 347944 0 1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_378
timestamp 1586364061
transform 1 0 349048 0 1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_3_3783
timestamp 1586364061
transform 1 0 349140 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_3795
timestamp 1586364061
transform 1 0 350244 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_3807
timestamp 1586364061
transform 1 0 351348 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_3819
timestamp 1586364061
transform 1 0 352452 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_3831
timestamp 1586364061
transform 1 0 353556 0 1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_379
timestamp 1586364061
transform 1 0 354660 0 1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_3_3844
timestamp 1586364061
transform 1 0 354752 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_3856
timestamp 1586364061
transform 1 0 355856 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_3868
timestamp 1586364061
transform 1 0 356960 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_3880
timestamp 1586364061
transform 1 0 358064 0 1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_380
timestamp 1586364061
transform 1 0 360272 0 1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_3_3892
timestamp 1586364061
transform 1 0 359168 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_3905
timestamp 1586364061
transform 1 0 360364 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_3917
timestamp 1586364061
transform 1 0 361468 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_3929
timestamp 1586364061
transform 1 0 362572 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_3941
timestamp 1586364061
transform 1 0 363676 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_3953
timestamp 1586364061
transform 1 0 364780 0 1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_381
timestamp 1586364061
transform 1 0 365884 0 1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_3_3966
timestamp 1586364061
transform 1 0 365976 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_3978
timestamp 1586364061
transform 1 0 367080 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_3990
timestamp 1586364061
transform 1 0 368184 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_4002
timestamp 1586364061
transform 1 0 369288 0 1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_382
timestamp 1586364061
transform 1 0 371496 0 1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_3_4014
timestamp 1586364061
transform 1 0 370392 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_4027
timestamp 1586364061
transform 1 0 371588 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_4039
timestamp 1586364061
transform 1 0 372692 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_4051
timestamp 1586364061
transform 1 0 373796 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_4063
timestamp 1586364061
transform 1 0 374900 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_4075
timestamp 1586364061
transform 1 0 376004 0 1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_383
timestamp 1586364061
transform 1 0 377108 0 1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_3_4088
timestamp 1586364061
transform 1 0 377200 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_4100
timestamp 1586364061
transform 1 0 378304 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_4112
timestamp 1586364061
transform 1 0 379408 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_4124
timestamp 1586364061
transform 1 0 380512 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_4136
timestamp 1586364061
transform 1 0 381616 0 1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_384
timestamp 1586364061
transform 1 0 382720 0 1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_3_4149
timestamp 1586364061
transform 1 0 382812 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_4161
timestamp 1586364061
transform 1 0 383916 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_4173
timestamp 1586364061
transform 1 0 385020 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_4185
timestamp 1586364061
transform 1 0 386124 0 1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_385
timestamp 1586364061
transform 1 0 388332 0 1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_3_4197
timestamp 1586364061
transform 1 0 387228 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_4210
timestamp 1586364061
transform 1 0 388424 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_4222
timestamp 1586364061
transform 1 0 389528 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_4234
timestamp 1586364061
transform 1 0 390632 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_4246
timestamp 1586364061
transform 1 0 391736 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_4258
timestamp 1586364061
transform 1 0 392840 0 1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_386
timestamp 1586364061
transform 1 0 393944 0 1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_3_4271
timestamp 1586364061
transform 1 0 394036 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_4283
timestamp 1586364061
transform 1 0 395140 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_4295
timestamp 1586364061
transform 1 0 396244 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_4307
timestamp 1586364061
transform 1 0 397348 0 1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_387
timestamp 1586364061
transform 1 0 399556 0 1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_3_4319
timestamp 1586364061
transform 1 0 398452 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_4332
timestamp 1586364061
transform 1 0 399648 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_4344
timestamp 1586364061
transform 1 0 400752 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_4356
timestamp 1586364061
transform 1 0 401856 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_4368
timestamp 1586364061
transform 1 0 402960 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_4380
timestamp 1586364061
transform 1 0 404064 0 1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_388
timestamp 1586364061
transform 1 0 405168 0 1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_3_4393
timestamp 1586364061
transform 1 0 405260 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_4405
timestamp 1586364061
transform 1 0 406364 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_4417
timestamp 1586364061
transform 1 0 407468 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_4429
timestamp 1586364061
transform 1 0 408572 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_4441
timestamp 1586364061
transform 1 0 409676 0 1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_389
timestamp 1586364061
transform 1 0 410780 0 1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_3_4454
timestamp 1586364061
transform 1 0 410872 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_4466
timestamp 1586364061
transform 1 0 411976 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_4478
timestamp 1586364061
transform 1 0 413080 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_4490
timestamp 1586364061
transform 1 0 414184 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_4502
timestamp 1586364061
transform 1 0 415288 0 1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_390
timestamp 1586364061
transform 1 0 416392 0 1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_3_4515
timestamp 1586364061
transform 1 0 416484 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_4527
timestamp 1586364061
transform 1 0 417588 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_4539
timestamp 1586364061
transform 1 0 418692 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_4551
timestamp 1586364061
transform 1 0 419796 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_4563
timestamp 1586364061
transform 1 0 420900 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_3  PHY_7
timestamp 1586364061
transform -1 0 422832 0 1 3808
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_391
timestamp 1586364061
transform 1 0 422004 0 1 3808
box -38 -48 130 592
use scs8hd_decap_4  FILLER_3_4576
timestamp 1586364061
transform 1 0 422096 0 1 3808
box -38 -48 406 592
use scs8hd_fill_1  FILLER_3_4580
timestamp 1586364061
transform 1 0 422464 0 1 3808
box -38 -48 130 592
use scs8hd_decap_3  PHY_8
timestamp 1586364061
transform 1 0 1104 0 -1 4896
box -38 -48 314 592
use scs8hd_decap_12  FILLER_4_3
timestamp 1586364061
transform 1 0 1380 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_15
timestamp 1586364061
transform 1 0 2484 0 -1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_392
timestamp 1586364061
transform 1 0 3956 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_4  FILLER_4_27
timestamp 1586364061
transform 1 0 3588 0 -1 4896
box -38 -48 406 592
use scs8hd_decap_12  FILLER_4_32
timestamp 1586364061
transform 1 0 4048 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_44
timestamp 1586364061
transform 1 0 5152 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_56
timestamp 1586364061
transform 1 0 6256 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_68
timestamp 1586364061
transform 1 0 7360 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_80
timestamp 1586364061
transform 1 0 8464 0 -1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_393
timestamp 1586364061
transform 1 0 9568 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_4_93
timestamp 1586364061
transform 1 0 9660 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_105
timestamp 1586364061
transform 1 0 10764 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_117
timestamp 1586364061
transform 1 0 11868 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_129
timestamp 1586364061
transform 1 0 12972 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_141
timestamp 1586364061
transform 1 0 14076 0 -1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_394
timestamp 1586364061
transform 1 0 15180 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_4_154
timestamp 1586364061
transform 1 0 15272 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_166
timestamp 1586364061
transform 1 0 16376 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_178
timestamp 1586364061
transform 1 0 17480 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_190
timestamp 1586364061
transform 1 0 18584 0 -1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_395
timestamp 1586364061
transform 1 0 20792 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_4_202
timestamp 1586364061
transform 1 0 19688 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_215
timestamp 1586364061
transform 1 0 20884 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_227
timestamp 1586364061
transform 1 0 21988 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_239
timestamp 1586364061
transform 1 0 23092 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_251
timestamp 1586364061
transform 1 0 24196 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_263
timestamp 1586364061
transform 1 0 25300 0 -1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_396
timestamp 1586364061
transform 1 0 26404 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_4_276
timestamp 1586364061
transform 1 0 26496 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_288
timestamp 1586364061
transform 1 0 27600 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_300
timestamp 1586364061
transform 1 0 28704 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_312
timestamp 1586364061
transform 1 0 29808 0 -1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_397
timestamp 1586364061
transform 1 0 32016 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_4_324
timestamp 1586364061
transform 1 0 30912 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_337
timestamp 1586364061
transform 1 0 32108 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_349
timestamp 1586364061
transform 1 0 33212 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_361
timestamp 1586364061
transform 1 0 34316 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_373
timestamp 1586364061
transform 1 0 35420 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_385
timestamp 1586364061
transform 1 0 36524 0 -1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_398
timestamp 1586364061
transform 1 0 37628 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_4_398
timestamp 1586364061
transform 1 0 37720 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_410
timestamp 1586364061
transform 1 0 38824 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_422
timestamp 1586364061
transform 1 0 39928 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_434
timestamp 1586364061
transform 1 0 41032 0 -1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_399
timestamp 1586364061
transform 1 0 43240 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_4_446
timestamp 1586364061
transform 1 0 42136 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_459
timestamp 1586364061
transform 1 0 43332 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_471
timestamp 1586364061
transform 1 0 44436 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_483
timestamp 1586364061
transform 1 0 45540 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_495
timestamp 1586364061
transform 1 0 46644 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_507
timestamp 1586364061
transform 1 0 47748 0 -1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_400
timestamp 1586364061
transform 1 0 48852 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_4_520
timestamp 1586364061
transform 1 0 48944 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_532
timestamp 1586364061
transform 1 0 50048 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_544
timestamp 1586364061
transform 1 0 51152 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_556
timestamp 1586364061
transform 1 0 52256 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_568
timestamp 1586364061
transform 1 0 53360 0 -1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_401
timestamp 1586364061
transform 1 0 54464 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_4_581
timestamp 1586364061
transform 1 0 54556 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_593
timestamp 1586364061
transform 1 0 55660 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_605
timestamp 1586364061
transform 1 0 56764 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_617
timestamp 1586364061
transform 1 0 57868 0 -1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_402
timestamp 1586364061
transform 1 0 60076 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_4_629
timestamp 1586364061
transform 1 0 58972 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_642
timestamp 1586364061
transform 1 0 60168 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_654
timestamp 1586364061
transform 1 0 61272 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_666
timestamp 1586364061
transform 1 0 62376 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_678
timestamp 1586364061
transform 1 0 63480 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_690
timestamp 1586364061
transform 1 0 64584 0 -1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_403
timestamp 1586364061
transform 1 0 65688 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_4_703
timestamp 1586364061
transform 1 0 65780 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_715
timestamp 1586364061
transform 1 0 66884 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_727
timestamp 1586364061
transform 1 0 67988 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_739
timestamp 1586364061
transform 1 0 69092 0 -1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_404
timestamp 1586364061
transform 1 0 71300 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_4_751
timestamp 1586364061
transform 1 0 70196 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_764
timestamp 1586364061
transform 1 0 71392 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_776
timestamp 1586364061
transform 1 0 72496 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_788
timestamp 1586364061
transform 1 0 73600 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_800
timestamp 1586364061
transform 1 0 74704 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_812
timestamp 1586364061
transform 1 0 75808 0 -1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_405
timestamp 1586364061
transform 1 0 76912 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_4_825
timestamp 1586364061
transform 1 0 77004 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_837
timestamp 1586364061
transform 1 0 78108 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_849
timestamp 1586364061
transform 1 0 79212 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_861
timestamp 1586364061
transform 1 0 80316 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_873
timestamp 1586364061
transform 1 0 81420 0 -1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_406
timestamp 1586364061
transform 1 0 82524 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_4_886
timestamp 1586364061
transform 1 0 82616 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_898
timestamp 1586364061
transform 1 0 83720 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_910
timestamp 1586364061
transform 1 0 84824 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_922
timestamp 1586364061
transform 1 0 85928 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_934
timestamp 1586364061
transform 1 0 87032 0 -1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_407
timestamp 1586364061
transform 1 0 88136 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_4_947
timestamp 1586364061
transform 1 0 88228 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_959
timestamp 1586364061
transform 1 0 89332 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_971
timestamp 1586364061
transform 1 0 90436 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_983
timestamp 1586364061
transform 1 0 91540 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_995
timestamp 1586364061
transform 1 0 92644 0 -1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_408
timestamp 1586364061
transform 1 0 93748 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_4_1008
timestamp 1586364061
transform 1 0 93840 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_1020
timestamp 1586364061
transform 1 0 94944 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_1032
timestamp 1586364061
transform 1 0 96048 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_1044
timestamp 1586364061
transform 1 0 97152 0 -1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_409
timestamp 1586364061
transform 1 0 99360 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_4_1056
timestamp 1586364061
transform 1 0 98256 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_1069
timestamp 1586364061
transform 1 0 99452 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_1081
timestamp 1586364061
transform 1 0 100556 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_1093
timestamp 1586364061
transform 1 0 101660 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_1105
timestamp 1586364061
transform 1 0 102764 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_1117
timestamp 1586364061
transform 1 0 103868 0 -1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_410
timestamp 1586364061
transform 1 0 104972 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_4_1130
timestamp 1586364061
transform 1 0 105064 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_1142
timestamp 1586364061
transform 1 0 106168 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_1154
timestamp 1586364061
transform 1 0 107272 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_1166
timestamp 1586364061
transform 1 0 108376 0 -1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_411
timestamp 1586364061
transform 1 0 110584 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_4_1178
timestamp 1586364061
transform 1 0 109480 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_1191
timestamp 1586364061
transform 1 0 110676 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_1203
timestamp 1586364061
transform 1 0 111780 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_1215
timestamp 1586364061
transform 1 0 112884 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_1227
timestamp 1586364061
transform 1 0 113988 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_1239
timestamp 1586364061
transform 1 0 115092 0 -1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_412
timestamp 1586364061
transform 1 0 116196 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_4_1252
timestamp 1586364061
transform 1 0 116288 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_1264
timestamp 1586364061
transform 1 0 117392 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_1276
timestamp 1586364061
transform 1 0 118496 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_1288
timestamp 1586364061
transform 1 0 119600 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_1300
timestamp 1586364061
transform 1 0 120704 0 -1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_413
timestamp 1586364061
transform 1 0 121808 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_4_1313
timestamp 1586364061
transform 1 0 121900 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_1325
timestamp 1586364061
transform 1 0 123004 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_1337
timestamp 1586364061
transform 1 0 124108 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_1349
timestamp 1586364061
transform 1 0 125212 0 -1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_414
timestamp 1586364061
transform 1 0 127420 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_4_1361
timestamp 1586364061
transform 1 0 126316 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_1374
timestamp 1586364061
transform 1 0 127512 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_1386
timestamp 1586364061
transform 1 0 128616 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_1398
timestamp 1586364061
transform 1 0 129720 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_1410
timestamp 1586364061
transform 1 0 130824 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_1422
timestamp 1586364061
transform 1 0 131928 0 -1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_415
timestamp 1586364061
transform 1 0 133032 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_4_1435
timestamp 1586364061
transform 1 0 133124 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_1447
timestamp 1586364061
transform 1 0 134228 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_1459
timestamp 1586364061
transform 1 0 135332 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_1471
timestamp 1586364061
transform 1 0 136436 0 -1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_416
timestamp 1586364061
transform 1 0 138644 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_4_1483
timestamp 1586364061
transform 1 0 137540 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_1496
timestamp 1586364061
transform 1 0 138736 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_1508
timestamp 1586364061
transform 1 0 139840 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_1520
timestamp 1586364061
transform 1 0 140944 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_1532
timestamp 1586364061
transform 1 0 142048 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_1544
timestamp 1586364061
transform 1 0 143152 0 -1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_417
timestamp 1586364061
transform 1 0 144256 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_4_1557
timestamp 1586364061
transform 1 0 144348 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_1569
timestamp 1586364061
transform 1 0 145452 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_1581
timestamp 1586364061
transform 1 0 146556 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_1593
timestamp 1586364061
transform 1 0 147660 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_1605
timestamp 1586364061
transform 1 0 148764 0 -1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_418
timestamp 1586364061
transform 1 0 149868 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_4_1618
timestamp 1586364061
transform 1 0 149960 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_1630
timestamp 1586364061
transform 1 0 151064 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_1642
timestamp 1586364061
transform 1 0 152168 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_1654
timestamp 1586364061
transform 1 0 153272 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_1666
timestamp 1586364061
transform 1 0 154376 0 -1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_419
timestamp 1586364061
transform 1 0 155480 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_4_1679
timestamp 1586364061
transform 1 0 155572 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_1691
timestamp 1586364061
transform 1 0 156676 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_1703
timestamp 1586364061
transform 1 0 157780 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_1715
timestamp 1586364061
transform 1 0 158884 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_1727
timestamp 1586364061
transform 1 0 159988 0 -1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_420
timestamp 1586364061
transform 1 0 161092 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_4_1740
timestamp 1586364061
transform 1 0 161184 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_1752
timestamp 1586364061
transform 1 0 162288 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_1764
timestamp 1586364061
transform 1 0 163392 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_1776
timestamp 1586364061
transform 1 0 164496 0 -1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_421
timestamp 1586364061
transform 1 0 166704 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_4_1788
timestamp 1586364061
transform 1 0 165600 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_1801
timestamp 1586364061
transform 1 0 166796 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_1813
timestamp 1586364061
transform 1 0 167900 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_1825
timestamp 1586364061
transform 1 0 169004 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_1837
timestamp 1586364061
transform 1 0 170108 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_1849
timestamp 1586364061
transform 1 0 171212 0 -1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_422
timestamp 1586364061
transform 1 0 172316 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_4_1862
timestamp 1586364061
transform 1 0 172408 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_1874
timestamp 1586364061
transform 1 0 173512 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_1886
timestamp 1586364061
transform 1 0 174616 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_1898
timestamp 1586364061
transform 1 0 175720 0 -1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_423
timestamp 1586364061
transform 1 0 177928 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_4_1910
timestamp 1586364061
transform 1 0 176824 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_1923
timestamp 1586364061
transform 1 0 178020 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_1935
timestamp 1586364061
transform 1 0 179124 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_1947
timestamp 1586364061
transform 1 0 180228 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_1959
timestamp 1586364061
transform 1 0 181332 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_1971
timestamp 1586364061
transform 1 0 182436 0 -1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_424
timestamp 1586364061
transform 1 0 183540 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_4_1984
timestamp 1586364061
transform 1 0 183632 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_1996
timestamp 1586364061
transform 1 0 184736 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_2008
timestamp 1586364061
transform 1 0 185840 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_2020
timestamp 1586364061
transform 1 0 186944 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_2032
timestamp 1586364061
transform 1 0 188048 0 -1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_425
timestamp 1586364061
transform 1 0 189152 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_4_2045
timestamp 1586364061
transform 1 0 189244 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_2057
timestamp 1586364061
transform 1 0 190348 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_2069
timestamp 1586364061
transform 1 0 191452 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_2081
timestamp 1586364061
transform 1 0 192556 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_2093
timestamp 1586364061
transform 1 0 193660 0 -1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_426
timestamp 1586364061
transform 1 0 194764 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_4_2106
timestamp 1586364061
transform 1 0 194856 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_2118
timestamp 1586364061
transform 1 0 195960 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_2130
timestamp 1586364061
transform 1 0 197064 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_2142
timestamp 1586364061
transform 1 0 198168 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_2154
timestamp 1586364061
transform 1 0 199272 0 -1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_427
timestamp 1586364061
transform 1 0 200376 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_4_2167
timestamp 1586364061
transform 1 0 200468 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_2179
timestamp 1586364061
transform 1 0 201572 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_2191
timestamp 1586364061
transform 1 0 202676 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_2203
timestamp 1586364061
transform 1 0 203780 0 -1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_428
timestamp 1586364061
transform 1 0 205988 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_4_2215
timestamp 1586364061
transform 1 0 204884 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_2228
timestamp 1586364061
transform 1 0 206080 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_2240
timestamp 1586364061
transform 1 0 207184 0 -1 4896
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA_logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer_TEB
timestamp 1586364061
transform 1 0 208840 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_6  FILLER_4_2252
timestamp 1586364061
transform 1 0 208288 0 -1 4896
box -38 -48 590 592
use scs8hd_decap_12  FILLER_4_2260
timestamp 1586364061
transform 1 0 209024 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_2272
timestamp 1586364061
transform 1 0 210128 0 -1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_429
timestamp 1586364061
transform 1 0 211600 0 -1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 212244 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_4_2284
timestamp 1586364061
transform 1 0 211232 0 -1 4896
box -38 -48 406 592
use scs8hd_decap_6  FILLER_4_2289
timestamp 1586364061
transform 1 0 211692 0 -1 4896
box -38 -48 590 592
use scs8hd_decap_4  FILLER_4_2297
timestamp 1586364061
transform 1 0 212428 0 -1 4896
box -38 -48 406 592
use scs8hd_inv_8  _06_
timestamp 1586364061
transform 1 0 213716 0 -1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__07__A
timestamp 1586364061
transform 1 0 212796 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_8  FILLER_4_2303
timestamp 1586364061
transform 1 0 212980 0 -1 4896
box -38 -48 774 592
use scs8hd_lpflow_inputisolatch_1  logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.LATCH_0_.latch
timestamp 1586364061
transform 1 0 215280 0 -1 4896
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA__11__A
timestamp 1586364061
transform 1 0 215096 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__13__B
timestamp 1586364061
transform 1 0 214728 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_2320
timestamp 1586364061
transform 1 0 214544 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_2324
timestamp 1586364061
transform 1 0 214912 0 -1 4896
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_430
timestamp 1586364061
transform 1 0 217212 0 -1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__10__B
timestamp 1586364061
transform 1 0 216752 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_4_2339
timestamp 1586364061
transform 1 0 216292 0 -1 4896
box -38 -48 406 592
use scs8hd_fill_1  FILLER_4_2343
timestamp 1586364061
transform 1 0 216660 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_3  FILLER_4_2346
timestamp 1586364061
transform 1 0 216936 0 -1 4896
box -38 -48 314 592
use scs8hd_decap_6  FILLER_4_2350
timestamp 1586364061
transform 1 0 217304 0 -1 4896
box -38 -48 590 592
use scs8hd_lpflow_inputisolatch_1  logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.LATCH_0_.latch
timestamp 1586364061
transform 1 0 217948 0 -1 4896
box -38 -48 1050 592
use scs8hd_fill_1  FILLER_4_2356
timestamp 1586364061
transform 1 0 217856 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_4_2368
timestamp 1586364061
transform 1 0 218960 0 -1 4896
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA_logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 220524 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_4_2380
timestamp 1586364061
transform 1 0 220064 0 -1 4896
box -38 -48 406 592
use scs8hd_fill_1  FILLER_4_2384
timestamp 1586364061
transform 1 0 220432 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_4_2387
timestamp 1586364061
transform 1 0 220708 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_4_2399
timestamp 1586364061
transform 1 0 221812 0 -1 4896
box -38 -48 774 592
use scs8hd_decap_3  FILLER_4_2407
timestamp 1586364061
transform 1 0 222548 0 -1 4896
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_431
timestamp 1586364061
transform 1 0 222824 0 -1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer_TEB
timestamp 1586364061
transform 1 0 224020 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_12  FILLER_4_2411
timestamp 1586364061
transform 1 0 222916 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_2425
timestamp 1586364061
transform 1 0 224204 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_2437
timestamp 1586364061
transform 1 0 225308 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_2449
timestamp 1586364061
transform 1 0 226412 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_4_2461
timestamp 1586364061
transform 1 0 227516 0 -1 4896
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_432
timestamp 1586364061
transform 1 0 228436 0 -1 4896
box -38 -48 130 592
use scs8hd_fill_2  FILLER_4_2469
timestamp 1586364061
transform 1 0 228252 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_12  FILLER_4_2472
timestamp 1586364061
transform 1 0 228528 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_2484
timestamp 1586364061
transform 1 0 229632 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_2496
timestamp 1586364061
transform 1 0 230736 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_2508
timestamp 1586364061
transform 1 0 231840 0 -1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_433
timestamp 1586364061
transform 1 0 234048 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_4_2520
timestamp 1586364061
transform 1 0 232944 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_2533
timestamp 1586364061
transform 1 0 234140 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_2545
timestamp 1586364061
transform 1 0 235244 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_2557
timestamp 1586364061
transform 1 0 236348 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_2569
timestamp 1586364061
transform 1 0 237452 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_2581
timestamp 1586364061
transform 1 0 238556 0 -1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_434
timestamp 1586364061
transform 1 0 239660 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_4_2594
timestamp 1586364061
transform 1 0 239752 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_2606
timestamp 1586364061
transform 1 0 240856 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_2618
timestamp 1586364061
transform 1 0 241960 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_2630
timestamp 1586364061
transform 1 0 243064 0 -1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_435
timestamp 1586364061
transform 1 0 245272 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_4_2642
timestamp 1586364061
transform 1 0 244168 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_2655
timestamp 1586364061
transform 1 0 245364 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_2667
timestamp 1586364061
transform 1 0 246468 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_2679
timestamp 1586364061
transform 1 0 247572 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_2691
timestamp 1586364061
transform 1 0 248676 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_2703
timestamp 1586364061
transform 1 0 249780 0 -1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_436
timestamp 1586364061
transform 1 0 250884 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_4_2716
timestamp 1586364061
transform 1 0 250976 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_2728
timestamp 1586364061
transform 1 0 252080 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_2740
timestamp 1586364061
transform 1 0 253184 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_2752
timestamp 1586364061
transform 1 0 254288 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_2764
timestamp 1586364061
transform 1 0 255392 0 -1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_437
timestamp 1586364061
transform 1 0 256496 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_4_2777
timestamp 1586364061
transform 1 0 256588 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_2789
timestamp 1586364061
transform 1 0 257692 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_2801
timestamp 1586364061
transform 1 0 258796 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_2813
timestamp 1586364061
transform 1 0 259900 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_2825
timestamp 1586364061
transform 1 0 261004 0 -1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_438
timestamp 1586364061
transform 1 0 262108 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_4_2838
timestamp 1586364061
transform 1 0 262200 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_2850
timestamp 1586364061
transform 1 0 263304 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_2862
timestamp 1586364061
transform 1 0 264408 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_2874
timestamp 1586364061
transform 1 0 265512 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_2886
timestamp 1586364061
transform 1 0 266616 0 -1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_439
timestamp 1586364061
transform 1 0 267720 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_4_2899
timestamp 1586364061
transform 1 0 267812 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_2911
timestamp 1586364061
transform 1 0 268916 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_2923
timestamp 1586364061
transform 1 0 270020 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_2935
timestamp 1586364061
transform 1 0 271124 0 -1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_440
timestamp 1586364061
transform 1 0 273332 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_4_2947
timestamp 1586364061
transform 1 0 272228 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_2960
timestamp 1586364061
transform 1 0 273424 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_2972
timestamp 1586364061
transform 1 0 274528 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_2984
timestamp 1586364061
transform 1 0 275632 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_2996
timestamp 1586364061
transform 1 0 276736 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_3008
timestamp 1586364061
transform 1 0 277840 0 -1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_441
timestamp 1586364061
transform 1 0 278944 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_4_3021
timestamp 1586364061
transform 1 0 279036 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_3033
timestamp 1586364061
transform 1 0 280140 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_3045
timestamp 1586364061
transform 1 0 281244 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_3057
timestamp 1586364061
transform 1 0 282348 0 -1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_442
timestamp 1586364061
transform 1 0 284556 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_4_3069
timestamp 1586364061
transform 1 0 283452 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_3082
timestamp 1586364061
transform 1 0 284648 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_3094
timestamp 1586364061
transform 1 0 285752 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_3106
timestamp 1586364061
transform 1 0 286856 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_3118
timestamp 1586364061
transform 1 0 287960 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_3130
timestamp 1586364061
transform 1 0 289064 0 -1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_443
timestamp 1586364061
transform 1 0 290168 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_4_3143
timestamp 1586364061
transform 1 0 290260 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_3155
timestamp 1586364061
transform 1 0 291364 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_3167
timestamp 1586364061
transform 1 0 292468 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_3179
timestamp 1586364061
transform 1 0 293572 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_3191
timestamp 1586364061
transform 1 0 294676 0 -1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_444
timestamp 1586364061
transform 1 0 295780 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_4_3204
timestamp 1586364061
transform 1 0 295872 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_3216
timestamp 1586364061
transform 1 0 296976 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_3228
timestamp 1586364061
transform 1 0 298080 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_3240
timestamp 1586364061
transform 1 0 299184 0 -1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_445
timestamp 1586364061
transform 1 0 301392 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_4_3252
timestamp 1586364061
transform 1 0 300288 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_3265
timestamp 1586364061
transform 1 0 301484 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_3277
timestamp 1586364061
transform 1 0 302588 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_3289
timestamp 1586364061
transform 1 0 303692 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_3301
timestamp 1586364061
transform 1 0 304796 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_3313
timestamp 1586364061
transform 1 0 305900 0 -1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_446
timestamp 1586364061
transform 1 0 307004 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_4_3326
timestamp 1586364061
transform 1 0 307096 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_3338
timestamp 1586364061
transform 1 0 308200 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_3350
timestamp 1586364061
transform 1 0 309304 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_3362
timestamp 1586364061
transform 1 0 310408 0 -1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_447
timestamp 1586364061
transform 1 0 312616 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_4_3374
timestamp 1586364061
transform 1 0 311512 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_3387
timestamp 1586364061
transform 1 0 312708 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_3399
timestamp 1586364061
transform 1 0 313812 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_3411
timestamp 1586364061
transform 1 0 314916 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_3423
timestamp 1586364061
transform 1 0 316020 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_3435
timestamp 1586364061
transform 1 0 317124 0 -1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_448
timestamp 1586364061
transform 1 0 318228 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_4_3448
timestamp 1586364061
transform 1 0 318320 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_3460
timestamp 1586364061
transform 1 0 319424 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_3472
timestamp 1586364061
transform 1 0 320528 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_3484
timestamp 1586364061
transform 1 0 321632 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_3496
timestamp 1586364061
transform 1 0 322736 0 -1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_449
timestamp 1586364061
transform 1 0 323840 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_4_3509
timestamp 1586364061
transform 1 0 323932 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_3521
timestamp 1586364061
transform 1 0 325036 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_3533
timestamp 1586364061
transform 1 0 326140 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_3545
timestamp 1586364061
transform 1 0 327244 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_3557
timestamp 1586364061
transform 1 0 328348 0 -1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_450
timestamp 1586364061
transform 1 0 329452 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_4_3570
timestamp 1586364061
transform 1 0 329544 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_3582
timestamp 1586364061
transform 1 0 330648 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_3594
timestamp 1586364061
transform 1 0 331752 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_3606
timestamp 1586364061
transform 1 0 332856 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_3618
timestamp 1586364061
transform 1 0 333960 0 -1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_451
timestamp 1586364061
transform 1 0 335064 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_4_3631
timestamp 1586364061
transform 1 0 335156 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_3643
timestamp 1586364061
transform 1 0 336260 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_3655
timestamp 1586364061
transform 1 0 337364 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_3667
timestamp 1586364061
transform 1 0 338468 0 -1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_452
timestamp 1586364061
transform 1 0 340676 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_4_3679
timestamp 1586364061
transform 1 0 339572 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_3692
timestamp 1586364061
transform 1 0 340768 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_3704
timestamp 1586364061
transform 1 0 341872 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_3716
timestamp 1586364061
transform 1 0 342976 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_3728
timestamp 1586364061
transform 1 0 344080 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_3740
timestamp 1586364061
transform 1 0 345184 0 -1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_453
timestamp 1586364061
transform 1 0 346288 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_4_3753
timestamp 1586364061
transform 1 0 346380 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_3765
timestamp 1586364061
transform 1 0 347484 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_3777
timestamp 1586364061
transform 1 0 348588 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_3789
timestamp 1586364061
transform 1 0 349692 0 -1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_454
timestamp 1586364061
transform 1 0 351900 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_4_3801
timestamp 1586364061
transform 1 0 350796 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_3814
timestamp 1586364061
transform 1 0 351992 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_3826
timestamp 1586364061
transform 1 0 353096 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_3838
timestamp 1586364061
transform 1 0 354200 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_3850
timestamp 1586364061
transform 1 0 355304 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_3862
timestamp 1586364061
transform 1 0 356408 0 -1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_455
timestamp 1586364061
transform 1 0 357512 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_4_3875
timestamp 1586364061
transform 1 0 357604 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_3887
timestamp 1586364061
transform 1 0 358708 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_3899
timestamp 1586364061
transform 1 0 359812 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_3911
timestamp 1586364061
transform 1 0 360916 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_3923
timestamp 1586364061
transform 1 0 362020 0 -1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_456
timestamp 1586364061
transform 1 0 363124 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_4_3936
timestamp 1586364061
transform 1 0 363216 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_3948
timestamp 1586364061
transform 1 0 364320 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_3960
timestamp 1586364061
transform 1 0 365424 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_3972
timestamp 1586364061
transform 1 0 366528 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_3984
timestamp 1586364061
transform 1 0 367632 0 -1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_457
timestamp 1586364061
transform 1 0 368736 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_4_3997
timestamp 1586364061
transform 1 0 368828 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_4009
timestamp 1586364061
transform 1 0 369932 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_4021
timestamp 1586364061
transform 1 0 371036 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_4033
timestamp 1586364061
transform 1 0 372140 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_4045
timestamp 1586364061
transform 1 0 373244 0 -1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_458
timestamp 1586364061
transform 1 0 374348 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_4_4058
timestamp 1586364061
transform 1 0 374440 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_4070
timestamp 1586364061
transform 1 0 375544 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_4082
timestamp 1586364061
transform 1 0 376648 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_4094
timestamp 1586364061
transform 1 0 377752 0 -1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_459
timestamp 1586364061
transform 1 0 379960 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_4_4106
timestamp 1586364061
transform 1 0 378856 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_4119
timestamp 1586364061
transform 1 0 380052 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_4131
timestamp 1586364061
transform 1 0 381156 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_4143
timestamp 1586364061
transform 1 0 382260 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_4155
timestamp 1586364061
transform 1 0 383364 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_4167
timestamp 1586364061
transform 1 0 384468 0 -1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_460
timestamp 1586364061
transform 1 0 385572 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_4_4180
timestamp 1586364061
transform 1 0 385664 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_4192
timestamp 1586364061
transform 1 0 386768 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_4204
timestamp 1586364061
transform 1 0 387872 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_4216
timestamp 1586364061
transform 1 0 388976 0 -1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_461
timestamp 1586364061
transform 1 0 391184 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_4_4228
timestamp 1586364061
transform 1 0 390080 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_4241
timestamp 1586364061
transform 1 0 391276 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_4253
timestamp 1586364061
transform 1 0 392380 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_4265
timestamp 1586364061
transform 1 0 393484 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_4277
timestamp 1586364061
transform 1 0 394588 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_4289
timestamp 1586364061
transform 1 0 395692 0 -1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_462
timestamp 1586364061
transform 1 0 396796 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_4_4302
timestamp 1586364061
transform 1 0 396888 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_4314
timestamp 1586364061
transform 1 0 397992 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_4326
timestamp 1586364061
transform 1 0 399096 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_4338
timestamp 1586364061
transform 1 0 400200 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_4350
timestamp 1586364061
transform 1 0 401304 0 -1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_463
timestamp 1586364061
transform 1 0 402408 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_4_4363
timestamp 1586364061
transform 1 0 402500 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_4375
timestamp 1586364061
transform 1 0 403604 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_4387
timestamp 1586364061
transform 1 0 404708 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_4399
timestamp 1586364061
transform 1 0 405812 0 -1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_464
timestamp 1586364061
transform 1 0 408020 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_4_4411
timestamp 1586364061
transform 1 0 406916 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_4424
timestamp 1586364061
transform 1 0 408112 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_4436
timestamp 1586364061
transform 1 0 409216 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_4448
timestamp 1586364061
transform 1 0 410320 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_4460
timestamp 1586364061
transform 1 0 411424 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_4472
timestamp 1586364061
transform 1 0 412528 0 -1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_465
timestamp 1586364061
transform 1 0 413632 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_4_4485
timestamp 1586364061
transform 1 0 413724 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_4497
timestamp 1586364061
transform 1 0 414828 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_4509
timestamp 1586364061
transform 1 0 415932 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_4521
timestamp 1586364061
transform 1 0 417036 0 -1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_466
timestamp 1586364061
transform 1 0 419244 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_4_4533
timestamp 1586364061
transform 1 0 418140 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_4546
timestamp 1586364061
transform 1 0 419336 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_4558
timestamp 1586364061
transform 1 0 420440 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_3  PHY_9
timestamp 1586364061
transform -1 0 422832 0 -1 4896
box -38 -48 314 592
use scs8hd_decap_8  FILLER_4_4570
timestamp 1586364061
transform 1 0 421544 0 -1 4896
box -38 -48 774 592
use scs8hd_decap_3  FILLER_4_4578
timestamp 1586364061
transform 1 0 422280 0 -1 4896
box -38 -48 314 592
use scs8hd_decap_3  PHY_10
timestamp 1586364061
transform 1 0 1104 0 1 4896
box -38 -48 314 592
use scs8hd_decap_12  FILLER_5_3
timestamp 1586364061
transform 1 0 1380 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_15
timestamp 1586364061
transform 1 0 2484 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_27
timestamp 1586364061
transform 1 0 3588 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_39
timestamp 1586364061
transform 1 0 4692 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_5_51
timestamp 1586364061
transform 1 0 5796 0 1 4896
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_467
timestamp 1586364061
transform 1 0 6716 0 1 4896
box -38 -48 130 592
use scs8hd_fill_2  FILLER_5_59
timestamp 1586364061
transform 1 0 6532 0 1 4896
box -38 -48 222 592
use scs8hd_decap_12  FILLER_5_62
timestamp 1586364061
transform 1 0 6808 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_74
timestamp 1586364061
transform 1 0 7912 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_86
timestamp 1586364061
transform 1 0 9016 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_98
timestamp 1586364061
transform 1 0 10120 0 1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_468
timestamp 1586364061
transform 1 0 12328 0 1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_5_110
timestamp 1586364061
transform 1 0 11224 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_123
timestamp 1586364061
transform 1 0 12420 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_135
timestamp 1586364061
transform 1 0 13524 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_147
timestamp 1586364061
transform 1 0 14628 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_159
timestamp 1586364061
transform 1 0 15732 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_171
timestamp 1586364061
transform 1 0 16836 0 1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_469
timestamp 1586364061
transform 1 0 17940 0 1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_5_184
timestamp 1586364061
transform 1 0 18032 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_196
timestamp 1586364061
transform 1 0 19136 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_208
timestamp 1586364061
transform 1 0 20240 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_220
timestamp 1586364061
transform 1 0 21344 0 1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_470
timestamp 1586364061
transform 1 0 23552 0 1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_5_232
timestamp 1586364061
transform 1 0 22448 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_245
timestamp 1586364061
transform 1 0 23644 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_257
timestamp 1586364061
transform 1 0 24748 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_269
timestamp 1586364061
transform 1 0 25852 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_281
timestamp 1586364061
transform 1 0 26956 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_293
timestamp 1586364061
transform 1 0 28060 0 1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_471
timestamp 1586364061
transform 1 0 29164 0 1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_5_306
timestamp 1586364061
transform 1 0 29256 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_318
timestamp 1586364061
transform 1 0 30360 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_330
timestamp 1586364061
transform 1 0 31464 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_342
timestamp 1586364061
transform 1 0 32568 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_354
timestamp 1586364061
transform 1 0 33672 0 1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_472
timestamp 1586364061
transform 1 0 34776 0 1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_5_367
timestamp 1586364061
transform 1 0 34868 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_379
timestamp 1586364061
transform 1 0 35972 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_391
timestamp 1586364061
transform 1 0 37076 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_403
timestamp 1586364061
transform 1 0 38180 0 1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_473
timestamp 1586364061
transform 1 0 40388 0 1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_5_415
timestamp 1586364061
transform 1 0 39284 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_428
timestamp 1586364061
transform 1 0 40480 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_440
timestamp 1586364061
transform 1 0 41584 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_452
timestamp 1586364061
transform 1 0 42688 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_464
timestamp 1586364061
transform 1 0 43792 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_476
timestamp 1586364061
transform 1 0 44896 0 1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_474
timestamp 1586364061
transform 1 0 46000 0 1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_5_489
timestamp 1586364061
transform 1 0 46092 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_501
timestamp 1586364061
transform 1 0 47196 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_513
timestamp 1586364061
transform 1 0 48300 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_525
timestamp 1586364061
transform 1 0 49404 0 1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_475
timestamp 1586364061
transform 1 0 51612 0 1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_5_537
timestamp 1586364061
transform 1 0 50508 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_550
timestamp 1586364061
transform 1 0 51704 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_562
timestamp 1586364061
transform 1 0 52808 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_574
timestamp 1586364061
transform 1 0 53912 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_586
timestamp 1586364061
transform 1 0 55016 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_598
timestamp 1586364061
transform 1 0 56120 0 1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_476
timestamp 1586364061
transform 1 0 57224 0 1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_5_611
timestamp 1586364061
transform 1 0 57316 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_623
timestamp 1586364061
transform 1 0 58420 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_635
timestamp 1586364061
transform 1 0 59524 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_647
timestamp 1586364061
transform 1 0 60628 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_659
timestamp 1586364061
transform 1 0 61732 0 1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_477
timestamp 1586364061
transform 1 0 62836 0 1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_5_672
timestamp 1586364061
transform 1 0 62928 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_684
timestamp 1586364061
transform 1 0 64032 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_696
timestamp 1586364061
transform 1 0 65136 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_708
timestamp 1586364061
transform 1 0 66240 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_720
timestamp 1586364061
transform 1 0 67344 0 1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_478
timestamp 1586364061
transform 1 0 68448 0 1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_5_733
timestamp 1586364061
transform 1 0 68540 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_745
timestamp 1586364061
transform 1 0 69644 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_757
timestamp 1586364061
transform 1 0 70748 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_769
timestamp 1586364061
transform 1 0 71852 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_781
timestamp 1586364061
transform 1 0 72956 0 1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_479
timestamp 1586364061
transform 1 0 74060 0 1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_5_794
timestamp 1586364061
transform 1 0 74152 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_806
timestamp 1586364061
transform 1 0 75256 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_818
timestamp 1586364061
transform 1 0 76360 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_830
timestamp 1586364061
transform 1 0 77464 0 1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_480
timestamp 1586364061
transform 1 0 79672 0 1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_5_842
timestamp 1586364061
transform 1 0 78568 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_855
timestamp 1586364061
transform 1 0 79764 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_867
timestamp 1586364061
transform 1 0 80868 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_879
timestamp 1586364061
transform 1 0 81972 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_891
timestamp 1586364061
transform 1 0 83076 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_903
timestamp 1586364061
transform 1 0 84180 0 1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_481
timestamp 1586364061
transform 1 0 85284 0 1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_5_916
timestamp 1586364061
transform 1 0 85376 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_928
timestamp 1586364061
transform 1 0 86480 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_940
timestamp 1586364061
transform 1 0 87584 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_952
timestamp 1586364061
transform 1 0 88688 0 1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_482
timestamp 1586364061
transform 1 0 90896 0 1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_5_964
timestamp 1586364061
transform 1 0 89792 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_977
timestamp 1586364061
transform 1 0 90988 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_5_989
timestamp 1586364061
transform 1 0 92092 0 1 4896
box -38 -48 774 592
use scs8hd_decap_3  FILLER_5_997
timestamp 1586364061
transform 1 0 92828 0 1 4896
box -38 -48 314 592
use scs8hd_buf_2  _16_
timestamp 1586364061
transform 1 0 93104 0 1 4896
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__16__A
timestamp 1586364061
transform 1 0 93656 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_1004
timestamp 1586364061
transform 1 0 93472 0 1 4896
box -38 -48 222 592
use scs8hd_decap_12  FILLER_5_1008
timestamp 1586364061
transform 1 0 93840 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_1020
timestamp 1586364061
transform 1 0 94944 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_5_1032
timestamp 1586364061
transform 1 0 96048 0 1 4896
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_483
timestamp 1586364061
transform 1 0 96508 0 1 4896
box -38 -48 130 592
use scs8hd_fill_1  FILLER_5_1036
timestamp 1586364061
transform 1 0 96416 0 1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_5_1038
timestamp 1586364061
transform 1 0 96600 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_1050
timestamp 1586364061
transform 1 0 97704 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_1062
timestamp 1586364061
transform 1 0 98808 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_1074
timestamp 1586364061
transform 1 0 99912 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_1086
timestamp 1586364061
transform 1 0 101016 0 1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_484
timestamp 1586364061
transform 1 0 102120 0 1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_5_1099
timestamp 1586364061
transform 1 0 102212 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_1111
timestamp 1586364061
transform 1 0 103316 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_1123
timestamp 1586364061
transform 1 0 104420 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_1135
timestamp 1586364061
transform 1 0 105524 0 1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_485
timestamp 1586364061
transform 1 0 107732 0 1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_5_1147
timestamp 1586364061
transform 1 0 106628 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_1160
timestamp 1586364061
transform 1 0 107824 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_1172
timestamp 1586364061
transform 1 0 108928 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_1184
timestamp 1586364061
transform 1 0 110032 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_1196
timestamp 1586364061
transform 1 0 111136 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_1208
timestamp 1586364061
transform 1 0 112240 0 1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_486
timestamp 1586364061
transform 1 0 113344 0 1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_5_1221
timestamp 1586364061
transform 1 0 113436 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_1233
timestamp 1586364061
transform 1 0 114540 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_1245
timestamp 1586364061
transform 1 0 115644 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_1257
timestamp 1586364061
transform 1 0 116748 0 1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_487
timestamp 1586364061
transform 1 0 118956 0 1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_5_1269
timestamp 1586364061
transform 1 0 117852 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_1282
timestamp 1586364061
transform 1 0 119048 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_1294
timestamp 1586364061
transform 1 0 120152 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_1306
timestamp 1586364061
transform 1 0 121256 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_1318
timestamp 1586364061
transform 1 0 122360 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_1330
timestamp 1586364061
transform 1 0 123464 0 1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_488
timestamp 1586364061
transform 1 0 124568 0 1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_5_1343
timestamp 1586364061
transform 1 0 124660 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_1355
timestamp 1586364061
transform 1 0 125764 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_1367
timestamp 1586364061
transform 1 0 126868 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_1379
timestamp 1586364061
transform 1 0 127972 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_1391
timestamp 1586364061
transform 1 0 129076 0 1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_489
timestamp 1586364061
transform 1 0 130180 0 1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_5_1404
timestamp 1586364061
transform 1 0 130272 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_1416
timestamp 1586364061
transform 1 0 131376 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_1428
timestamp 1586364061
transform 1 0 132480 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_1440
timestamp 1586364061
transform 1 0 133584 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_1452
timestamp 1586364061
transform 1 0 134688 0 1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_490
timestamp 1586364061
transform 1 0 135792 0 1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_5_1465
timestamp 1586364061
transform 1 0 135884 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_1477
timestamp 1586364061
transform 1 0 136988 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_1489
timestamp 1586364061
transform 1 0 138092 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_1501
timestamp 1586364061
transform 1 0 139196 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_1513
timestamp 1586364061
transform 1 0 140300 0 1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_491
timestamp 1586364061
transform 1 0 141404 0 1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_5_1526
timestamp 1586364061
transform 1 0 141496 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_1538
timestamp 1586364061
transform 1 0 142600 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_1550
timestamp 1586364061
transform 1 0 143704 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_1562
timestamp 1586364061
transform 1 0 144808 0 1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_492
timestamp 1586364061
transform 1 0 147016 0 1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_5_1574
timestamp 1586364061
transform 1 0 145912 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_1587
timestamp 1586364061
transform 1 0 147108 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_1599
timestamp 1586364061
transform 1 0 148212 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_1611
timestamp 1586364061
transform 1 0 149316 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_1623
timestamp 1586364061
transform 1 0 150420 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_1635
timestamp 1586364061
transform 1 0 151524 0 1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_493
timestamp 1586364061
transform 1 0 152628 0 1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_5_1648
timestamp 1586364061
transform 1 0 152720 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_1660
timestamp 1586364061
transform 1 0 153824 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_1672
timestamp 1586364061
transform 1 0 154928 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_1684
timestamp 1586364061
transform 1 0 156032 0 1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_494
timestamp 1586364061
transform 1 0 158240 0 1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_5_1696
timestamp 1586364061
transform 1 0 157136 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_1709
timestamp 1586364061
transform 1 0 158332 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_1721
timestamp 1586364061
transform 1 0 159436 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_1733
timestamp 1586364061
transform 1 0 160540 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_1745
timestamp 1586364061
transform 1 0 161644 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_1757
timestamp 1586364061
transform 1 0 162748 0 1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_495
timestamp 1586364061
transform 1 0 163852 0 1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_5_1770
timestamp 1586364061
transform 1 0 163944 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_1782
timestamp 1586364061
transform 1 0 165048 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_1794
timestamp 1586364061
transform 1 0 166152 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_1806
timestamp 1586364061
transform 1 0 167256 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_1818
timestamp 1586364061
transform 1 0 168360 0 1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_496
timestamp 1586364061
transform 1 0 169464 0 1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_5_1831
timestamp 1586364061
transform 1 0 169556 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_1843
timestamp 1586364061
transform 1 0 170660 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_1855
timestamp 1586364061
transform 1 0 171764 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_1867
timestamp 1586364061
transform 1 0 172868 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_1879
timestamp 1586364061
transform 1 0 173972 0 1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_497
timestamp 1586364061
transform 1 0 175076 0 1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_5_1892
timestamp 1586364061
transform 1 0 175168 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_1904
timestamp 1586364061
transform 1 0 176272 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_1916
timestamp 1586364061
transform 1 0 177376 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_1928
timestamp 1586364061
transform 1 0 178480 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_1940
timestamp 1586364061
transform 1 0 179584 0 1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_498
timestamp 1586364061
transform 1 0 180688 0 1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_5_1953
timestamp 1586364061
transform 1 0 180780 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_1965
timestamp 1586364061
transform 1 0 181884 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_1977
timestamp 1586364061
transform 1 0 182988 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_1989
timestamp 1586364061
transform 1 0 184092 0 1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_499
timestamp 1586364061
transform 1 0 186300 0 1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_5_2001
timestamp 1586364061
transform 1 0 185196 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_2014
timestamp 1586364061
transform 1 0 186392 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_2026
timestamp 1586364061
transform 1 0 187496 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_2038
timestamp 1586364061
transform 1 0 188600 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_2050
timestamp 1586364061
transform 1 0 189704 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_2062
timestamp 1586364061
transform 1 0 190808 0 1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_500
timestamp 1586364061
transform 1 0 191912 0 1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_5_2075
timestamp 1586364061
transform 1 0 192004 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_2087
timestamp 1586364061
transform 1 0 193108 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_2099
timestamp 1586364061
transform 1 0 194212 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_2111
timestamp 1586364061
transform 1 0 195316 0 1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_501
timestamp 1586364061
transform 1 0 197524 0 1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_5_2123
timestamp 1586364061
transform 1 0 196420 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_2136
timestamp 1586364061
transform 1 0 197616 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_2148
timestamp 1586364061
transform 1 0 198720 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_2160
timestamp 1586364061
transform 1 0 199824 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_2172
timestamp 1586364061
transform 1 0 200928 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_2184
timestamp 1586364061
transform 1 0 202032 0 1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_502
timestamp 1586364061
transform 1 0 203136 0 1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_5_2197
timestamp 1586364061
transform 1 0 203228 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_2209
timestamp 1586364061
transform 1 0 204332 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_2221
timestamp 1586364061
transform 1 0 205436 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_2233
timestamp 1586364061
transform 1 0 206540 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_5_2245
timestamp 1586364061
transform 1 0 207644 0 1 4896
box -38 -48 774 592
use scs8hd_ebufn_1  logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer
timestamp 1586364061
transform 1 0 208840 0 1 4896
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_503
timestamp 1586364061
transform 1 0 208748 0 1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer_A
timestamp 1586364061
transform 1 0 208564 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_2253
timestamp 1586364061
transform 1 0 208380 0 1 4896
box -38 -48 222 592
use scs8hd_decap_12  FILLER_5_2266
timestamp 1586364061
transform 1 0 209576 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_2278
timestamp 1586364061
transform 1 0 210680 0 1 4896
box -38 -48 1142 592
use scs8hd_lpflow_inputisolatch_1  logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.LATCH_0_.latch
timestamp 1586364061
transform 1 0 212244 0 1 4896
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 212060 0 1 4896
box -38 -48 222 592
use scs8hd_decap_3  FILLER_5_2290
timestamp 1586364061
transform 1 0 211784 0 1 4896
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_504
timestamp 1586364061
transform 1 0 214360 0 1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 214176 0 1 4896
box -38 -48 222 592
use scs8hd_decap_8  FILLER_5_2306
timestamp 1586364061
transform 1 0 213256 0 1 4896
box -38 -48 774 592
use scs8hd_fill_2  FILLER_5_2314
timestamp 1586364061
transform 1 0 213992 0 1 4896
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.LATCH_0_.latch
timestamp 1586364061
transform 1 0 215004 0 1 4896
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 214820 0 1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_5_2319
timestamp 1586364061
transform 1 0 214452 0 1 4896
box -38 -48 406 592
use scs8hd_fill_2  FILLER_5_2336
timestamp 1586364061
transform 1 0 216016 0 1 4896
box -38 -48 222 592
use scs8hd_and4_4  _10_
timestamp 1586364061
transform 1 0 216752 0 1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__10__C
timestamp 1586364061
transform 1 0 216568 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__10__D
timestamp 1586364061
transform 1 0 216200 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_2340
timestamp 1586364061
transform 1 0 216384 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_2353
timestamp 1586364061
transform 1 0 217580 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer_A
timestamp 1586364061
transform 1 0 217764 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer_TEB
timestamp 1586364061
transform 1 0 218132 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_2357
timestamp 1586364061
transform 1 0 217948 0 1 4896
box -38 -48 222 592
use scs8hd_decap_12  FILLER_5_2361
timestamp 1586364061
transform 1 0 218316 0 1 4896
box -38 -48 1142 592
use scs8hd_lpflow_inputisolatch_1  logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.LATCH_0_.latch
timestamp 1586364061
transform 1 0 220524 0 1 4896
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_505
timestamp 1586364061
transform 1 0 219972 0 1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 220340 0 1 4896
box -38 -48 222 592
use scs8hd_decap_6  FILLER_5_2373
timestamp 1586364061
transform 1 0 219420 0 1 4896
box -38 -48 590 592
use scs8hd_decap_3  FILLER_5_2380
timestamp 1586364061
transform 1 0 220064 0 1 4896
box -38 -48 314 592
use scs8hd_decap_12  FILLER_5_2396
timestamp 1586364061
transform 1 0 221536 0 1 4896
box -38 -48 1142 592
use scs8hd_ebufn_1  logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer
timestamp 1586364061
transform 1 0 224020 0 1 4896
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA_logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer_A
timestamp 1586364061
transform 1 0 223836 0 1 4896
box -38 -48 222 592
use scs8hd_decap_12  FILLER_5_2408
timestamp 1586364061
transform 1 0 222640 0 1 4896
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_5_2420
timestamp 1586364061
transform 1 0 223744 0 1 4896
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_506
timestamp 1586364061
transform 1 0 225584 0 1 4896
box -38 -48 130 592
use scs8hd_decap_8  FILLER_5_2431
timestamp 1586364061
transform 1 0 224756 0 1 4896
box -38 -48 774 592
use scs8hd_fill_1  FILLER_5_2439
timestamp 1586364061
transform 1 0 225492 0 1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_5_2441
timestamp 1586364061
transform 1 0 225676 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_2453
timestamp 1586364061
transform 1 0 226780 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_2465
timestamp 1586364061
transform 1 0 227884 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_2477
timestamp 1586364061
transform 1 0 228988 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_2489
timestamp 1586364061
transform 1 0 230092 0 1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_507
timestamp 1586364061
transform 1 0 231196 0 1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_5_2502
timestamp 1586364061
transform 1 0 231288 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_2514
timestamp 1586364061
transform 1 0 232392 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_2526
timestamp 1586364061
transform 1 0 233496 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_2538
timestamp 1586364061
transform 1 0 234600 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_2550
timestamp 1586364061
transform 1 0 235704 0 1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_508
timestamp 1586364061
transform 1 0 236808 0 1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_5_2563
timestamp 1586364061
transform 1 0 236900 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_2575
timestamp 1586364061
transform 1 0 238004 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_2587
timestamp 1586364061
transform 1 0 239108 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_2599
timestamp 1586364061
transform 1 0 240212 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_2611
timestamp 1586364061
transform 1 0 241316 0 1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_509
timestamp 1586364061
transform 1 0 242420 0 1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_5_2624
timestamp 1586364061
transform 1 0 242512 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_2636
timestamp 1586364061
transform 1 0 243616 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_2648
timestamp 1586364061
transform 1 0 244720 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_2660
timestamp 1586364061
transform 1 0 245824 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_2672
timestamp 1586364061
transform 1 0 246928 0 1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_510
timestamp 1586364061
transform 1 0 248032 0 1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_5_2685
timestamp 1586364061
transform 1 0 248124 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_2697
timestamp 1586364061
transform 1 0 249228 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_2709
timestamp 1586364061
transform 1 0 250332 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_2721
timestamp 1586364061
transform 1 0 251436 0 1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_511
timestamp 1586364061
transform 1 0 253644 0 1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_5_2733
timestamp 1586364061
transform 1 0 252540 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_2746
timestamp 1586364061
transform 1 0 253736 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_2758
timestamp 1586364061
transform 1 0 254840 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_2770
timestamp 1586364061
transform 1 0 255944 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_2782
timestamp 1586364061
transform 1 0 257048 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_2794
timestamp 1586364061
transform 1 0 258152 0 1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_512
timestamp 1586364061
transform 1 0 259256 0 1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_5_2807
timestamp 1586364061
transform 1 0 259348 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_2819
timestamp 1586364061
transform 1 0 260452 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_2831
timestamp 1586364061
transform 1 0 261556 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_2843
timestamp 1586364061
transform 1 0 262660 0 1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_513
timestamp 1586364061
transform 1 0 264868 0 1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_5_2855
timestamp 1586364061
transform 1 0 263764 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_2868
timestamp 1586364061
transform 1 0 264960 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_2880
timestamp 1586364061
transform 1 0 266064 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_2892
timestamp 1586364061
transform 1 0 267168 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_2904
timestamp 1586364061
transform 1 0 268272 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_2916
timestamp 1586364061
transform 1 0 269376 0 1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_514
timestamp 1586364061
transform 1 0 270480 0 1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_5_2929
timestamp 1586364061
transform 1 0 270572 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_2941
timestamp 1586364061
transform 1 0 271676 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_2953
timestamp 1586364061
transform 1 0 272780 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_2965
timestamp 1586364061
transform 1 0 273884 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_2977
timestamp 1586364061
transform 1 0 274988 0 1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_515
timestamp 1586364061
transform 1 0 276092 0 1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_5_2990
timestamp 1586364061
transform 1 0 276184 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_3002
timestamp 1586364061
transform 1 0 277288 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_3014
timestamp 1586364061
transform 1 0 278392 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_3026
timestamp 1586364061
transform 1 0 279496 0 1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_516
timestamp 1586364061
transform 1 0 281704 0 1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_5_3038
timestamp 1586364061
transform 1 0 280600 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_3051
timestamp 1586364061
transform 1 0 281796 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_3063
timestamp 1586364061
transform 1 0 282900 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_3075
timestamp 1586364061
transform 1 0 284004 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_3087
timestamp 1586364061
transform 1 0 285108 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_3099
timestamp 1586364061
transform 1 0 286212 0 1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_517
timestamp 1586364061
transform 1 0 287316 0 1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_5_3112
timestamp 1586364061
transform 1 0 287408 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_3124
timestamp 1586364061
transform 1 0 288512 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_3136
timestamp 1586364061
transform 1 0 289616 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_3148
timestamp 1586364061
transform 1 0 290720 0 1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_518
timestamp 1586364061
transform 1 0 292928 0 1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_5_3160
timestamp 1586364061
transform 1 0 291824 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_3173
timestamp 1586364061
transform 1 0 293020 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_3185
timestamp 1586364061
transform 1 0 294124 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_3197
timestamp 1586364061
transform 1 0 295228 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_3209
timestamp 1586364061
transform 1 0 296332 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_3221
timestamp 1586364061
transform 1 0 297436 0 1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_519
timestamp 1586364061
transform 1 0 298540 0 1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_5_3234
timestamp 1586364061
transform 1 0 298632 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_3246
timestamp 1586364061
transform 1 0 299736 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_3258
timestamp 1586364061
transform 1 0 300840 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_3270
timestamp 1586364061
transform 1 0 301944 0 1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_520
timestamp 1586364061
transform 1 0 304152 0 1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_5_3282
timestamp 1586364061
transform 1 0 303048 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_3295
timestamp 1586364061
transform 1 0 304244 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_3307
timestamp 1586364061
transform 1 0 305348 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_3319
timestamp 1586364061
transform 1 0 306452 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_3331
timestamp 1586364061
transform 1 0 307556 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_3343
timestamp 1586364061
transform 1 0 308660 0 1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_521
timestamp 1586364061
transform 1 0 309764 0 1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_5_3356
timestamp 1586364061
transform 1 0 309856 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_3368
timestamp 1586364061
transform 1 0 310960 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_3380
timestamp 1586364061
transform 1 0 312064 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_3392
timestamp 1586364061
transform 1 0 313168 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_3404
timestamp 1586364061
transform 1 0 314272 0 1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_522
timestamp 1586364061
transform 1 0 315376 0 1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_5_3417
timestamp 1586364061
transform 1 0 315468 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_3429
timestamp 1586364061
transform 1 0 316572 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_3441
timestamp 1586364061
transform 1 0 317676 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_3453
timestamp 1586364061
transform 1 0 318780 0 1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_523
timestamp 1586364061
transform 1 0 320988 0 1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_5_3465
timestamp 1586364061
transform 1 0 319884 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_3478
timestamp 1586364061
transform 1 0 321080 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_3490
timestamp 1586364061
transform 1 0 322184 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_3502
timestamp 1586364061
transform 1 0 323288 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_3514
timestamp 1586364061
transform 1 0 324392 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_3526
timestamp 1586364061
transform 1 0 325496 0 1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_524
timestamp 1586364061
transform 1 0 326600 0 1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_5_3539
timestamp 1586364061
transform 1 0 326692 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_3551
timestamp 1586364061
transform 1 0 327796 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_3563
timestamp 1586364061
transform 1 0 328900 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_3575
timestamp 1586364061
transform 1 0 330004 0 1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_525
timestamp 1586364061
transform 1 0 332212 0 1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_5_3587
timestamp 1586364061
transform 1 0 331108 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_3600
timestamp 1586364061
transform 1 0 332304 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_3612
timestamp 1586364061
transform 1 0 333408 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_3624
timestamp 1586364061
transform 1 0 334512 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_3636
timestamp 1586364061
transform 1 0 335616 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_3648
timestamp 1586364061
transform 1 0 336720 0 1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_526
timestamp 1586364061
transform 1 0 337824 0 1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_5_3661
timestamp 1586364061
transform 1 0 337916 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_3673
timestamp 1586364061
transform 1 0 339020 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_3685
timestamp 1586364061
transform 1 0 340124 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_3697
timestamp 1586364061
transform 1 0 341228 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_3709
timestamp 1586364061
transform 1 0 342332 0 1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_527
timestamp 1586364061
transform 1 0 343436 0 1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_5_3722
timestamp 1586364061
transform 1 0 343528 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_3734
timestamp 1586364061
transform 1 0 344632 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_3746
timestamp 1586364061
transform 1 0 345736 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_3758
timestamp 1586364061
transform 1 0 346840 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_3770
timestamp 1586364061
transform 1 0 347944 0 1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_528
timestamp 1586364061
transform 1 0 349048 0 1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_5_3783
timestamp 1586364061
transform 1 0 349140 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_3795
timestamp 1586364061
transform 1 0 350244 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_3807
timestamp 1586364061
transform 1 0 351348 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_3819
timestamp 1586364061
transform 1 0 352452 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_3831
timestamp 1586364061
transform 1 0 353556 0 1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_529
timestamp 1586364061
transform 1 0 354660 0 1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_5_3844
timestamp 1586364061
transform 1 0 354752 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_3856
timestamp 1586364061
transform 1 0 355856 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_3868
timestamp 1586364061
transform 1 0 356960 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_3880
timestamp 1586364061
transform 1 0 358064 0 1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_530
timestamp 1586364061
transform 1 0 360272 0 1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_5_3892
timestamp 1586364061
transform 1 0 359168 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_3905
timestamp 1586364061
transform 1 0 360364 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_3917
timestamp 1586364061
transform 1 0 361468 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_3929
timestamp 1586364061
transform 1 0 362572 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_3941
timestamp 1586364061
transform 1 0 363676 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_3953
timestamp 1586364061
transform 1 0 364780 0 1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_531
timestamp 1586364061
transform 1 0 365884 0 1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_5_3966
timestamp 1586364061
transform 1 0 365976 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_3978
timestamp 1586364061
transform 1 0 367080 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_3990
timestamp 1586364061
transform 1 0 368184 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_4002
timestamp 1586364061
transform 1 0 369288 0 1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_532
timestamp 1586364061
transform 1 0 371496 0 1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_5_4014
timestamp 1586364061
transform 1 0 370392 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_4027
timestamp 1586364061
transform 1 0 371588 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_4039
timestamp 1586364061
transform 1 0 372692 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_4051
timestamp 1586364061
transform 1 0 373796 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_4063
timestamp 1586364061
transform 1 0 374900 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_4075
timestamp 1586364061
transform 1 0 376004 0 1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_533
timestamp 1586364061
transform 1 0 377108 0 1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_5_4088
timestamp 1586364061
transform 1 0 377200 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_4100
timestamp 1586364061
transform 1 0 378304 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_4112
timestamp 1586364061
transform 1 0 379408 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_4124
timestamp 1586364061
transform 1 0 380512 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_4136
timestamp 1586364061
transform 1 0 381616 0 1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_534
timestamp 1586364061
transform 1 0 382720 0 1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_5_4149
timestamp 1586364061
transform 1 0 382812 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_4161
timestamp 1586364061
transform 1 0 383916 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_4173
timestamp 1586364061
transform 1 0 385020 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_4185
timestamp 1586364061
transform 1 0 386124 0 1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_535
timestamp 1586364061
transform 1 0 388332 0 1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_5_4197
timestamp 1586364061
transform 1 0 387228 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_4210
timestamp 1586364061
transform 1 0 388424 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_4222
timestamp 1586364061
transform 1 0 389528 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_4234
timestamp 1586364061
transform 1 0 390632 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_4246
timestamp 1586364061
transform 1 0 391736 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_4258
timestamp 1586364061
transform 1 0 392840 0 1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_536
timestamp 1586364061
transform 1 0 393944 0 1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_5_4271
timestamp 1586364061
transform 1 0 394036 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_4283
timestamp 1586364061
transform 1 0 395140 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_4295
timestamp 1586364061
transform 1 0 396244 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_4307
timestamp 1586364061
transform 1 0 397348 0 1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_537
timestamp 1586364061
transform 1 0 399556 0 1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_5_4319
timestamp 1586364061
transform 1 0 398452 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_4332
timestamp 1586364061
transform 1 0 399648 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_4344
timestamp 1586364061
transform 1 0 400752 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_4356
timestamp 1586364061
transform 1 0 401856 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_4368
timestamp 1586364061
transform 1 0 402960 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_4380
timestamp 1586364061
transform 1 0 404064 0 1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_538
timestamp 1586364061
transform 1 0 405168 0 1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_5_4393
timestamp 1586364061
transform 1 0 405260 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_4405
timestamp 1586364061
transform 1 0 406364 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_4417
timestamp 1586364061
transform 1 0 407468 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_4429
timestamp 1586364061
transform 1 0 408572 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_4441
timestamp 1586364061
transform 1 0 409676 0 1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_539
timestamp 1586364061
transform 1 0 410780 0 1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_5_4454
timestamp 1586364061
transform 1 0 410872 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_4466
timestamp 1586364061
transform 1 0 411976 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_4478
timestamp 1586364061
transform 1 0 413080 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_4490
timestamp 1586364061
transform 1 0 414184 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_4502
timestamp 1586364061
transform 1 0 415288 0 1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_540
timestamp 1586364061
transform 1 0 416392 0 1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_5_4515
timestamp 1586364061
transform 1 0 416484 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_4527
timestamp 1586364061
transform 1 0 417588 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_4539
timestamp 1586364061
transform 1 0 418692 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_4551
timestamp 1586364061
transform 1 0 419796 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_4563
timestamp 1586364061
transform 1 0 420900 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_3  PHY_11
timestamp 1586364061
transform -1 0 422832 0 1 4896
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_541
timestamp 1586364061
transform 1 0 422004 0 1 4896
box -38 -48 130 592
use scs8hd_decap_4  FILLER_5_4576
timestamp 1586364061
transform 1 0 422096 0 1 4896
box -38 -48 406 592
use scs8hd_fill_1  FILLER_5_4580
timestamp 1586364061
transform 1 0 422464 0 1 4896
box -38 -48 130 592
use scs8hd_decap_3  PHY_12
timestamp 1586364061
transform 1 0 1104 0 -1 5984
box -38 -48 314 592
use scs8hd_decap_3  PHY_14
timestamp 1586364061
transform 1 0 1104 0 1 5984
box -38 -48 314 592
use scs8hd_decap_12  FILLER_6_3
timestamp 1586364061
transform 1 0 1380 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_15
timestamp 1586364061
transform 1 0 2484 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_3
timestamp 1586364061
transform 1 0 1380 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_15
timestamp 1586364061
transform 1 0 2484 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_542
timestamp 1586364061
transform 1 0 3956 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_4  FILLER_6_27
timestamp 1586364061
transform 1 0 3588 0 -1 5984
box -38 -48 406 592
use scs8hd_decap_12  FILLER_6_32
timestamp 1586364061
transform 1 0 4048 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_27
timestamp 1586364061
transform 1 0 3588 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_44
timestamp 1586364061
transform 1 0 5152 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_39
timestamp 1586364061
transform 1 0 4692 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_7_51
timestamp 1586364061
transform 1 0 5796 0 1 5984
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_617
timestamp 1586364061
transform 1 0 6716 0 1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_56
timestamp 1586364061
transform 1 0 6256 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_68
timestamp 1586364061
transform 1 0 7360 0 -1 5984
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_7_59
timestamp 1586364061
transform 1 0 6532 0 1 5984
box -38 -48 222 592
use scs8hd_decap_12  FILLER_7_62
timestamp 1586364061
transform 1 0 6808 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_80
timestamp 1586364061
transform 1 0 8464 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_74
timestamp 1586364061
transform 1 0 7912 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_86
timestamp 1586364061
transform 1 0 9016 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_543
timestamp 1586364061
transform 1 0 9568 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_93
timestamp 1586364061
transform 1 0 9660 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_105
timestamp 1586364061
transform 1 0 10764 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_98
timestamp 1586364061
transform 1 0 10120 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_618
timestamp 1586364061
transform 1 0 12328 0 1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_117
timestamp 1586364061
transform 1 0 11868 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_110
timestamp 1586364061
transform 1 0 11224 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_123
timestamp 1586364061
transform 1 0 12420 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_129
timestamp 1586364061
transform 1 0 12972 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_141
timestamp 1586364061
transform 1 0 14076 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_135
timestamp 1586364061
transform 1 0 13524 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_544
timestamp 1586364061
transform 1 0 15180 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_154
timestamp 1586364061
transform 1 0 15272 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_147
timestamp 1586364061
transform 1 0 14628 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_159
timestamp 1586364061
transform 1 0 15732 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_166
timestamp 1586364061
transform 1 0 16376 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_178
timestamp 1586364061
transform 1 0 17480 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_171
timestamp 1586364061
transform 1 0 16836 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_619
timestamp 1586364061
transform 1 0 17940 0 1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_190
timestamp 1586364061
transform 1 0 18584 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_184
timestamp 1586364061
transform 1 0 18032 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_196
timestamp 1586364061
transform 1 0 19136 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_545
timestamp 1586364061
transform 1 0 20792 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_202
timestamp 1586364061
transform 1 0 19688 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_208
timestamp 1586364061
transform 1 0 20240 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_215
timestamp 1586364061
transform 1 0 20884 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_227
timestamp 1586364061
transform 1 0 21988 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_220
timestamp 1586364061
transform 1 0 21344 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_620
timestamp 1586364061
transform 1 0 23552 0 1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_239
timestamp 1586364061
transform 1 0 23092 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_232
timestamp 1586364061
transform 1 0 22448 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_245
timestamp 1586364061
transform 1 0 23644 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_251
timestamp 1586364061
transform 1 0 24196 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_263
timestamp 1586364061
transform 1 0 25300 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_257
timestamp 1586364061
transform 1 0 24748 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_546
timestamp 1586364061
transform 1 0 26404 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_276
timestamp 1586364061
transform 1 0 26496 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_269
timestamp 1586364061
transform 1 0 25852 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_281
timestamp 1586364061
transform 1 0 26956 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_288
timestamp 1586364061
transform 1 0 27600 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_300
timestamp 1586364061
transform 1 0 28704 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_293
timestamp 1586364061
transform 1 0 28060 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_621
timestamp 1586364061
transform 1 0 29164 0 1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_312
timestamp 1586364061
transform 1 0 29808 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_306
timestamp 1586364061
transform 1 0 29256 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_318
timestamp 1586364061
transform 1 0 30360 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_547
timestamp 1586364061
transform 1 0 32016 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_324
timestamp 1586364061
transform 1 0 30912 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_337
timestamp 1586364061
transform 1 0 32108 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_330
timestamp 1586364061
transform 1 0 31464 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_349
timestamp 1586364061
transform 1 0 33212 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_342
timestamp 1586364061
transform 1 0 32568 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_354
timestamp 1586364061
transform 1 0 33672 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_622
timestamp 1586364061
transform 1 0 34776 0 1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_361
timestamp 1586364061
transform 1 0 34316 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_373
timestamp 1586364061
transform 1 0 35420 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_367
timestamp 1586364061
transform 1 0 34868 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_385
timestamp 1586364061
transform 1 0 36524 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_379
timestamp 1586364061
transform 1 0 35972 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_391
timestamp 1586364061
transform 1 0 37076 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_548
timestamp 1586364061
transform 1 0 37628 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_398
timestamp 1586364061
transform 1 0 37720 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_410
timestamp 1586364061
transform 1 0 38824 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_403
timestamp 1586364061
transform 1 0 38180 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_623
timestamp 1586364061
transform 1 0 40388 0 1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_422
timestamp 1586364061
transform 1 0 39928 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_415
timestamp 1586364061
transform 1 0 39284 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_428
timestamp 1586364061
transform 1 0 40480 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_434
timestamp 1586364061
transform 1 0 41032 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_440
timestamp 1586364061
transform 1 0 41584 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_549
timestamp 1586364061
transform 1 0 43240 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_446
timestamp 1586364061
transform 1 0 42136 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_459
timestamp 1586364061
transform 1 0 43332 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_452
timestamp 1586364061
transform 1 0 42688 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_471
timestamp 1586364061
transform 1 0 44436 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_464
timestamp 1586364061
transform 1 0 43792 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_476
timestamp 1586364061
transform 1 0 44896 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_624
timestamp 1586364061
transform 1 0 46000 0 1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_483
timestamp 1586364061
transform 1 0 45540 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_495
timestamp 1586364061
transform 1 0 46644 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_489
timestamp 1586364061
transform 1 0 46092 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_507
timestamp 1586364061
transform 1 0 47748 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_501
timestamp 1586364061
transform 1 0 47196 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_513
timestamp 1586364061
transform 1 0 48300 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_550
timestamp 1586364061
transform 1 0 48852 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_520
timestamp 1586364061
transform 1 0 48944 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_532
timestamp 1586364061
transform 1 0 50048 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_525
timestamp 1586364061
transform 1 0 49404 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_625
timestamp 1586364061
transform 1 0 51612 0 1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_544
timestamp 1586364061
transform 1 0 51152 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_537
timestamp 1586364061
transform 1 0 50508 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_550
timestamp 1586364061
transform 1 0 51704 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_556
timestamp 1586364061
transform 1 0 52256 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_568
timestamp 1586364061
transform 1 0 53360 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_562
timestamp 1586364061
transform 1 0 52808 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_551
timestamp 1586364061
transform 1 0 54464 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_581
timestamp 1586364061
transform 1 0 54556 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_574
timestamp 1586364061
transform 1 0 53912 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_586
timestamp 1586364061
transform 1 0 55016 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_593
timestamp 1586364061
transform 1 0 55660 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_605
timestamp 1586364061
transform 1 0 56764 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_598
timestamp 1586364061
transform 1 0 56120 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_626
timestamp 1586364061
transform 1 0 57224 0 1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_617
timestamp 1586364061
transform 1 0 57868 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_611
timestamp 1586364061
transform 1 0 57316 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_623
timestamp 1586364061
transform 1 0 58420 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_552
timestamp 1586364061
transform 1 0 60076 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_629
timestamp 1586364061
transform 1 0 58972 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_642
timestamp 1586364061
transform 1 0 60168 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_635
timestamp 1586364061
transform 1 0 59524 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_654
timestamp 1586364061
transform 1 0 61272 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_647
timestamp 1586364061
transform 1 0 60628 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_659
timestamp 1586364061
transform 1 0 61732 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_627
timestamp 1586364061
transform 1 0 62836 0 1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_666
timestamp 1586364061
transform 1 0 62376 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_672
timestamp 1586364061
transform 1 0 62928 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_678
timestamp 1586364061
transform 1 0 63480 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_690
timestamp 1586364061
transform 1 0 64584 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_684
timestamp 1586364061
transform 1 0 64032 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_553
timestamp 1586364061
transform 1 0 65688 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_703
timestamp 1586364061
transform 1 0 65780 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_696
timestamp 1586364061
transform 1 0 65136 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_708
timestamp 1586364061
transform 1 0 66240 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_715
timestamp 1586364061
transform 1 0 66884 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_727
timestamp 1586364061
transform 1 0 67988 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_720
timestamp 1586364061
transform 1 0 67344 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_628
timestamp 1586364061
transform 1 0 68448 0 1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_739
timestamp 1586364061
transform 1 0 69092 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_733
timestamp 1586364061
transform 1 0 68540 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_745
timestamp 1586364061
transform 1 0 69644 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_554
timestamp 1586364061
transform 1 0 71300 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_751
timestamp 1586364061
transform 1 0 70196 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_764
timestamp 1586364061
transform 1 0 71392 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_757
timestamp 1586364061
transform 1 0 70748 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_776
timestamp 1586364061
transform 1 0 72496 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_769
timestamp 1586364061
transform 1 0 71852 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_781
timestamp 1586364061
transform 1 0 72956 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_629
timestamp 1586364061
transform 1 0 74060 0 1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_788
timestamp 1586364061
transform 1 0 73600 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_800
timestamp 1586364061
transform 1 0 74704 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_794
timestamp 1586364061
transform 1 0 74152 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_812
timestamp 1586364061
transform 1 0 75808 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_806
timestamp 1586364061
transform 1 0 75256 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_818
timestamp 1586364061
transform 1 0 76360 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_555
timestamp 1586364061
transform 1 0 76912 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_825
timestamp 1586364061
transform 1 0 77004 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_837
timestamp 1586364061
transform 1 0 78108 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_830
timestamp 1586364061
transform 1 0 77464 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_630
timestamp 1586364061
transform 1 0 79672 0 1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_849
timestamp 1586364061
transform 1 0 79212 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_842
timestamp 1586364061
transform 1 0 78568 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_855
timestamp 1586364061
transform 1 0 79764 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_861
timestamp 1586364061
transform 1 0 80316 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_873
timestamp 1586364061
transform 1 0 81420 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_867
timestamp 1586364061
transform 1 0 80868 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_556
timestamp 1586364061
transform 1 0 82524 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_886
timestamp 1586364061
transform 1 0 82616 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_879
timestamp 1586364061
transform 1 0 81972 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_891
timestamp 1586364061
transform 1 0 83076 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_898
timestamp 1586364061
transform 1 0 83720 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_903
timestamp 1586364061
transform 1 0 84180 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_631
timestamp 1586364061
transform 1 0 85284 0 1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_910
timestamp 1586364061
transform 1 0 84824 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_922
timestamp 1586364061
transform 1 0 85928 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_916
timestamp 1586364061
transform 1 0 85376 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_934
timestamp 1586364061
transform 1 0 87032 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_928
timestamp 1586364061
transform 1 0 86480 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_7_940
timestamp 1586364061
transform 1 0 87584 0 1 5984
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_557
timestamp 1586364061
transform 1 0 88136 0 -1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer_A
timestamp 1586364061
transform 1 0 88228 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer_TEB
timestamp 1586364061
transform 1 0 88596 0 1 5984
box -38 -48 222 592
use scs8hd_decap_12  FILLER_6_947
timestamp 1586364061
transform 1 0 88228 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_959
timestamp 1586364061
transform 1 0 89332 0 -1 5984
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_7_946
timestamp 1586364061
transform 1 0 88136 0 1 5984
box -38 -48 130 592
use scs8hd_fill_2  FILLER_7_949
timestamp 1586364061
transform 1 0 88412 0 1 5984
box -38 -48 222 592
use scs8hd_decap_12  FILLER_7_953
timestamp 1586364061
transform 1 0 88780 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_632
timestamp 1586364061
transform 1 0 90896 0 1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_971
timestamp 1586364061
transform 1 0 90436 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_7_965
timestamp 1586364061
transform 1 0 89884 0 1 5984
box -38 -48 774 592
use scs8hd_decap_3  FILLER_7_973
timestamp 1586364061
transform 1 0 90620 0 1 5984
box -38 -48 314 592
use scs8hd_decap_12  FILLER_7_977
timestamp 1586364061
transform 1 0 90988 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_983
timestamp 1586364061
transform 1 0 91540 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_995
timestamp 1586364061
transform 1 0 92644 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_989
timestamp 1586364061
transform 1 0 92092 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_558
timestamp 1586364061
transform 1 0 93748 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_1008
timestamp 1586364061
transform 1 0 93840 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_1001
timestamp 1586364061
transform 1 0 93196 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_1013
timestamp 1586364061
transform 1 0 94300 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_1020
timestamp 1586364061
transform 1 0 94944 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_1032
timestamp 1586364061
transform 1 0 96048 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_1025
timestamp 1586364061
transform 1 0 95404 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_633
timestamp 1586364061
transform 1 0 96508 0 1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_1044
timestamp 1586364061
transform 1 0 97152 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_1038
timestamp 1586364061
transform 1 0 96600 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_1050
timestamp 1586364061
transform 1 0 97704 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_559
timestamp 1586364061
transform 1 0 99360 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_1056
timestamp 1586364061
transform 1 0 98256 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_1069
timestamp 1586364061
transform 1 0 99452 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_1062
timestamp 1586364061
transform 1 0 98808 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_1081
timestamp 1586364061
transform 1 0 100556 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_1074
timestamp 1586364061
transform 1 0 99912 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_1086
timestamp 1586364061
transform 1 0 101016 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_634
timestamp 1586364061
transform 1 0 102120 0 1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_1093
timestamp 1586364061
transform 1 0 101660 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_1105
timestamp 1586364061
transform 1 0 102764 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_1099
timestamp 1586364061
transform 1 0 102212 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_1117
timestamp 1586364061
transform 1 0 103868 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_1111
timestamp 1586364061
transform 1 0 103316 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_1123
timestamp 1586364061
transform 1 0 104420 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_560
timestamp 1586364061
transform 1 0 104972 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_1130
timestamp 1586364061
transform 1 0 105064 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_1135
timestamp 1586364061
transform 1 0 105524 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_635
timestamp 1586364061
transform 1 0 107732 0 1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_1142
timestamp 1586364061
transform 1 0 106168 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_1154
timestamp 1586364061
transform 1 0 107272 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_1147
timestamp 1586364061
transform 1 0 106628 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_1166
timestamp 1586364061
transform 1 0 108376 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_1160
timestamp 1586364061
transform 1 0 107824 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_1172
timestamp 1586364061
transform 1 0 108928 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_561
timestamp 1586364061
transform 1 0 110584 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_1178
timestamp 1586364061
transform 1 0 109480 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_1191
timestamp 1586364061
transform 1 0 110676 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_1184
timestamp 1586364061
transform 1 0 110032 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_1203
timestamp 1586364061
transform 1 0 111780 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_1196
timestamp 1586364061
transform 1 0 111136 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_1208
timestamp 1586364061
transform 1 0 112240 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_636
timestamp 1586364061
transform 1 0 113344 0 1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_1215
timestamp 1586364061
transform 1 0 112884 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_1227
timestamp 1586364061
transform 1 0 113988 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_1221
timestamp 1586364061
transform 1 0 113436 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_1239
timestamp 1586364061
transform 1 0 115092 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_1233
timestamp 1586364061
transform 1 0 114540 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_1245
timestamp 1586364061
transform 1 0 115644 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_562
timestamp 1586364061
transform 1 0 116196 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_1252
timestamp 1586364061
transform 1 0 116288 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_1264
timestamp 1586364061
transform 1 0 117392 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_1257
timestamp 1586364061
transform 1 0 116748 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_637
timestamp 1586364061
transform 1 0 118956 0 1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_1276
timestamp 1586364061
transform 1 0 118496 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_1269
timestamp 1586364061
transform 1 0 117852 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_1282
timestamp 1586364061
transform 1 0 119048 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_1288
timestamp 1586364061
transform 1 0 119600 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_1300
timestamp 1586364061
transform 1 0 120704 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_1294
timestamp 1586364061
transform 1 0 120152 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_563
timestamp 1586364061
transform 1 0 121808 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_1313
timestamp 1586364061
transform 1 0 121900 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_1306
timestamp 1586364061
transform 1 0 121256 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_1318
timestamp 1586364061
transform 1 0 122360 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_1325
timestamp 1586364061
transform 1 0 123004 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_1337
timestamp 1586364061
transform 1 0 124108 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_1330
timestamp 1586364061
transform 1 0 123464 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_638
timestamp 1586364061
transform 1 0 124568 0 1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_1349
timestamp 1586364061
transform 1 0 125212 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_1343
timestamp 1586364061
transform 1 0 124660 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_1355
timestamp 1586364061
transform 1 0 125764 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_564
timestamp 1586364061
transform 1 0 127420 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_1361
timestamp 1586364061
transform 1 0 126316 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_1367
timestamp 1586364061
transform 1 0 126868 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_1374
timestamp 1586364061
transform 1 0 127512 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_1386
timestamp 1586364061
transform 1 0 128616 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_1379
timestamp 1586364061
transform 1 0 127972 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_1391
timestamp 1586364061
transform 1 0 129076 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_639
timestamp 1586364061
transform 1 0 130180 0 1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_1398
timestamp 1586364061
transform 1 0 129720 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_1404
timestamp 1586364061
transform 1 0 130272 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_1410
timestamp 1586364061
transform 1 0 130824 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_1422
timestamp 1586364061
transform 1 0 131928 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_1416
timestamp 1586364061
transform 1 0 131376 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_565
timestamp 1586364061
transform 1 0 133032 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_1435
timestamp 1586364061
transform 1 0 133124 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_1428
timestamp 1586364061
transform 1 0 132480 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_1440
timestamp 1586364061
transform 1 0 133584 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_1447
timestamp 1586364061
transform 1 0 134228 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_1459
timestamp 1586364061
transform 1 0 135332 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_1452
timestamp 1586364061
transform 1 0 134688 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_640
timestamp 1586364061
transform 1 0 135792 0 1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_1471
timestamp 1586364061
transform 1 0 136436 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_1465
timestamp 1586364061
transform 1 0 135884 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_1477
timestamp 1586364061
transform 1 0 136988 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_566
timestamp 1586364061
transform 1 0 138644 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_1483
timestamp 1586364061
transform 1 0 137540 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_1496
timestamp 1586364061
transform 1 0 138736 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_1489
timestamp 1586364061
transform 1 0 138092 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_1508
timestamp 1586364061
transform 1 0 139840 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_1501
timestamp 1586364061
transform 1 0 139196 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_1513
timestamp 1586364061
transform 1 0 140300 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_641
timestamp 1586364061
transform 1 0 141404 0 1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_1520
timestamp 1586364061
transform 1 0 140944 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_1532
timestamp 1586364061
transform 1 0 142048 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_1526
timestamp 1586364061
transform 1 0 141496 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_1544
timestamp 1586364061
transform 1 0 143152 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_1538
timestamp 1586364061
transform 1 0 142600 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_1550
timestamp 1586364061
transform 1 0 143704 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_567
timestamp 1586364061
transform 1 0 144256 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_1557
timestamp 1586364061
transform 1 0 144348 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_1569
timestamp 1586364061
transform 1 0 145452 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_1562
timestamp 1586364061
transform 1 0 144808 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_642
timestamp 1586364061
transform 1 0 147016 0 1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_1581
timestamp 1586364061
transform 1 0 146556 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_1574
timestamp 1586364061
transform 1 0 145912 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_1587
timestamp 1586364061
transform 1 0 147108 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_1593
timestamp 1586364061
transform 1 0 147660 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_1605
timestamp 1586364061
transform 1 0 148764 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_1599
timestamp 1586364061
transform 1 0 148212 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_568
timestamp 1586364061
transform 1 0 149868 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_1618
timestamp 1586364061
transform 1 0 149960 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_1611
timestamp 1586364061
transform 1 0 149316 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_1623
timestamp 1586364061
transform 1 0 150420 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_1630
timestamp 1586364061
transform 1 0 151064 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_1635
timestamp 1586364061
transform 1 0 151524 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_643
timestamp 1586364061
transform 1 0 152628 0 1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_1642
timestamp 1586364061
transform 1 0 152168 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_1654
timestamp 1586364061
transform 1 0 153272 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_1648
timestamp 1586364061
transform 1 0 152720 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_1666
timestamp 1586364061
transform 1 0 154376 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_1660
timestamp 1586364061
transform 1 0 153824 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_1672
timestamp 1586364061
transform 1 0 154928 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_569
timestamp 1586364061
transform 1 0 155480 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_1679
timestamp 1586364061
transform 1 0 155572 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_1691
timestamp 1586364061
transform 1 0 156676 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_1684
timestamp 1586364061
transform 1 0 156032 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_644
timestamp 1586364061
transform 1 0 158240 0 1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_1703
timestamp 1586364061
transform 1 0 157780 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_1696
timestamp 1586364061
transform 1 0 157136 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_1709
timestamp 1586364061
transform 1 0 158332 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_1715
timestamp 1586364061
transform 1 0 158884 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_1727
timestamp 1586364061
transform 1 0 159988 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_1721
timestamp 1586364061
transform 1 0 159436 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_570
timestamp 1586364061
transform 1 0 161092 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_1740
timestamp 1586364061
transform 1 0 161184 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_1733
timestamp 1586364061
transform 1 0 160540 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_1745
timestamp 1586364061
transform 1 0 161644 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_1752
timestamp 1586364061
transform 1 0 162288 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_1764
timestamp 1586364061
transform 1 0 163392 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_1757
timestamp 1586364061
transform 1 0 162748 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_645
timestamp 1586364061
transform 1 0 163852 0 1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_1776
timestamp 1586364061
transform 1 0 164496 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_1770
timestamp 1586364061
transform 1 0 163944 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_1782
timestamp 1586364061
transform 1 0 165048 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_571
timestamp 1586364061
transform 1 0 166704 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_1788
timestamp 1586364061
transform 1 0 165600 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_1801
timestamp 1586364061
transform 1 0 166796 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_1794
timestamp 1586364061
transform 1 0 166152 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_1813
timestamp 1586364061
transform 1 0 167900 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_1806
timestamp 1586364061
transform 1 0 167256 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_1818
timestamp 1586364061
transform 1 0 168360 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_646
timestamp 1586364061
transform 1 0 169464 0 1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_1825
timestamp 1586364061
transform 1 0 169004 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_1837
timestamp 1586364061
transform 1 0 170108 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_7_1831
timestamp 1586364061
transform 1 0 169556 0 1 5984
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA__20__A
timestamp 1586364061
transform 1 0 170568 0 1 5984
box -38 -48 222 592
use scs8hd_decap_12  FILLER_6_1849
timestamp 1586364061
transform 1 0 171212 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_7_1839
timestamp 1586364061
transform 1 0 170292 0 1 5984
box -38 -48 314 592
use scs8hd_decap_12  FILLER_7_1844
timestamp 1586364061
transform 1 0 170752 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_572
timestamp 1586364061
transform 1 0 172316 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_1862
timestamp 1586364061
transform 1 0 172408 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_1856
timestamp 1586364061
transform 1 0 171856 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_1868
timestamp 1586364061
transform 1 0 172960 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_1874
timestamp 1586364061
transform 1 0 173512 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_1886
timestamp 1586364061
transform 1 0 174616 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_7_1880
timestamp 1586364061
transform 1 0 174064 0 1 5984
box -38 -48 774 592
use scs8hd_decap_3  FILLER_7_1888
timestamp 1586364061
transform 1 0 174800 0 1 5984
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_647
timestamp 1586364061
transform 1 0 175076 0 1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_1898
timestamp 1586364061
transform 1 0 175720 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_1892
timestamp 1586364061
transform 1 0 175168 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_1904
timestamp 1586364061
transform 1 0 176272 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_573
timestamp 1586364061
transform 1 0 177928 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_1910
timestamp 1586364061
transform 1 0 176824 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_1923
timestamp 1586364061
transform 1 0 178020 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_1916
timestamp 1586364061
transform 1 0 177376 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_1935
timestamp 1586364061
transform 1 0 179124 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_1928
timestamp 1586364061
transform 1 0 178480 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_1940
timestamp 1586364061
transform 1 0 179584 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_648
timestamp 1586364061
transform 1 0 180688 0 1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_1947
timestamp 1586364061
transform 1 0 180228 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_1959
timestamp 1586364061
transform 1 0 181332 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_1953
timestamp 1586364061
transform 1 0 180780 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_1971
timestamp 1586364061
transform 1 0 182436 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_1965
timestamp 1586364061
transform 1 0 181884 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_1977
timestamp 1586364061
transform 1 0 182988 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_574
timestamp 1586364061
transform 1 0 183540 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_1984
timestamp 1586364061
transform 1 0 183632 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_1996
timestamp 1586364061
transform 1 0 184736 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_1989
timestamp 1586364061
transform 1 0 184092 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_649
timestamp 1586364061
transform 1 0 186300 0 1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_2008
timestamp 1586364061
transform 1 0 185840 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_2001
timestamp 1586364061
transform 1 0 185196 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_2014
timestamp 1586364061
transform 1 0 186392 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_2020
timestamp 1586364061
transform 1 0 186944 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_2032
timestamp 1586364061
transform 1 0 188048 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_2026
timestamp 1586364061
transform 1 0 187496 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_575
timestamp 1586364061
transform 1 0 189152 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_2045
timestamp 1586364061
transform 1 0 189244 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_2038
timestamp 1586364061
transform 1 0 188600 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_2050
timestamp 1586364061
transform 1 0 189704 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_2057
timestamp 1586364061
transform 1 0 190348 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_2069
timestamp 1586364061
transform 1 0 191452 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_2062
timestamp 1586364061
transform 1 0 190808 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_650
timestamp 1586364061
transform 1 0 191912 0 1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_2081
timestamp 1586364061
transform 1 0 192556 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_2075
timestamp 1586364061
transform 1 0 192004 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_2093
timestamp 1586364061
transform 1 0 193660 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_2087
timestamp 1586364061
transform 1 0 193108 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_2099
timestamp 1586364061
transform 1 0 194212 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_576
timestamp 1586364061
transform 1 0 194764 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_2106
timestamp 1586364061
transform 1 0 194856 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_2118
timestamp 1586364061
transform 1 0 195960 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_2111
timestamp 1586364061
transform 1 0 195316 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_651
timestamp 1586364061
transform 1 0 197524 0 1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_2130
timestamp 1586364061
transform 1 0 197064 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_2123
timestamp 1586364061
transform 1 0 196420 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_2136
timestamp 1586364061
transform 1 0 197616 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_2142
timestamp 1586364061
transform 1 0 198168 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_2154
timestamp 1586364061
transform 1 0 199272 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_2148
timestamp 1586364061
transform 1 0 198720 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_577
timestamp 1586364061
transform 1 0 200376 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_2167
timestamp 1586364061
transform 1 0 200468 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_2160
timestamp 1586364061
transform 1 0 199824 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_2172
timestamp 1586364061
transform 1 0 200928 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_2179
timestamp 1586364061
transform 1 0 201572 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_2191
timestamp 1586364061
transform 1 0 202676 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_2184
timestamp 1586364061
transform 1 0 202032 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_652
timestamp 1586364061
transform 1 0 203136 0 1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_2203
timestamp 1586364061
transform 1 0 203780 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_2197
timestamp 1586364061
transform 1 0 203228 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_2209
timestamp 1586364061
transform 1 0 204332 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_578
timestamp 1586364061
transform 1 0 205988 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_2215
timestamp 1586364061
transform 1 0 204884 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_2228
timestamp 1586364061
transform 1 0 206080 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_2221
timestamp 1586364061
transform 1 0 205436 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_2240
timestamp 1586364061
transform 1 0 207184 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_2233
timestamp 1586364061
transform 1 0 206540 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_2245
timestamp 1586364061
transform 1 0 207644 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_653
timestamp 1586364061
transform 1 0 208748 0 1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_2252
timestamp 1586364061
transform 1 0 208288 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_2264
timestamp 1586364061
transform 1 0 209392 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_2258
timestamp 1586364061
transform 1 0 208840 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_2276
timestamp 1586364061
transform 1 0 210496 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_2270
timestamp 1586364061
transform 1 0 209944 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_2282
timestamp 1586364061
transform 1 0 211048 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_579
timestamp 1586364061
transform 1 0 211600 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_2289
timestamp 1586364061
transform 1 0 211692 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_2294
timestamp 1586364061
transform 1 0 212152 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_654
timestamp 1586364061
transform 1 0 214360 0 1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_2301
timestamp 1586364061
transform 1 0 212796 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_2313
timestamp 1586364061
transform 1 0 213900 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_2306
timestamp 1586364061
transform 1 0 213256 0 1 5984
box -38 -48 1142 592
use scs8hd_inv_8  _11_
timestamp 1586364061
transform 1 0 215096 0 -1 5984
box -38 -48 866 592
use scs8hd_ebufn_1  logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer
timestamp 1586364061
transform 1 0 215556 0 1 5984
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA_logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer_A
timestamp 1586364061
transform 1 0 215372 0 1 5984
box -38 -48 222 592
use scs8hd_fill_1  FILLER_6_2325
timestamp 1586364061
transform 1 0 215004 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_8  FILLER_6_2335
timestamp 1586364061
transform 1 0 215924 0 -1 5984
box -38 -48 774 592
use scs8hd_decap_8  FILLER_7_2319
timestamp 1586364061
transform 1 0 214452 0 1 5984
box -38 -48 774 592
use scs8hd_fill_2  FILLER_7_2327
timestamp 1586364061
transform 1 0 215188 0 1 5984
box -38 -48 222 592
use scs8hd_ebufn_1  logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer
timestamp 1586364061
transform 1 0 217304 0 -1 5984
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_580
timestamp 1586364061
transform 1 0 217212 0 -1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__10__A
timestamp 1586364061
transform 1 0 216752 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_1  FILLER_6_2343
timestamp 1586364061
transform 1 0 216660 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_3  FILLER_6_2346
timestamp 1586364061
transform 1 0 216936 0 -1 5984
box -38 -48 314 592
use scs8hd_decap_12  FILLER_7_2339
timestamp 1586364061
transform 1 0 216292 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_2351
timestamp 1586364061
transform 1 0 217396 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_2358
timestamp 1586364061
transform 1 0 218040 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_2370
timestamp 1586364061
transform 1 0 219144 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_2363
timestamp 1586364061
transform 1 0 218500 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_655
timestamp 1586364061
transform 1 0 219972 0 1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_2382
timestamp 1586364061
transform 1 0 220248 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_7_2375
timestamp 1586364061
transform 1 0 219604 0 1 5984
box -38 -48 406 592
use scs8hd_decap_12  FILLER_7_2380
timestamp 1586364061
transform 1 0 220064 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_2394
timestamp 1586364061
transform 1 0 221352 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_6_2406
timestamp 1586364061
transform 1 0 222456 0 -1 5984
box -38 -48 406 592
use scs8hd_decap_12  FILLER_7_2392
timestamp 1586364061
transform 1 0 221168 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_2404
timestamp 1586364061
transform 1 0 222272 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_581
timestamp 1586364061
transform 1 0 222824 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_2411
timestamp 1586364061
transform 1 0 222916 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_2423
timestamp 1586364061
transform 1 0 224020 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_2416
timestamp 1586364061
transform 1 0 223376 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_656
timestamp 1586364061
transform 1 0 225584 0 1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer_A
timestamp 1586364061
transform 1 0 225308 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer_TEB
timestamp 1586364061
transform 1 0 225860 0 1 5984
box -38 -48 222 592
use scs8hd_decap_12  FILLER_6_2435
timestamp 1586364061
transform 1 0 225124 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_7_2428
timestamp 1586364061
transform 1 0 224480 0 1 5984
box -38 -48 774 592
use scs8hd_fill_1  FILLER_7_2436
timestamp 1586364061
transform 1 0 225216 0 1 5984
box -38 -48 130 592
use scs8hd_fill_1  FILLER_7_2439
timestamp 1586364061
transform 1 0 225492 0 1 5984
box -38 -48 130 592
use scs8hd_fill_2  FILLER_7_2441
timestamp 1586364061
transform 1 0 225676 0 1 5984
box -38 -48 222 592
use scs8hd_decap_12  FILLER_6_2447
timestamp 1586364061
transform 1 0 226228 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_2459
timestamp 1586364061
transform 1 0 227332 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_2445
timestamp 1586364061
transform 1 0 226044 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_2457
timestamp 1586364061
transform 1 0 227148 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_582
timestamp 1586364061
transform 1 0 228436 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_2472
timestamp 1586364061
transform 1 0 228528 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_2469
timestamp 1586364061
transform 1 0 228252 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_2484
timestamp 1586364061
transform 1 0 229632 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_2496
timestamp 1586364061
transform 1 0 230736 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_2481
timestamp 1586364061
transform 1 0 229356 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_7_2493
timestamp 1586364061
transform 1 0 230460 0 1 5984
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_657
timestamp 1586364061
transform 1 0 231196 0 1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_2508
timestamp 1586364061
transform 1 0 231840 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_2502
timestamp 1586364061
transform 1 0 231288 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_2514
timestamp 1586364061
transform 1 0 232392 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_583
timestamp 1586364061
transform 1 0 234048 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_2520
timestamp 1586364061
transform 1 0 232944 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_2526
timestamp 1586364061
transform 1 0 233496 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_2533
timestamp 1586364061
transform 1 0 234140 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_2545
timestamp 1586364061
transform 1 0 235244 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_2538
timestamp 1586364061
transform 1 0 234600 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_2550
timestamp 1586364061
transform 1 0 235704 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_658
timestamp 1586364061
transform 1 0 236808 0 1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_2557
timestamp 1586364061
transform 1 0 236348 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_2563
timestamp 1586364061
transform 1 0 236900 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_2569
timestamp 1586364061
transform 1 0 237452 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_2581
timestamp 1586364061
transform 1 0 238556 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_2575
timestamp 1586364061
transform 1 0 238004 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_584
timestamp 1586364061
transform 1 0 239660 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_2594
timestamp 1586364061
transform 1 0 239752 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_2587
timestamp 1586364061
transform 1 0 239108 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_2599
timestamp 1586364061
transform 1 0 240212 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_2606
timestamp 1586364061
transform 1 0 240856 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_2618
timestamp 1586364061
transform 1 0 241960 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_2611
timestamp 1586364061
transform 1 0 241316 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_659
timestamp 1586364061
transform 1 0 242420 0 1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_2630
timestamp 1586364061
transform 1 0 243064 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_2624
timestamp 1586364061
transform 1 0 242512 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_2636
timestamp 1586364061
transform 1 0 243616 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_585
timestamp 1586364061
transform 1 0 245272 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_2642
timestamp 1586364061
transform 1 0 244168 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_2655
timestamp 1586364061
transform 1 0 245364 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_2648
timestamp 1586364061
transform 1 0 244720 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_2667
timestamp 1586364061
transform 1 0 246468 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_2660
timestamp 1586364061
transform 1 0 245824 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_2672
timestamp 1586364061
transform 1 0 246928 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_660
timestamp 1586364061
transform 1 0 248032 0 1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_2679
timestamp 1586364061
transform 1 0 247572 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_2691
timestamp 1586364061
transform 1 0 248676 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_2685
timestamp 1586364061
transform 1 0 248124 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_2703
timestamp 1586364061
transform 1 0 249780 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_2697
timestamp 1586364061
transform 1 0 249228 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_2709
timestamp 1586364061
transform 1 0 250332 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_586
timestamp 1586364061
transform 1 0 250884 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_2716
timestamp 1586364061
transform 1 0 250976 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_2728
timestamp 1586364061
transform 1 0 252080 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_2721
timestamp 1586364061
transform 1 0 251436 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_661
timestamp 1586364061
transform 1 0 253644 0 1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_2740
timestamp 1586364061
transform 1 0 253184 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_2733
timestamp 1586364061
transform 1 0 252540 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_2746
timestamp 1586364061
transform 1 0 253736 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_2752
timestamp 1586364061
transform 1 0 254288 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_2764
timestamp 1586364061
transform 1 0 255392 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_2758
timestamp 1586364061
transform 1 0 254840 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_587
timestamp 1586364061
transform 1 0 256496 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_2777
timestamp 1586364061
transform 1 0 256588 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_2770
timestamp 1586364061
transform 1 0 255944 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_2782
timestamp 1586364061
transform 1 0 257048 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_2789
timestamp 1586364061
transform 1 0 257692 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_2794
timestamp 1586364061
transform 1 0 258152 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_662
timestamp 1586364061
transform 1 0 259256 0 1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_2801
timestamp 1586364061
transform 1 0 258796 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_2813
timestamp 1586364061
transform 1 0 259900 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_2807
timestamp 1586364061
transform 1 0 259348 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_2825
timestamp 1586364061
transform 1 0 261004 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_2819
timestamp 1586364061
transform 1 0 260452 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_2831
timestamp 1586364061
transform 1 0 261556 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_588
timestamp 1586364061
transform 1 0 262108 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_2838
timestamp 1586364061
transform 1 0 262200 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_2850
timestamp 1586364061
transform 1 0 263304 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_2843
timestamp 1586364061
transform 1 0 262660 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_663
timestamp 1586364061
transform 1 0 264868 0 1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_2862
timestamp 1586364061
transform 1 0 264408 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_2855
timestamp 1586364061
transform 1 0 263764 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_2868
timestamp 1586364061
transform 1 0 264960 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_2874
timestamp 1586364061
transform 1 0 265512 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_2886
timestamp 1586364061
transform 1 0 266616 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_2880
timestamp 1586364061
transform 1 0 266064 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_589
timestamp 1586364061
transform 1 0 267720 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_2899
timestamp 1586364061
transform 1 0 267812 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_2892
timestamp 1586364061
transform 1 0 267168 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_2904
timestamp 1586364061
transform 1 0 268272 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_2911
timestamp 1586364061
transform 1 0 268916 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_2923
timestamp 1586364061
transform 1 0 270020 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_2916
timestamp 1586364061
transform 1 0 269376 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_664
timestamp 1586364061
transform 1 0 270480 0 1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_2935
timestamp 1586364061
transform 1 0 271124 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_2929
timestamp 1586364061
transform 1 0 270572 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_2941
timestamp 1586364061
transform 1 0 271676 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_590
timestamp 1586364061
transform 1 0 273332 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_2947
timestamp 1586364061
transform 1 0 272228 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_2960
timestamp 1586364061
transform 1 0 273424 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_2953
timestamp 1586364061
transform 1 0 272780 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_2972
timestamp 1586364061
transform 1 0 274528 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_2965
timestamp 1586364061
transform 1 0 273884 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_2977
timestamp 1586364061
transform 1 0 274988 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_665
timestamp 1586364061
transform 1 0 276092 0 1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_2984
timestamp 1586364061
transform 1 0 275632 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_2996
timestamp 1586364061
transform 1 0 276736 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_2990
timestamp 1586364061
transform 1 0 276184 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_3008
timestamp 1586364061
transform 1 0 277840 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_3002
timestamp 1586364061
transform 1 0 277288 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_3014
timestamp 1586364061
transform 1 0 278392 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_591
timestamp 1586364061
transform 1 0 278944 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_3021
timestamp 1586364061
transform 1 0 279036 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_3026
timestamp 1586364061
transform 1 0 279496 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_666
timestamp 1586364061
transform 1 0 281704 0 1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_3033
timestamp 1586364061
transform 1 0 280140 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_3045
timestamp 1586364061
transform 1 0 281244 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_3038
timestamp 1586364061
transform 1 0 280600 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_3057
timestamp 1586364061
transform 1 0 282348 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_3051
timestamp 1586364061
transform 1 0 281796 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_3063
timestamp 1586364061
transform 1 0 282900 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_592
timestamp 1586364061
transform 1 0 284556 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_3069
timestamp 1586364061
transform 1 0 283452 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_3082
timestamp 1586364061
transform 1 0 284648 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_3075
timestamp 1586364061
transform 1 0 284004 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_3094
timestamp 1586364061
transform 1 0 285752 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_3087
timestamp 1586364061
transform 1 0 285108 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_3099
timestamp 1586364061
transform 1 0 286212 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_667
timestamp 1586364061
transform 1 0 287316 0 1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_3106
timestamp 1586364061
transform 1 0 286856 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_3118
timestamp 1586364061
transform 1 0 287960 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_3112
timestamp 1586364061
transform 1 0 287408 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_3130
timestamp 1586364061
transform 1 0 289064 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_3124
timestamp 1586364061
transform 1 0 288512 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_3136
timestamp 1586364061
transform 1 0 289616 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_593
timestamp 1586364061
transform 1 0 290168 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_3143
timestamp 1586364061
transform 1 0 290260 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_3155
timestamp 1586364061
transform 1 0 291364 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_3148
timestamp 1586364061
transform 1 0 290720 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_668
timestamp 1586364061
transform 1 0 292928 0 1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_3167
timestamp 1586364061
transform 1 0 292468 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_3160
timestamp 1586364061
transform 1 0 291824 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_3173
timestamp 1586364061
transform 1 0 293020 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_3179
timestamp 1586364061
transform 1 0 293572 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_3191
timestamp 1586364061
transform 1 0 294676 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_3185
timestamp 1586364061
transform 1 0 294124 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_594
timestamp 1586364061
transform 1 0 295780 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_3204
timestamp 1586364061
transform 1 0 295872 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_3197
timestamp 1586364061
transform 1 0 295228 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_3209
timestamp 1586364061
transform 1 0 296332 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_3216
timestamp 1586364061
transform 1 0 296976 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_3228
timestamp 1586364061
transform 1 0 298080 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_3221
timestamp 1586364061
transform 1 0 297436 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_669
timestamp 1586364061
transform 1 0 298540 0 1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_3240
timestamp 1586364061
transform 1 0 299184 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_3234
timestamp 1586364061
transform 1 0 298632 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_3246
timestamp 1586364061
transform 1 0 299736 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_595
timestamp 1586364061
transform 1 0 301392 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_3252
timestamp 1586364061
transform 1 0 300288 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_3258
timestamp 1586364061
transform 1 0 300840 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_3265
timestamp 1586364061
transform 1 0 301484 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_3277
timestamp 1586364061
transform 1 0 302588 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_3270
timestamp 1586364061
transform 1 0 301944 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_670
timestamp 1586364061
transform 1 0 304152 0 1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_3289
timestamp 1586364061
transform 1 0 303692 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_3282
timestamp 1586364061
transform 1 0 303048 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_3295
timestamp 1586364061
transform 1 0 304244 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_3301
timestamp 1586364061
transform 1 0 304796 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_3313
timestamp 1586364061
transform 1 0 305900 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_3307
timestamp 1586364061
transform 1 0 305348 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_596
timestamp 1586364061
transform 1 0 307004 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_3326
timestamp 1586364061
transform 1 0 307096 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_3319
timestamp 1586364061
transform 1 0 306452 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_3331
timestamp 1586364061
transform 1 0 307556 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_3338
timestamp 1586364061
transform 1 0 308200 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_3350
timestamp 1586364061
transform 1 0 309304 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_3343
timestamp 1586364061
transform 1 0 308660 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_671
timestamp 1586364061
transform 1 0 309764 0 1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_3362
timestamp 1586364061
transform 1 0 310408 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_3356
timestamp 1586364061
transform 1 0 309856 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_3368
timestamp 1586364061
transform 1 0 310960 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_597
timestamp 1586364061
transform 1 0 312616 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_3374
timestamp 1586364061
transform 1 0 311512 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_3387
timestamp 1586364061
transform 1 0 312708 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_3380
timestamp 1586364061
transform 1 0 312064 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_3399
timestamp 1586364061
transform 1 0 313812 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_3392
timestamp 1586364061
transform 1 0 313168 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_3404
timestamp 1586364061
transform 1 0 314272 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_672
timestamp 1586364061
transform 1 0 315376 0 1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_3411
timestamp 1586364061
transform 1 0 314916 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_3423
timestamp 1586364061
transform 1 0 316020 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_3417
timestamp 1586364061
transform 1 0 315468 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_3435
timestamp 1586364061
transform 1 0 317124 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_3429
timestamp 1586364061
transform 1 0 316572 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_3441
timestamp 1586364061
transform 1 0 317676 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_598
timestamp 1586364061
transform 1 0 318228 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_3448
timestamp 1586364061
transform 1 0 318320 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_3460
timestamp 1586364061
transform 1 0 319424 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_3453
timestamp 1586364061
transform 1 0 318780 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_673
timestamp 1586364061
transform 1 0 320988 0 1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_3472
timestamp 1586364061
transform 1 0 320528 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_3465
timestamp 1586364061
transform 1 0 319884 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_3478
timestamp 1586364061
transform 1 0 321080 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_3484
timestamp 1586364061
transform 1 0 321632 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_3496
timestamp 1586364061
transform 1 0 322736 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_3490
timestamp 1586364061
transform 1 0 322184 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_599
timestamp 1586364061
transform 1 0 323840 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_3509
timestamp 1586364061
transform 1 0 323932 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_3502
timestamp 1586364061
transform 1 0 323288 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_3521
timestamp 1586364061
transform 1 0 325036 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_3514
timestamp 1586364061
transform 1 0 324392 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_3526
timestamp 1586364061
transform 1 0 325496 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_674
timestamp 1586364061
transform 1 0 326600 0 1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_3533
timestamp 1586364061
transform 1 0 326140 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_3545
timestamp 1586364061
transform 1 0 327244 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_3539
timestamp 1586364061
transform 1 0 326692 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_3557
timestamp 1586364061
transform 1 0 328348 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_3551
timestamp 1586364061
transform 1 0 327796 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_3563
timestamp 1586364061
transform 1 0 328900 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_600
timestamp 1586364061
transform 1 0 329452 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_3570
timestamp 1586364061
transform 1 0 329544 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_3582
timestamp 1586364061
transform 1 0 330648 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_3575
timestamp 1586364061
transform 1 0 330004 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_675
timestamp 1586364061
transform 1 0 332212 0 1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_3594
timestamp 1586364061
transform 1 0 331752 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_3587
timestamp 1586364061
transform 1 0 331108 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_3600
timestamp 1586364061
transform 1 0 332304 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_3606
timestamp 1586364061
transform 1 0 332856 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_3618
timestamp 1586364061
transform 1 0 333960 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_3612
timestamp 1586364061
transform 1 0 333408 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_601
timestamp 1586364061
transform 1 0 335064 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_3631
timestamp 1586364061
transform 1 0 335156 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_3624
timestamp 1586364061
transform 1 0 334512 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_3636
timestamp 1586364061
transform 1 0 335616 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_3643
timestamp 1586364061
transform 1 0 336260 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_3655
timestamp 1586364061
transform 1 0 337364 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_3648
timestamp 1586364061
transform 1 0 336720 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_676
timestamp 1586364061
transform 1 0 337824 0 1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_3667
timestamp 1586364061
transform 1 0 338468 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_3661
timestamp 1586364061
transform 1 0 337916 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_3673
timestamp 1586364061
transform 1 0 339020 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_602
timestamp 1586364061
transform 1 0 340676 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_3679
timestamp 1586364061
transform 1 0 339572 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_3692
timestamp 1586364061
transform 1 0 340768 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_3685
timestamp 1586364061
transform 1 0 340124 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_3704
timestamp 1586364061
transform 1 0 341872 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_3697
timestamp 1586364061
transform 1 0 341228 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_3709
timestamp 1586364061
transform 1 0 342332 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_677
timestamp 1586364061
transform 1 0 343436 0 1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_3716
timestamp 1586364061
transform 1 0 342976 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_3722
timestamp 1586364061
transform 1 0 343528 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_3728
timestamp 1586364061
transform 1 0 344080 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_3740
timestamp 1586364061
transform 1 0 345184 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_3734
timestamp 1586364061
transform 1 0 344632 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_603
timestamp 1586364061
transform 1 0 346288 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_3753
timestamp 1586364061
transform 1 0 346380 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_3746
timestamp 1586364061
transform 1 0 345736 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_3758
timestamp 1586364061
transform 1 0 346840 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_3765
timestamp 1586364061
transform 1 0 347484 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_3777
timestamp 1586364061
transform 1 0 348588 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_3770
timestamp 1586364061
transform 1 0 347944 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_678
timestamp 1586364061
transform 1 0 349048 0 1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_3789
timestamp 1586364061
transform 1 0 349692 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_3783
timestamp 1586364061
transform 1 0 349140 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_3795
timestamp 1586364061
transform 1 0 350244 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_604
timestamp 1586364061
transform 1 0 351900 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_3801
timestamp 1586364061
transform 1 0 350796 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_3814
timestamp 1586364061
transform 1 0 351992 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_3807
timestamp 1586364061
transform 1 0 351348 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_3826
timestamp 1586364061
transform 1 0 353096 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_3819
timestamp 1586364061
transform 1 0 352452 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_3831
timestamp 1586364061
transform 1 0 353556 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_679
timestamp 1586364061
transform 1 0 354660 0 1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_3838
timestamp 1586364061
transform 1 0 354200 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_3850
timestamp 1586364061
transform 1 0 355304 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_3844
timestamp 1586364061
transform 1 0 354752 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_3862
timestamp 1586364061
transform 1 0 356408 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_3856
timestamp 1586364061
transform 1 0 355856 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_3868
timestamp 1586364061
transform 1 0 356960 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_605
timestamp 1586364061
transform 1 0 357512 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_3875
timestamp 1586364061
transform 1 0 357604 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_3887
timestamp 1586364061
transform 1 0 358708 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_3880
timestamp 1586364061
transform 1 0 358064 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_680
timestamp 1586364061
transform 1 0 360272 0 1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_3899
timestamp 1586364061
transform 1 0 359812 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_3892
timestamp 1586364061
transform 1 0 359168 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_3905
timestamp 1586364061
transform 1 0 360364 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_3911
timestamp 1586364061
transform 1 0 360916 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_3923
timestamp 1586364061
transform 1 0 362020 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_3917
timestamp 1586364061
transform 1 0 361468 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_606
timestamp 1586364061
transform 1 0 363124 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_3936
timestamp 1586364061
transform 1 0 363216 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_3929
timestamp 1586364061
transform 1 0 362572 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_3941
timestamp 1586364061
transform 1 0 363676 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_3948
timestamp 1586364061
transform 1 0 364320 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_3953
timestamp 1586364061
transform 1 0 364780 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_681
timestamp 1586364061
transform 1 0 365884 0 1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_3960
timestamp 1586364061
transform 1 0 365424 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_3972
timestamp 1586364061
transform 1 0 366528 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_3966
timestamp 1586364061
transform 1 0 365976 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_3984
timestamp 1586364061
transform 1 0 367632 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_3978
timestamp 1586364061
transform 1 0 367080 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_3990
timestamp 1586364061
transform 1 0 368184 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_607
timestamp 1586364061
transform 1 0 368736 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_3997
timestamp 1586364061
transform 1 0 368828 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_4009
timestamp 1586364061
transform 1 0 369932 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_4002
timestamp 1586364061
transform 1 0 369288 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_682
timestamp 1586364061
transform 1 0 371496 0 1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_4021
timestamp 1586364061
transform 1 0 371036 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_4014
timestamp 1586364061
transform 1 0 370392 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_4027
timestamp 1586364061
transform 1 0 371588 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_4033
timestamp 1586364061
transform 1 0 372140 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_4045
timestamp 1586364061
transform 1 0 373244 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_4039
timestamp 1586364061
transform 1 0 372692 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_608
timestamp 1586364061
transform 1 0 374348 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_4058
timestamp 1586364061
transform 1 0 374440 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_4051
timestamp 1586364061
transform 1 0 373796 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_4063
timestamp 1586364061
transform 1 0 374900 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_4070
timestamp 1586364061
transform 1 0 375544 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_4082
timestamp 1586364061
transform 1 0 376648 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_4075
timestamp 1586364061
transform 1 0 376004 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_683
timestamp 1586364061
transform 1 0 377108 0 1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_4094
timestamp 1586364061
transform 1 0 377752 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_4088
timestamp 1586364061
transform 1 0 377200 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_4100
timestamp 1586364061
transform 1 0 378304 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_609
timestamp 1586364061
transform 1 0 379960 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_4106
timestamp 1586364061
transform 1 0 378856 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_4119
timestamp 1586364061
transform 1 0 380052 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_4112
timestamp 1586364061
transform 1 0 379408 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_4131
timestamp 1586364061
transform 1 0 381156 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_4124
timestamp 1586364061
transform 1 0 380512 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_4136
timestamp 1586364061
transform 1 0 381616 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_684
timestamp 1586364061
transform 1 0 382720 0 1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_4143
timestamp 1586364061
transform 1 0 382260 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_4155
timestamp 1586364061
transform 1 0 383364 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_4149
timestamp 1586364061
transform 1 0 382812 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_4167
timestamp 1586364061
transform 1 0 384468 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_4161
timestamp 1586364061
transform 1 0 383916 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_4173
timestamp 1586364061
transform 1 0 385020 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_610
timestamp 1586364061
transform 1 0 385572 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_4180
timestamp 1586364061
transform 1 0 385664 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_4185
timestamp 1586364061
transform 1 0 386124 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_685
timestamp 1586364061
transform 1 0 388332 0 1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_4192
timestamp 1586364061
transform 1 0 386768 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_4204
timestamp 1586364061
transform 1 0 387872 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_4197
timestamp 1586364061
transform 1 0 387228 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_4216
timestamp 1586364061
transform 1 0 388976 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_4210
timestamp 1586364061
transform 1 0 388424 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_4222
timestamp 1586364061
transform 1 0 389528 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_611
timestamp 1586364061
transform 1 0 391184 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_4228
timestamp 1586364061
transform 1 0 390080 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_4241
timestamp 1586364061
transform 1 0 391276 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_4234
timestamp 1586364061
transform 1 0 390632 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_4253
timestamp 1586364061
transform 1 0 392380 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_4246
timestamp 1586364061
transform 1 0 391736 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_4258
timestamp 1586364061
transform 1 0 392840 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_686
timestamp 1586364061
transform 1 0 393944 0 1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_4265
timestamp 1586364061
transform 1 0 393484 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_4277
timestamp 1586364061
transform 1 0 394588 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_4271
timestamp 1586364061
transform 1 0 394036 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_4289
timestamp 1586364061
transform 1 0 395692 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_4283
timestamp 1586364061
transform 1 0 395140 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_4295
timestamp 1586364061
transform 1 0 396244 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_612
timestamp 1586364061
transform 1 0 396796 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_4302
timestamp 1586364061
transform 1 0 396888 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_4314
timestamp 1586364061
transform 1 0 397992 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_4307
timestamp 1586364061
transform 1 0 397348 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_687
timestamp 1586364061
transform 1 0 399556 0 1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_4326
timestamp 1586364061
transform 1 0 399096 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_4319
timestamp 1586364061
transform 1 0 398452 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_4332
timestamp 1586364061
transform 1 0 399648 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_4338
timestamp 1586364061
transform 1 0 400200 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_4350
timestamp 1586364061
transform 1 0 401304 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_4344
timestamp 1586364061
transform 1 0 400752 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_613
timestamp 1586364061
transform 1 0 402408 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_4363
timestamp 1586364061
transform 1 0 402500 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_4356
timestamp 1586364061
transform 1 0 401856 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_4368
timestamp 1586364061
transform 1 0 402960 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_4375
timestamp 1586364061
transform 1 0 403604 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_4387
timestamp 1586364061
transform 1 0 404708 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_4380
timestamp 1586364061
transform 1 0 404064 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_688
timestamp 1586364061
transform 1 0 405168 0 1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_4399
timestamp 1586364061
transform 1 0 405812 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_4393
timestamp 1586364061
transform 1 0 405260 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_4405
timestamp 1586364061
transform 1 0 406364 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_614
timestamp 1586364061
transform 1 0 408020 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_4411
timestamp 1586364061
transform 1 0 406916 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_4417
timestamp 1586364061
transform 1 0 407468 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_4424
timestamp 1586364061
transform 1 0 408112 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_4436
timestamp 1586364061
transform 1 0 409216 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_4429
timestamp 1586364061
transform 1 0 408572 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_4441
timestamp 1586364061
transform 1 0 409676 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_689
timestamp 1586364061
transform 1 0 410780 0 1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_4448
timestamp 1586364061
transform 1 0 410320 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_4454
timestamp 1586364061
transform 1 0 410872 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_4460
timestamp 1586364061
transform 1 0 411424 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_4472
timestamp 1586364061
transform 1 0 412528 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_4466
timestamp 1586364061
transform 1 0 411976 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_615
timestamp 1586364061
transform 1 0 413632 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_4485
timestamp 1586364061
transform 1 0 413724 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_4478
timestamp 1586364061
transform 1 0 413080 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_4490
timestamp 1586364061
transform 1 0 414184 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_4497
timestamp 1586364061
transform 1 0 414828 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_4509
timestamp 1586364061
transform 1 0 415932 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_4502
timestamp 1586364061
transform 1 0 415288 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_690
timestamp 1586364061
transform 1 0 416392 0 1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_4521
timestamp 1586364061
transform 1 0 417036 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_4515
timestamp 1586364061
transform 1 0 416484 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_4527
timestamp 1586364061
transform 1 0 417588 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_616
timestamp 1586364061
transform 1 0 419244 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_4533
timestamp 1586364061
transform 1 0 418140 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_4546
timestamp 1586364061
transform 1 0 419336 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_4539
timestamp 1586364061
transform 1 0 418692 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_4558
timestamp 1586364061
transform 1 0 420440 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_4551
timestamp 1586364061
transform 1 0 419796 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_4563
timestamp 1586364061
transform 1 0 420900 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_3  PHY_13
timestamp 1586364061
transform -1 0 422832 0 -1 5984
box -38 -48 314 592
use scs8hd_decap_3  PHY_15
timestamp 1586364061
transform -1 0 422832 0 1 5984
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_691
timestamp 1586364061
transform 1 0 422004 0 1 5984
box -38 -48 130 592
use scs8hd_decap_8  FILLER_6_4570
timestamp 1586364061
transform 1 0 421544 0 -1 5984
box -38 -48 774 592
use scs8hd_decap_3  FILLER_6_4578
timestamp 1586364061
transform 1 0 422280 0 -1 5984
box -38 -48 314 592
use scs8hd_decap_4  FILLER_7_4576
timestamp 1586364061
transform 1 0 422096 0 1 5984
box -38 -48 406 592
use scs8hd_fill_1  FILLER_7_4580
timestamp 1586364061
transform 1 0 422464 0 1 5984
box -38 -48 130 592
use scs8hd_decap_3  PHY_16
timestamp 1586364061
transform 1 0 1104 0 -1 7072
box -38 -48 314 592
use scs8hd_decap_12  FILLER_8_3
timestamp 1586364061
transform 1 0 1380 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_15
timestamp 1586364061
transform 1 0 2484 0 -1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_692
timestamp 1586364061
transform 1 0 3956 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_4  FILLER_8_27
timestamp 1586364061
transform 1 0 3588 0 -1 7072
box -38 -48 406 592
use scs8hd_decap_12  FILLER_8_32
timestamp 1586364061
transform 1 0 4048 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_44
timestamp 1586364061
transform 1 0 5152 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_56
timestamp 1586364061
transform 1 0 6256 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_68
timestamp 1586364061
transform 1 0 7360 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_80
timestamp 1586364061
transform 1 0 8464 0 -1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_693
timestamp 1586364061
transform 1 0 9568 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_8_93
timestamp 1586364061
transform 1 0 9660 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_105
timestamp 1586364061
transform 1 0 10764 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_117
timestamp 1586364061
transform 1 0 11868 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_129
timestamp 1586364061
transform 1 0 12972 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_141
timestamp 1586364061
transform 1 0 14076 0 -1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_694
timestamp 1586364061
transform 1 0 15180 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_8_154
timestamp 1586364061
transform 1 0 15272 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_166
timestamp 1586364061
transform 1 0 16376 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_178
timestamp 1586364061
transform 1 0 17480 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_190
timestamp 1586364061
transform 1 0 18584 0 -1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_695
timestamp 1586364061
transform 1 0 20792 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_8_202
timestamp 1586364061
transform 1 0 19688 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_215
timestamp 1586364061
transform 1 0 20884 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_227
timestamp 1586364061
transform 1 0 21988 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_239
timestamp 1586364061
transform 1 0 23092 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_251
timestamp 1586364061
transform 1 0 24196 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_263
timestamp 1586364061
transform 1 0 25300 0 -1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_696
timestamp 1586364061
transform 1 0 26404 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_8_276
timestamp 1586364061
transform 1 0 26496 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_288
timestamp 1586364061
transform 1 0 27600 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_300
timestamp 1586364061
transform 1 0 28704 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_312
timestamp 1586364061
transform 1 0 29808 0 -1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_697
timestamp 1586364061
transform 1 0 32016 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_8_324
timestamp 1586364061
transform 1 0 30912 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_337
timestamp 1586364061
transform 1 0 32108 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_349
timestamp 1586364061
transform 1 0 33212 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_361
timestamp 1586364061
transform 1 0 34316 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_373
timestamp 1586364061
transform 1 0 35420 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_385
timestamp 1586364061
transform 1 0 36524 0 -1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_698
timestamp 1586364061
transform 1 0 37628 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_8_398
timestamp 1586364061
transform 1 0 37720 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_410
timestamp 1586364061
transform 1 0 38824 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_422
timestamp 1586364061
transform 1 0 39928 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_434
timestamp 1586364061
transform 1 0 41032 0 -1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_699
timestamp 1586364061
transform 1 0 43240 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_8_446
timestamp 1586364061
transform 1 0 42136 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_459
timestamp 1586364061
transform 1 0 43332 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_471
timestamp 1586364061
transform 1 0 44436 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_483
timestamp 1586364061
transform 1 0 45540 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_495
timestamp 1586364061
transform 1 0 46644 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_507
timestamp 1586364061
transform 1 0 47748 0 -1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_700
timestamp 1586364061
transform 1 0 48852 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_8_520
timestamp 1586364061
transform 1 0 48944 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_532
timestamp 1586364061
transform 1 0 50048 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_544
timestamp 1586364061
transform 1 0 51152 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_556
timestamp 1586364061
transform 1 0 52256 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_568
timestamp 1586364061
transform 1 0 53360 0 -1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_701
timestamp 1586364061
transform 1 0 54464 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_8_581
timestamp 1586364061
transform 1 0 54556 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_593
timestamp 1586364061
transform 1 0 55660 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_605
timestamp 1586364061
transform 1 0 56764 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_617
timestamp 1586364061
transform 1 0 57868 0 -1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_702
timestamp 1586364061
transform 1 0 60076 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_8_629
timestamp 1586364061
transform 1 0 58972 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_642
timestamp 1586364061
transform 1 0 60168 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_654
timestamp 1586364061
transform 1 0 61272 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_666
timestamp 1586364061
transform 1 0 62376 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_678
timestamp 1586364061
transform 1 0 63480 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_690
timestamp 1586364061
transform 1 0 64584 0 -1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_703
timestamp 1586364061
transform 1 0 65688 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_8_703
timestamp 1586364061
transform 1 0 65780 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_715
timestamp 1586364061
transform 1 0 66884 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_727
timestamp 1586364061
transform 1 0 67988 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_739
timestamp 1586364061
transform 1 0 69092 0 -1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_704
timestamp 1586364061
transform 1 0 71300 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_8_751
timestamp 1586364061
transform 1 0 70196 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_764
timestamp 1586364061
transform 1 0 71392 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_776
timestamp 1586364061
transform 1 0 72496 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_788
timestamp 1586364061
transform 1 0 73600 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_800
timestamp 1586364061
transform 1 0 74704 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_812
timestamp 1586364061
transform 1 0 75808 0 -1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_705
timestamp 1586364061
transform 1 0 76912 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_8_825
timestamp 1586364061
transform 1 0 77004 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_837
timestamp 1586364061
transform 1 0 78108 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_849
timestamp 1586364061
transform 1 0 79212 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_861
timestamp 1586364061
transform 1 0 80316 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_873
timestamp 1586364061
transform 1 0 81420 0 -1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_706
timestamp 1586364061
transform 1 0 82524 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_8_886
timestamp 1586364061
transform 1 0 82616 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_898
timestamp 1586364061
transform 1 0 83720 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_910
timestamp 1586364061
transform 1 0 84824 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_922
timestamp 1586364061
transform 1 0 85928 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_934
timestamp 1586364061
transform 1 0 87032 0 -1 7072
box -38 -48 1142 592
use scs8hd_ebufn_1  logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer
timestamp 1586364061
transform 1 0 88228 0 -1 7072
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_707
timestamp 1586364061
transform 1 0 88136 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_8_955
timestamp 1586364061
transform 1 0 88964 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_967
timestamp 1586364061
transform 1 0 90068 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_979
timestamp 1586364061
transform 1 0 91172 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_991
timestamp 1586364061
transform 1 0 92276 0 -1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_708
timestamp 1586364061
transform 1 0 93748 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_4  FILLER_8_1003
timestamp 1586364061
transform 1 0 93380 0 -1 7072
box -38 -48 406 592
use scs8hd_decap_12  FILLER_8_1008
timestamp 1586364061
transform 1 0 93840 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_1020
timestamp 1586364061
transform 1 0 94944 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_1032
timestamp 1586364061
transform 1 0 96048 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_1044
timestamp 1586364061
transform 1 0 97152 0 -1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_709
timestamp 1586364061
transform 1 0 99360 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_8_1056
timestamp 1586364061
transform 1 0 98256 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_1069
timestamp 1586364061
transform 1 0 99452 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_1081
timestamp 1586364061
transform 1 0 100556 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_1093
timestamp 1586364061
transform 1 0 101660 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_1105
timestamp 1586364061
transform 1 0 102764 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_1117
timestamp 1586364061
transform 1 0 103868 0 -1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_710
timestamp 1586364061
transform 1 0 104972 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_8_1130
timestamp 1586364061
transform 1 0 105064 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_1142
timestamp 1586364061
transform 1 0 106168 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_1154
timestamp 1586364061
transform 1 0 107272 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_1166
timestamp 1586364061
transform 1 0 108376 0 -1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_711
timestamp 1586364061
transform 1 0 110584 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_8_1178
timestamp 1586364061
transform 1 0 109480 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_1191
timestamp 1586364061
transform 1 0 110676 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_1203
timestamp 1586364061
transform 1 0 111780 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_1215
timestamp 1586364061
transform 1 0 112884 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_1227
timestamp 1586364061
transform 1 0 113988 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_1239
timestamp 1586364061
transform 1 0 115092 0 -1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_712
timestamp 1586364061
transform 1 0 116196 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_8_1252
timestamp 1586364061
transform 1 0 116288 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_1264
timestamp 1586364061
transform 1 0 117392 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_1276
timestamp 1586364061
transform 1 0 118496 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_1288
timestamp 1586364061
transform 1 0 119600 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_1300
timestamp 1586364061
transform 1 0 120704 0 -1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_713
timestamp 1586364061
transform 1 0 121808 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_8_1313
timestamp 1586364061
transform 1 0 121900 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_1325
timestamp 1586364061
transform 1 0 123004 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_1337
timestamp 1586364061
transform 1 0 124108 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_1349
timestamp 1586364061
transform 1 0 125212 0 -1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_714
timestamp 1586364061
transform 1 0 127420 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_8_1361
timestamp 1586364061
transform 1 0 126316 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_1374
timestamp 1586364061
transform 1 0 127512 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_1386
timestamp 1586364061
transform 1 0 128616 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_1398
timestamp 1586364061
transform 1 0 129720 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_1410
timestamp 1586364061
transform 1 0 130824 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_1422
timestamp 1586364061
transform 1 0 131928 0 -1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_715
timestamp 1586364061
transform 1 0 133032 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_8_1435
timestamp 1586364061
transform 1 0 133124 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_1447
timestamp 1586364061
transform 1 0 134228 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_1459
timestamp 1586364061
transform 1 0 135332 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_1471
timestamp 1586364061
transform 1 0 136436 0 -1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_716
timestamp 1586364061
transform 1 0 138644 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_8_1483
timestamp 1586364061
transform 1 0 137540 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_1496
timestamp 1586364061
transform 1 0 138736 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_1508
timestamp 1586364061
transform 1 0 139840 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_1520
timestamp 1586364061
transform 1 0 140944 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_1532
timestamp 1586364061
transform 1 0 142048 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_1544
timestamp 1586364061
transform 1 0 143152 0 -1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_717
timestamp 1586364061
transform 1 0 144256 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_8_1557
timestamp 1586364061
transform 1 0 144348 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_1569
timestamp 1586364061
transform 1 0 145452 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_1581
timestamp 1586364061
transform 1 0 146556 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_1593
timestamp 1586364061
transform 1 0 147660 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_1605
timestamp 1586364061
transform 1 0 148764 0 -1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_718
timestamp 1586364061
transform 1 0 149868 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_8_1618
timestamp 1586364061
transform 1 0 149960 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_1630
timestamp 1586364061
transform 1 0 151064 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_1642
timestamp 1586364061
transform 1 0 152168 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_1654
timestamp 1586364061
transform 1 0 153272 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_1666
timestamp 1586364061
transform 1 0 154376 0 -1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_719
timestamp 1586364061
transform 1 0 155480 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_8_1679
timestamp 1586364061
transform 1 0 155572 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_1691
timestamp 1586364061
transform 1 0 156676 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_1703
timestamp 1586364061
transform 1 0 157780 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_1715
timestamp 1586364061
transform 1 0 158884 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_1727
timestamp 1586364061
transform 1 0 159988 0 -1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_720
timestamp 1586364061
transform 1 0 161092 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_8_1740
timestamp 1586364061
transform 1 0 161184 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_1752
timestamp 1586364061
transform 1 0 162288 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_1764
timestamp 1586364061
transform 1 0 163392 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_1776
timestamp 1586364061
transform 1 0 164496 0 -1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_721
timestamp 1586364061
transform 1 0 166704 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_8_1788
timestamp 1586364061
transform 1 0 165600 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_1801
timestamp 1586364061
transform 1 0 166796 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_1813
timestamp 1586364061
transform 1 0 167900 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_1825
timestamp 1586364061
transform 1 0 169004 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_8_1837
timestamp 1586364061
transform 1 0 170108 0 -1 7072
box -38 -48 406 592
use scs8hd_buf_2  _20_
timestamp 1586364061
transform 1 0 170568 0 -1 7072
box -38 -48 406 592
use scs8hd_fill_1  FILLER_8_1841
timestamp 1586364061
transform 1 0 170476 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_8_1846
timestamp 1586364061
transform 1 0 170936 0 -1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_722
timestamp 1586364061
transform 1 0 172316 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_3  FILLER_8_1858
timestamp 1586364061
transform 1 0 172040 0 -1 7072
box -38 -48 314 592
use scs8hd_decap_12  FILLER_8_1862
timestamp 1586364061
transform 1 0 172408 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_1874
timestamp 1586364061
transform 1 0 173512 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_1886
timestamp 1586364061
transform 1 0 174616 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_1898
timestamp 1586364061
transform 1 0 175720 0 -1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_723
timestamp 1586364061
transform 1 0 177928 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_8_1910
timestamp 1586364061
transform 1 0 176824 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_1923
timestamp 1586364061
transform 1 0 178020 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_1935
timestamp 1586364061
transform 1 0 179124 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_1947
timestamp 1586364061
transform 1 0 180228 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_1959
timestamp 1586364061
transform 1 0 181332 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_1971
timestamp 1586364061
transform 1 0 182436 0 -1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_724
timestamp 1586364061
transform 1 0 183540 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_8_1984
timestamp 1586364061
transform 1 0 183632 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_1996
timestamp 1586364061
transform 1 0 184736 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_2008
timestamp 1586364061
transform 1 0 185840 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_2020
timestamp 1586364061
transform 1 0 186944 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_2032
timestamp 1586364061
transform 1 0 188048 0 -1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_725
timestamp 1586364061
transform 1 0 189152 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_8_2045
timestamp 1586364061
transform 1 0 189244 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_2057
timestamp 1586364061
transform 1 0 190348 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_2069
timestamp 1586364061
transform 1 0 191452 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_2081
timestamp 1586364061
transform 1 0 192556 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_2093
timestamp 1586364061
transform 1 0 193660 0 -1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_726
timestamp 1586364061
transform 1 0 194764 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_8_2106
timestamp 1586364061
transform 1 0 194856 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_2118
timestamp 1586364061
transform 1 0 195960 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_2130
timestamp 1586364061
transform 1 0 197064 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_2142
timestamp 1586364061
transform 1 0 198168 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_2154
timestamp 1586364061
transform 1 0 199272 0 -1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_727
timestamp 1586364061
transform 1 0 200376 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_8_2167
timestamp 1586364061
transform 1 0 200468 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_2179
timestamp 1586364061
transform 1 0 201572 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_2191
timestamp 1586364061
transform 1 0 202676 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_2203
timestamp 1586364061
transform 1 0 203780 0 -1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_728
timestamp 1586364061
transform 1 0 205988 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_8_2215
timestamp 1586364061
transform 1 0 204884 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_2228
timestamp 1586364061
transform 1 0 206080 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_2240
timestamp 1586364061
transform 1 0 207184 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_2252
timestamp 1586364061
transform 1 0 208288 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_2264
timestamp 1586364061
transform 1 0 209392 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_2276
timestamp 1586364061
transform 1 0 210496 0 -1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_729
timestamp 1586364061
transform 1 0 211600 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_8_2289
timestamp 1586364061
transform 1 0 211692 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_2301
timestamp 1586364061
transform 1 0 212796 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_2313
timestamp 1586364061
transform 1 0 213900 0 -1 7072
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA_logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer_TEB
timestamp 1586364061
transform 1 0 215556 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_6  FILLER_8_2325
timestamp 1586364061
transform 1 0 215004 0 -1 7072
box -38 -48 590 592
use scs8hd_decap_12  FILLER_8_2333
timestamp 1586364061
transform 1 0 215740 0 -1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_730
timestamp 1586364061
transform 1 0 217212 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_4  FILLER_8_2345
timestamp 1586364061
transform 1 0 216844 0 -1 7072
box -38 -48 406 592
use scs8hd_decap_12  FILLER_8_2350
timestamp 1586364061
transform 1 0 217304 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_2362
timestamp 1586364061
transform 1 0 218408 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_2374
timestamp 1586364061
transform 1 0 219512 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_2386
timestamp 1586364061
transform 1 0 220616 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_2398
timestamp 1586364061
transform 1 0 221720 0 -1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_731
timestamp 1586364061
transform 1 0 222824 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_8_2411
timestamp 1586364061
transform 1 0 222916 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_2423
timestamp 1586364061
transform 1 0 224020 0 -1 7072
box -38 -48 1142 592
use scs8hd_ebufn_1  logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer
timestamp 1586364061
transform 1 0 225308 0 -1 7072
box -38 -48 774 592
use scs8hd_fill_2  FILLER_8_2435
timestamp 1586364061
transform 1 0 225124 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_12  FILLER_8_2445
timestamp 1586364061
transform 1 0 226044 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_2457
timestamp 1586364061
transform 1 0 227148 0 -1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_732
timestamp 1586364061
transform 1 0 228436 0 -1 7072
box -38 -48 130 592
use scs8hd_fill_2  FILLER_8_2469
timestamp 1586364061
transform 1 0 228252 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_12  FILLER_8_2472
timestamp 1586364061
transform 1 0 228528 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_2484
timestamp 1586364061
transform 1 0 229632 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_2496
timestamp 1586364061
transform 1 0 230736 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_2508
timestamp 1586364061
transform 1 0 231840 0 -1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_733
timestamp 1586364061
transform 1 0 234048 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_8_2520
timestamp 1586364061
transform 1 0 232944 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_2533
timestamp 1586364061
transform 1 0 234140 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_2545
timestamp 1586364061
transform 1 0 235244 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_2557
timestamp 1586364061
transform 1 0 236348 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_2569
timestamp 1586364061
transform 1 0 237452 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_2581
timestamp 1586364061
transform 1 0 238556 0 -1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_734
timestamp 1586364061
transform 1 0 239660 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_8_2594
timestamp 1586364061
transform 1 0 239752 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_2606
timestamp 1586364061
transform 1 0 240856 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_2618
timestamp 1586364061
transform 1 0 241960 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_2630
timestamp 1586364061
transform 1 0 243064 0 -1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_735
timestamp 1586364061
transform 1 0 245272 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_8_2642
timestamp 1586364061
transform 1 0 244168 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_2655
timestamp 1586364061
transform 1 0 245364 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_2667
timestamp 1586364061
transform 1 0 246468 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_2679
timestamp 1586364061
transform 1 0 247572 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_2691
timestamp 1586364061
transform 1 0 248676 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_2703
timestamp 1586364061
transform 1 0 249780 0 -1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_736
timestamp 1586364061
transform 1 0 250884 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_8_2716
timestamp 1586364061
transform 1 0 250976 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_2728
timestamp 1586364061
transform 1 0 252080 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_2740
timestamp 1586364061
transform 1 0 253184 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_2752
timestamp 1586364061
transform 1 0 254288 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_2764
timestamp 1586364061
transform 1 0 255392 0 -1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_737
timestamp 1586364061
transform 1 0 256496 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_8_2777
timestamp 1586364061
transform 1 0 256588 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_2789
timestamp 1586364061
transform 1 0 257692 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_2801
timestamp 1586364061
transform 1 0 258796 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_2813
timestamp 1586364061
transform 1 0 259900 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_2825
timestamp 1586364061
transform 1 0 261004 0 -1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_738
timestamp 1586364061
transform 1 0 262108 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_8_2838
timestamp 1586364061
transform 1 0 262200 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_2850
timestamp 1586364061
transform 1 0 263304 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_2862
timestamp 1586364061
transform 1 0 264408 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_2874
timestamp 1586364061
transform 1 0 265512 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_2886
timestamp 1586364061
transform 1 0 266616 0 -1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_739
timestamp 1586364061
transform 1 0 267720 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_8_2899
timestamp 1586364061
transform 1 0 267812 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_2911
timestamp 1586364061
transform 1 0 268916 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_2923
timestamp 1586364061
transform 1 0 270020 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_2935
timestamp 1586364061
transform 1 0 271124 0 -1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_740
timestamp 1586364061
transform 1 0 273332 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_8_2947
timestamp 1586364061
transform 1 0 272228 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_2960
timestamp 1586364061
transform 1 0 273424 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_2972
timestamp 1586364061
transform 1 0 274528 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_2984
timestamp 1586364061
transform 1 0 275632 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_2996
timestamp 1586364061
transform 1 0 276736 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_3008
timestamp 1586364061
transform 1 0 277840 0 -1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_741
timestamp 1586364061
transform 1 0 278944 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_8_3021
timestamp 1586364061
transform 1 0 279036 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_3033
timestamp 1586364061
transform 1 0 280140 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_3045
timestamp 1586364061
transform 1 0 281244 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_3057
timestamp 1586364061
transform 1 0 282348 0 -1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_742
timestamp 1586364061
transform 1 0 284556 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_8_3069
timestamp 1586364061
transform 1 0 283452 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_3082
timestamp 1586364061
transform 1 0 284648 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_3094
timestamp 1586364061
transform 1 0 285752 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_3106
timestamp 1586364061
transform 1 0 286856 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_3118
timestamp 1586364061
transform 1 0 287960 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_3130
timestamp 1586364061
transform 1 0 289064 0 -1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_743
timestamp 1586364061
transform 1 0 290168 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_8_3143
timestamp 1586364061
transform 1 0 290260 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_3155
timestamp 1586364061
transform 1 0 291364 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_3167
timestamp 1586364061
transform 1 0 292468 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_3179
timestamp 1586364061
transform 1 0 293572 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_3191
timestamp 1586364061
transform 1 0 294676 0 -1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_744
timestamp 1586364061
transform 1 0 295780 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_8_3204
timestamp 1586364061
transform 1 0 295872 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_3216
timestamp 1586364061
transform 1 0 296976 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_3228
timestamp 1586364061
transform 1 0 298080 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_3240
timestamp 1586364061
transform 1 0 299184 0 -1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_745
timestamp 1586364061
transform 1 0 301392 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_8_3252
timestamp 1586364061
transform 1 0 300288 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_3265
timestamp 1586364061
transform 1 0 301484 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_3277
timestamp 1586364061
transform 1 0 302588 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_3289
timestamp 1586364061
transform 1 0 303692 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_3301
timestamp 1586364061
transform 1 0 304796 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_3313
timestamp 1586364061
transform 1 0 305900 0 -1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_746
timestamp 1586364061
transform 1 0 307004 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_8_3326
timestamp 1586364061
transform 1 0 307096 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_3338
timestamp 1586364061
transform 1 0 308200 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_3350
timestamp 1586364061
transform 1 0 309304 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_3362
timestamp 1586364061
transform 1 0 310408 0 -1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_747
timestamp 1586364061
transform 1 0 312616 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_8_3374
timestamp 1586364061
transform 1 0 311512 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_3387
timestamp 1586364061
transform 1 0 312708 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_3399
timestamp 1586364061
transform 1 0 313812 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_3411
timestamp 1586364061
transform 1 0 314916 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_3423
timestamp 1586364061
transform 1 0 316020 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_3435
timestamp 1586364061
transform 1 0 317124 0 -1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_748
timestamp 1586364061
transform 1 0 318228 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_8_3448
timestamp 1586364061
transform 1 0 318320 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_3460
timestamp 1586364061
transform 1 0 319424 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_3472
timestamp 1586364061
transform 1 0 320528 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_3484
timestamp 1586364061
transform 1 0 321632 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_3496
timestamp 1586364061
transform 1 0 322736 0 -1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_749
timestamp 1586364061
transform 1 0 323840 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_8_3509
timestamp 1586364061
transform 1 0 323932 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_3521
timestamp 1586364061
transform 1 0 325036 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_3533
timestamp 1586364061
transform 1 0 326140 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_3545
timestamp 1586364061
transform 1 0 327244 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_3557
timestamp 1586364061
transform 1 0 328348 0 -1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_750
timestamp 1586364061
transform 1 0 329452 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_8_3570
timestamp 1586364061
transform 1 0 329544 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_3582
timestamp 1586364061
transform 1 0 330648 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_3594
timestamp 1586364061
transform 1 0 331752 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_3606
timestamp 1586364061
transform 1 0 332856 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_3618
timestamp 1586364061
transform 1 0 333960 0 -1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_751
timestamp 1586364061
transform 1 0 335064 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_8_3631
timestamp 1586364061
transform 1 0 335156 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_3643
timestamp 1586364061
transform 1 0 336260 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_3655
timestamp 1586364061
transform 1 0 337364 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_3667
timestamp 1586364061
transform 1 0 338468 0 -1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_752
timestamp 1586364061
transform 1 0 340676 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_8_3679
timestamp 1586364061
transform 1 0 339572 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_3692
timestamp 1586364061
transform 1 0 340768 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_3704
timestamp 1586364061
transform 1 0 341872 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_3716
timestamp 1586364061
transform 1 0 342976 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_3728
timestamp 1586364061
transform 1 0 344080 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_3740
timestamp 1586364061
transform 1 0 345184 0 -1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_753
timestamp 1586364061
transform 1 0 346288 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_8_3753
timestamp 1586364061
transform 1 0 346380 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_3765
timestamp 1586364061
transform 1 0 347484 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_3777
timestamp 1586364061
transform 1 0 348588 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_3789
timestamp 1586364061
transform 1 0 349692 0 -1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_754
timestamp 1586364061
transform 1 0 351900 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_8_3801
timestamp 1586364061
transform 1 0 350796 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_3814
timestamp 1586364061
transform 1 0 351992 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_3826
timestamp 1586364061
transform 1 0 353096 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_3838
timestamp 1586364061
transform 1 0 354200 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_3850
timestamp 1586364061
transform 1 0 355304 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_3862
timestamp 1586364061
transform 1 0 356408 0 -1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_755
timestamp 1586364061
transform 1 0 357512 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_8_3875
timestamp 1586364061
transform 1 0 357604 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_3887
timestamp 1586364061
transform 1 0 358708 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_3899
timestamp 1586364061
transform 1 0 359812 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_3911
timestamp 1586364061
transform 1 0 360916 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_3923
timestamp 1586364061
transform 1 0 362020 0 -1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_756
timestamp 1586364061
transform 1 0 363124 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_8_3936
timestamp 1586364061
transform 1 0 363216 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_3948
timestamp 1586364061
transform 1 0 364320 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_3960
timestamp 1586364061
transform 1 0 365424 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_3972
timestamp 1586364061
transform 1 0 366528 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_3984
timestamp 1586364061
transform 1 0 367632 0 -1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_757
timestamp 1586364061
transform 1 0 368736 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_8_3997
timestamp 1586364061
transform 1 0 368828 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_4009
timestamp 1586364061
transform 1 0 369932 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_4021
timestamp 1586364061
transform 1 0 371036 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_4033
timestamp 1586364061
transform 1 0 372140 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_4045
timestamp 1586364061
transform 1 0 373244 0 -1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_758
timestamp 1586364061
transform 1 0 374348 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_8_4058
timestamp 1586364061
transform 1 0 374440 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_4070
timestamp 1586364061
transform 1 0 375544 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_4082
timestamp 1586364061
transform 1 0 376648 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_4094
timestamp 1586364061
transform 1 0 377752 0 -1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_759
timestamp 1586364061
transform 1 0 379960 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_8_4106
timestamp 1586364061
transform 1 0 378856 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_4119
timestamp 1586364061
transform 1 0 380052 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_4131
timestamp 1586364061
transform 1 0 381156 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_4143
timestamp 1586364061
transform 1 0 382260 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_4155
timestamp 1586364061
transform 1 0 383364 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_4167
timestamp 1586364061
transform 1 0 384468 0 -1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_760
timestamp 1586364061
transform 1 0 385572 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_8_4180
timestamp 1586364061
transform 1 0 385664 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_4192
timestamp 1586364061
transform 1 0 386768 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_4204
timestamp 1586364061
transform 1 0 387872 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_4216
timestamp 1586364061
transform 1 0 388976 0 -1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_761
timestamp 1586364061
transform 1 0 391184 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_8_4228
timestamp 1586364061
transform 1 0 390080 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_4241
timestamp 1586364061
transform 1 0 391276 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_4253
timestamp 1586364061
transform 1 0 392380 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_4265
timestamp 1586364061
transform 1 0 393484 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_4277
timestamp 1586364061
transform 1 0 394588 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_4289
timestamp 1586364061
transform 1 0 395692 0 -1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_762
timestamp 1586364061
transform 1 0 396796 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_8_4302
timestamp 1586364061
transform 1 0 396888 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_4314
timestamp 1586364061
transform 1 0 397992 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_4326
timestamp 1586364061
transform 1 0 399096 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_4338
timestamp 1586364061
transform 1 0 400200 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_4350
timestamp 1586364061
transform 1 0 401304 0 -1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_763
timestamp 1586364061
transform 1 0 402408 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_8_4363
timestamp 1586364061
transform 1 0 402500 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_4375
timestamp 1586364061
transform 1 0 403604 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_4387
timestamp 1586364061
transform 1 0 404708 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_4399
timestamp 1586364061
transform 1 0 405812 0 -1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_764
timestamp 1586364061
transform 1 0 408020 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_8_4411
timestamp 1586364061
transform 1 0 406916 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_4424
timestamp 1586364061
transform 1 0 408112 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_4436
timestamp 1586364061
transform 1 0 409216 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_4448
timestamp 1586364061
transform 1 0 410320 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_4460
timestamp 1586364061
transform 1 0 411424 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_4472
timestamp 1586364061
transform 1 0 412528 0 -1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_765
timestamp 1586364061
transform 1 0 413632 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_8_4485
timestamp 1586364061
transform 1 0 413724 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_4497
timestamp 1586364061
transform 1 0 414828 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_4509
timestamp 1586364061
transform 1 0 415932 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_4521
timestamp 1586364061
transform 1 0 417036 0 -1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_766
timestamp 1586364061
transform 1 0 419244 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_8_4533
timestamp 1586364061
transform 1 0 418140 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_4546
timestamp 1586364061
transform 1 0 419336 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_4558
timestamp 1586364061
transform 1 0 420440 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_3  PHY_17
timestamp 1586364061
transform -1 0 422832 0 -1 7072
box -38 -48 314 592
use scs8hd_decap_8  FILLER_8_4570
timestamp 1586364061
transform 1 0 421544 0 -1 7072
box -38 -48 774 592
use scs8hd_decap_3  FILLER_8_4578
timestamp 1586364061
transform 1 0 422280 0 -1 7072
box -38 -48 314 592
use scs8hd_decap_3  PHY_18
timestamp 1586364061
transform 1 0 1104 0 1 7072
box -38 -48 314 592
use scs8hd_decap_12  FILLER_9_3
timestamp 1586364061
transform 1 0 1380 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_15
timestamp 1586364061
transform 1 0 2484 0 1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_767
timestamp 1586364061
transform 1 0 3956 0 1 7072
box -38 -48 130 592
use scs8hd_decap_4  FILLER_9_27
timestamp 1586364061
transform 1 0 3588 0 1 7072
box -38 -48 406 592
use scs8hd_decap_12  FILLER_9_32
timestamp 1586364061
transform 1 0 4048 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_44
timestamp 1586364061
transform 1 0 5152 0 1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_768
timestamp 1586364061
transform 1 0 6808 0 1 7072
box -38 -48 130 592
use scs8hd_decap_6  FILLER_9_56
timestamp 1586364061
transform 1 0 6256 0 1 7072
box -38 -48 590 592
use scs8hd_decap_12  FILLER_9_63
timestamp 1586364061
transform 1 0 6900 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_75
timestamp 1586364061
transform 1 0 8004 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_9_87
timestamp 1586364061
transform 1 0 9108 0 1 7072
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_769
timestamp 1586364061
transform 1 0 9660 0 1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_9_94
timestamp 1586364061
transform 1 0 9752 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_106
timestamp 1586364061
transform 1 0 10856 0 1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_770
timestamp 1586364061
transform 1 0 12512 0 1 7072
box -38 -48 130 592
use scs8hd_decap_6  FILLER_9_118
timestamp 1586364061
transform 1 0 11960 0 1 7072
box -38 -48 590 592
use scs8hd_decap_12  FILLER_9_125
timestamp 1586364061
transform 1 0 12604 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_137
timestamp 1586364061
transform 1 0 13708 0 1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_771
timestamp 1586364061
transform 1 0 15364 0 1 7072
box -38 -48 130 592
use scs8hd_decap_6  FILLER_9_149
timestamp 1586364061
transform 1 0 14812 0 1 7072
box -38 -48 590 592
use scs8hd_decap_12  FILLER_9_156
timestamp 1586364061
transform 1 0 15456 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_168
timestamp 1586364061
transform 1 0 16560 0 1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_772
timestamp 1586364061
transform 1 0 18216 0 1 7072
box -38 -48 130 592
use scs8hd_decap_6  FILLER_9_180
timestamp 1586364061
transform 1 0 17664 0 1 7072
box -38 -48 590 592
use scs8hd_decap_12  FILLER_9_187
timestamp 1586364061
transform 1 0 18308 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_199
timestamp 1586364061
transform 1 0 19412 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_9_211
timestamp 1586364061
transform 1 0 20516 0 1 7072
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_773
timestamp 1586364061
transform 1 0 21068 0 1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_9_218
timestamp 1586364061
transform 1 0 21160 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_230
timestamp 1586364061
transform 1 0 22264 0 1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_774
timestamp 1586364061
transform 1 0 23920 0 1 7072
box -38 -48 130 592
use scs8hd_decap_6  FILLER_9_242
timestamp 1586364061
transform 1 0 23368 0 1 7072
box -38 -48 590 592
use scs8hd_decap_12  FILLER_9_249
timestamp 1586364061
transform 1 0 24012 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_261
timestamp 1586364061
transform 1 0 25116 0 1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_775
timestamp 1586364061
transform 1 0 26772 0 1 7072
box -38 -48 130 592
use scs8hd_decap_6  FILLER_9_273
timestamp 1586364061
transform 1 0 26220 0 1 7072
box -38 -48 590 592
use scs8hd_decap_12  FILLER_9_280
timestamp 1586364061
transform 1 0 26864 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_292
timestamp 1586364061
transform 1 0 27968 0 1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_776
timestamp 1586364061
transform 1 0 29624 0 1 7072
box -38 -48 130 592
use scs8hd_decap_6  FILLER_9_304
timestamp 1586364061
transform 1 0 29072 0 1 7072
box -38 -48 590 592
use scs8hd_decap_12  FILLER_9_311
timestamp 1586364061
transform 1 0 29716 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_323
timestamp 1586364061
transform 1 0 30820 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_9_335
timestamp 1586364061
transform 1 0 31924 0 1 7072
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_777
timestamp 1586364061
transform 1 0 32476 0 1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_9_342
timestamp 1586364061
transform 1 0 32568 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_354
timestamp 1586364061
transform 1 0 33672 0 1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_778
timestamp 1586364061
transform 1 0 35328 0 1 7072
box -38 -48 130 592
use scs8hd_decap_6  FILLER_9_366
timestamp 1586364061
transform 1 0 34776 0 1 7072
box -38 -48 590 592
use scs8hd_decap_12  FILLER_9_373
timestamp 1586364061
transform 1 0 35420 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_385
timestamp 1586364061
transform 1 0 36524 0 1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_779
timestamp 1586364061
transform 1 0 38180 0 1 7072
box -38 -48 130 592
use scs8hd_decap_6  FILLER_9_397
timestamp 1586364061
transform 1 0 37628 0 1 7072
box -38 -48 590 592
use scs8hd_decap_12  FILLER_9_404
timestamp 1586364061
transform 1 0 38272 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_416
timestamp 1586364061
transform 1 0 39376 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_9_428
timestamp 1586364061
transform 1 0 40480 0 1 7072
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_780
timestamp 1586364061
transform 1 0 41032 0 1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_9_435
timestamp 1586364061
transform 1 0 41124 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_447
timestamp 1586364061
transform 1 0 42228 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_9_459
timestamp 1586364061
transform 1 0 43332 0 1 7072
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_781
timestamp 1586364061
transform 1 0 43884 0 1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_9_466
timestamp 1586364061
transform 1 0 43976 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_478
timestamp 1586364061
transform 1 0 45080 0 1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_782
timestamp 1586364061
transform 1 0 46736 0 1 7072
box -38 -48 130 592
use scs8hd_decap_6  FILLER_9_490
timestamp 1586364061
transform 1 0 46184 0 1 7072
box -38 -48 590 592
use scs8hd_decap_12  FILLER_9_497
timestamp 1586364061
transform 1 0 46828 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_509
timestamp 1586364061
transform 1 0 47932 0 1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_783
timestamp 1586364061
transform 1 0 49588 0 1 7072
box -38 -48 130 592
use scs8hd_decap_6  FILLER_9_521
timestamp 1586364061
transform 1 0 49036 0 1 7072
box -38 -48 590 592
use scs8hd_decap_12  FILLER_9_528
timestamp 1586364061
transform 1 0 49680 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_540
timestamp 1586364061
transform 1 0 50784 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_9_552
timestamp 1586364061
transform 1 0 51888 0 1 7072
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_784
timestamp 1586364061
transform 1 0 52440 0 1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_9_559
timestamp 1586364061
transform 1 0 52532 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_571
timestamp 1586364061
transform 1 0 53636 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_9_583
timestamp 1586364061
transform 1 0 54740 0 1 7072
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_785
timestamp 1586364061
transform 1 0 55292 0 1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_9_590
timestamp 1586364061
transform 1 0 55384 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_602
timestamp 1586364061
transform 1 0 56488 0 1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_786
timestamp 1586364061
transform 1 0 58144 0 1 7072
box -38 -48 130 592
use scs8hd_decap_6  FILLER_9_614
timestamp 1586364061
transform 1 0 57592 0 1 7072
box -38 -48 590 592
use scs8hd_decap_12  FILLER_9_621
timestamp 1586364061
transform 1 0 58236 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_633
timestamp 1586364061
transform 1 0 59340 0 1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_787
timestamp 1586364061
transform 1 0 60996 0 1 7072
box -38 -48 130 592
use scs8hd_decap_6  FILLER_9_645
timestamp 1586364061
transform 1 0 60444 0 1 7072
box -38 -48 590 592
use scs8hd_decap_12  FILLER_9_652
timestamp 1586364061
transform 1 0 61088 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_664
timestamp 1586364061
transform 1 0 62192 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_9_676
timestamp 1586364061
transform 1 0 63296 0 1 7072
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_788
timestamp 1586364061
transform 1 0 63848 0 1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_9_683
timestamp 1586364061
transform 1 0 63940 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_695
timestamp 1586364061
transform 1 0 65044 0 1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_789
timestamp 1586364061
transform 1 0 66700 0 1 7072
box -38 -48 130 592
use scs8hd_decap_6  FILLER_9_707
timestamp 1586364061
transform 1 0 66148 0 1 7072
box -38 -48 590 592
use scs8hd_decap_12  FILLER_9_714
timestamp 1586364061
transform 1 0 66792 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_726
timestamp 1586364061
transform 1 0 67896 0 1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_790
timestamp 1586364061
transform 1 0 69552 0 1 7072
box -38 -48 130 592
use scs8hd_decap_6  FILLER_9_738
timestamp 1586364061
transform 1 0 69000 0 1 7072
box -38 -48 590 592
use scs8hd_decap_12  FILLER_9_745
timestamp 1586364061
transform 1 0 69644 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_757
timestamp 1586364061
transform 1 0 70748 0 1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_791
timestamp 1586364061
transform 1 0 72404 0 1 7072
box -38 -48 130 592
use scs8hd_decap_6  FILLER_9_769
timestamp 1586364061
transform 1 0 71852 0 1 7072
box -38 -48 590 592
use scs8hd_decap_12  FILLER_9_776
timestamp 1586364061
transform 1 0 72496 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_788
timestamp 1586364061
transform 1 0 73600 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_9_800
timestamp 1586364061
transform 1 0 74704 0 1 7072
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_792
timestamp 1586364061
transform 1 0 75256 0 1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_9_807
timestamp 1586364061
transform 1 0 75348 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_819
timestamp 1586364061
transform 1 0 76452 0 1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_793
timestamp 1586364061
transform 1 0 78108 0 1 7072
box -38 -48 130 592
use scs8hd_decap_6  FILLER_9_831
timestamp 1586364061
transform 1 0 77556 0 1 7072
box -38 -48 590 592
use scs8hd_decap_12  FILLER_9_838
timestamp 1586364061
transform 1 0 78200 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_850
timestamp 1586364061
transform 1 0 79304 0 1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_794
timestamp 1586364061
transform 1 0 80960 0 1 7072
box -38 -48 130 592
use scs8hd_decap_6  FILLER_9_862
timestamp 1586364061
transform 1 0 80408 0 1 7072
box -38 -48 590 592
use scs8hd_decap_12  FILLER_9_869
timestamp 1586364061
transform 1 0 81052 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_881
timestamp 1586364061
transform 1 0 82156 0 1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_795
timestamp 1586364061
transform 1 0 83812 0 1 7072
box -38 -48 130 592
use scs8hd_decap_6  FILLER_9_893
timestamp 1586364061
transform 1 0 83260 0 1 7072
box -38 -48 590 592
use scs8hd_decap_12  FILLER_9_900
timestamp 1586364061
transform 1 0 83904 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_912
timestamp 1586364061
transform 1 0 85008 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_9_924
timestamp 1586364061
transform 1 0 86112 0 1 7072
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_796
timestamp 1586364061
transform 1 0 86664 0 1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_9_931
timestamp 1586364061
transform 1 0 86756 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_943
timestamp 1586364061
transform 1 0 87860 0 1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_797
timestamp 1586364061
transform 1 0 89516 0 1 7072
box -38 -48 130 592
use scs8hd_decap_6  FILLER_9_955
timestamp 1586364061
transform 1 0 88964 0 1 7072
box -38 -48 590 592
use scs8hd_decap_12  FILLER_9_962
timestamp 1586364061
transform 1 0 89608 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_974
timestamp 1586364061
transform 1 0 90712 0 1 7072
box -38 -48 1142 592
use scs8hd_buf_2  _19_
timestamp 1586364061
transform 1 0 92736 0 1 7072
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_798
timestamp 1586364061
transform 1 0 92368 0 1 7072
box -38 -48 130 592
use scs8hd_decap_6  FILLER_9_986
timestamp 1586364061
transform 1 0 91816 0 1 7072
box -38 -48 590 592
use scs8hd_decap_3  FILLER_9_993
timestamp 1586364061
transform 1 0 92460 0 1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__19__A
timestamp 1586364061
transform 1 0 93288 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_1000
timestamp 1586364061
transform 1 0 93104 0 1 7072
box -38 -48 222 592
use scs8hd_decap_12  FILLER_9_1004
timestamp 1586364061
transform 1 0 93472 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_9_1016
timestamp 1586364061
transform 1 0 94576 0 1 7072
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_799
timestamp 1586364061
transform 1 0 95220 0 1 7072
box -38 -48 130 592
use scs8hd_fill_1  FILLER_9_1022
timestamp 1586364061
transform 1 0 95128 0 1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_9_1024
timestamp 1586364061
transform 1 0 95312 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_1036
timestamp 1586364061
transform 1 0 96416 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_9_1048
timestamp 1586364061
transform 1 0 97520 0 1 7072
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_800
timestamp 1586364061
transform 1 0 98072 0 1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_9_1055
timestamp 1586364061
transform 1 0 98164 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_1067
timestamp 1586364061
transform 1 0 99268 0 1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_801
timestamp 1586364061
transform 1 0 100924 0 1 7072
box -38 -48 130 592
use scs8hd_decap_6  FILLER_9_1079
timestamp 1586364061
transform 1 0 100372 0 1 7072
box -38 -48 590 592
use scs8hd_decap_12  FILLER_9_1086
timestamp 1586364061
transform 1 0 101016 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_1098
timestamp 1586364061
transform 1 0 102120 0 1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_802
timestamp 1586364061
transform 1 0 103776 0 1 7072
box -38 -48 130 592
use scs8hd_decap_6  FILLER_9_1110
timestamp 1586364061
transform 1 0 103224 0 1 7072
box -38 -48 590 592
use scs8hd_decap_12  FILLER_9_1117
timestamp 1586364061
transform 1 0 103868 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_1129
timestamp 1586364061
transform 1 0 104972 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_9_1141
timestamp 1586364061
transform 1 0 106076 0 1 7072
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_803
timestamp 1586364061
transform 1 0 106628 0 1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_9_1148
timestamp 1586364061
transform 1 0 106720 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_1160
timestamp 1586364061
transform 1 0 107824 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_9_1172
timestamp 1586364061
transform 1 0 108928 0 1 7072
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_804
timestamp 1586364061
transform 1 0 109480 0 1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_9_1179
timestamp 1586364061
transform 1 0 109572 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_1191
timestamp 1586364061
transform 1 0 110676 0 1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_805
timestamp 1586364061
transform 1 0 112332 0 1 7072
box -38 -48 130 592
use scs8hd_decap_6  FILLER_9_1203
timestamp 1586364061
transform 1 0 111780 0 1 7072
box -38 -48 590 592
use scs8hd_decap_12  FILLER_9_1210
timestamp 1586364061
transform 1 0 112424 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_1222
timestamp 1586364061
transform 1 0 113528 0 1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_806
timestamp 1586364061
transform 1 0 115184 0 1 7072
box -38 -48 130 592
use scs8hd_decap_6  FILLER_9_1234
timestamp 1586364061
transform 1 0 114632 0 1 7072
box -38 -48 590 592
use scs8hd_decap_12  FILLER_9_1241
timestamp 1586364061
transform 1 0 115276 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_1253
timestamp 1586364061
transform 1 0 116380 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_9_1265
timestamp 1586364061
transform 1 0 117484 0 1 7072
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_807
timestamp 1586364061
transform 1 0 118036 0 1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_9_1272
timestamp 1586364061
transform 1 0 118128 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_1284
timestamp 1586364061
transform 1 0 119232 0 1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_808
timestamp 1586364061
transform 1 0 120888 0 1 7072
box -38 -48 130 592
use scs8hd_decap_6  FILLER_9_1296
timestamp 1586364061
transform 1 0 120336 0 1 7072
box -38 -48 590 592
use scs8hd_decap_12  FILLER_9_1303
timestamp 1586364061
transform 1 0 120980 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_1315
timestamp 1586364061
transform 1 0 122084 0 1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_809
timestamp 1586364061
transform 1 0 123740 0 1 7072
box -38 -48 130 592
use scs8hd_decap_6  FILLER_9_1327
timestamp 1586364061
transform 1 0 123188 0 1 7072
box -38 -48 590 592
use scs8hd_decap_12  FILLER_9_1334
timestamp 1586364061
transform 1 0 123832 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_1346
timestamp 1586364061
transform 1 0 124936 0 1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_810
timestamp 1586364061
transform 1 0 126592 0 1 7072
box -38 -48 130 592
use scs8hd_decap_6  FILLER_9_1358
timestamp 1586364061
transform 1 0 126040 0 1 7072
box -38 -48 590 592
use scs8hd_decap_12  FILLER_9_1365
timestamp 1586364061
transform 1 0 126684 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_1377
timestamp 1586364061
transform 1 0 127788 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_9_1389
timestamp 1586364061
transform 1 0 128892 0 1 7072
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_811
timestamp 1586364061
transform 1 0 129444 0 1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_9_1396
timestamp 1586364061
transform 1 0 129536 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_1408
timestamp 1586364061
transform 1 0 130640 0 1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_812
timestamp 1586364061
transform 1 0 132296 0 1 7072
box -38 -48 130 592
use scs8hd_decap_6  FILLER_9_1420
timestamp 1586364061
transform 1 0 131744 0 1 7072
box -38 -48 590 592
use scs8hd_decap_12  FILLER_9_1427
timestamp 1586364061
transform 1 0 132388 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_1439
timestamp 1586364061
transform 1 0 133492 0 1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_813
timestamp 1586364061
transform 1 0 135148 0 1 7072
box -38 -48 130 592
use scs8hd_decap_6  FILLER_9_1451
timestamp 1586364061
transform 1 0 134596 0 1 7072
box -38 -48 590 592
use scs8hd_decap_12  FILLER_9_1458
timestamp 1586364061
transform 1 0 135240 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_1470
timestamp 1586364061
transform 1 0 136344 0 1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_814
timestamp 1586364061
transform 1 0 138000 0 1 7072
box -38 -48 130 592
use scs8hd_decap_6  FILLER_9_1482
timestamp 1586364061
transform 1 0 137448 0 1 7072
box -38 -48 590 592
use scs8hd_decap_12  FILLER_9_1489
timestamp 1586364061
transform 1 0 138092 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_1501
timestamp 1586364061
transform 1 0 139196 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_9_1513
timestamp 1586364061
transform 1 0 140300 0 1 7072
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_815
timestamp 1586364061
transform 1 0 140852 0 1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_9_1520
timestamp 1586364061
transform 1 0 140944 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_1532
timestamp 1586364061
transform 1 0 142048 0 1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_816
timestamp 1586364061
transform 1 0 143704 0 1 7072
box -38 -48 130 592
use scs8hd_decap_6  FILLER_9_1544
timestamp 1586364061
transform 1 0 143152 0 1 7072
box -38 -48 590 592
use scs8hd_decap_12  FILLER_9_1551
timestamp 1586364061
transform 1 0 143796 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_1563
timestamp 1586364061
transform 1 0 144900 0 1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_817
timestamp 1586364061
transform 1 0 146556 0 1 7072
box -38 -48 130 592
use scs8hd_decap_6  FILLER_9_1575
timestamp 1586364061
transform 1 0 146004 0 1 7072
box -38 -48 590 592
use scs8hd_decap_12  FILLER_9_1582
timestamp 1586364061
transform 1 0 146648 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_1594
timestamp 1586364061
transform 1 0 147752 0 1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_818
timestamp 1586364061
transform 1 0 149408 0 1 7072
box -38 -48 130 592
use scs8hd_decap_6  FILLER_9_1606
timestamp 1586364061
transform 1 0 148856 0 1 7072
box -38 -48 590 592
use scs8hd_decap_12  FILLER_9_1613
timestamp 1586364061
transform 1 0 149500 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_1625
timestamp 1586364061
transform 1 0 150604 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_9_1637
timestamp 1586364061
transform 1 0 151708 0 1 7072
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_819
timestamp 1586364061
transform 1 0 152260 0 1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_9_1644
timestamp 1586364061
transform 1 0 152352 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_1656
timestamp 1586364061
transform 1 0 153456 0 1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_820
timestamp 1586364061
transform 1 0 155112 0 1 7072
box -38 -48 130 592
use scs8hd_decap_6  FILLER_9_1668
timestamp 1586364061
transform 1 0 154560 0 1 7072
box -38 -48 590 592
use scs8hd_decap_12  FILLER_9_1675
timestamp 1586364061
transform 1 0 155204 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_1687
timestamp 1586364061
transform 1 0 156308 0 1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_821
timestamp 1586364061
transform 1 0 157964 0 1 7072
box -38 -48 130 592
use scs8hd_decap_6  FILLER_9_1699
timestamp 1586364061
transform 1 0 157412 0 1 7072
box -38 -48 590 592
use scs8hd_decap_12  FILLER_9_1706
timestamp 1586364061
transform 1 0 158056 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_1718
timestamp 1586364061
transform 1 0 159160 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_9_1730
timestamp 1586364061
transform 1 0 160264 0 1 7072
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_822
timestamp 1586364061
transform 1 0 160816 0 1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_9_1737
timestamp 1586364061
transform 1 0 160908 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_1749
timestamp 1586364061
transform 1 0 162012 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_9_1761
timestamp 1586364061
transform 1 0 163116 0 1 7072
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_823
timestamp 1586364061
transform 1 0 163668 0 1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_9_1768
timestamp 1586364061
transform 1 0 163760 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_1780
timestamp 1586364061
transform 1 0 164864 0 1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_824
timestamp 1586364061
transform 1 0 166520 0 1 7072
box -38 -48 130 592
use scs8hd_decap_6  FILLER_9_1792
timestamp 1586364061
transform 1 0 165968 0 1 7072
box -38 -48 590 592
use scs8hd_decap_12  FILLER_9_1799
timestamp 1586364061
transform 1 0 166612 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_1811
timestamp 1586364061
transform 1 0 167716 0 1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_825
timestamp 1586364061
transform 1 0 169372 0 1 7072
box -38 -48 130 592
use scs8hd_decap_6  FILLER_9_1823
timestamp 1586364061
transform 1 0 168820 0 1 7072
box -38 -48 590 592
use scs8hd_decap_12  FILLER_9_1830
timestamp 1586364061
transform 1 0 169464 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_1842
timestamp 1586364061
transform 1 0 170568 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_9_1854
timestamp 1586364061
transform 1 0 171672 0 1 7072
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_826
timestamp 1586364061
transform 1 0 172224 0 1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_9_1861
timestamp 1586364061
transform 1 0 172316 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_1873
timestamp 1586364061
transform 1 0 173420 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_9_1885
timestamp 1586364061
transform 1 0 174524 0 1 7072
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_827
timestamp 1586364061
transform 1 0 175076 0 1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_9_1892
timestamp 1586364061
transform 1 0 175168 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_1904
timestamp 1586364061
transform 1 0 176272 0 1 7072
box -38 -48 1142 592
use scs8hd_buf_2  _18_
timestamp 1586364061
transform 1 0 178020 0 1 7072
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_828
timestamp 1586364061
transform 1 0 177928 0 1 7072
box -38 -48 130 592
use scs8hd_decap_6  FILLER_9_1916
timestamp 1586364061
transform 1 0 177376 0 1 7072
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA__18__A
timestamp 1586364061
transform 1 0 178572 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_1927
timestamp 1586364061
transform 1 0 178388 0 1 7072
box -38 -48 222 592
use scs8hd_decap_12  FILLER_9_1931
timestamp 1586364061
transform 1 0 178756 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_9_1943
timestamp 1586364061
transform 1 0 179860 0 1 7072
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_829
timestamp 1586364061
transform 1 0 180780 0 1 7072
box -38 -48 130 592
use scs8hd_fill_2  FILLER_9_1951
timestamp 1586364061
transform 1 0 180596 0 1 7072
box -38 -48 222 592
use scs8hd_decap_12  FILLER_9_1954
timestamp 1586364061
transform 1 0 180872 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_1966
timestamp 1586364061
transform 1 0 181976 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_9_1978
timestamp 1586364061
transform 1 0 183080 0 1 7072
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_830
timestamp 1586364061
transform 1 0 183632 0 1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_9_1985
timestamp 1586364061
transform 1 0 183724 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_1997
timestamp 1586364061
transform 1 0 184828 0 1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_831
timestamp 1586364061
transform 1 0 186484 0 1 7072
box -38 -48 130 592
use scs8hd_decap_6  FILLER_9_2009
timestamp 1586364061
transform 1 0 185932 0 1 7072
box -38 -48 590 592
use scs8hd_decap_12  FILLER_9_2016
timestamp 1586364061
transform 1 0 186576 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_2028
timestamp 1586364061
transform 1 0 187680 0 1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_832
timestamp 1586364061
transform 1 0 189336 0 1 7072
box -38 -48 130 592
use scs8hd_decap_6  FILLER_9_2040
timestamp 1586364061
transform 1 0 188784 0 1 7072
box -38 -48 590 592
use scs8hd_decap_12  FILLER_9_2047
timestamp 1586364061
transform 1 0 189428 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_2059
timestamp 1586364061
transform 1 0 190532 0 1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_833
timestamp 1586364061
transform 1 0 192188 0 1 7072
box -38 -48 130 592
use scs8hd_decap_6  FILLER_9_2071
timestamp 1586364061
transform 1 0 191636 0 1 7072
box -38 -48 590 592
use scs8hd_decap_12  FILLER_9_2078
timestamp 1586364061
transform 1 0 192280 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_2090
timestamp 1586364061
transform 1 0 193384 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_9_2102
timestamp 1586364061
transform 1 0 194488 0 1 7072
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_834
timestamp 1586364061
transform 1 0 195040 0 1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_9_2109
timestamp 1586364061
transform 1 0 195132 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_2121
timestamp 1586364061
transform 1 0 196236 0 1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_835
timestamp 1586364061
transform 1 0 197892 0 1 7072
box -38 -48 130 592
use scs8hd_decap_6  FILLER_9_2133
timestamp 1586364061
transform 1 0 197340 0 1 7072
box -38 -48 590 592
use scs8hd_decap_12  FILLER_9_2140
timestamp 1586364061
transform 1 0 197984 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_2152
timestamp 1586364061
transform 1 0 199088 0 1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_836
timestamp 1586364061
transform 1 0 200744 0 1 7072
box -38 -48 130 592
use scs8hd_decap_6  FILLER_9_2164
timestamp 1586364061
transform 1 0 200192 0 1 7072
box -38 -48 590 592
use scs8hd_decap_12  FILLER_9_2171
timestamp 1586364061
transform 1 0 200836 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_2183
timestamp 1586364061
transform 1 0 201940 0 1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_837
timestamp 1586364061
transform 1 0 203596 0 1 7072
box -38 -48 130 592
use scs8hd_decap_6  FILLER_9_2195
timestamp 1586364061
transform 1 0 203044 0 1 7072
box -38 -48 590 592
use scs8hd_decap_12  FILLER_9_2202
timestamp 1586364061
transform 1 0 203688 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_2214
timestamp 1586364061
transform 1 0 204792 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_9_2226
timestamp 1586364061
transform 1 0 205896 0 1 7072
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_838
timestamp 1586364061
transform 1 0 206448 0 1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_9_2233
timestamp 1586364061
transform 1 0 206540 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_2245
timestamp 1586364061
transform 1 0 207644 0 1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_839
timestamp 1586364061
transform 1 0 209300 0 1 7072
box -38 -48 130 592
use scs8hd_decap_6  FILLER_9_2257
timestamp 1586364061
transform 1 0 208748 0 1 7072
box -38 -48 590 592
use scs8hd_decap_12  FILLER_9_2264
timestamp 1586364061
transform 1 0 209392 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_2276
timestamp 1586364061
transform 1 0 210496 0 1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_840
timestamp 1586364061
transform 1 0 212152 0 1 7072
box -38 -48 130 592
use scs8hd_decap_6  FILLER_9_2288
timestamp 1586364061
transform 1 0 211600 0 1 7072
box -38 -48 590 592
use scs8hd_decap_12  FILLER_9_2295
timestamp 1586364061
transform 1 0 212244 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_2307
timestamp 1586364061
transform 1 0 213348 0 1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_841
timestamp 1586364061
transform 1 0 215004 0 1 7072
box -38 -48 130 592
use scs8hd_decap_6  FILLER_9_2319
timestamp 1586364061
transform 1 0 214452 0 1 7072
box -38 -48 590 592
use scs8hd_decap_12  FILLER_9_2326
timestamp 1586364061
transform 1 0 215096 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_2338
timestamp 1586364061
transform 1 0 216200 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_9_2350
timestamp 1586364061
transform 1 0 217304 0 1 7072
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_842
timestamp 1586364061
transform 1 0 217856 0 1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_9_2357
timestamp 1586364061
transform 1 0 217948 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_2369
timestamp 1586364061
transform 1 0 219052 0 1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_843
timestamp 1586364061
transform 1 0 220708 0 1 7072
box -38 -48 130 592
use scs8hd_decap_6  FILLER_9_2381
timestamp 1586364061
transform 1 0 220156 0 1 7072
box -38 -48 590 592
use scs8hd_decap_12  FILLER_9_2388
timestamp 1586364061
transform 1 0 220800 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_2400
timestamp 1586364061
transform 1 0 221904 0 1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_844
timestamp 1586364061
transform 1 0 223560 0 1 7072
box -38 -48 130 592
use scs8hd_decap_6  FILLER_9_2412
timestamp 1586364061
transform 1 0 223008 0 1 7072
box -38 -48 590 592
use scs8hd_decap_12  FILLER_9_2419
timestamp 1586364061
transform 1 0 223652 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_2431
timestamp 1586364061
transform 1 0 224756 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_9_2443
timestamp 1586364061
transform 1 0 225860 0 1 7072
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_845
timestamp 1586364061
transform 1 0 226412 0 1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_9_2450
timestamp 1586364061
transform 1 0 226504 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_2462
timestamp 1586364061
transform 1 0 227608 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_9_2474
timestamp 1586364061
transform 1 0 228712 0 1 7072
box -38 -48 590 592
use scs8hd_buf_2  _23_
timestamp 1586364061
transform 1 0 229356 0 1 7072
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_846
timestamp 1586364061
transform 1 0 229264 0 1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__23__A
timestamp 1586364061
transform 1 0 229908 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_2485
timestamp 1586364061
transform 1 0 229724 0 1 7072
box -38 -48 222 592
use scs8hd_decap_12  FILLER_9_2489
timestamp 1586364061
transform 1 0 230092 0 1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_847
timestamp 1586364061
transform 1 0 232116 0 1 7072
box -38 -48 130 592
use scs8hd_decap_8  FILLER_9_2501
timestamp 1586364061
transform 1 0 231196 0 1 7072
box -38 -48 774 592
use scs8hd_fill_2  FILLER_9_2509
timestamp 1586364061
transform 1 0 231932 0 1 7072
box -38 -48 222 592
use scs8hd_decap_12  FILLER_9_2512
timestamp 1586364061
transform 1 0 232208 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_2524
timestamp 1586364061
transform 1 0 233312 0 1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_848
timestamp 1586364061
transform 1 0 234968 0 1 7072
box -38 -48 130 592
use scs8hd_decap_6  FILLER_9_2536
timestamp 1586364061
transform 1 0 234416 0 1 7072
box -38 -48 590 592
use scs8hd_decap_12  FILLER_9_2543
timestamp 1586364061
transform 1 0 235060 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_2555
timestamp 1586364061
transform 1 0 236164 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_9_2567
timestamp 1586364061
transform 1 0 237268 0 1 7072
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_849
timestamp 1586364061
transform 1 0 237820 0 1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_9_2574
timestamp 1586364061
transform 1 0 237912 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_2586
timestamp 1586364061
transform 1 0 239016 0 1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_850
timestamp 1586364061
transform 1 0 240672 0 1 7072
box -38 -48 130 592
use scs8hd_decap_6  FILLER_9_2598
timestamp 1586364061
transform 1 0 240120 0 1 7072
box -38 -48 590 592
use scs8hd_decap_12  FILLER_9_2605
timestamp 1586364061
transform 1 0 240764 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_2617
timestamp 1586364061
transform 1 0 241868 0 1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_851
timestamp 1586364061
transform 1 0 243524 0 1 7072
box -38 -48 130 592
use scs8hd_decap_6  FILLER_9_2629
timestamp 1586364061
transform 1 0 242972 0 1 7072
box -38 -48 590 592
use scs8hd_decap_12  FILLER_9_2636
timestamp 1586364061
transform 1 0 243616 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_2648
timestamp 1586364061
transform 1 0 244720 0 1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_852
timestamp 1586364061
transform 1 0 246376 0 1 7072
box -38 -48 130 592
use scs8hd_decap_6  FILLER_9_2660
timestamp 1586364061
transform 1 0 245824 0 1 7072
box -38 -48 590 592
use scs8hd_decap_12  FILLER_9_2667
timestamp 1586364061
transform 1 0 246468 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_2679
timestamp 1586364061
transform 1 0 247572 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_9_2691
timestamp 1586364061
transform 1 0 248676 0 1 7072
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_853
timestamp 1586364061
transform 1 0 249228 0 1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_9_2698
timestamp 1586364061
transform 1 0 249320 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_2710
timestamp 1586364061
transform 1 0 250424 0 1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_854
timestamp 1586364061
transform 1 0 252080 0 1 7072
box -38 -48 130 592
use scs8hd_decap_6  FILLER_9_2722
timestamp 1586364061
transform 1 0 251528 0 1 7072
box -38 -48 590 592
use scs8hd_decap_12  FILLER_9_2729
timestamp 1586364061
transform 1 0 252172 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_2741
timestamp 1586364061
transform 1 0 253276 0 1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_855
timestamp 1586364061
transform 1 0 254932 0 1 7072
box -38 -48 130 592
use scs8hd_decap_6  FILLER_9_2753
timestamp 1586364061
transform 1 0 254380 0 1 7072
box -38 -48 590 592
use scs8hd_decap_12  FILLER_9_2760
timestamp 1586364061
transform 1 0 255024 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_2772
timestamp 1586364061
transform 1 0 256128 0 1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_856
timestamp 1586364061
transform 1 0 257784 0 1 7072
box -38 -48 130 592
use scs8hd_decap_6  FILLER_9_2784
timestamp 1586364061
transform 1 0 257232 0 1 7072
box -38 -48 590 592
use scs8hd_decap_12  FILLER_9_2791
timestamp 1586364061
transform 1 0 257876 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_2803
timestamp 1586364061
transform 1 0 258980 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_9_2815
timestamp 1586364061
transform 1 0 260084 0 1 7072
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_857
timestamp 1586364061
transform 1 0 260636 0 1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_9_2822
timestamp 1586364061
transform 1 0 260728 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_2834
timestamp 1586364061
transform 1 0 261832 0 1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_858
timestamp 1586364061
transform 1 0 263488 0 1 7072
box -38 -48 130 592
use scs8hd_decap_6  FILLER_9_2846
timestamp 1586364061
transform 1 0 262936 0 1 7072
box -38 -48 590 592
use scs8hd_decap_12  FILLER_9_2853
timestamp 1586364061
transform 1 0 263580 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_2865
timestamp 1586364061
transform 1 0 264684 0 1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_859
timestamp 1586364061
transform 1 0 266340 0 1 7072
box -38 -48 130 592
use scs8hd_decap_6  FILLER_9_2877
timestamp 1586364061
transform 1 0 265788 0 1 7072
box -38 -48 590 592
use scs8hd_decap_12  FILLER_9_2884
timestamp 1586364061
transform 1 0 266432 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_2896
timestamp 1586364061
transform 1 0 267536 0 1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_860
timestamp 1586364061
transform 1 0 269192 0 1 7072
box -38 -48 130 592
use scs8hd_decap_6  FILLER_9_2908
timestamp 1586364061
transform 1 0 268640 0 1 7072
box -38 -48 590 592
use scs8hd_decap_12  FILLER_9_2915
timestamp 1586364061
transform 1 0 269284 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_2927
timestamp 1586364061
transform 1 0 270388 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_9_2939
timestamp 1586364061
transform 1 0 271492 0 1 7072
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_861
timestamp 1586364061
transform 1 0 272044 0 1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_9_2946
timestamp 1586364061
transform 1 0 272136 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_2958
timestamp 1586364061
transform 1 0 273240 0 1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_862
timestamp 1586364061
transform 1 0 274896 0 1 7072
box -38 -48 130 592
use scs8hd_decap_6  FILLER_9_2970
timestamp 1586364061
transform 1 0 274344 0 1 7072
box -38 -48 590 592
use scs8hd_decap_12  FILLER_9_2977
timestamp 1586364061
transform 1 0 274988 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_2989
timestamp 1586364061
transform 1 0 276092 0 1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_863
timestamp 1586364061
transform 1 0 277748 0 1 7072
box -38 -48 130 592
use scs8hd_decap_6  FILLER_9_3001
timestamp 1586364061
transform 1 0 277196 0 1 7072
box -38 -48 590 592
use scs8hd_decap_12  FILLER_9_3008
timestamp 1586364061
transform 1 0 277840 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_3020
timestamp 1586364061
transform 1 0 278944 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_9_3032
timestamp 1586364061
transform 1 0 280048 0 1 7072
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_864
timestamp 1586364061
transform 1 0 280600 0 1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_9_3039
timestamp 1586364061
transform 1 0 280692 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_3051
timestamp 1586364061
transform 1 0 281796 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_9_3063
timestamp 1586364061
transform 1 0 282900 0 1 7072
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_865
timestamp 1586364061
transform 1 0 283452 0 1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_9_3070
timestamp 1586364061
transform 1 0 283544 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_3082
timestamp 1586364061
transform 1 0 284648 0 1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_866
timestamp 1586364061
transform 1 0 286304 0 1 7072
box -38 -48 130 592
use scs8hd_decap_6  FILLER_9_3094
timestamp 1586364061
transform 1 0 285752 0 1 7072
box -38 -48 590 592
use scs8hd_decap_12  FILLER_9_3101
timestamp 1586364061
transform 1 0 286396 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_3113
timestamp 1586364061
transform 1 0 287500 0 1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_867
timestamp 1586364061
transform 1 0 289156 0 1 7072
box -38 -48 130 592
use scs8hd_decap_6  FILLER_9_3125
timestamp 1586364061
transform 1 0 288604 0 1 7072
box -38 -48 590 592
use scs8hd_decap_12  FILLER_9_3132
timestamp 1586364061
transform 1 0 289248 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_3144
timestamp 1586364061
transform 1 0 290352 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_9_3156
timestamp 1586364061
transform 1 0 291456 0 1 7072
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_868
timestamp 1586364061
transform 1 0 292008 0 1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_9_3163
timestamp 1586364061
transform 1 0 292100 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_3175
timestamp 1586364061
transform 1 0 293204 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_9_3187
timestamp 1586364061
transform 1 0 294308 0 1 7072
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_869
timestamp 1586364061
transform 1 0 294860 0 1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_9_3194
timestamp 1586364061
transform 1 0 294952 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_3206
timestamp 1586364061
transform 1 0 296056 0 1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_870
timestamp 1586364061
transform 1 0 297712 0 1 7072
box -38 -48 130 592
use scs8hd_decap_6  FILLER_9_3218
timestamp 1586364061
transform 1 0 297160 0 1 7072
box -38 -48 590 592
use scs8hd_decap_12  FILLER_9_3225
timestamp 1586364061
transform 1 0 297804 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_3237
timestamp 1586364061
transform 1 0 298908 0 1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_871
timestamp 1586364061
transform 1 0 300564 0 1 7072
box -38 -48 130 592
use scs8hd_decap_6  FILLER_9_3249
timestamp 1586364061
transform 1 0 300012 0 1 7072
box -38 -48 590 592
use scs8hd_decap_12  FILLER_9_3256
timestamp 1586364061
transform 1 0 300656 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_3268
timestamp 1586364061
transform 1 0 301760 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_9_3280
timestamp 1586364061
transform 1 0 302864 0 1 7072
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_872
timestamp 1586364061
transform 1 0 303416 0 1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_9_3287
timestamp 1586364061
transform 1 0 303508 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_3299
timestamp 1586364061
transform 1 0 304612 0 1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_873
timestamp 1586364061
transform 1 0 306268 0 1 7072
box -38 -48 130 592
use scs8hd_decap_6  FILLER_9_3311
timestamp 1586364061
transform 1 0 305716 0 1 7072
box -38 -48 590 592
use scs8hd_decap_12  FILLER_9_3318
timestamp 1586364061
transform 1 0 306360 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_3330
timestamp 1586364061
transform 1 0 307464 0 1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_874
timestamp 1586364061
transform 1 0 309120 0 1 7072
box -38 -48 130 592
use scs8hd_decap_6  FILLER_9_3342
timestamp 1586364061
transform 1 0 308568 0 1 7072
box -38 -48 590 592
use scs8hd_decap_12  FILLER_9_3349
timestamp 1586364061
transform 1 0 309212 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_3361
timestamp 1586364061
transform 1 0 310316 0 1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_875
timestamp 1586364061
transform 1 0 311972 0 1 7072
box -38 -48 130 592
use scs8hd_decap_6  FILLER_9_3373
timestamp 1586364061
transform 1 0 311420 0 1 7072
box -38 -48 590 592
use scs8hd_decap_12  FILLER_9_3380
timestamp 1586364061
transform 1 0 312064 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_3392
timestamp 1586364061
transform 1 0 313168 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_9_3404
timestamp 1586364061
transform 1 0 314272 0 1 7072
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_876
timestamp 1586364061
transform 1 0 314824 0 1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_9_3411
timestamp 1586364061
transform 1 0 314916 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_3423
timestamp 1586364061
transform 1 0 316020 0 1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_877
timestamp 1586364061
transform 1 0 317676 0 1 7072
box -38 -48 130 592
use scs8hd_decap_6  FILLER_9_3435
timestamp 1586364061
transform 1 0 317124 0 1 7072
box -38 -48 590 592
use scs8hd_decap_12  FILLER_9_3442
timestamp 1586364061
transform 1 0 317768 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_3454
timestamp 1586364061
transform 1 0 318872 0 1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_878
timestamp 1586364061
transform 1 0 320528 0 1 7072
box -38 -48 130 592
use scs8hd_decap_6  FILLER_9_3466
timestamp 1586364061
transform 1 0 319976 0 1 7072
box -38 -48 590 592
use scs8hd_decap_12  FILLER_9_3473
timestamp 1586364061
transform 1 0 320620 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_3485
timestamp 1586364061
transform 1 0 321724 0 1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_879
timestamp 1586364061
transform 1 0 323380 0 1 7072
box -38 -48 130 592
use scs8hd_decap_6  FILLER_9_3497
timestamp 1586364061
transform 1 0 322828 0 1 7072
box -38 -48 590 592
use scs8hd_decap_12  FILLER_9_3504
timestamp 1586364061
transform 1 0 323472 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_3516
timestamp 1586364061
transform 1 0 324576 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_9_3528
timestamp 1586364061
transform 1 0 325680 0 1 7072
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_880
timestamp 1586364061
transform 1 0 326232 0 1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_9_3535
timestamp 1586364061
transform 1 0 326324 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_3547
timestamp 1586364061
transform 1 0 327428 0 1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_881
timestamp 1586364061
transform 1 0 329084 0 1 7072
box -38 -48 130 592
use scs8hd_decap_6  FILLER_9_3559
timestamp 1586364061
transform 1 0 328532 0 1 7072
box -38 -48 590 592
use scs8hd_decap_12  FILLER_9_3566
timestamp 1586364061
transform 1 0 329176 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_3578
timestamp 1586364061
transform 1 0 330280 0 1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_882
timestamp 1586364061
transform 1 0 331936 0 1 7072
box -38 -48 130 592
use scs8hd_decap_6  FILLER_9_3590
timestamp 1586364061
transform 1 0 331384 0 1 7072
box -38 -48 590 592
use scs8hd_decap_12  FILLER_9_3597
timestamp 1586364061
transform 1 0 332028 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_3609
timestamp 1586364061
transform 1 0 333132 0 1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_883
timestamp 1586364061
transform 1 0 334788 0 1 7072
box -38 -48 130 592
use scs8hd_decap_6  FILLER_9_3621
timestamp 1586364061
transform 1 0 334236 0 1 7072
box -38 -48 590 592
use scs8hd_decap_12  FILLER_9_3628
timestamp 1586364061
transform 1 0 334880 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_3640
timestamp 1586364061
transform 1 0 335984 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_9_3652
timestamp 1586364061
transform 1 0 337088 0 1 7072
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_884
timestamp 1586364061
transform 1 0 337640 0 1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_9_3659
timestamp 1586364061
transform 1 0 337732 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_3671
timestamp 1586364061
transform 1 0 338836 0 1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_885
timestamp 1586364061
transform 1 0 340492 0 1 7072
box -38 -48 130 592
use scs8hd_decap_6  FILLER_9_3683
timestamp 1586364061
transform 1 0 339940 0 1 7072
box -38 -48 590 592
use scs8hd_decap_12  FILLER_9_3690
timestamp 1586364061
transform 1 0 340584 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_3702
timestamp 1586364061
transform 1 0 341688 0 1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_886
timestamp 1586364061
transform 1 0 343344 0 1 7072
box -38 -48 130 592
use scs8hd_decap_6  FILLER_9_3714
timestamp 1586364061
transform 1 0 342792 0 1 7072
box -38 -48 590 592
use scs8hd_decap_12  FILLER_9_3721
timestamp 1586364061
transform 1 0 343436 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_3733
timestamp 1586364061
transform 1 0 344540 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_9_3745
timestamp 1586364061
transform 1 0 345644 0 1 7072
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_887
timestamp 1586364061
transform 1 0 346196 0 1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_9_3752
timestamp 1586364061
transform 1 0 346288 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_3764
timestamp 1586364061
transform 1 0 347392 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_9_3776
timestamp 1586364061
transform 1 0 348496 0 1 7072
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_888
timestamp 1586364061
transform 1 0 349048 0 1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_9_3783
timestamp 1586364061
transform 1 0 349140 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_3795
timestamp 1586364061
transform 1 0 350244 0 1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_889
timestamp 1586364061
transform 1 0 351900 0 1 7072
box -38 -48 130 592
use scs8hd_decap_6  FILLER_9_3807
timestamp 1586364061
transform 1 0 351348 0 1 7072
box -38 -48 590 592
use scs8hd_decap_12  FILLER_9_3814
timestamp 1586364061
transform 1 0 351992 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_3826
timestamp 1586364061
transform 1 0 353096 0 1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_890
timestamp 1586364061
transform 1 0 354752 0 1 7072
box -38 -48 130 592
use scs8hd_decap_6  FILLER_9_3838
timestamp 1586364061
transform 1 0 354200 0 1 7072
box -38 -48 590 592
use scs8hd_decap_12  FILLER_9_3845
timestamp 1586364061
transform 1 0 354844 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_3857
timestamp 1586364061
transform 1 0 355948 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_9_3869
timestamp 1586364061
transform 1 0 357052 0 1 7072
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_891
timestamp 1586364061
transform 1 0 357604 0 1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_9_3876
timestamp 1586364061
transform 1 0 357696 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_3888
timestamp 1586364061
transform 1 0 358800 0 1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_892
timestamp 1586364061
transform 1 0 360456 0 1 7072
box -38 -48 130 592
use scs8hd_decap_6  FILLER_9_3900
timestamp 1586364061
transform 1 0 359904 0 1 7072
box -38 -48 590 592
use scs8hd_decap_12  FILLER_9_3907
timestamp 1586364061
transform 1 0 360548 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_3919
timestamp 1586364061
transform 1 0 361652 0 1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_893
timestamp 1586364061
transform 1 0 363308 0 1 7072
box -38 -48 130 592
use scs8hd_decap_6  FILLER_9_3931
timestamp 1586364061
transform 1 0 362756 0 1 7072
box -38 -48 590 592
use scs8hd_decap_12  FILLER_9_3938
timestamp 1586364061
transform 1 0 363400 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_3950
timestamp 1586364061
transform 1 0 364504 0 1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_894
timestamp 1586364061
transform 1 0 366160 0 1 7072
box -38 -48 130 592
use scs8hd_decap_6  FILLER_9_3962
timestamp 1586364061
transform 1 0 365608 0 1 7072
box -38 -48 590 592
use scs8hd_decap_12  FILLER_9_3969
timestamp 1586364061
transform 1 0 366252 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_3981
timestamp 1586364061
transform 1 0 367356 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_9_3993
timestamp 1586364061
transform 1 0 368460 0 1 7072
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_895
timestamp 1586364061
transform 1 0 369012 0 1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_9_4000
timestamp 1586364061
transform 1 0 369104 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_4012
timestamp 1586364061
transform 1 0 370208 0 1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_896
timestamp 1586364061
transform 1 0 371864 0 1 7072
box -38 -48 130 592
use scs8hd_decap_6  FILLER_9_4024
timestamp 1586364061
transform 1 0 371312 0 1 7072
box -38 -48 590 592
use scs8hd_decap_12  FILLER_9_4031
timestamp 1586364061
transform 1 0 371956 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_4043
timestamp 1586364061
transform 1 0 373060 0 1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_897
timestamp 1586364061
transform 1 0 374716 0 1 7072
box -38 -48 130 592
use scs8hd_decap_6  FILLER_9_4055
timestamp 1586364061
transform 1 0 374164 0 1 7072
box -38 -48 590 592
use scs8hd_decap_12  FILLER_9_4062
timestamp 1586364061
transform 1 0 374808 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_4074
timestamp 1586364061
transform 1 0 375912 0 1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_898
timestamp 1586364061
transform 1 0 377568 0 1 7072
box -38 -48 130 592
use scs8hd_decap_6  FILLER_9_4086
timestamp 1586364061
transform 1 0 377016 0 1 7072
box -38 -48 590 592
use scs8hd_decap_12  FILLER_9_4093
timestamp 1586364061
transform 1 0 377660 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_4105
timestamp 1586364061
transform 1 0 378764 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_9_4117
timestamp 1586364061
transform 1 0 379868 0 1 7072
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_899
timestamp 1586364061
transform 1 0 380420 0 1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_9_4124
timestamp 1586364061
transform 1 0 380512 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_4136
timestamp 1586364061
transform 1 0 381616 0 1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_900
timestamp 1586364061
transform 1 0 383272 0 1 7072
box -38 -48 130 592
use scs8hd_decap_6  FILLER_9_4148
timestamp 1586364061
transform 1 0 382720 0 1 7072
box -38 -48 590 592
use scs8hd_decap_12  FILLER_9_4155
timestamp 1586364061
transform 1 0 383364 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_4167
timestamp 1586364061
transform 1 0 384468 0 1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_901
timestamp 1586364061
transform 1 0 386124 0 1 7072
box -38 -48 130 592
use scs8hd_decap_6  FILLER_9_4179
timestamp 1586364061
transform 1 0 385572 0 1 7072
box -38 -48 590 592
use scs8hd_decap_12  FILLER_9_4186
timestamp 1586364061
transform 1 0 386216 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_4198
timestamp 1586364061
transform 1 0 387320 0 1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_902
timestamp 1586364061
transform 1 0 388976 0 1 7072
box -38 -48 130 592
use scs8hd_decap_6  FILLER_9_4210
timestamp 1586364061
transform 1 0 388424 0 1 7072
box -38 -48 590 592
use scs8hd_decap_12  FILLER_9_4217
timestamp 1586364061
transform 1 0 389068 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_4229
timestamp 1586364061
transform 1 0 390172 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_9_4241
timestamp 1586364061
transform 1 0 391276 0 1 7072
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_903
timestamp 1586364061
transform 1 0 391828 0 1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_9_4248
timestamp 1586364061
transform 1 0 391920 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_4260
timestamp 1586364061
transform 1 0 393024 0 1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_904
timestamp 1586364061
transform 1 0 394680 0 1 7072
box -38 -48 130 592
use scs8hd_decap_6  FILLER_9_4272
timestamp 1586364061
transform 1 0 394128 0 1 7072
box -38 -48 590 592
use scs8hd_decap_12  FILLER_9_4279
timestamp 1586364061
transform 1 0 394772 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_4291
timestamp 1586364061
transform 1 0 395876 0 1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_905
timestamp 1586364061
transform 1 0 397532 0 1 7072
box -38 -48 130 592
use scs8hd_decap_6  FILLER_9_4303
timestamp 1586364061
transform 1 0 396980 0 1 7072
box -38 -48 590 592
use scs8hd_decap_12  FILLER_9_4310
timestamp 1586364061
transform 1 0 397624 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_4322
timestamp 1586364061
transform 1 0 398728 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_9_4334
timestamp 1586364061
transform 1 0 399832 0 1 7072
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_906
timestamp 1586364061
transform 1 0 400384 0 1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_9_4341
timestamp 1586364061
transform 1 0 400476 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_4353
timestamp 1586364061
transform 1 0 401580 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_9_4365
timestamp 1586364061
transform 1 0 402684 0 1 7072
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_907
timestamp 1586364061
transform 1 0 403236 0 1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_9_4372
timestamp 1586364061
transform 1 0 403328 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_4384
timestamp 1586364061
transform 1 0 404432 0 1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_908
timestamp 1586364061
transform 1 0 406088 0 1 7072
box -38 -48 130 592
use scs8hd_decap_6  FILLER_9_4396
timestamp 1586364061
transform 1 0 405536 0 1 7072
box -38 -48 590 592
use scs8hd_decap_12  FILLER_9_4403
timestamp 1586364061
transform 1 0 406180 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_4415
timestamp 1586364061
transform 1 0 407284 0 1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_909
timestamp 1586364061
transform 1 0 408940 0 1 7072
box -38 -48 130 592
use scs8hd_decap_6  FILLER_9_4427
timestamp 1586364061
transform 1 0 408388 0 1 7072
box -38 -48 590 592
use scs8hd_decap_12  FILLER_9_4434
timestamp 1586364061
transform 1 0 409032 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_4446
timestamp 1586364061
transform 1 0 410136 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_9_4458
timestamp 1586364061
transform 1 0 411240 0 1 7072
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_910
timestamp 1586364061
transform 1 0 411792 0 1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_9_4465
timestamp 1586364061
transform 1 0 411884 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_4477
timestamp 1586364061
transform 1 0 412988 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_9_4489
timestamp 1586364061
transform 1 0 414092 0 1 7072
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_911
timestamp 1586364061
transform 1 0 414644 0 1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_9_4496
timestamp 1586364061
transform 1 0 414736 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_4508
timestamp 1586364061
transform 1 0 415840 0 1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_912
timestamp 1586364061
transform 1 0 417496 0 1 7072
box -38 -48 130 592
use scs8hd_decap_6  FILLER_9_4520
timestamp 1586364061
transform 1 0 416944 0 1 7072
box -38 -48 590 592
use scs8hd_decap_12  FILLER_9_4527
timestamp 1586364061
transform 1 0 417588 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_4539
timestamp 1586364061
transform 1 0 418692 0 1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_913
timestamp 1586364061
transform 1 0 420348 0 1 7072
box -38 -48 130 592
use scs8hd_decap_6  FILLER_9_4551
timestamp 1586364061
transform 1 0 419796 0 1 7072
box -38 -48 590 592
use scs8hd_decap_12  FILLER_9_4558
timestamp 1586364061
transform 1 0 420440 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_3  PHY_19
timestamp 1586364061
transform -1 0 422832 0 1 7072
box -38 -48 314 592
use scs8hd_decap_8  FILLER_9_4570
timestamp 1586364061
transform 1 0 421544 0 1 7072
box -38 -48 774 592
use scs8hd_decap_3  FILLER_9_4578
timestamp 1586364061
transform 1 0 422280 0 1 7072
box -38 -48 314 592
<< labels >>
rlabel metal3 s 0 552 480 672 6 address[0]
port 0 nsew default input
rlabel metal3 s 0 1776 480 1896 6 address[1]
port 1 nsew default input
rlabel metal3 s 0 3000 480 3120 6 address[2]
port 2 nsew default input
rlabel metal2 s 21178 0 21234 480 6 address[3]
port 3 nsew default input
rlabel metal3 s 423520 2456 424000 2576 6 data_in
port 4 nsew default input
rlabel metal3 s 423520 824 424000 944 6 enable
port 5 nsew default input
rlabel metal3 s 0 4224 480 4344 6 gfpga_pad_GPIO_PAD[0]
port 6 nsew default bidirectional
rlabel metal3 s 423520 4088 424000 4208 6 gfpga_pad_GPIO_PAD[1]
port 7 nsew default bidirectional
rlabel metal2 s 63498 0 63554 480 6 gfpga_pad_GPIO_PAD[2]
port 8 nsew default bidirectional
rlabel metal3 s 423520 5856 424000 5976 6 gfpga_pad_GPIO_PAD[3]
port 9 nsew default bidirectional
rlabel metal3 s 0 5584 480 5704 6 gfpga_pad_GPIO_PAD[4]
port 10 nsew default bidirectional
rlabel metal2 s 105910 0 105966 480 6 gfpga_pad_GPIO_PAD[5]
port 11 nsew default bidirectional
rlabel metal2 s 148322 0 148378 480 6 gfpga_pad_GPIO_PAD[6]
port 12 nsew default bidirectional
rlabel metal2 s 190734 0 190790 480 6 gfpga_pad_GPIO_PAD[7]
port 13 nsew default bidirectional
rlabel metal2 s 35346 9520 35402 10000 6 top_width_0_height_0__pin_0_
port 14 nsew default input
rlabel metal3 s 423520 9120 424000 9240 6 top_width_0_height_0__pin_10_
port 15 nsew default input
rlabel metal3 s 0 6808 480 6928 6 top_width_0_height_0__pin_11_
port 16 nsew default tristate
rlabel metal3 s 0 8032 480 8152 6 top_width_0_height_0__pin_12_
port 17 nsew default input
rlabel metal2 s 402794 0 402850 480 6 top_width_0_height_0__pin_13_
port 18 nsew default tristate
rlabel metal2 s 388626 9520 388682 10000 6 top_width_0_height_0__pin_14_
port 19 nsew default input
rlabel metal3 s 0 9256 480 9376 6 top_width_0_height_0__pin_15_
port 20 nsew default tristate
rlabel metal2 s 106002 9520 106058 10000 6 top_width_0_height_0__pin_1_
port 21 nsew default tristate
rlabel metal2 s 233146 0 233202 480 6 top_width_0_height_0__pin_2_
port 22 nsew default input
rlabel metal2 s 176658 9520 176714 10000 6 top_width_0_height_0__pin_3_
port 23 nsew default tristate
rlabel metal3 s 423520 7488 424000 7608 6 top_width_0_height_0__pin_4_
port 24 nsew default input
rlabel metal2 s 275558 0 275614 480 6 top_width_0_height_0__pin_5_
port 25 nsew default tristate
rlabel metal2 s 317970 0 318026 480 6 top_width_0_height_0__pin_6_
port 26 nsew default input
rlabel metal2 s 360382 0 360438 480 6 top_width_0_height_0__pin_7_
port 27 nsew default tristate
rlabel metal2 s 247314 9520 247370 10000 6 top_width_0_height_0__pin_8_
port 28 nsew default input
rlabel metal2 s 317970 9520 318026 10000 6 top_width_0_height_0__pin_9_
port 29 nsew default tristate
rlabel metal4 s 71611 2128 71931 7664 6 vpwr
port 30 nsew default input
rlabel metal4 s 142277 2128 142597 7664 6 vgnd
port 31 nsew default input
<< end >>
