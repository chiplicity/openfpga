magic
tech EFS8A
magscale 1 2
timestamp 1602269676
<< locali >>
rect 18613 19159 18647 19261
rect 18647 18785 18682 18819
rect 13823 15657 13829 15691
rect 18883 15657 18889 15691
rect 13823 15589 13857 15657
rect 18883 15589 18917 15657
rect 6779 14909 6871 14943
rect 12391 14909 12518 14943
rect 19763 14025 19901 14059
rect 6469 13719 6503 13957
rect 7199 13719 7233 13787
rect 7199 13685 7205 13719
rect 2881 13379 2915 13481
rect 2881 13345 3042 13379
rect 2881 13175 2915 13345
rect 17503 12393 17509 12427
rect 6503 12325 6548 12359
rect 17503 12325 17537 12393
rect 1995 12257 2030 12291
rect 2743 11781 2881 11815
rect 6009 11747 6043 11781
rect 5917 11713 6043 11747
rect 11713 11679 11747 11781
rect 13921 11679 13955 11781
rect 8217 10999 8251 11101
rect 3007 10081 3042 10115
rect 4905 9571 4939 9673
rect 13001 9367 13035 9469
rect 16951 9129 16957 9163
rect 1995 8993 2030 9027
rect 3801 8891 3835 9129
rect 8723 9061 8769 9095
rect 16951 9061 16985 9129
rect 8527 8993 8654 9027
rect 9539 8313 9584 8347
rect 13639 8041 13645 8075
rect 13639 7973 13673 8041
rect 3617 7735 3651 7973
rect 5733 7803 5767 7973
rect 9873 7327 9907 7497
rect 2881 6307 2915 6409
rect 4537 6103 4571 6205
rect 7843 5865 7849 5899
rect 7843 5797 7877 5865
rect 9045 5559 9079 5661
rect 14013 5559 14047 5865
rect 2639 5117 2674 5151
rect 13277 5015 13311 5253
rect 13737 5151 13771 5321
rect 6469 3995 6503 4165
rect 7475 3927 7509 3995
rect 7475 3893 7481 3927
rect 7941 2907 7975 3077
rect 11621 3043 11655 3145
rect 4203 2465 4330 2499
rect 9413 2431 9447 2601
rect 4997 2295 5031 2397
<< viali >>
rect 15623 19465 15657 19499
rect 13921 19329 13955 19363
rect 13436 19261 13470 19295
rect 14448 19261 14482 19295
rect 15520 19261 15554 19295
rect 15945 19261 15979 19295
rect 17300 19261 17334 19295
rect 18404 19261 18438 19295
rect 18613 19261 18647 19295
rect 19384 19261 19418 19295
rect 19809 19261 19843 19295
rect 19487 19193 19521 19227
rect 13507 19125 13541 19159
rect 14519 19125 14553 19159
rect 14841 19125 14875 19159
rect 17371 19125 17405 19159
rect 17785 19125 17819 19159
rect 18475 19125 18509 19159
rect 18613 19125 18647 19159
rect 18889 19125 18923 19159
rect 14335 18921 14369 18955
rect 12311 18853 12345 18887
rect 12208 18785 12242 18819
rect 13252 18785 13286 18819
rect 14264 18785 14298 18819
rect 16037 18785 16071 18819
rect 16313 18785 16347 18819
rect 17636 18785 17670 18819
rect 18613 18785 18647 18819
rect 19692 18785 19726 18819
rect 16497 18717 16531 18751
rect 18751 18649 18785 18683
rect 12633 18581 12667 18615
rect 13323 18581 13357 18615
rect 15577 18581 15611 18615
rect 17739 18581 17773 18615
rect 19763 18581 19797 18615
rect 1593 18377 1627 18411
rect 2053 18377 2087 18411
rect 8125 18377 8159 18411
rect 13553 18377 13587 18411
rect 14565 18377 14599 18411
rect 18245 18377 18279 18411
rect 19993 18377 20027 18411
rect 18981 18309 19015 18343
rect 1409 18173 1443 18207
rect 7941 18173 7975 18207
rect 10492 18173 10526 18207
rect 12541 18173 12575 18207
rect 13001 18173 13035 18207
rect 14381 18173 14415 18207
rect 14933 18173 14967 18207
rect 15761 18173 15795 18207
rect 16037 18173 16071 18207
rect 18061 18173 18095 18207
rect 19232 18173 19266 18207
rect 8585 18105 8619 18139
rect 13277 18105 13311 18139
rect 16221 18105 16255 18139
rect 17601 18105 17635 18139
rect 10563 18037 10597 18071
rect 10977 18037 11011 18071
rect 11897 18037 11931 18071
rect 12265 18037 12299 18071
rect 14289 18037 14323 18071
rect 15393 18037 15427 18071
rect 16497 18037 16531 18071
rect 18613 18037 18647 18071
rect 19303 18037 19337 18071
rect 19625 18037 19659 18071
rect 15393 17833 15427 17867
rect 16957 17833 16991 17867
rect 18521 17833 18555 17867
rect 10517 17697 10551 17731
rect 10701 17697 10735 17731
rect 12817 17697 12851 17731
rect 13185 17697 13219 17731
rect 14232 17697 14266 17731
rect 15301 17697 15335 17731
rect 15761 17697 15795 17731
rect 16865 17697 16899 17731
rect 17325 17697 17359 17731
rect 18705 17697 18739 17731
rect 18889 17697 18923 17731
rect 10793 17629 10827 17663
rect 13369 17629 13403 17663
rect 16313 17561 16347 17595
rect 12541 17493 12575 17527
rect 14335 17493 14369 17527
rect 18061 17493 18095 17527
rect 17233 17289 17267 17323
rect 19763 17221 19797 17255
rect 8539 17153 8573 17187
rect 14381 17153 14415 17187
rect 8452 17085 8486 17119
rect 9505 17085 9539 17119
rect 9873 17085 9907 17119
rect 12725 17085 12759 17119
rect 12909 17085 12943 17119
rect 13461 17085 13495 17119
rect 15853 17085 15887 17119
rect 16313 17085 16347 17119
rect 16865 17085 16899 17119
rect 18061 17085 18095 17119
rect 18521 17085 18555 17119
rect 19073 17085 19107 17119
rect 19692 17085 19726 17119
rect 20085 17085 20119 17119
rect 10149 17017 10183 17051
rect 10793 17017 10827 17051
rect 14473 17017 14507 17051
rect 15025 17017 15059 17051
rect 16589 17017 16623 17051
rect 8861 16949 8895 16983
rect 9321 16949 9355 16983
rect 10425 16949 10459 16983
rect 11069 16949 11103 16983
rect 12265 16949 12299 16983
rect 12725 16949 12759 16983
rect 14105 16949 14139 16983
rect 15301 16949 15335 16983
rect 15669 16949 15703 16983
rect 17785 16949 17819 16983
rect 18153 16949 18187 16983
rect 10793 16745 10827 16779
rect 13277 16745 13311 16779
rect 15393 16745 15427 16779
rect 16313 16745 16347 16779
rect 18889 16745 18923 16779
rect 19625 16745 19659 16779
rect 11805 16677 11839 16711
rect 17969 16677 18003 16711
rect 18061 16677 18095 16711
rect 8309 16609 8343 16643
rect 8493 16609 8527 16643
rect 9689 16609 9723 16643
rect 10149 16609 10183 16643
rect 13185 16609 13219 16643
rect 13645 16609 13679 16643
rect 15577 16609 15611 16643
rect 15761 16609 15795 16643
rect 19441 16609 19475 16643
rect 8769 16541 8803 16575
rect 10425 16541 10459 16575
rect 11713 16541 11747 16575
rect 11989 16541 12023 16575
rect 16865 16541 16899 16575
rect 18613 16541 18647 16575
rect 7941 16405 7975 16439
rect 9505 16405 9539 16439
rect 12633 16405 12667 16439
rect 14381 16405 14415 16439
rect 14657 16405 14691 16439
rect 15025 16405 15059 16439
rect 1593 16201 1627 16235
rect 11897 16201 11931 16235
rect 14105 16201 14139 16235
rect 14841 16201 14875 16235
rect 17509 16201 17543 16235
rect 17785 16201 17819 16235
rect 11529 16133 11563 16167
rect 12173 16133 12207 16167
rect 18705 16133 18739 16167
rect 10609 16065 10643 16099
rect 12633 16065 12667 16099
rect 13185 16065 13219 16099
rect 14381 16065 14415 16099
rect 14933 16065 14967 16099
rect 15485 16065 15519 16099
rect 18153 16065 18187 16099
rect 19763 16065 19797 16099
rect 1409 15997 1443 16031
rect 6964 15997 6998 16031
rect 7389 15997 7423 16031
rect 9632 15997 9666 16031
rect 10057 15997 10091 16031
rect 16221 15997 16255 16031
rect 16405 15997 16439 16031
rect 17141 15997 17175 16031
rect 19660 15997 19694 16031
rect 20085 15997 20119 16031
rect 7067 15929 7101 15963
rect 8033 15929 8067 15963
rect 8125 15929 8159 15963
rect 8677 15929 8711 15963
rect 9505 15929 9539 15963
rect 10517 15929 10551 15963
rect 10971 15929 11005 15963
rect 13547 15929 13581 15963
rect 16681 15929 16715 15963
rect 18245 15929 18279 15963
rect 2053 15861 2087 15895
rect 7757 15861 7791 15895
rect 9045 15861 9079 15895
rect 9735 15861 9769 15895
rect 13093 15861 13127 15895
rect 15761 15861 15795 15895
rect 19441 15861 19475 15895
rect 6285 15657 6319 15691
rect 8217 15657 8251 15691
rect 10701 15657 10735 15691
rect 13829 15657 13863 15691
rect 16037 15657 16071 15691
rect 17693 15657 17727 15691
rect 18153 15657 18187 15691
rect 18889 15657 18923 15691
rect 7659 15589 7693 15623
rect 8493 15589 8527 15623
rect 10143 15589 10177 15623
rect 11713 15589 11747 15623
rect 17135 15589 17169 15623
rect 9781 15521 9815 15555
rect 13461 15521 13495 15555
rect 15336 15521 15370 15555
rect 16773 15521 16807 15555
rect 18521 15521 18555 15555
rect 7297 15453 7331 15487
rect 11621 15453 11655 15487
rect 11897 15453 11931 15487
rect 9413 15385 9447 15419
rect 6929 15317 6963 15351
rect 8953 15317 8987 15351
rect 13185 15317 13219 15351
rect 14381 15317 14415 15351
rect 15439 15317 15473 15351
rect 19441 15317 19475 15351
rect 6285 15113 6319 15147
rect 7941 15113 7975 15147
rect 9873 15113 9907 15147
rect 11713 15113 11747 15147
rect 13369 15113 13403 15147
rect 16405 15113 16439 15147
rect 17049 15113 17083 15147
rect 19441 15113 19475 15147
rect 14749 15045 14783 15079
rect 16773 15045 16807 15079
rect 18337 15045 18371 15079
rect 19073 15045 19107 15079
rect 7573 14977 7607 15011
rect 8217 14977 8251 15011
rect 8585 14977 8619 15011
rect 10057 14977 10091 15011
rect 11253 14977 11287 15011
rect 13461 14977 13495 15011
rect 15577 14977 15611 15011
rect 18521 14977 18555 15011
rect 19809 14977 19843 15011
rect 5800 14909 5834 14943
rect 6653 14909 6687 14943
rect 6745 14909 6779 14943
rect 7297 14909 7331 14943
rect 12357 14909 12391 14943
rect 12909 14909 12943 14943
rect 14381 14909 14415 14943
rect 16865 14909 16899 14943
rect 17417 14909 17451 14943
rect 8677 14841 8711 14875
rect 9229 14841 9263 14875
rect 10378 14841 10412 14875
rect 11989 14841 12023 14875
rect 13823 14841 13857 14875
rect 15301 14841 15335 14875
rect 15393 14841 15427 14875
rect 17877 14841 17911 14875
rect 18613 14841 18647 14875
rect 5871 14773 5905 14807
rect 10977 14773 11011 14807
rect 12587 14773 12621 14807
rect 15025 14773 15059 14807
rect 9229 14569 9263 14603
rect 9873 14569 9907 14603
rect 10517 14569 10551 14603
rect 10885 14569 10919 14603
rect 12541 14569 12575 14603
rect 13277 14569 13311 14603
rect 15117 14569 15151 14603
rect 15485 14569 15519 14603
rect 15853 14569 15887 14603
rect 17693 14569 17727 14603
rect 7291 14501 7325 14535
rect 11253 14501 11287 14535
rect 11805 14501 11839 14535
rect 13553 14501 13587 14535
rect 14105 14501 14139 14535
rect 17135 14501 17169 14535
rect 18613 14501 18647 14535
rect 18705 14501 18739 14535
rect 19257 14501 19291 14535
rect 4420 14433 4454 14467
rect 5273 14433 5307 14467
rect 5641 14433 5675 14467
rect 5917 14433 5951 14467
rect 10124 14433 10158 14467
rect 15669 14433 15703 14467
rect 16773 14433 16807 14467
rect 6101 14365 6135 14399
rect 6929 14365 6963 14399
rect 11161 14365 11195 14399
rect 13461 14365 13495 14399
rect 16313 14365 16347 14399
rect 4491 14297 4525 14331
rect 4813 14229 4847 14263
rect 7849 14229 7883 14263
rect 8769 14229 8803 14263
rect 10195 14229 10229 14263
rect 12909 14229 12943 14263
rect 14381 14229 14415 14263
rect 4721 14025 4755 14059
rect 5089 14025 5123 14059
rect 8033 14025 8067 14059
rect 14197 14025 14231 14059
rect 15669 14025 15703 14059
rect 17141 14025 17175 14059
rect 17785 14025 17819 14059
rect 19073 14025 19107 14059
rect 19901 14025 19935 14059
rect 6469 13957 6503 13991
rect 17417 13957 17451 13991
rect 20085 13957 20119 13991
rect 5917 13889 5951 13923
rect 4220 13821 4254 13855
rect 5457 13821 5491 13855
rect 5641 13821 5675 13855
rect 8769 13889 8803 13923
rect 10517 13889 10551 13923
rect 11713 13889 11747 13923
rect 12449 13889 12483 13923
rect 15025 13889 15059 13923
rect 16221 13889 16255 13923
rect 18153 13889 18187 13923
rect 6837 13821 6871 13855
rect 9689 13821 9723 13855
rect 10057 13821 10091 13855
rect 16129 13821 16163 13855
rect 19660 13821 19694 13855
rect 8585 13753 8619 13787
rect 9090 13753 9124 13787
rect 10879 13753 10913 13787
rect 12770 13753 12804 13787
rect 14381 13753 14415 13787
rect 14473 13753 14507 13787
rect 16583 13753 16617 13787
rect 18245 13753 18279 13787
rect 18797 13753 18831 13787
rect 4307 13685 4341 13719
rect 6285 13685 6319 13719
rect 6469 13685 6503 13719
rect 6561 13685 6595 13719
rect 7205 13685 7239 13719
rect 7757 13685 7791 13719
rect 11437 13685 11471 13719
rect 12265 13685 12299 13719
rect 13369 13685 13403 13719
rect 13645 13685 13679 13719
rect 19441 13685 19475 13719
rect 2881 13481 2915 13515
rect 11529 13481 11563 13515
rect 13461 13481 13495 13515
rect 16221 13481 16255 13515
rect 17509 13481 17543 13515
rect 18153 13481 18187 13515
rect 6561 13413 6595 13447
rect 7389 13413 7423 13447
rect 8125 13413 8159 13447
rect 10701 13413 10735 13447
rect 12265 13413 12299 13447
rect 13829 13413 13863 13447
rect 16634 13413 16668 13447
rect 18429 13413 18463 13447
rect 5089 13345 5123 13379
rect 5365 13345 5399 13379
rect 5549 13345 5583 13379
rect 15368 13345 15402 13379
rect 6469 13277 6503 13311
rect 7113 13277 7147 13311
rect 8033 13277 8067 13311
rect 8677 13277 8711 13311
rect 10609 13277 10643 13311
rect 12173 13277 12207 13311
rect 13737 13277 13771 13311
rect 14381 13277 14415 13311
rect 16313 13277 16347 13311
rect 18337 13277 18371 13311
rect 18613 13277 18647 13311
rect 11161 13209 11195 13243
rect 12725 13209 12759 13243
rect 2881 13141 2915 13175
rect 3111 13141 3145 13175
rect 5825 13141 5859 13175
rect 6285 13141 6319 13175
rect 7757 13141 7791 13175
rect 10333 13141 10367 13175
rect 11897 13141 11931 13175
rect 15439 13141 15473 13175
rect 17233 13141 17267 13175
rect 2697 12937 2731 12971
rect 2973 12937 3007 12971
rect 3985 12937 4019 12971
rect 4307 12937 4341 12971
rect 11437 12937 11471 12971
rect 13645 12937 13679 12971
rect 13921 12937 13955 12971
rect 14289 12937 14323 12971
rect 15485 12937 15519 12971
rect 11897 12869 11931 12903
rect 7113 12801 7147 12835
rect 9137 12801 9171 12835
rect 10425 12801 10459 12835
rect 12265 12801 12299 12835
rect 12725 12801 12759 12835
rect 14565 12801 14599 12835
rect 14841 12801 14875 12835
rect 16129 12801 16163 12835
rect 18613 12801 18647 12835
rect 18889 12801 18923 12835
rect 2212 12733 2246 12767
rect 3192 12733 3226 12767
rect 3617 12733 3651 12767
rect 4236 12733 4270 12767
rect 5089 12733 5123 12767
rect 5457 12733 5491 12767
rect 5733 12733 5767 12767
rect 5917 12733 5951 12767
rect 17049 12733 17083 12767
rect 17785 12733 17819 12767
rect 18337 12733 18371 12767
rect 7205 12665 7239 12699
rect 7757 12665 7791 12699
rect 8861 12665 8895 12699
rect 8953 12665 8987 12699
rect 10517 12665 10551 12699
rect 11069 12665 11103 12699
rect 13046 12665 13080 12699
rect 14657 12665 14691 12699
rect 16450 12665 16484 12699
rect 18705 12665 18739 12699
rect 2283 12597 2317 12631
rect 3295 12597 3329 12631
rect 4721 12597 4755 12631
rect 6285 12597 6319 12631
rect 6653 12597 6687 12631
rect 8033 12597 8067 12631
rect 8677 12597 8711 12631
rect 10241 12597 10275 12631
rect 15945 12597 15979 12631
rect 3111 12393 3145 12427
rect 6009 12393 6043 12427
rect 7389 12393 7423 12427
rect 7849 12393 7883 12427
rect 8953 12393 8987 12427
rect 10701 12393 10735 12427
rect 12357 12393 12391 12427
rect 13461 12393 13495 12427
rect 14657 12393 14691 12427
rect 16681 12393 16715 12427
rect 17509 12393 17543 12427
rect 18337 12393 18371 12427
rect 18797 12393 18831 12427
rect 6469 12325 6503 12359
rect 8125 12325 8159 12359
rect 9873 12325 9907 12359
rect 10425 12325 10459 12359
rect 11437 12325 11471 12359
rect 13829 12325 13863 12359
rect 14381 12325 14415 12359
rect 15485 12325 15519 12359
rect 16037 12325 16071 12359
rect 19073 12325 19107 12359
rect 1961 12257 1995 12291
rect 3008 12257 3042 12291
rect 4905 12257 4939 12291
rect 5181 12257 5215 12291
rect 7113 12257 7147 12291
rect 17141 12257 17175 12291
rect 3709 12189 3743 12223
rect 5365 12189 5399 12223
rect 6193 12189 6227 12223
rect 8033 12189 8067 12223
rect 8309 12189 8343 12223
rect 9781 12189 9815 12223
rect 11345 12189 11379 12223
rect 11621 12189 11655 12223
rect 13737 12189 13771 12223
rect 15393 12189 15427 12223
rect 18981 12189 19015 12223
rect 19257 12189 19291 12223
rect 18061 12121 18095 12155
rect 2099 12053 2133 12087
rect 5733 12053 5767 12087
rect 12725 12053 12759 12087
rect 15025 12053 15059 12087
rect 16313 12053 16347 12087
rect 3065 11849 3099 11883
rect 4721 11849 4755 11883
rect 8125 11849 8159 11883
rect 9045 11849 9079 11883
rect 10701 11849 10735 11883
rect 13829 11849 13863 11883
rect 14197 11849 14231 11883
rect 15853 11849 15887 11883
rect 17785 11849 17819 11883
rect 19625 11849 19659 11883
rect 2881 11781 2915 11815
rect 6009 11781 6043 11815
rect 11713 11781 11747 11815
rect 5089 11713 5123 11747
rect 6837 11713 6871 11747
rect 11483 11713 11517 11747
rect 13921 11781 13955 11815
rect 19993 11781 20027 11815
rect 14933 11713 14967 11747
rect 15577 11713 15611 11747
rect 16497 11713 16531 11747
rect 17141 11713 17175 11747
rect 19349 11713 19383 11747
rect 1644 11645 1678 11679
rect 2672 11645 2706 11679
rect 3433 11645 3467 11679
rect 3893 11645 3927 11679
rect 4169 11645 4203 11679
rect 5181 11645 5215 11679
rect 5733 11645 5767 11679
rect 8585 11645 8619 11679
rect 9505 11645 9539 11679
rect 10425 11645 10459 11679
rect 11380 11645 11414 11679
rect 11713 11645 11747 11679
rect 12909 11645 12943 11679
rect 13921 11645 13955 11679
rect 1731 11577 1765 11611
rect 4353 11577 4387 11611
rect 7199 11577 7233 11611
rect 9867 11577 9901 11611
rect 11805 11577 11839 11611
rect 13271 11577 13305 11611
rect 14749 11577 14783 11611
rect 15025 11577 15059 11611
rect 16313 11577 16347 11611
rect 16589 11577 16623 11611
rect 18521 11577 18555 11611
rect 18705 11577 18739 11611
rect 18797 11577 18831 11611
rect 2053 11509 2087 11543
rect 2513 11509 2547 11543
rect 6285 11509 6319 11543
rect 6653 11509 6687 11543
rect 7757 11509 7791 11543
rect 9413 11509 9447 11543
rect 11253 11509 11287 11543
rect 12817 11509 12851 11543
rect 17417 11509 17451 11543
rect 1593 11305 1627 11339
rect 5181 11305 5215 11339
rect 5549 11305 5583 11339
rect 6745 11305 6779 11339
rect 7113 11305 7147 11339
rect 10701 11305 10735 11339
rect 11253 11305 11287 11339
rect 12909 11305 12943 11339
rect 14933 11305 14967 11339
rect 16865 11305 16899 11339
rect 18705 11305 18739 11339
rect 4905 11237 4939 11271
rect 7481 11237 7515 11271
rect 8033 11237 8067 11271
rect 8677 11237 8711 11271
rect 10143 11237 10177 11271
rect 11713 11237 11747 11271
rect 13461 11237 13495 11271
rect 15939 11237 15973 11271
rect 17646 11237 17680 11271
rect 19257 11237 19291 11271
rect 1409 11169 1443 11203
rect 3040 11169 3074 11203
rect 4169 11169 4203 11203
rect 4721 11169 4755 11203
rect 5733 11169 5767 11203
rect 6193 11169 6227 11203
rect 9781 11169 9815 11203
rect 15577 11169 15611 11203
rect 18245 11169 18279 11203
rect 3709 11101 3743 11135
rect 6469 11101 6503 11135
rect 7389 11101 7423 11135
rect 8217 11101 8251 11135
rect 11621 11101 11655 11135
rect 11897 11101 11931 11135
rect 13369 11101 13403 11135
rect 14013 11101 14047 11135
rect 17141 11101 17175 11135
rect 17325 11101 17359 11135
rect 19165 11101 19199 11135
rect 19533 11101 19567 11135
rect 3111 11033 3145 11067
rect 12541 11033 12575 11067
rect 8217 10965 8251 10999
rect 8401 10965 8435 10999
rect 14289 10965 14323 10999
rect 16497 10965 16531 10999
rect 2145 10761 2179 10795
rect 4721 10761 4755 10795
rect 6561 10761 6595 10795
rect 9459 10761 9493 10795
rect 11621 10761 11655 10795
rect 16313 10761 16347 10795
rect 19625 10761 19659 10795
rect 2513 10693 2547 10727
rect 7849 10625 7883 10659
rect 8493 10625 8527 10659
rect 10609 10625 10643 10659
rect 11253 10625 11287 10659
rect 12817 10625 12851 10659
rect 14381 10625 14415 10659
rect 14657 10625 14691 10659
rect 16497 10625 16531 10659
rect 19257 10625 19291 10659
rect 1660 10557 1694 10591
rect 2672 10557 2706 10591
rect 3893 10557 3927 10591
rect 4077 10557 4111 10591
rect 5457 10557 5491 10591
rect 5733 10557 5767 10591
rect 5917 10557 5951 10591
rect 9388 10557 9422 10591
rect 9781 10557 9815 10591
rect 7389 10489 7423 10523
rect 7941 10489 7975 10523
rect 9137 10489 9171 10523
rect 10701 10489 10735 10523
rect 12909 10489 12943 10523
rect 13461 10489 13495 10523
rect 14473 10489 14507 10523
rect 16589 10489 16623 10523
rect 17141 10489 17175 10523
rect 18613 10489 18647 10523
rect 18705 10489 18739 10523
rect 1731 10421 1765 10455
rect 2743 10421 2777 10455
rect 3065 10421 3099 10455
rect 3433 10421 3467 10455
rect 3893 10421 3927 10455
rect 5089 10421 5123 10455
rect 6193 10421 6227 10455
rect 8769 10421 8803 10455
rect 10241 10421 10275 10455
rect 12265 10421 12299 10455
rect 13737 10421 13771 10455
rect 14197 10421 14231 10455
rect 15669 10421 15703 10455
rect 17417 10421 17451 10455
rect 17785 10421 17819 10455
rect 18337 10421 18371 10455
rect 19901 10421 19935 10455
rect 1685 10217 1719 10251
rect 5457 10217 5491 10251
rect 5825 10217 5859 10251
rect 7389 10217 7423 10251
rect 9873 10217 9907 10251
rect 10885 10217 10919 10251
rect 13553 10217 13587 10251
rect 14289 10217 14323 10251
rect 15853 10217 15887 10251
rect 17325 10217 17359 10251
rect 19349 10217 19383 10251
rect 2099 10149 2133 10183
rect 6101 10149 6135 10183
rect 7665 10149 7699 10183
rect 10195 10149 10229 10183
rect 11253 10149 11287 10183
rect 12081 10149 12115 10183
rect 12995 10149 13029 10183
rect 16767 10149 16801 10183
rect 18521 10149 18555 10183
rect 1996 10081 2030 10115
rect 2973 10081 3007 10115
rect 4537 10081 4571 10115
rect 4813 10081 4847 10115
rect 10092 10081 10126 10115
rect 12449 10081 12483 10115
rect 12633 10081 12667 10115
rect 15301 10081 15335 10115
rect 5089 10013 5123 10047
rect 6009 10013 6043 10047
rect 7573 10013 7607 10047
rect 7849 10013 7883 10047
rect 11161 10013 11195 10047
rect 16405 10013 16439 10047
rect 18429 10013 18463 10047
rect 18797 10013 18831 10047
rect 3111 9945 3145 9979
rect 6561 9945 6595 9979
rect 11713 9945 11747 9979
rect 15485 9945 15519 9979
rect 3617 9877 3651 9911
rect 6929 9877 6963 9911
rect 8677 9877 8711 9911
rect 10609 9877 10643 9911
rect 13829 9877 13863 9911
rect 16313 9877 16347 9911
rect 2329 9673 2363 9707
rect 4905 9673 4939 9707
rect 5089 9673 5123 9707
rect 6193 9673 6227 9707
rect 12817 9673 12851 9707
rect 14657 9673 14691 9707
rect 15301 9673 15335 9707
rect 17417 9673 17451 9707
rect 19073 9673 19107 9707
rect 1593 9605 1627 9639
rect 2743 9605 2777 9639
rect 9689 9605 9723 9639
rect 15945 9605 15979 9639
rect 4905 9537 4939 9571
rect 6837 9537 6871 9571
rect 8677 9537 8711 9571
rect 8953 9537 8987 9571
rect 10517 9537 10551 9571
rect 13737 9537 13771 9571
rect 16313 9537 16347 9571
rect 17141 9537 17175 9571
rect 18153 9537 18187 9571
rect 18429 9537 18463 9571
rect 19625 9537 19659 9571
rect 1409 9469 1443 9503
rect 1961 9469 1995 9503
rect 2640 9469 2674 9503
rect 3433 9469 3467 9503
rect 3617 9469 3651 9503
rect 4077 9469 4111 9503
rect 4629 9469 4663 9503
rect 7757 9469 7791 9503
rect 8033 9469 8067 9503
rect 12633 9469 12667 9503
rect 13001 9469 13035 9503
rect 5273 9401 5307 9435
rect 5365 9401 5399 9435
rect 5917 9401 5951 9435
rect 7158 9401 7192 9435
rect 8769 9401 8803 9435
rect 10879 9401 10913 9435
rect 12173 9401 12207 9435
rect 13553 9401 13587 9435
rect 14058 9401 14092 9435
rect 16497 9401 16531 9435
rect 16589 9401 16623 9435
rect 18245 9401 18279 9435
rect 3065 9333 3099 9367
rect 3893 9333 3927 9367
rect 6561 9333 6595 9367
rect 8401 9333 8435 9367
rect 10057 9333 10091 9367
rect 11437 9333 11471 9367
rect 11805 9333 11839 9367
rect 13001 9333 13035 9367
rect 13277 9333 13311 9367
rect 17877 9333 17911 9367
rect 19533 9333 19567 9367
rect 3111 9129 3145 9163
rect 3801 9129 3835 9163
rect 4629 9129 4663 9163
rect 5089 9129 5123 9163
rect 6193 9129 6227 9163
rect 8309 9129 8343 9163
rect 10609 9129 10643 9163
rect 12633 9129 12667 9163
rect 16037 9129 16071 9163
rect 16957 9129 16991 9163
rect 17509 9129 17543 9163
rect 18153 9129 18187 9163
rect 19257 9129 19291 9163
rect 2099 9061 2133 9095
rect 1961 8993 1995 9027
rect 2881 8993 2915 9027
rect 3040 8993 3074 9027
rect 7107 9061 7141 9095
rect 7941 9061 7975 9095
rect 8769 9061 8803 9095
rect 11345 9061 11379 9095
rect 13829 9061 13863 9095
rect 14381 9061 14415 9095
rect 18658 9061 18692 9095
rect 5365 8993 5399 9027
rect 5641 8993 5675 9027
rect 7665 8993 7699 9027
rect 8493 8993 8527 9027
rect 10057 8993 10091 9027
rect 15485 8993 15519 9027
rect 4169 8925 4203 8959
rect 5917 8925 5951 8959
rect 6745 8925 6779 8959
rect 11253 8925 11287 8959
rect 11897 8925 11931 8959
rect 13461 8925 13495 8959
rect 13737 8925 13771 8959
rect 16589 8925 16623 8959
rect 18337 8925 18371 8959
rect 3801 8857 3835 8891
rect 10241 8857 10275 8891
rect 15669 8857 15703 8891
rect 3709 8789 3743 8823
rect 6561 8789 6595 8823
rect 10977 8789 11011 8823
rect 16405 8789 16439 8823
rect 1961 8585 1995 8619
rect 6285 8585 6319 8619
rect 7389 8585 7423 8619
rect 9045 8585 9079 8619
rect 10425 8585 10459 8619
rect 11253 8585 11287 8619
rect 13737 8585 13771 8619
rect 15485 8585 15519 8619
rect 17785 8585 17819 8619
rect 19165 8585 19199 8619
rect 4077 8517 4111 8551
rect 4537 8517 4571 8551
rect 7021 8517 7055 8551
rect 12173 8517 12207 8551
rect 13093 8517 13127 8551
rect 18797 8517 18831 8551
rect 4629 8449 4663 8483
rect 7757 8449 7791 8483
rect 8033 8449 8067 8483
rect 9229 8449 9263 8483
rect 12541 8449 12575 8483
rect 14749 8449 14783 8483
rect 16681 8449 16715 8483
rect 18245 8449 18279 8483
rect 2099 8381 2133 8415
rect 3341 8381 3375 8415
rect 3617 8381 3651 8415
rect 3801 8381 3835 8415
rect 11161 8381 11195 8415
rect 11805 8381 11839 8415
rect 15945 8381 15979 8415
rect 16405 8381 16439 8415
rect 2191 8313 2225 8347
rect 4991 8313 5025 8347
rect 7858 8313 7892 8347
rect 9505 8313 9539 8347
rect 10885 8313 10919 8347
rect 10977 8313 11011 8347
rect 12633 8313 12667 8347
rect 14197 8313 14231 8347
rect 14473 8313 14507 8347
rect 14565 8313 14599 8347
rect 18337 8313 18371 8347
rect 2605 8245 2639 8279
rect 2973 8245 3007 8279
rect 5549 8245 5583 8279
rect 5825 8245 5859 8279
rect 8677 8245 8711 8279
rect 10149 8245 10183 8279
rect 16957 8245 16991 8279
rect 17417 8245 17451 8279
rect 19625 8245 19659 8279
rect 2513 8041 2547 8075
rect 2881 8041 2915 8075
rect 3433 8041 3467 8075
rect 4721 8041 4755 8075
rect 5917 8041 5951 8075
rect 8861 8041 8895 8075
rect 9229 8041 9263 8075
rect 9873 8041 9907 8075
rect 13645 8041 13679 8075
rect 14197 8041 14231 8075
rect 18981 8041 19015 8075
rect 3617 7973 3651 8007
rect 4261 7973 4295 8007
rect 4997 7973 5031 8007
rect 5089 7973 5123 8007
rect 5733 7973 5767 8007
rect 8033 7973 8067 8007
rect 11247 7973 11281 8007
rect 16865 7973 16899 8007
rect 17509 7973 17543 8007
rect 18705 7973 18739 8007
rect 2012 7905 2046 7939
rect 3040 7905 3074 7939
rect 2099 7837 2133 7871
rect 1869 7769 1903 7803
rect 3111 7769 3145 7803
rect 6904 7905 6938 7939
rect 7665 7905 7699 7939
rect 13277 7905 13311 7939
rect 15761 7905 15795 7939
rect 16313 7905 16347 7939
rect 18889 7905 18923 7939
rect 19349 7905 19383 7939
rect 7941 7837 7975 7871
rect 8217 7837 8251 7871
rect 10885 7837 10919 7871
rect 16497 7837 16531 7871
rect 17417 7837 17451 7871
rect 18337 7837 18371 7871
rect 5549 7769 5583 7803
rect 5733 7769 5767 7803
rect 6975 7769 7009 7803
rect 17969 7769 18003 7803
rect 3617 7701 3651 7735
rect 3893 7701 3927 7735
rect 7297 7701 7331 7735
rect 11805 7701 11839 7735
rect 12449 7701 12483 7735
rect 12817 7701 12851 7735
rect 14565 7701 14599 7735
rect 17141 7701 17175 7735
rect 1961 7497 1995 7531
rect 3157 7497 3191 7531
rect 4629 7497 4663 7531
rect 6653 7497 6687 7531
rect 9873 7497 9907 7531
rect 11621 7497 11655 7531
rect 14657 7497 14691 7531
rect 15393 7497 15427 7531
rect 16129 7497 16163 7531
rect 17509 7497 17543 7531
rect 19763 7497 19797 7531
rect 3525 7429 3559 7463
rect 4353 7361 4387 7395
rect 6929 7361 6963 7395
rect 10057 7429 10091 7463
rect 14933 7429 14967 7463
rect 15853 7429 15887 7463
rect 17049 7429 17083 7463
rect 18705 7429 18739 7463
rect 10333 7361 10367 7395
rect 10609 7361 10643 7395
rect 13737 7361 13771 7395
rect 19441 7361 19475 7395
rect 2237 7293 2271 7327
rect 2605 7293 2639 7327
rect 3801 7293 3835 7327
rect 4077 7293 4111 7327
rect 5181 7293 5215 7327
rect 5641 7293 5675 7327
rect 5917 7293 5951 7327
rect 7849 7293 7883 7327
rect 8493 7293 8527 7327
rect 9413 7293 9447 7327
rect 9781 7293 9815 7327
rect 9873 7293 9907 7327
rect 12633 7293 12667 7327
rect 13185 7293 13219 7327
rect 19692 7293 19726 7327
rect 2789 7225 2823 7259
rect 7250 7225 7284 7259
rect 8769 7225 8803 7259
rect 8861 7225 8895 7259
rect 10425 7225 10459 7259
rect 11345 7225 11379 7259
rect 14058 7225 14092 7259
rect 16497 7225 16531 7259
rect 16589 7225 16623 7259
rect 18153 7225 18187 7259
rect 18245 7225 18279 7259
rect 5089 7157 5123 7191
rect 6285 7157 6319 7191
rect 8125 7157 8159 7191
rect 12817 7157 12851 7191
rect 13553 7157 13587 7191
rect 17877 7157 17911 7191
rect 19073 7157 19107 7191
rect 20085 7157 20119 7191
rect 1547 6953 1581 6987
rect 7481 6953 7515 6987
rect 8723 6953 8757 6987
rect 16773 6953 16807 6987
rect 17049 6953 17083 6987
rect 19533 6953 19567 6987
rect 2329 6885 2363 6919
rect 3709 6885 3743 6919
rect 6009 6885 6043 6919
rect 6882 6885 6916 6919
rect 9045 6885 9079 6919
rect 11621 6885 11655 6919
rect 11713 6885 11747 6919
rect 12265 6885 12299 6919
rect 14381 6885 14415 6919
rect 16215 6885 16249 6919
rect 17922 6885 17956 6919
rect 1476 6817 1510 6851
rect 2513 6817 2547 6851
rect 2881 6817 2915 6851
rect 5273 6817 5307 6851
rect 5549 6817 5583 6851
rect 5733 6817 5767 6851
rect 8652 6817 8686 6851
rect 9965 6817 9999 6851
rect 10241 6817 10275 6851
rect 13645 6817 13679 6851
rect 13921 6817 13955 6851
rect 19349 6817 19383 6851
rect 3157 6749 3191 6783
rect 6561 6749 6595 6783
rect 7941 6749 7975 6783
rect 10517 6749 10551 6783
rect 15853 6749 15887 6783
rect 17601 6749 17635 6783
rect 9413 6681 9447 6715
rect 10057 6681 10091 6715
rect 13737 6681 13771 6715
rect 1869 6613 1903 6647
rect 4261 6613 4295 6647
rect 4629 6613 4663 6647
rect 10977 6613 11011 6647
rect 13369 6613 13403 6647
rect 17417 6613 17451 6647
rect 18521 6613 18555 6647
rect 2881 6409 2915 6443
rect 3525 6409 3559 6443
rect 8033 6409 8067 6443
rect 11529 6409 11563 6443
rect 11805 6409 11839 6443
rect 14381 6409 14415 6443
rect 15485 6409 15519 6443
rect 19349 6409 19383 6443
rect 19763 6409 19797 6443
rect 1961 6341 1995 6375
rect 2145 6341 2179 6375
rect 12173 6341 12207 6375
rect 20085 6341 20119 6375
rect 2881 6273 2915 6307
rect 4353 6273 4387 6307
rect 10793 6273 10827 6307
rect 15025 6273 15059 6307
rect 16313 6273 16347 6307
rect 18429 6273 18463 6307
rect 2053 6205 2087 6239
rect 2329 6205 2363 6239
rect 3893 6205 3927 6239
rect 4077 6205 4111 6239
rect 4537 6205 4571 6239
rect 5089 6205 5123 6239
rect 5825 6205 5859 6239
rect 6193 6205 6227 6239
rect 6837 6205 6871 6239
rect 7297 6205 7331 6239
rect 10057 6205 10091 6239
rect 13277 6205 13311 6239
rect 14013 6205 14047 6239
rect 15577 6205 15611 6239
rect 16037 6205 16071 6239
rect 19676 6205 19710 6239
rect 3157 6137 3191 6171
rect 7573 6137 7607 6171
rect 8953 6137 8987 6171
rect 9054 6137 9088 6171
rect 9597 6137 9631 6171
rect 10517 6137 10551 6171
rect 10609 6137 10643 6171
rect 13369 6137 13403 6171
rect 17325 6137 17359 6171
rect 18153 6137 18187 6171
rect 18245 6137 18279 6171
rect 2513 6069 2547 6103
rect 4537 6069 4571 6103
rect 4629 6069 4663 6103
rect 5457 6069 5491 6103
rect 6653 6069 6687 6103
rect 8677 6069 8711 6103
rect 12909 6069 12943 6103
rect 16589 6069 16623 6103
rect 17601 6069 17635 6103
rect 4813 5865 4847 5899
rect 5733 5865 5767 5899
rect 6561 5865 6595 5899
rect 7021 5865 7055 5899
rect 7389 5865 7423 5899
rect 7849 5865 7883 5899
rect 9229 5865 9263 5899
rect 10701 5865 10735 5899
rect 14013 5865 14047 5899
rect 14197 5865 14231 5899
rect 19533 5865 19567 5899
rect 1547 5797 1581 5831
rect 9873 5797 9907 5831
rect 12081 5797 12115 5831
rect 13185 5797 13219 5831
rect 1460 5729 1494 5763
rect 1869 5729 1903 5763
rect 2421 5729 2455 5763
rect 2697 5729 2731 5763
rect 3617 5729 3651 5763
rect 4353 5729 4387 5763
rect 4629 5729 4663 5763
rect 5917 5729 5951 5763
rect 11437 5729 11471 5763
rect 12541 5729 12575 5763
rect 13461 5729 13495 5763
rect 3157 5661 3191 5695
rect 6285 5661 6319 5695
rect 7481 5661 7515 5695
rect 8953 5661 8987 5695
rect 9045 5661 9079 5695
rect 9781 5661 9815 5695
rect 10425 5661 10459 5695
rect 11069 5661 11103 5695
rect 2513 5593 2547 5627
rect 4445 5593 4479 5627
rect 6193 5593 6227 5627
rect 16129 5797 16163 5831
rect 16681 5797 16715 5831
rect 17693 5797 17727 5831
rect 18245 5797 18279 5831
rect 19073 5729 19107 5763
rect 19349 5729 19383 5763
rect 16037 5661 16071 5695
rect 17417 5661 17451 5695
rect 17601 5661 17635 5695
rect 15577 5593 15611 5627
rect 19165 5593 19199 5627
rect 2329 5525 2363 5559
rect 5365 5525 5399 5559
rect 6082 5525 6116 5559
rect 8401 5525 8435 5559
rect 9045 5525 9079 5559
rect 12817 5525 12851 5559
rect 14013 5525 14047 5559
rect 18521 5525 18555 5559
rect 1731 5321 1765 5355
rect 3065 5321 3099 5355
rect 4997 5321 5031 5355
rect 8585 5321 8619 5355
rect 11805 5321 11839 5355
rect 13737 5321 13771 5355
rect 13829 5321 13863 5355
rect 15301 5321 15335 5355
rect 16681 5321 16715 5355
rect 17509 5321 17543 5355
rect 19441 5321 19475 5355
rect 19763 5321 19797 5355
rect 5273 5253 5307 5287
rect 6653 5253 6687 5287
rect 13277 5253 13311 5287
rect 2513 5185 2547 5219
rect 3525 5185 3559 5219
rect 4077 5185 4111 5219
rect 5641 5185 5675 5219
rect 6285 5185 6319 5219
rect 9229 5185 9263 5219
rect 9873 5185 9907 5219
rect 12265 5185 12299 5219
rect 12541 5185 12575 5219
rect 1660 5117 1694 5151
rect 2605 5117 2639 5151
rect 3617 5117 3651 5151
rect 3709 5117 3743 5151
rect 3893 5117 3927 5151
rect 5181 5117 5215 5151
rect 5457 5117 5491 5151
rect 7389 5117 7423 5151
rect 10333 5117 10367 5151
rect 10793 5117 10827 5151
rect 10885 5117 10919 5151
rect 11069 5117 11103 5151
rect 12449 5117 12483 5151
rect 12725 5117 12759 5151
rect 4721 5049 4755 5083
rect 7710 5049 7744 5083
rect 9321 5049 9355 5083
rect 10609 5049 10643 5083
rect 16957 5253 16991 5287
rect 18153 5185 18187 5219
rect 13737 5117 13771 5151
rect 14105 5117 14139 5151
rect 15761 5117 15795 5151
rect 19676 5117 19710 5151
rect 20085 5117 20119 5151
rect 14013 5049 14047 5083
rect 15669 5049 15703 5083
rect 16123 5049 16157 5083
rect 18245 5049 18279 5083
rect 18797 5049 18831 5083
rect 2145 4981 2179 5015
rect 2743 4981 2777 5015
rect 7297 4981 7331 5015
rect 8309 4981 8343 5015
rect 9045 4981 9079 5015
rect 11253 4981 11287 5015
rect 12909 4981 12943 5015
rect 13277 4981 13311 5015
rect 13461 4981 13495 5015
rect 19073 4981 19107 5015
rect 3525 4777 3559 4811
rect 4445 4777 4479 4811
rect 6009 4777 6043 4811
rect 6285 4777 6319 4811
rect 9229 4777 9263 4811
rect 13001 4777 13035 4811
rect 17785 4777 17819 4811
rect 18153 4777 18187 4811
rect 18429 4777 18463 4811
rect 19625 4777 19659 4811
rect 3157 4709 3191 4743
rect 7205 4709 7239 4743
rect 7849 4709 7883 4743
rect 8217 4709 8251 4743
rect 9873 4709 9907 4743
rect 15485 4709 15519 4743
rect 17186 4709 17220 4743
rect 18797 4709 18831 4743
rect 1444 4641 1478 4675
rect 2421 4641 2455 4675
rect 2697 4641 2731 4675
rect 3801 4641 3835 4675
rect 4721 4641 4755 4675
rect 5181 4641 5215 4675
rect 5365 4641 5399 4675
rect 6469 4641 6503 4675
rect 7021 4641 7055 4675
rect 11805 4641 11839 4675
rect 11989 4641 12023 4675
rect 12265 4641 12299 4675
rect 13553 4641 13587 4675
rect 13737 4641 13771 4675
rect 5641 4573 5675 4607
rect 8125 4573 8159 4607
rect 8769 4573 8803 4607
rect 9781 4573 9815 4607
rect 10057 4573 10091 4607
rect 12449 4573 12483 4607
rect 14381 4573 14415 4607
rect 15393 4573 15427 4607
rect 16037 4573 16071 4607
rect 16865 4573 16899 4607
rect 18705 4573 18739 4607
rect 18981 4573 19015 4607
rect 2145 4505 2179 4539
rect 2513 4505 2547 4539
rect 12081 4505 12115 4539
rect 16313 4505 16347 4539
rect 1547 4437 1581 4471
rect 7481 4437 7515 4471
rect 10793 4437 10827 4471
rect 11437 4437 11471 4471
rect 9137 4233 9171 4267
rect 10517 4233 10551 4267
rect 11483 4233 11517 4267
rect 15485 4233 15519 4267
rect 18981 4233 19015 4267
rect 19257 4233 19291 4267
rect 2145 4165 2179 4199
rect 4721 4165 4755 4199
rect 6469 4165 6503 4199
rect 11253 4165 11287 4199
rect 12081 4165 12115 4199
rect 14841 4165 14875 4199
rect 15117 4165 15151 4199
rect 1961 4097 1995 4131
rect 2789 4097 2823 4131
rect 5089 4097 5123 4131
rect 5917 4097 5951 4131
rect 2053 4029 2087 4063
rect 2329 4029 2363 4063
rect 3433 4029 3467 4063
rect 3893 4029 3927 4063
rect 4169 4029 4203 4063
rect 4353 4029 4387 4063
rect 5181 4029 5215 4063
rect 5641 4029 5675 4063
rect 6193 4029 6227 4063
rect 9597 4097 9631 4131
rect 10793 4097 10827 4131
rect 13737 4097 13771 4131
rect 7113 4029 7147 4063
rect 8033 4029 8067 4063
rect 11380 4029 11414 4063
rect 12725 4029 12759 4063
rect 13461 4029 13495 4063
rect 13921 4029 13955 4063
rect 18061 4029 18095 4063
rect 6469 3961 6503 3995
rect 9918 3961 9952 3995
rect 12541 3961 12575 3995
rect 14242 3961 14276 3995
rect 15761 3961 15795 3995
rect 15853 3961 15887 3995
rect 16405 3961 16439 3995
rect 17785 3961 17819 3995
rect 18382 3961 18416 3995
rect 3065 3893 3099 3927
rect 6653 3893 6687 3927
rect 7481 3893 7515 3927
rect 8309 3893 8343 3927
rect 8769 3893 8803 3927
rect 9413 3893 9447 3927
rect 12817 3893 12851 3927
rect 16957 3893 16991 3927
rect 17233 3893 17267 3927
rect 2881 3689 2915 3723
rect 3525 3689 3559 3723
rect 3801 3689 3835 3723
rect 4261 3689 4295 3723
rect 5917 3689 5951 3723
rect 11897 3689 11931 3723
rect 12541 3689 12575 3723
rect 14197 3689 14231 3723
rect 14657 3689 14691 3723
rect 15485 3689 15519 3723
rect 16681 3689 16715 3723
rect 18613 3689 18647 3723
rect 19073 3689 19107 3723
rect 1409 3621 1443 3655
rect 4813 3621 4847 3655
rect 6285 3621 6319 3655
rect 7205 3621 7239 3655
rect 7849 3621 7883 3655
rect 8125 3621 8159 3655
rect 8217 3621 8251 3655
rect 9873 3621 9907 3655
rect 11161 3621 11195 3655
rect 15761 3621 15795 3655
rect 15853 3621 15887 3655
rect 2421 3553 2455 3587
rect 2697 3553 2731 3587
rect 5549 3553 5583 3587
rect 6469 3553 6503 3587
rect 6929 3553 6963 3587
rect 7481 3553 7515 3587
rect 11437 3553 11471 3587
rect 11713 3553 11747 3587
rect 13093 3553 13127 3587
rect 13277 3553 13311 3587
rect 14105 3553 14139 3587
rect 14289 3553 14323 3587
rect 16405 3553 16439 3587
rect 17325 3553 17359 3587
rect 18797 3553 18831 3587
rect 19257 3553 19291 3587
rect 5641 3485 5675 3519
rect 8769 3485 8803 3519
rect 9781 3485 9815 3519
rect 17233 3485 17267 3519
rect 2513 3417 2547 3451
rect 10333 3417 10367 3451
rect 10885 3417 10919 3451
rect 11529 3417 11563 3451
rect 2145 3349 2179 3383
rect 9045 3349 9079 3383
rect 9413 3349 9447 3383
rect 15025 3349 15059 3383
rect 18245 3349 18279 3383
rect 3065 3145 3099 3179
rect 3433 3145 3467 3179
rect 4997 3145 5031 3179
rect 6469 3145 6503 3179
rect 9137 3145 9171 3179
rect 9873 3145 9907 3179
rect 10149 3145 10183 3179
rect 11621 3145 11655 3179
rect 12265 3145 12299 3179
rect 12633 3145 12667 3179
rect 14565 3145 14599 3179
rect 17049 3145 17083 3179
rect 17417 3145 17451 3179
rect 19165 3145 19199 3179
rect 7941 3077 7975 3111
rect 9413 3077 9447 3111
rect 10885 3077 10919 3111
rect 2789 3009 2823 3043
rect 2329 2941 2363 2975
rect 2605 2941 2639 2975
rect 3801 2941 3835 2975
rect 4169 2941 4203 2975
rect 5181 2941 5215 2975
rect 5733 2941 5767 2975
rect 5917 2941 5951 2975
rect 7113 2941 7147 2975
rect 7665 2941 7699 2975
rect 13001 3077 13035 3111
rect 15025 3077 15059 3111
rect 19763 3077 19797 3111
rect 8217 3009 8251 3043
rect 11529 3009 11563 3043
rect 11621 3009 11655 3043
rect 16405 3009 16439 3043
rect 18061 3009 18095 3043
rect 19441 3009 19475 3043
rect 10793 2941 10827 2975
rect 11069 2941 11103 2975
rect 13185 2941 13219 2975
rect 13645 2941 13679 2975
rect 14013 2941 14047 2975
rect 17877 2941 17911 2975
rect 18705 2941 18739 2975
rect 19692 2941 19726 2975
rect 20085 2941 20119 2975
rect 4353 2873 4387 2907
rect 7941 2873 7975 2907
rect 8579 2873 8613 2907
rect 15485 2873 15519 2907
rect 16129 2873 16163 2907
rect 16221 2873 16255 2907
rect 1869 2805 1903 2839
rect 7297 2805 7331 2839
rect 8033 2805 8067 2839
rect 10609 2805 10643 2839
rect 11897 2805 11931 2839
rect 14289 2805 14323 2839
rect 15945 2805 15979 2839
rect 1869 2601 1903 2635
rect 2329 2601 2363 2635
rect 3433 2601 3467 2635
rect 3801 2601 3835 2635
rect 4813 2601 4847 2635
rect 6469 2601 6503 2635
rect 6929 2601 6963 2635
rect 9413 2601 9447 2635
rect 9505 2601 9539 2635
rect 10885 2601 10919 2635
rect 11253 2601 11287 2635
rect 13185 2601 13219 2635
rect 13553 2601 13587 2635
rect 14841 2601 14875 2635
rect 15623 2601 15657 2635
rect 4399 2533 4433 2567
rect 6009 2533 6043 2567
rect 7481 2533 7515 2567
rect 8262 2533 8296 2567
rect 9229 2533 9263 2567
rect 2697 2465 2731 2499
rect 2973 2465 3007 2499
rect 4169 2465 4203 2499
rect 5181 2465 5215 2499
rect 5365 2465 5399 2499
rect 8861 2465 8895 2499
rect 9965 2533 9999 2567
rect 13966 2533 14000 2567
rect 16818 2533 16852 2567
rect 17785 2533 17819 2567
rect 18521 2533 18555 2567
rect 11437 2465 11471 2499
rect 11989 2465 12023 2499
rect 12449 2465 12483 2499
rect 12668 2465 12702 2499
rect 13645 2465 13679 2499
rect 15552 2465 15586 2499
rect 15945 2465 15979 2499
rect 17417 2465 17451 2499
rect 1409 2397 1443 2431
rect 3157 2397 3191 2431
rect 4997 2397 5031 2431
rect 7941 2397 7975 2431
rect 9413 2397 9447 2431
rect 9873 2397 9907 2431
rect 10333 2397 10367 2431
rect 12771 2397 12805 2431
rect 16497 2397 16531 2431
rect 18429 2397 18463 2431
rect 18705 2397 18739 2431
rect 11621 2329 11655 2363
rect 16313 2329 16347 2363
rect 4997 2261 5031 2295
rect 7757 2261 7791 2295
rect 14565 2261 14599 2295
rect 15209 2261 15243 2295
rect 18061 2261 18095 2295
<< metal1 >>
rect 1104 19610 20884 19632
rect 1104 19558 4648 19610
rect 4700 19558 4712 19610
rect 4764 19558 4776 19610
rect 4828 19558 4840 19610
rect 4892 19558 11982 19610
rect 12034 19558 12046 19610
rect 12098 19558 12110 19610
rect 12162 19558 12174 19610
rect 12226 19558 19315 19610
rect 19367 19558 19379 19610
rect 19431 19558 19443 19610
rect 19495 19558 19507 19610
rect 19559 19558 20884 19610
rect 1104 19536 20884 19558
rect 15611 19499 15669 19505
rect 15611 19465 15623 19499
rect 15657 19496 15669 19499
rect 15746 19496 15752 19508
rect 15657 19468 15752 19496
rect 15657 19465 15669 19468
rect 15611 19459 15669 19465
rect 15746 19456 15752 19468
rect 15804 19456 15810 19508
rect 13909 19363 13967 19369
rect 13909 19360 13921 19363
rect 13786 19332 13921 19360
rect 13786 19304 13814 19332
rect 13909 19329 13921 19332
rect 13955 19360 13967 19363
rect 13955 19332 16620 19360
rect 13955 19329 13967 19332
rect 13909 19323 13967 19329
rect 13424 19295 13482 19301
rect 13424 19261 13436 19295
rect 13470 19292 13482 19295
rect 13786 19292 13820 19304
rect 13470 19264 13820 19292
rect 13470 19261 13482 19264
rect 13424 19255 13482 19261
rect 13814 19252 13820 19264
rect 13872 19252 13878 19304
rect 14436 19295 14494 19301
rect 14436 19261 14448 19295
rect 14482 19292 14494 19295
rect 14482 19264 14872 19292
rect 14482 19261 14494 19264
rect 14436 19255 14494 19261
rect 13998 19224 14004 19236
rect 13786 19196 14004 19224
rect 13495 19159 13553 19165
rect 13495 19125 13507 19159
rect 13541 19156 13553 19159
rect 13786 19156 13814 19196
rect 13998 19184 14004 19196
rect 14056 19184 14062 19236
rect 14844 19168 14872 19264
rect 15102 19252 15108 19304
rect 15160 19292 15166 19304
rect 15508 19295 15566 19301
rect 15508 19292 15520 19295
rect 15160 19264 15520 19292
rect 15160 19252 15166 19264
rect 15508 19261 15520 19264
rect 15554 19292 15566 19295
rect 15933 19295 15991 19301
rect 15933 19292 15945 19295
rect 15554 19264 15945 19292
rect 15554 19261 15566 19264
rect 15508 19255 15566 19261
rect 15933 19261 15945 19264
rect 15979 19261 15991 19295
rect 16592 19292 16620 19332
rect 17288 19295 17346 19301
rect 17288 19292 17300 19295
rect 16592 19264 17300 19292
rect 15933 19255 15991 19261
rect 17288 19261 17300 19264
rect 17334 19292 17346 19295
rect 17862 19292 17868 19304
rect 17334 19264 17868 19292
rect 17334 19261 17346 19264
rect 17288 19255 17346 19261
rect 17862 19252 17868 19264
rect 17920 19252 17926 19304
rect 18392 19295 18450 19301
rect 18392 19261 18404 19295
rect 18438 19292 18450 19295
rect 18601 19295 18659 19301
rect 18601 19292 18613 19295
rect 18438 19264 18613 19292
rect 18438 19261 18450 19264
rect 18392 19255 18450 19261
rect 18601 19261 18613 19264
rect 18647 19261 18659 19295
rect 19372 19295 19430 19301
rect 19372 19292 19384 19295
rect 18601 19255 18659 19261
rect 18845 19264 19384 19292
rect 17126 19184 17132 19236
rect 17184 19224 17190 19236
rect 18845 19224 18873 19264
rect 19372 19261 19384 19264
rect 19418 19292 19430 19295
rect 19797 19295 19855 19301
rect 19797 19292 19809 19295
rect 19418 19264 19809 19292
rect 19418 19261 19430 19264
rect 19372 19255 19430 19261
rect 19797 19261 19809 19264
rect 19843 19261 19855 19295
rect 19797 19255 19855 19261
rect 17184 19196 18873 19224
rect 19475 19227 19533 19233
rect 17184 19184 17190 19196
rect 19475 19193 19487 19227
rect 19521 19224 19533 19227
rect 20622 19224 20628 19236
rect 19521 19196 20628 19224
rect 19521 19193 19533 19196
rect 19475 19187 19533 19193
rect 20622 19184 20628 19196
rect 20680 19184 20686 19236
rect 13541 19128 13814 19156
rect 13541 19125 13553 19128
rect 13495 19119 13553 19125
rect 14274 19116 14280 19168
rect 14332 19156 14338 19168
rect 14507 19159 14565 19165
rect 14507 19156 14519 19159
rect 14332 19128 14519 19156
rect 14332 19116 14338 19128
rect 14507 19125 14519 19128
rect 14553 19125 14565 19159
rect 14826 19156 14832 19168
rect 14787 19128 14832 19156
rect 14507 19119 14565 19125
rect 14826 19116 14832 19128
rect 14884 19116 14890 19168
rect 17359 19159 17417 19165
rect 17359 19125 17371 19159
rect 17405 19156 17417 19159
rect 17586 19156 17592 19168
rect 17405 19128 17592 19156
rect 17405 19125 17417 19128
rect 17359 19119 17417 19125
rect 17586 19116 17592 19128
rect 17644 19116 17650 19168
rect 17773 19159 17831 19165
rect 17773 19125 17785 19159
rect 17819 19156 17831 19159
rect 17862 19156 17868 19168
rect 17819 19128 17868 19156
rect 17819 19125 17831 19128
rect 17773 19119 17831 19125
rect 17862 19116 17868 19128
rect 17920 19116 17926 19168
rect 18138 19116 18144 19168
rect 18196 19156 18202 19168
rect 18463 19159 18521 19165
rect 18463 19156 18475 19159
rect 18196 19128 18475 19156
rect 18196 19116 18202 19128
rect 18463 19125 18475 19128
rect 18509 19125 18521 19159
rect 18463 19119 18521 19125
rect 18601 19159 18659 19165
rect 18601 19125 18613 19159
rect 18647 19156 18659 19159
rect 18877 19159 18935 19165
rect 18877 19156 18889 19159
rect 18647 19128 18889 19156
rect 18647 19125 18659 19128
rect 18601 19119 18659 19125
rect 18877 19125 18889 19128
rect 18923 19156 18935 19159
rect 19794 19156 19800 19168
rect 18923 19128 19800 19156
rect 18923 19125 18935 19128
rect 18877 19119 18935 19125
rect 19794 19116 19800 19128
rect 19852 19116 19858 19168
rect 1104 19066 20884 19088
rect 1104 19014 8315 19066
rect 8367 19014 8379 19066
rect 8431 19014 8443 19066
rect 8495 19014 8507 19066
rect 8559 19014 15648 19066
rect 15700 19014 15712 19066
rect 15764 19014 15776 19066
rect 15828 19014 15840 19066
rect 15892 19014 20884 19066
rect 1104 18992 20884 19014
rect 14323 18955 14381 18961
rect 14323 18921 14335 18955
rect 14369 18952 14381 18955
rect 14458 18952 14464 18964
rect 14369 18924 14464 18952
rect 14369 18921 14381 18924
rect 14323 18915 14381 18921
rect 14458 18912 14464 18924
rect 14516 18912 14522 18964
rect 12299 18887 12357 18893
rect 12299 18853 12311 18887
rect 12345 18884 12357 18887
rect 21634 18884 21640 18896
rect 12345 18856 21640 18884
rect 12345 18853 12357 18856
rect 12299 18847 12357 18853
rect 21634 18844 21640 18856
rect 21692 18844 21698 18896
rect 11882 18776 11888 18828
rect 11940 18816 11946 18828
rect 12196 18819 12254 18825
rect 12196 18816 12208 18819
rect 11940 18788 12208 18816
rect 11940 18776 11946 18788
rect 12196 18785 12208 18788
rect 12242 18785 12254 18819
rect 12196 18779 12254 18785
rect 13240 18819 13298 18825
rect 13240 18785 13252 18819
rect 13286 18816 13298 18819
rect 13446 18816 13452 18828
rect 13286 18788 13452 18816
rect 13286 18785 13298 18788
rect 13240 18779 13298 18785
rect 13446 18776 13452 18788
rect 13504 18776 13510 18828
rect 14252 18819 14310 18825
rect 14252 18785 14264 18819
rect 14298 18816 14310 18819
rect 14550 18816 14556 18828
rect 14298 18788 14556 18816
rect 14298 18785 14310 18788
rect 14252 18779 14310 18785
rect 14550 18776 14556 18788
rect 14608 18776 14614 18828
rect 16022 18816 16028 18828
rect 15983 18788 16028 18816
rect 16022 18776 16028 18788
rect 16080 18776 16086 18828
rect 16298 18816 16304 18828
rect 16259 18788 16304 18816
rect 16298 18776 16304 18788
rect 16356 18776 16362 18828
rect 17494 18776 17500 18828
rect 17552 18816 17558 18828
rect 17624 18819 17682 18825
rect 17624 18816 17636 18819
rect 17552 18788 17636 18816
rect 17552 18776 17558 18788
rect 17624 18785 17636 18788
rect 17670 18785 17682 18819
rect 18598 18816 18604 18828
rect 18559 18788 18604 18816
rect 17624 18779 17682 18785
rect 18598 18776 18604 18788
rect 18656 18776 18662 18828
rect 19680 18819 19738 18825
rect 19680 18785 19692 18819
rect 19726 18816 19738 18819
rect 19978 18816 19984 18828
rect 19726 18788 19984 18816
rect 19726 18785 19738 18788
rect 19680 18779 19738 18785
rect 19978 18776 19984 18788
rect 20036 18776 20042 18828
rect 16482 18748 16488 18760
rect 16443 18720 16488 18748
rect 16482 18708 16488 18720
rect 16540 18708 16546 18760
rect 16942 18640 16948 18692
rect 17000 18680 17006 18692
rect 18739 18683 18797 18689
rect 18739 18680 18751 18683
rect 17000 18652 18751 18680
rect 17000 18640 17006 18652
rect 18739 18649 18751 18652
rect 18785 18649 18797 18683
rect 18739 18643 18797 18649
rect 12618 18612 12624 18624
rect 12579 18584 12624 18612
rect 12618 18572 12624 18584
rect 12676 18572 12682 18624
rect 13311 18615 13369 18621
rect 13311 18581 13323 18615
rect 13357 18612 13369 18615
rect 13630 18612 13636 18624
rect 13357 18584 13636 18612
rect 13357 18581 13369 18584
rect 13311 18575 13369 18581
rect 13630 18572 13636 18584
rect 13688 18572 13694 18624
rect 15562 18612 15568 18624
rect 15523 18584 15568 18612
rect 15562 18572 15568 18584
rect 15620 18572 15626 18624
rect 17727 18615 17785 18621
rect 17727 18581 17739 18615
rect 17773 18612 17785 18615
rect 17954 18612 17960 18624
rect 17773 18584 17960 18612
rect 17773 18581 17785 18584
rect 17727 18575 17785 18581
rect 17954 18572 17960 18584
rect 18012 18572 18018 18624
rect 19751 18615 19809 18621
rect 19751 18581 19763 18615
rect 19797 18612 19809 18615
rect 21542 18612 21548 18624
rect 19797 18584 21548 18612
rect 19797 18581 19809 18584
rect 19751 18575 19809 18581
rect 21542 18572 21548 18584
rect 21600 18572 21606 18624
rect 1104 18522 20884 18544
rect 1104 18470 4648 18522
rect 4700 18470 4712 18522
rect 4764 18470 4776 18522
rect 4828 18470 4840 18522
rect 4892 18470 11982 18522
rect 12034 18470 12046 18522
rect 12098 18470 12110 18522
rect 12162 18470 12174 18522
rect 12226 18470 19315 18522
rect 19367 18470 19379 18522
rect 19431 18470 19443 18522
rect 19495 18470 19507 18522
rect 19559 18470 20884 18522
rect 1104 18448 20884 18470
rect 1578 18408 1584 18420
rect 1539 18380 1584 18408
rect 1578 18368 1584 18380
rect 1636 18368 1642 18420
rect 2041 18411 2099 18417
rect 2041 18377 2053 18411
rect 2087 18408 2099 18411
rect 2774 18408 2780 18420
rect 2087 18380 2780 18408
rect 2087 18377 2099 18380
rect 2041 18371 2099 18377
rect 1397 18207 1455 18213
rect 1397 18173 1409 18207
rect 1443 18204 1455 18207
rect 2056 18204 2084 18371
rect 2774 18368 2780 18380
rect 2832 18408 2838 18420
rect 3326 18408 3332 18420
rect 2832 18380 3332 18408
rect 2832 18368 2838 18380
rect 3326 18368 3332 18380
rect 3384 18368 3390 18420
rect 8113 18411 8171 18417
rect 8113 18377 8125 18411
rect 8159 18408 8171 18411
rect 8202 18408 8208 18420
rect 8159 18380 8208 18408
rect 8159 18377 8171 18380
rect 8113 18371 8171 18377
rect 8202 18368 8208 18380
rect 8260 18368 8266 18420
rect 13446 18408 13452 18420
rect 9646 18380 13452 18408
rect 7374 18300 7380 18352
rect 7432 18340 7438 18352
rect 9646 18340 9674 18380
rect 13446 18368 13452 18380
rect 13504 18408 13510 18420
rect 13541 18411 13599 18417
rect 13541 18408 13553 18411
rect 13504 18380 13553 18408
rect 13504 18368 13510 18380
rect 13541 18377 13553 18380
rect 13587 18377 13599 18411
rect 13541 18371 13599 18377
rect 14553 18411 14611 18417
rect 14553 18377 14565 18411
rect 14599 18408 14611 18411
rect 15930 18408 15936 18420
rect 14599 18380 15936 18408
rect 14599 18377 14611 18380
rect 14553 18371 14611 18377
rect 15930 18368 15936 18380
rect 15988 18368 15994 18420
rect 18233 18411 18291 18417
rect 18233 18377 18245 18411
rect 18279 18408 18291 18411
rect 18322 18408 18328 18420
rect 18279 18380 18328 18408
rect 18279 18377 18291 18380
rect 18233 18371 18291 18377
rect 18322 18368 18328 18380
rect 18380 18368 18386 18420
rect 19978 18408 19984 18420
rect 19939 18380 19984 18408
rect 19978 18368 19984 18380
rect 20036 18368 20042 18420
rect 7432 18312 9674 18340
rect 7432 18300 7438 18312
rect 10870 18300 10876 18352
rect 10928 18340 10934 18352
rect 18598 18340 18604 18352
rect 10928 18312 18604 18340
rect 10928 18300 10934 18312
rect 18598 18300 18604 18312
rect 18656 18340 18662 18352
rect 18969 18343 19027 18349
rect 18969 18340 18981 18343
rect 18656 18312 18981 18340
rect 18656 18300 18662 18312
rect 18969 18309 18981 18312
rect 19015 18309 19027 18343
rect 18969 18303 19027 18309
rect 1443 18176 2084 18204
rect 7929 18207 7987 18213
rect 1443 18173 1455 18176
rect 1397 18167 1455 18173
rect 7929 18173 7941 18207
rect 7975 18173 7987 18207
rect 7929 18167 7987 18173
rect 10480 18207 10538 18213
rect 10480 18173 10492 18207
rect 10526 18173 10538 18207
rect 10480 18167 10538 18173
rect 7944 18136 7972 18167
rect 8573 18139 8631 18145
rect 8573 18136 8585 18139
rect 7944 18108 8585 18136
rect 8573 18105 8585 18108
rect 8619 18136 8631 18139
rect 9582 18136 9588 18148
rect 8619 18108 9588 18136
rect 8619 18105 8631 18108
rect 8573 18099 8631 18105
rect 9582 18096 9588 18108
rect 9640 18096 9646 18148
rect 10495 18136 10523 18167
rect 10594 18164 10600 18216
rect 10652 18204 10658 18216
rect 12529 18207 12587 18213
rect 12529 18204 12541 18207
rect 10652 18176 12541 18204
rect 10652 18164 10658 18176
rect 12529 18173 12541 18176
rect 12575 18204 12587 18207
rect 12618 18204 12624 18216
rect 12575 18176 12624 18204
rect 12575 18173 12587 18176
rect 12529 18167 12587 18173
rect 12618 18164 12624 18176
rect 12676 18164 12682 18216
rect 12989 18207 13047 18213
rect 12989 18173 13001 18207
rect 13035 18204 13047 18207
rect 13170 18204 13176 18216
rect 13035 18176 13176 18204
rect 13035 18173 13047 18176
rect 12989 18167 13047 18173
rect 13170 18164 13176 18176
rect 13228 18164 13234 18216
rect 14366 18204 14372 18216
rect 14327 18176 14372 18204
rect 14366 18164 14372 18176
rect 14424 18204 14430 18216
rect 14826 18204 14832 18216
rect 14424 18176 14832 18204
rect 14424 18164 14430 18176
rect 14826 18164 14832 18176
rect 14884 18204 14890 18216
rect 14921 18207 14979 18213
rect 14921 18204 14933 18207
rect 14884 18176 14933 18204
rect 14884 18164 14890 18176
rect 14921 18173 14933 18176
rect 14967 18173 14979 18207
rect 14921 18167 14979 18173
rect 15562 18164 15568 18216
rect 15620 18204 15626 18216
rect 15749 18207 15807 18213
rect 15749 18204 15761 18207
rect 15620 18176 15761 18204
rect 15620 18164 15626 18176
rect 15749 18173 15761 18176
rect 15795 18204 15807 18207
rect 15930 18204 15936 18216
rect 15795 18176 15936 18204
rect 15795 18173 15807 18176
rect 15749 18167 15807 18173
rect 15930 18164 15936 18176
rect 15988 18164 15994 18216
rect 16025 18207 16083 18213
rect 16025 18173 16037 18207
rect 16071 18173 16083 18207
rect 16025 18167 16083 18173
rect 18049 18207 18107 18213
rect 18049 18173 18061 18207
rect 18095 18204 18107 18207
rect 19220 18207 19278 18213
rect 18095 18176 18460 18204
rect 18095 18173 18107 18176
rect 18049 18167 18107 18173
rect 13262 18136 13268 18148
rect 10495 18108 11008 18136
rect 13223 18108 13268 18136
rect 10980 18080 11008 18108
rect 13262 18096 13268 18108
rect 13320 18096 13326 18148
rect 9306 18028 9312 18080
rect 9364 18068 9370 18080
rect 10551 18071 10609 18077
rect 10551 18068 10563 18071
rect 9364 18040 10563 18068
rect 9364 18028 9370 18040
rect 10551 18037 10563 18040
rect 10597 18037 10609 18071
rect 10962 18068 10968 18080
rect 10923 18040 10968 18068
rect 10551 18031 10609 18037
rect 10962 18028 10968 18040
rect 11020 18028 11026 18080
rect 11882 18068 11888 18080
rect 11843 18040 11888 18068
rect 11882 18028 11888 18040
rect 11940 18028 11946 18080
rect 12253 18071 12311 18077
rect 12253 18037 12265 18071
rect 12299 18068 12311 18071
rect 12342 18068 12348 18080
rect 12299 18040 12348 18068
rect 12299 18037 12311 18040
rect 12253 18031 12311 18037
rect 12342 18028 12348 18040
rect 12400 18028 12406 18080
rect 14277 18071 14335 18077
rect 14277 18037 14289 18071
rect 14323 18068 14335 18071
rect 14550 18068 14556 18080
rect 14323 18040 14556 18068
rect 14323 18037 14335 18040
rect 14277 18031 14335 18037
rect 14550 18028 14556 18040
rect 14608 18028 14614 18080
rect 15381 18071 15439 18077
rect 15381 18037 15393 18071
rect 15427 18068 15439 18071
rect 15470 18068 15476 18080
rect 15427 18040 15476 18068
rect 15427 18037 15439 18040
rect 15381 18031 15439 18037
rect 15470 18028 15476 18040
rect 15528 18068 15534 18080
rect 16040 18068 16068 18167
rect 16114 18096 16120 18148
rect 16172 18136 16178 18148
rect 16209 18139 16267 18145
rect 16209 18136 16221 18139
rect 16172 18108 16221 18136
rect 16172 18096 16178 18108
rect 16209 18105 16221 18108
rect 16255 18105 16267 18139
rect 16209 18099 16267 18105
rect 16390 18096 16396 18148
rect 16448 18136 16454 18148
rect 17494 18136 17500 18148
rect 16448 18108 17500 18136
rect 16448 18096 16454 18108
rect 17494 18096 17500 18108
rect 17552 18136 17558 18148
rect 17589 18139 17647 18145
rect 17589 18136 17601 18139
rect 17552 18108 17601 18136
rect 17552 18096 17558 18108
rect 17589 18105 17601 18108
rect 17635 18105 17647 18139
rect 17589 18099 17647 18105
rect 18432 18080 18460 18176
rect 19220 18173 19232 18207
rect 19266 18204 19278 18207
rect 19266 18176 19656 18204
rect 19266 18173 19278 18176
rect 19220 18167 19278 18173
rect 19628 18080 19656 18176
rect 16298 18068 16304 18080
rect 15528 18040 16304 18068
rect 15528 18028 15534 18040
rect 16298 18028 16304 18040
rect 16356 18068 16362 18080
rect 16485 18071 16543 18077
rect 16485 18068 16497 18071
rect 16356 18040 16497 18068
rect 16356 18028 16362 18040
rect 16485 18037 16497 18040
rect 16531 18037 16543 18071
rect 16485 18031 16543 18037
rect 18414 18028 18420 18080
rect 18472 18068 18478 18080
rect 18601 18071 18659 18077
rect 18601 18068 18613 18071
rect 18472 18040 18613 18068
rect 18472 18028 18478 18040
rect 18601 18037 18613 18040
rect 18647 18037 18659 18071
rect 18601 18031 18659 18037
rect 19150 18028 19156 18080
rect 19208 18068 19214 18080
rect 19291 18071 19349 18077
rect 19291 18068 19303 18071
rect 19208 18040 19303 18068
rect 19208 18028 19214 18040
rect 19291 18037 19303 18040
rect 19337 18037 19349 18071
rect 19610 18068 19616 18080
rect 19571 18040 19616 18068
rect 19291 18031 19349 18037
rect 19610 18028 19616 18040
rect 19668 18028 19674 18080
rect 1104 17978 20884 18000
rect 1104 17926 8315 17978
rect 8367 17926 8379 17978
rect 8431 17926 8443 17978
rect 8495 17926 8507 17978
rect 8559 17926 15648 17978
rect 15700 17926 15712 17978
rect 15764 17926 15776 17978
rect 15828 17926 15840 17978
rect 15892 17926 20884 17978
rect 1104 17904 20884 17926
rect 15378 17864 15384 17876
rect 15339 17836 15384 17864
rect 15378 17824 15384 17836
rect 15436 17824 15442 17876
rect 16298 17824 16304 17876
rect 16356 17864 16362 17876
rect 16945 17867 17003 17873
rect 16945 17864 16957 17867
rect 16356 17836 16957 17864
rect 16356 17824 16362 17836
rect 16945 17833 16957 17836
rect 16991 17833 17003 17867
rect 18506 17864 18512 17876
rect 18467 17836 18512 17864
rect 16945 17827 17003 17833
rect 18506 17824 18512 17836
rect 18564 17824 18570 17876
rect 13538 17756 13544 17808
rect 13596 17796 13602 17808
rect 14090 17796 14096 17808
rect 13596 17768 14096 17796
rect 13596 17756 13602 17768
rect 14090 17756 14096 17768
rect 14148 17756 14154 17808
rect 15304 17768 16896 17796
rect 10505 17731 10563 17737
rect 10505 17697 10517 17731
rect 10551 17697 10563 17731
rect 10686 17728 10692 17740
rect 10647 17700 10692 17728
rect 10505 17691 10563 17697
rect 10520 17660 10548 17691
rect 10686 17688 10692 17700
rect 10744 17688 10750 17740
rect 12802 17728 12808 17740
rect 12763 17700 12808 17728
rect 12802 17688 12808 17700
rect 12860 17688 12866 17740
rect 13170 17728 13176 17740
rect 13131 17700 13176 17728
rect 13170 17688 13176 17700
rect 13228 17688 13234 17740
rect 14108 17728 14136 17756
rect 14220 17731 14278 17737
rect 14220 17728 14232 17731
rect 14108 17700 14232 17728
rect 14220 17697 14232 17700
rect 14266 17697 14278 17731
rect 14220 17691 14278 17697
rect 14918 17688 14924 17740
rect 14976 17728 14982 17740
rect 15304 17737 15332 17768
rect 16868 17737 16896 17768
rect 15289 17731 15347 17737
rect 15289 17728 15301 17731
rect 14976 17700 15301 17728
rect 14976 17688 14982 17700
rect 15289 17697 15301 17700
rect 15335 17697 15347 17731
rect 15289 17691 15347 17697
rect 15749 17731 15807 17737
rect 15749 17697 15761 17731
rect 15795 17697 15807 17731
rect 15749 17691 15807 17697
rect 16853 17731 16911 17737
rect 16853 17697 16865 17731
rect 16899 17728 16911 17731
rect 17218 17728 17224 17740
rect 16899 17700 17224 17728
rect 16899 17697 16911 17700
rect 16853 17691 16911 17697
rect 10594 17660 10600 17672
rect 10520 17632 10600 17660
rect 10594 17620 10600 17632
rect 10652 17620 10658 17672
rect 10778 17660 10784 17672
rect 10739 17632 10784 17660
rect 10778 17620 10784 17632
rect 10836 17620 10842 17672
rect 13354 17660 13360 17672
rect 13315 17632 13360 17660
rect 13354 17620 13360 17632
rect 13412 17620 13418 17672
rect 15194 17620 15200 17672
rect 15252 17660 15258 17672
rect 15764 17660 15792 17691
rect 17218 17688 17224 17700
rect 17276 17688 17282 17740
rect 17310 17688 17316 17740
rect 17368 17728 17374 17740
rect 18690 17728 18696 17740
rect 17368 17700 17413 17728
rect 18651 17700 18696 17728
rect 17368 17688 17374 17700
rect 18690 17688 18696 17700
rect 18748 17688 18754 17740
rect 18874 17728 18880 17740
rect 18835 17700 18880 17728
rect 18874 17688 18880 17700
rect 18932 17688 18938 17740
rect 15252 17632 15792 17660
rect 15252 17620 15258 17632
rect 12802 17552 12808 17604
rect 12860 17592 12866 17604
rect 16022 17592 16028 17604
rect 12860 17564 16028 17592
rect 12860 17552 12866 17564
rect 16022 17552 16028 17564
rect 16080 17592 16086 17604
rect 16301 17595 16359 17601
rect 16301 17592 16313 17595
rect 16080 17564 16313 17592
rect 16080 17552 16086 17564
rect 16301 17561 16313 17564
rect 16347 17561 16359 17595
rect 16301 17555 16359 17561
rect 12529 17527 12587 17533
rect 12529 17493 12541 17527
rect 12575 17524 12587 17527
rect 12710 17524 12716 17536
rect 12575 17496 12716 17524
rect 12575 17493 12587 17496
rect 12529 17487 12587 17493
rect 12710 17484 12716 17496
rect 12768 17484 12774 17536
rect 13722 17484 13728 17536
rect 13780 17524 13786 17536
rect 14323 17527 14381 17533
rect 14323 17524 14335 17527
rect 13780 17496 14335 17524
rect 13780 17484 13786 17496
rect 14323 17493 14335 17496
rect 14369 17493 14381 17527
rect 14323 17487 14381 17493
rect 17770 17484 17776 17536
rect 17828 17524 17834 17536
rect 18049 17527 18107 17533
rect 18049 17524 18061 17527
rect 17828 17496 18061 17524
rect 17828 17484 17834 17496
rect 18049 17493 18061 17496
rect 18095 17493 18107 17527
rect 18049 17487 18107 17493
rect 1104 17434 20884 17456
rect 1104 17382 4648 17434
rect 4700 17382 4712 17434
rect 4764 17382 4776 17434
rect 4828 17382 4840 17434
rect 4892 17382 11982 17434
rect 12034 17382 12046 17434
rect 12098 17382 12110 17434
rect 12162 17382 12174 17434
rect 12226 17382 19315 17434
rect 19367 17382 19379 17434
rect 19431 17382 19443 17434
rect 19495 17382 19507 17434
rect 19559 17382 20884 17434
rect 1104 17360 20884 17382
rect 15194 17280 15200 17332
rect 15252 17320 15258 17332
rect 17218 17320 17224 17332
rect 15252 17292 16252 17320
rect 17179 17292 17224 17320
rect 15252 17280 15258 17292
rect 12618 17212 12624 17264
rect 12676 17252 12682 17264
rect 16224 17252 16252 17292
rect 17218 17280 17224 17292
rect 17276 17280 17282 17332
rect 19751 17255 19809 17261
rect 19751 17252 19763 17255
rect 12676 17224 15884 17252
rect 16224 17224 19763 17252
rect 12676 17212 12682 17224
rect 8527 17187 8585 17193
rect 8527 17153 8539 17187
rect 8573 17184 8585 17187
rect 11054 17184 11060 17196
rect 8573 17156 11060 17184
rect 8573 17153 8585 17156
rect 8527 17147 8585 17153
rect 11054 17144 11060 17156
rect 11112 17144 11118 17196
rect 12342 17144 12348 17196
rect 12400 17184 12406 17196
rect 14369 17187 14427 17193
rect 12400 17156 12940 17184
rect 12400 17144 12406 17156
rect 8440 17119 8498 17125
rect 8440 17085 8452 17119
rect 8486 17116 8498 17119
rect 9490 17116 9496 17128
rect 8486 17088 8708 17116
rect 9451 17088 9496 17116
rect 8486 17085 8498 17088
rect 8440 17079 8498 17085
rect 8680 16992 8708 17088
rect 9490 17076 9496 17088
rect 9548 17076 9554 17128
rect 9861 17119 9919 17125
rect 9861 17085 9873 17119
rect 9907 17085 9919 17119
rect 12710 17116 12716 17128
rect 12671 17088 12716 17116
rect 9861 17079 9919 17085
rect 9876 16992 9904 17079
rect 12710 17076 12716 17088
rect 12768 17076 12774 17128
rect 12912 17125 12940 17156
rect 14369 17153 14381 17187
rect 14415 17184 14427 17187
rect 14458 17184 14464 17196
rect 14415 17156 14464 17184
rect 14415 17153 14427 17156
rect 14369 17147 14427 17153
rect 14458 17144 14464 17156
rect 14516 17144 14522 17196
rect 12897 17119 12955 17125
rect 12897 17085 12909 17119
rect 12943 17116 12955 17119
rect 13170 17116 13176 17128
rect 12943 17088 13176 17116
rect 12943 17085 12955 17088
rect 12897 17079 12955 17085
rect 13170 17076 13176 17088
rect 13228 17116 13234 17128
rect 13449 17119 13507 17125
rect 13449 17116 13461 17119
rect 13228 17088 13461 17116
rect 13228 17076 13234 17088
rect 13449 17085 13461 17088
rect 13495 17116 13507 17119
rect 13538 17116 13544 17128
rect 13495 17088 13544 17116
rect 13495 17085 13507 17088
rect 13449 17079 13507 17085
rect 13538 17076 13544 17088
rect 13596 17076 13602 17128
rect 15856 17125 15884 17224
rect 19751 17221 19763 17224
rect 19797 17221 19809 17255
rect 19751 17215 19809 17221
rect 17862 17144 17868 17196
rect 17920 17184 17926 17196
rect 17920 17156 19723 17184
rect 17920 17144 17926 17156
rect 15841 17119 15899 17125
rect 15841 17085 15853 17119
rect 15887 17116 15899 17119
rect 16206 17116 16212 17128
rect 15887 17088 16212 17116
rect 15887 17085 15899 17088
rect 15841 17079 15899 17085
rect 16206 17076 16212 17088
rect 16264 17076 16270 17128
rect 16301 17119 16359 17125
rect 16301 17085 16313 17119
rect 16347 17116 16359 17119
rect 16853 17119 16911 17125
rect 16853 17116 16865 17119
rect 16347 17088 16865 17116
rect 16347 17085 16359 17088
rect 16301 17079 16359 17085
rect 16853 17085 16865 17088
rect 16899 17085 16911 17119
rect 16853 17079 16911 17085
rect 10134 17048 10140 17060
rect 10095 17020 10140 17048
rect 10134 17008 10140 17020
rect 10192 17008 10198 17060
rect 10594 17008 10600 17060
rect 10652 17048 10658 17060
rect 10781 17051 10839 17057
rect 10781 17048 10793 17051
rect 10652 17020 10793 17048
rect 10652 17008 10658 17020
rect 10781 17017 10793 17020
rect 10827 17017 10839 17051
rect 10781 17011 10839 17017
rect 14461 17051 14519 17057
rect 14461 17017 14473 17051
rect 14507 17048 14519 17051
rect 14642 17048 14648 17060
rect 14507 17020 14648 17048
rect 14507 17017 14519 17020
rect 14461 17011 14519 17017
rect 14642 17008 14648 17020
rect 14700 17008 14706 17060
rect 15013 17051 15071 17057
rect 15013 17017 15025 17051
rect 15059 17048 15071 17051
rect 15102 17048 15108 17060
rect 15059 17020 15108 17048
rect 15059 17017 15071 17020
rect 15013 17011 15071 17017
rect 15102 17008 15108 17020
rect 15160 17008 15166 17060
rect 16316 17048 16344 17079
rect 16574 17048 16580 17060
rect 15672 17020 16344 17048
rect 16535 17020 16580 17048
rect 8662 16940 8668 16992
rect 8720 16980 8726 16992
rect 8849 16983 8907 16989
rect 8849 16980 8861 16983
rect 8720 16952 8861 16980
rect 8720 16940 8726 16952
rect 8849 16949 8861 16952
rect 8895 16949 8907 16983
rect 8849 16943 8907 16949
rect 9309 16983 9367 16989
rect 9309 16949 9321 16983
rect 9355 16980 9367 16983
rect 9858 16980 9864 16992
rect 9355 16952 9864 16980
rect 9355 16949 9367 16952
rect 9309 16943 9367 16949
rect 9858 16940 9864 16952
rect 9916 16980 9922 16992
rect 10413 16983 10471 16989
rect 10413 16980 10425 16983
rect 9916 16952 10425 16980
rect 9916 16940 9922 16952
rect 10413 16949 10425 16952
rect 10459 16980 10471 16983
rect 10686 16980 10692 16992
rect 10459 16952 10692 16980
rect 10459 16949 10471 16952
rect 10413 16943 10471 16949
rect 10686 16940 10692 16952
rect 10744 16940 10750 16992
rect 11057 16983 11115 16989
rect 11057 16949 11069 16983
rect 11103 16980 11115 16983
rect 11698 16980 11704 16992
rect 11103 16952 11704 16980
rect 11103 16949 11115 16952
rect 11057 16943 11115 16949
rect 11698 16940 11704 16952
rect 11756 16940 11762 16992
rect 12253 16983 12311 16989
rect 12253 16949 12265 16983
rect 12299 16980 12311 16983
rect 12342 16980 12348 16992
rect 12299 16952 12348 16980
rect 12299 16949 12311 16952
rect 12253 16943 12311 16949
rect 12342 16940 12348 16952
rect 12400 16940 12406 16992
rect 12710 16980 12716 16992
rect 12671 16952 12716 16980
rect 12710 16940 12716 16952
rect 12768 16940 12774 16992
rect 14090 16980 14096 16992
rect 14051 16952 14096 16980
rect 14090 16940 14096 16952
rect 14148 16940 14154 16992
rect 15286 16980 15292 16992
rect 15247 16952 15292 16980
rect 15286 16940 15292 16952
rect 15344 16940 15350 16992
rect 15470 16940 15476 16992
rect 15528 16980 15534 16992
rect 15672 16989 15700 17020
rect 16574 17008 16580 17020
rect 16632 17008 16638 17060
rect 15657 16983 15715 16989
rect 15657 16980 15669 16983
rect 15528 16952 15669 16980
rect 15528 16940 15534 16952
rect 15657 16949 15669 16952
rect 15703 16949 15715 16983
rect 16868 16980 16896 17079
rect 17770 17076 17776 17128
rect 17828 17116 17834 17128
rect 18049 17119 18107 17125
rect 18049 17116 18061 17119
rect 17828 17088 18061 17116
rect 17828 17076 17834 17088
rect 18049 17085 18061 17088
rect 18095 17085 18107 17119
rect 18049 17079 18107 17085
rect 18509 17119 18567 17125
rect 18509 17085 18521 17119
rect 18555 17116 18567 17119
rect 18874 17116 18880 17128
rect 18555 17088 18880 17116
rect 18555 17085 18567 17088
rect 18509 17079 18567 17085
rect 18524 17048 18552 17079
rect 18874 17076 18880 17088
rect 18932 17116 18938 17128
rect 19695 17125 19723 17156
rect 19061 17119 19119 17125
rect 19061 17116 19073 17119
rect 18932 17088 19073 17116
rect 18932 17076 18938 17088
rect 19061 17085 19073 17088
rect 19107 17085 19119 17119
rect 19061 17079 19119 17085
rect 19680 17119 19738 17125
rect 19680 17085 19692 17119
rect 19726 17116 19738 17119
rect 20073 17119 20131 17125
rect 20073 17116 20085 17119
rect 19726 17088 20085 17116
rect 19726 17085 19738 17088
rect 19680 17079 19738 17085
rect 20073 17085 20085 17088
rect 20119 17085 20131 17119
rect 20073 17079 20131 17085
rect 17788 17020 18552 17048
rect 17310 16980 17316 16992
rect 16868 16952 17316 16980
rect 15657 16943 15715 16949
rect 17310 16940 17316 16952
rect 17368 16980 17374 16992
rect 17788 16989 17816 17020
rect 17773 16983 17831 16989
rect 17773 16980 17785 16983
rect 17368 16952 17785 16980
rect 17368 16940 17374 16952
rect 17773 16949 17785 16952
rect 17819 16949 17831 16983
rect 17773 16943 17831 16949
rect 17862 16940 17868 16992
rect 17920 16980 17926 16992
rect 18141 16983 18199 16989
rect 18141 16980 18153 16983
rect 17920 16952 18153 16980
rect 17920 16940 17926 16952
rect 18141 16949 18153 16952
rect 18187 16949 18199 16983
rect 18141 16943 18199 16949
rect 1104 16890 20884 16912
rect 1104 16838 8315 16890
rect 8367 16838 8379 16890
rect 8431 16838 8443 16890
rect 8495 16838 8507 16890
rect 8559 16838 15648 16890
rect 15700 16838 15712 16890
rect 15764 16838 15776 16890
rect 15828 16838 15840 16890
rect 15892 16838 20884 16890
rect 1104 16816 20884 16838
rect 10778 16776 10784 16788
rect 10739 16748 10784 16776
rect 10778 16736 10784 16748
rect 10836 16736 10842 16788
rect 12526 16736 12532 16788
rect 12584 16776 12590 16788
rect 13265 16779 13323 16785
rect 13265 16776 13277 16779
rect 12584 16748 13277 16776
rect 12584 16736 12590 16748
rect 13265 16745 13277 16748
rect 13311 16745 13323 16779
rect 13265 16739 13323 16745
rect 13446 16736 13452 16788
rect 13504 16776 13510 16788
rect 15381 16779 15439 16785
rect 15381 16776 15393 16779
rect 13504 16748 15393 16776
rect 13504 16736 13510 16748
rect 15381 16745 15393 16748
rect 15427 16745 15439 16779
rect 15381 16739 15439 16745
rect 16206 16736 16212 16788
rect 16264 16776 16270 16788
rect 16301 16779 16359 16785
rect 16301 16776 16313 16779
rect 16264 16748 16313 16776
rect 16264 16736 16270 16748
rect 16301 16745 16313 16748
rect 16347 16745 16359 16779
rect 16301 16739 16359 16745
rect 17494 16736 17500 16788
rect 17552 16776 17558 16788
rect 17552 16748 18092 16776
rect 17552 16736 17558 16748
rect 9030 16708 9036 16720
rect 8312 16680 9036 16708
rect 1486 16600 1492 16652
rect 1544 16640 1550 16652
rect 2866 16640 2872 16652
rect 1544 16612 2872 16640
rect 1544 16600 1550 16612
rect 2866 16600 2872 16612
rect 2924 16600 2930 16652
rect 8312 16649 8340 16680
rect 9030 16668 9036 16680
rect 9088 16668 9094 16720
rect 11790 16708 11796 16720
rect 11751 16680 11796 16708
rect 11790 16668 11796 16680
rect 11848 16668 11854 16720
rect 17770 16708 17776 16720
rect 13188 16680 17776 16708
rect 8297 16643 8355 16649
rect 8297 16609 8309 16643
rect 8343 16609 8355 16643
rect 8478 16640 8484 16652
rect 8439 16612 8484 16640
rect 8297 16603 8355 16609
rect 8478 16600 8484 16612
rect 8536 16600 8542 16652
rect 9674 16640 9680 16652
rect 9635 16612 9680 16640
rect 9674 16600 9680 16612
rect 9732 16600 9738 16652
rect 9858 16600 9864 16652
rect 9916 16640 9922 16652
rect 10137 16643 10195 16649
rect 10137 16640 10149 16643
rect 9916 16612 10149 16640
rect 9916 16600 9922 16612
rect 10137 16609 10149 16612
rect 10183 16609 10195 16643
rect 10137 16603 10195 16609
rect 12618 16600 12624 16652
rect 12676 16640 12682 16652
rect 13188 16649 13216 16680
rect 17770 16668 17776 16680
rect 17828 16668 17834 16720
rect 17954 16708 17960 16720
rect 17915 16680 17960 16708
rect 17954 16668 17960 16680
rect 18012 16668 18018 16720
rect 18064 16717 18092 16748
rect 18690 16736 18696 16788
rect 18748 16776 18754 16788
rect 18877 16779 18935 16785
rect 18877 16776 18889 16779
rect 18748 16748 18889 16776
rect 18748 16736 18754 16748
rect 18877 16745 18889 16748
rect 18923 16745 18935 16779
rect 18877 16739 18935 16745
rect 19613 16779 19671 16785
rect 19613 16745 19625 16779
rect 19659 16776 19671 16779
rect 21542 16776 21548 16788
rect 19659 16748 21548 16776
rect 19659 16745 19671 16748
rect 19613 16739 19671 16745
rect 21542 16736 21548 16748
rect 21600 16736 21606 16788
rect 18049 16711 18107 16717
rect 18049 16677 18061 16711
rect 18095 16677 18107 16711
rect 18049 16671 18107 16677
rect 13173 16643 13231 16649
rect 13173 16640 13185 16643
rect 12676 16612 13185 16640
rect 12676 16600 12682 16612
rect 13173 16609 13185 16612
rect 13219 16609 13231 16643
rect 13173 16603 13231 16609
rect 13538 16600 13544 16652
rect 13596 16640 13602 16652
rect 13633 16643 13691 16649
rect 13633 16640 13645 16643
rect 13596 16612 13645 16640
rect 13596 16600 13602 16612
rect 13633 16609 13645 16612
rect 13679 16640 13691 16643
rect 15562 16640 15568 16652
rect 13679 16612 13814 16640
rect 15523 16612 15568 16640
rect 13679 16609 13691 16612
rect 13633 16603 13691 16609
rect 8754 16572 8760 16584
rect 8715 16544 8760 16572
rect 8754 16532 8760 16544
rect 8812 16532 8818 16584
rect 10413 16575 10471 16581
rect 10413 16541 10425 16575
rect 10459 16572 10471 16575
rect 10502 16572 10508 16584
rect 10459 16544 10508 16572
rect 10459 16541 10471 16544
rect 10413 16535 10471 16541
rect 10502 16532 10508 16544
rect 10560 16532 10566 16584
rect 11698 16572 11704 16584
rect 11659 16544 11704 16572
rect 11698 16532 11704 16544
rect 11756 16532 11762 16584
rect 11882 16532 11888 16584
rect 11940 16572 11946 16584
rect 11977 16575 12035 16581
rect 11977 16572 11989 16575
rect 11940 16544 11989 16572
rect 11940 16532 11946 16544
rect 11977 16541 11989 16544
rect 12023 16541 12035 16575
rect 13786 16572 13814 16612
rect 15562 16600 15568 16612
rect 15620 16600 15626 16652
rect 15746 16640 15752 16652
rect 15707 16612 15752 16640
rect 15746 16600 15752 16612
rect 15804 16600 15810 16652
rect 19429 16643 19487 16649
rect 19429 16609 19441 16643
rect 19475 16640 19487 16643
rect 19610 16640 19616 16652
rect 19475 16612 19616 16640
rect 19475 16609 19487 16612
rect 19429 16603 19487 16609
rect 19610 16600 19616 16612
rect 19668 16600 19674 16652
rect 15764 16572 15792 16600
rect 13786 16544 15792 16572
rect 16853 16575 16911 16581
rect 11977 16535 12035 16541
rect 16853 16541 16865 16575
rect 16899 16572 16911 16575
rect 17770 16572 17776 16584
rect 16899 16544 17776 16572
rect 16899 16541 16911 16544
rect 16853 16535 16911 16541
rect 17770 16532 17776 16544
rect 17828 16532 17834 16584
rect 18598 16572 18604 16584
rect 18559 16544 18604 16572
rect 18598 16532 18604 16544
rect 18656 16532 18662 16584
rect 15562 16464 15568 16516
rect 15620 16504 15626 16516
rect 18690 16504 18696 16516
rect 15620 16476 18696 16504
rect 15620 16464 15626 16476
rect 18690 16464 18696 16476
rect 18748 16464 18754 16516
rect 7929 16439 7987 16445
rect 7929 16405 7941 16439
rect 7975 16436 7987 16439
rect 8110 16436 8116 16448
rect 7975 16408 8116 16436
rect 7975 16405 7987 16408
rect 7929 16399 7987 16405
rect 8110 16396 8116 16408
rect 8168 16396 8174 16448
rect 9490 16436 9496 16448
rect 9451 16408 9496 16436
rect 9490 16396 9496 16408
rect 9548 16436 9554 16448
rect 12621 16439 12679 16445
rect 12621 16436 12633 16439
rect 9548 16408 12633 16436
rect 9548 16396 9554 16408
rect 12621 16405 12633 16408
rect 12667 16436 12679 16439
rect 12802 16436 12808 16448
rect 12667 16408 12808 16436
rect 12667 16405 12679 16408
rect 12621 16399 12679 16405
rect 12802 16396 12808 16408
rect 12860 16396 12866 16448
rect 14369 16439 14427 16445
rect 14369 16405 14381 16439
rect 14415 16436 14427 16439
rect 14458 16436 14464 16448
rect 14415 16408 14464 16436
rect 14415 16405 14427 16408
rect 14369 16399 14427 16405
rect 14458 16396 14464 16408
rect 14516 16396 14522 16448
rect 14642 16436 14648 16448
rect 14603 16408 14648 16436
rect 14642 16396 14648 16408
rect 14700 16396 14706 16448
rect 14918 16396 14924 16448
rect 14976 16436 14982 16448
rect 15013 16439 15071 16445
rect 15013 16436 15025 16439
rect 14976 16408 15025 16436
rect 14976 16396 14982 16408
rect 15013 16405 15025 16408
rect 15059 16405 15071 16439
rect 15013 16399 15071 16405
rect 1104 16346 20884 16368
rect 1104 16294 4648 16346
rect 4700 16294 4712 16346
rect 4764 16294 4776 16346
rect 4828 16294 4840 16346
rect 4892 16294 11982 16346
rect 12034 16294 12046 16346
rect 12098 16294 12110 16346
rect 12162 16294 12174 16346
rect 12226 16294 19315 16346
rect 19367 16294 19379 16346
rect 19431 16294 19443 16346
rect 19495 16294 19507 16346
rect 19559 16294 20884 16346
rect 1104 16272 20884 16294
rect 1578 16232 1584 16244
rect 1539 16204 1584 16232
rect 1578 16192 1584 16204
rect 1636 16192 1642 16244
rect 11698 16192 11704 16244
rect 11756 16232 11762 16244
rect 11885 16235 11943 16241
rect 11885 16232 11897 16235
rect 11756 16204 11897 16232
rect 11756 16192 11762 16204
rect 11885 16201 11897 16204
rect 11931 16201 11943 16235
rect 11885 16195 11943 16201
rect 14093 16235 14151 16241
rect 14093 16201 14105 16235
rect 14139 16232 14151 16235
rect 14642 16232 14648 16244
rect 14139 16204 14648 16232
rect 14139 16201 14151 16204
rect 14093 16195 14151 16201
rect 14642 16192 14648 16204
rect 14700 16192 14706 16244
rect 14826 16232 14832 16244
rect 14739 16204 14832 16232
rect 14826 16192 14832 16204
rect 14884 16232 14890 16244
rect 15562 16232 15568 16244
rect 14884 16204 15568 16232
rect 14884 16192 14890 16204
rect 15562 16192 15568 16204
rect 15620 16192 15626 16244
rect 17494 16232 17500 16244
rect 17455 16204 17500 16232
rect 17494 16192 17500 16204
rect 17552 16192 17558 16244
rect 17770 16232 17776 16244
rect 17731 16204 17776 16232
rect 17770 16192 17776 16204
rect 17828 16192 17834 16244
rect 9674 16124 9680 16176
rect 9732 16164 9738 16176
rect 11517 16167 11575 16173
rect 9732 16136 11002 16164
rect 9732 16124 9738 16136
rect 1302 16056 1308 16108
rect 1360 16096 1366 16108
rect 10597 16099 10655 16105
rect 1360 16068 6913 16096
rect 1360 16056 1366 16068
rect 1397 16031 1455 16037
rect 1397 15997 1409 16031
rect 1443 16028 1455 16031
rect 6885 16028 6913 16068
rect 10597 16065 10609 16099
rect 10643 16096 10655 16099
rect 10778 16096 10784 16108
rect 10643 16068 10784 16096
rect 10643 16065 10655 16068
rect 10597 16059 10655 16065
rect 10778 16056 10784 16068
rect 10836 16056 10842 16108
rect 10974 16096 11002 16136
rect 11517 16133 11529 16167
rect 11563 16164 11575 16167
rect 11790 16164 11796 16176
rect 11563 16136 11796 16164
rect 11563 16133 11575 16136
rect 11517 16127 11575 16133
rect 11790 16124 11796 16136
rect 11848 16164 11854 16176
rect 12161 16167 12219 16173
rect 12161 16164 12173 16167
rect 11848 16136 12173 16164
rect 11848 16124 11854 16136
rect 12161 16133 12173 16136
rect 12207 16133 12219 16167
rect 12161 16127 12219 16133
rect 12618 16096 12624 16108
rect 10974 16068 12624 16096
rect 12618 16056 12624 16068
rect 12676 16056 12682 16108
rect 13173 16099 13231 16105
rect 13173 16065 13185 16099
rect 13219 16096 13231 16099
rect 13262 16096 13268 16108
rect 13219 16068 13268 16096
rect 13219 16065 13231 16068
rect 13173 16059 13231 16065
rect 13262 16056 13268 16068
rect 13320 16096 13326 16108
rect 14369 16099 14427 16105
rect 14369 16096 14381 16099
rect 13320 16068 14381 16096
rect 13320 16056 13326 16068
rect 14369 16065 14381 16068
rect 14415 16065 14427 16099
rect 14369 16059 14427 16065
rect 14458 16056 14464 16108
rect 14516 16096 14522 16108
rect 14921 16099 14979 16105
rect 14921 16096 14933 16099
rect 14516 16068 14933 16096
rect 14516 16056 14522 16068
rect 14921 16065 14933 16068
rect 14967 16065 14979 16099
rect 14921 16059 14979 16065
rect 15473 16099 15531 16105
rect 15473 16065 15485 16099
rect 15519 16096 15531 16099
rect 15746 16096 15752 16108
rect 15519 16068 15752 16096
rect 15519 16065 15531 16068
rect 15473 16059 15531 16065
rect 15746 16056 15752 16068
rect 15804 16096 15810 16108
rect 17310 16096 17316 16108
rect 15804 16068 17316 16096
rect 15804 16056 15810 16068
rect 17310 16056 17316 16068
rect 17368 16056 17374 16108
rect 17788 16096 17816 16192
rect 18693 16167 18751 16173
rect 18693 16133 18705 16167
rect 18739 16164 18751 16167
rect 19058 16164 19064 16176
rect 18739 16136 19064 16164
rect 18739 16133 18751 16136
rect 18693 16127 18751 16133
rect 19058 16124 19064 16136
rect 19116 16164 19122 16176
rect 19978 16164 19984 16176
rect 19116 16136 19984 16164
rect 19116 16124 19122 16136
rect 19978 16124 19984 16136
rect 20036 16124 20042 16176
rect 18141 16099 18199 16105
rect 18141 16096 18153 16099
rect 17788 16068 18153 16096
rect 18141 16065 18153 16068
rect 18187 16065 18199 16099
rect 18141 16059 18199 16065
rect 18322 16056 18328 16108
rect 18380 16096 18386 16108
rect 19751 16099 19809 16105
rect 19751 16096 19763 16099
rect 18380 16068 19763 16096
rect 18380 16056 18386 16068
rect 19751 16065 19763 16068
rect 19797 16065 19809 16099
rect 19751 16059 19809 16065
rect 6952 16031 7010 16037
rect 6952 16028 6964 16031
rect 1443 16000 2084 16028
rect 6885 16000 6964 16028
rect 1443 15997 1455 16000
rect 1397 15991 1455 15997
rect 2056 15901 2084 16000
rect 6952 15997 6964 16000
rect 6998 16028 7010 16031
rect 7374 16028 7380 16040
rect 6998 16000 7380 16028
rect 6998 15997 7010 16000
rect 6952 15991 7010 15997
rect 7374 15988 7380 16000
rect 7432 15988 7438 16040
rect 9582 16028 9588 16040
rect 9640 16037 9646 16040
rect 9640 16031 9678 16037
rect 9530 16000 9588 16028
rect 9582 15988 9588 16000
rect 9666 16028 9678 16031
rect 10045 16031 10103 16037
rect 10045 16028 10057 16031
rect 9666 16000 10057 16028
rect 9666 15997 9678 16000
rect 9640 15991 9678 15997
rect 10045 15997 10057 16000
rect 10091 15997 10103 16031
rect 12636 16028 12664 16056
rect 13906 16028 13912 16040
rect 12636 16000 13912 16028
rect 10045 15991 10103 15997
rect 9640 15988 9646 15991
rect 13906 15988 13912 16000
rect 13964 15988 13970 16040
rect 16206 16028 16212 16040
rect 16167 16000 16212 16028
rect 16206 15988 16212 16000
rect 16264 15988 16270 16040
rect 16393 16031 16451 16037
rect 16393 15997 16405 16031
rect 16439 15997 16451 16031
rect 16393 15991 16451 15997
rect 17129 16031 17187 16037
rect 17129 15997 17141 16031
rect 17175 16028 17187 16031
rect 17954 16028 17960 16040
rect 17175 16000 17960 16028
rect 17175 15997 17187 16000
rect 17129 15991 17187 15997
rect 7055 15963 7113 15969
rect 7055 15929 7067 15963
rect 7101 15960 7113 15963
rect 7466 15960 7472 15972
rect 7101 15932 7472 15960
rect 7101 15929 7113 15932
rect 7055 15923 7113 15929
rect 7466 15920 7472 15932
rect 7524 15920 7530 15972
rect 8018 15960 8024 15972
rect 7979 15932 8024 15960
rect 8018 15920 8024 15932
rect 8076 15920 8082 15972
rect 8110 15920 8116 15972
rect 8168 15960 8174 15972
rect 8168 15932 8213 15960
rect 8168 15920 8174 15932
rect 8478 15920 8484 15972
rect 8536 15920 8542 15972
rect 8662 15960 8668 15972
rect 8623 15932 8668 15960
rect 8662 15920 8668 15932
rect 8720 15920 8726 15972
rect 9493 15963 9551 15969
rect 9493 15960 9505 15963
rect 8864 15932 9505 15960
rect 2041 15895 2099 15901
rect 2041 15861 2053 15895
rect 2087 15892 2099 15895
rect 2958 15892 2964 15904
rect 2087 15864 2964 15892
rect 2087 15861 2099 15864
rect 2041 15855 2099 15861
rect 2958 15852 2964 15864
rect 3016 15852 3022 15904
rect 7742 15892 7748 15904
rect 7703 15864 7748 15892
rect 7742 15852 7748 15864
rect 7800 15892 7806 15904
rect 8496 15892 8524 15920
rect 8864 15892 8892 15932
rect 9493 15929 9505 15932
rect 9539 15960 9551 15963
rect 9858 15960 9864 15972
rect 9539 15932 9864 15960
rect 9539 15929 9551 15932
rect 9493 15923 9551 15929
rect 9858 15920 9864 15932
rect 9916 15920 9922 15972
rect 10226 15920 10232 15972
rect 10284 15960 10290 15972
rect 10505 15963 10563 15969
rect 10505 15960 10517 15963
rect 10284 15932 10517 15960
rect 10284 15920 10290 15932
rect 10505 15929 10517 15932
rect 10551 15960 10563 15963
rect 10959 15963 11017 15969
rect 10959 15960 10971 15963
rect 10551 15932 10971 15960
rect 10551 15929 10563 15932
rect 10505 15923 10563 15929
rect 10959 15929 10971 15932
rect 11005 15960 11017 15963
rect 13535 15963 13593 15969
rect 11005 15932 13124 15960
rect 11005 15929 11017 15932
rect 10959 15923 11017 15929
rect 9030 15892 9036 15904
rect 7800 15864 8892 15892
rect 8991 15864 9036 15892
rect 7800 15852 7806 15864
rect 9030 15852 9036 15864
rect 9088 15852 9094 15904
rect 9723 15895 9781 15901
rect 9723 15861 9735 15895
rect 9769 15892 9781 15895
rect 9950 15892 9956 15904
rect 9769 15864 9956 15892
rect 9769 15861 9781 15864
rect 9723 15855 9781 15861
rect 9950 15852 9956 15864
rect 10008 15852 10014 15904
rect 13096 15901 13124 15932
rect 13535 15929 13547 15963
rect 13581 15929 13593 15963
rect 16408 15960 16436 15991
rect 17954 15988 17960 16000
rect 18012 15988 18018 16040
rect 18874 15988 18880 16040
rect 18932 16028 18938 16040
rect 19648 16031 19706 16037
rect 19648 16028 19660 16031
rect 18932 16000 19660 16028
rect 18932 15988 18938 16000
rect 19648 15997 19660 16000
rect 19694 16028 19706 16031
rect 20073 16031 20131 16037
rect 20073 16028 20085 16031
rect 19694 16000 20085 16028
rect 19694 15997 19706 16000
rect 19648 15991 19706 15997
rect 20073 15997 20085 16000
rect 20119 15997 20131 16031
rect 20073 15991 20131 15997
rect 16666 15960 16672 15972
rect 13535 15923 13593 15929
rect 15764 15932 16436 15960
rect 16627 15932 16672 15960
rect 13081 15895 13139 15901
rect 13081 15861 13093 15895
rect 13127 15892 13139 15895
rect 13550 15892 13578 15923
rect 13814 15892 13820 15904
rect 13127 15864 13820 15892
rect 13127 15861 13139 15864
rect 13081 15855 13139 15861
rect 13814 15852 13820 15864
rect 13872 15852 13878 15904
rect 15010 15852 15016 15904
rect 15068 15892 15074 15904
rect 15286 15892 15292 15904
rect 15068 15864 15292 15892
rect 15068 15852 15074 15864
rect 15286 15852 15292 15864
rect 15344 15892 15350 15904
rect 15764 15901 15792 15932
rect 16666 15920 16672 15932
rect 16724 15920 16730 15972
rect 18230 15920 18236 15972
rect 18288 15960 18294 15972
rect 18288 15932 18333 15960
rect 18288 15920 18294 15932
rect 15749 15895 15807 15901
rect 15749 15892 15761 15895
rect 15344 15864 15761 15892
rect 15344 15852 15350 15864
rect 15749 15861 15761 15864
rect 15795 15861 15807 15895
rect 15749 15855 15807 15861
rect 17402 15852 17408 15904
rect 17460 15892 17466 15904
rect 19429 15895 19487 15901
rect 19429 15892 19441 15895
rect 17460 15864 19441 15892
rect 17460 15852 17466 15864
rect 19429 15861 19441 15864
rect 19475 15892 19487 15895
rect 19610 15892 19616 15904
rect 19475 15864 19616 15892
rect 19475 15861 19487 15864
rect 19429 15855 19487 15861
rect 19610 15852 19616 15864
rect 19668 15852 19674 15904
rect 1104 15802 20884 15824
rect 1104 15750 8315 15802
rect 8367 15750 8379 15802
rect 8431 15750 8443 15802
rect 8495 15750 8507 15802
rect 8559 15750 15648 15802
rect 15700 15750 15712 15802
rect 15764 15750 15776 15802
rect 15828 15750 15840 15802
rect 15892 15750 20884 15802
rect 1104 15728 20884 15750
rect 6273 15691 6331 15697
rect 6273 15657 6285 15691
rect 6319 15688 6331 15691
rect 8018 15688 8024 15700
rect 6319 15660 8024 15688
rect 6319 15657 6331 15660
rect 6273 15651 6331 15657
rect 8018 15648 8024 15660
rect 8076 15648 8082 15700
rect 8110 15648 8116 15700
rect 8168 15688 8174 15700
rect 8205 15691 8263 15697
rect 8205 15688 8217 15691
rect 8168 15660 8217 15688
rect 8168 15648 8174 15660
rect 8205 15657 8217 15660
rect 8251 15657 8263 15691
rect 8205 15651 8263 15657
rect 10689 15691 10747 15697
rect 10689 15657 10701 15691
rect 10735 15688 10747 15691
rect 10735 15660 11744 15688
rect 10735 15657 10747 15660
rect 10689 15651 10747 15657
rect 7647 15623 7705 15629
rect 7647 15589 7659 15623
rect 7693 15620 7705 15623
rect 7926 15620 7932 15632
rect 7693 15592 7932 15620
rect 7693 15589 7705 15592
rect 7647 15583 7705 15589
rect 7926 15580 7932 15592
rect 7984 15580 7990 15632
rect 8036 15620 8064 15648
rect 11716 15632 11744 15660
rect 13814 15648 13820 15700
rect 13872 15688 13878 15700
rect 16025 15691 16083 15697
rect 13872 15660 13917 15688
rect 13872 15648 13878 15660
rect 16025 15657 16037 15691
rect 16071 15688 16083 15691
rect 16206 15688 16212 15700
rect 16071 15660 16212 15688
rect 16071 15657 16083 15660
rect 16025 15651 16083 15657
rect 16206 15648 16212 15660
rect 16264 15648 16270 15700
rect 17681 15691 17739 15697
rect 17681 15657 17693 15691
rect 17727 15688 17739 15691
rect 18141 15691 18199 15697
rect 18141 15688 18153 15691
rect 17727 15660 18153 15688
rect 17727 15657 17739 15660
rect 17681 15651 17739 15657
rect 18141 15657 18153 15660
rect 18187 15688 18199 15691
rect 18230 15688 18236 15700
rect 18187 15660 18236 15688
rect 18187 15657 18199 15660
rect 18141 15651 18199 15657
rect 18230 15648 18236 15660
rect 18288 15648 18294 15700
rect 18782 15648 18788 15700
rect 18840 15688 18846 15700
rect 18877 15691 18935 15697
rect 18877 15688 18889 15691
rect 18840 15660 18889 15688
rect 18840 15648 18846 15660
rect 18877 15657 18889 15660
rect 18923 15657 18935 15691
rect 18877 15651 18935 15657
rect 8481 15623 8539 15629
rect 8481 15620 8493 15623
rect 8036 15592 8493 15620
rect 8481 15589 8493 15592
rect 8527 15589 8539 15623
rect 8481 15583 8539 15589
rect 10131 15623 10189 15629
rect 10131 15589 10143 15623
rect 10177 15620 10189 15623
rect 10226 15620 10232 15632
rect 10177 15592 10232 15620
rect 10177 15589 10189 15592
rect 10131 15583 10189 15589
rect 10226 15580 10232 15592
rect 10284 15580 10290 15632
rect 11698 15620 11704 15632
rect 11611 15592 11704 15620
rect 11698 15580 11704 15592
rect 11756 15580 11762 15632
rect 17123 15623 17181 15629
rect 17123 15589 17135 15623
rect 17169 15620 17181 15623
rect 18800 15620 18828 15648
rect 17169 15592 18828 15620
rect 17169 15589 17181 15592
rect 17123 15583 17181 15589
rect 8754 15512 8760 15564
rect 8812 15552 8818 15564
rect 9769 15555 9827 15561
rect 9769 15552 9781 15555
rect 8812 15524 9781 15552
rect 8812 15512 8818 15524
rect 9769 15521 9781 15524
rect 9815 15552 9827 15555
rect 9858 15552 9864 15564
rect 9815 15524 9864 15552
rect 9815 15521 9827 15524
rect 9769 15515 9827 15521
rect 9858 15512 9864 15524
rect 9916 15512 9922 15564
rect 13354 15512 13360 15564
rect 13412 15552 13418 15564
rect 13449 15555 13507 15561
rect 13449 15552 13461 15555
rect 13412 15524 13461 15552
rect 13412 15512 13418 15524
rect 13449 15521 13461 15524
rect 13495 15521 13507 15555
rect 13449 15515 13507 15521
rect 14734 15512 14740 15564
rect 14792 15552 14798 15564
rect 15324 15555 15382 15561
rect 15324 15552 15336 15555
rect 14792 15524 15336 15552
rect 14792 15512 14798 15524
rect 15324 15521 15336 15524
rect 15370 15521 15382 15555
rect 15324 15515 15382 15521
rect 16574 15512 16580 15564
rect 16632 15552 16638 15564
rect 16761 15555 16819 15561
rect 16761 15552 16773 15555
rect 16632 15524 16773 15552
rect 16632 15512 16638 15524
rect 16761 15521 16773 15524
rect 16807 15521 16819 15555
rect 18506 15552 18512 15564
rect 18467 15524 18512 15552
rect 16761 15515 16819 15521
rect 18506 15512 18512 15524
rect 18564 15512 18570 15564
rect 7285 15487 7343 15493
rect 7285 15453 7297 15487
rect 7331 15484 7343 15487
rect 7558 15484 7564 15496
rect 7331 15456 7564 15484
rect 7331 15453 7343 15456
rect 7285 15447 7343 15453
rect 7558 15444 7564 15456
rect 7616 15444 7622 15496
rect 11606 15484 11612 15496
rect 11567 15456 11612 15484
rect 11606 15444 11612 15456
rect 11664 15444 11670 15496
rect 11882 15484 11888 15496
rect 11843 15456 11888 15484
rect 11882 15444 11888 15456
rect 11940 15444 11946 15496
rect 5350 15376 5356 15428
rect 5408 15416 5414 15428
rect 9401 15419 9459 15425
rect 9401 15416 9413 15419
rect 5408 15388 9413 15416
rect 5408 15376 5414 15388
rect 9401 15385 9413 15388
rect 9447 15416 9459 15419
rect 9674 15416 9680 15428
rect 9447 15388 9680 15416
rect 9447 15385 9459 15388
rect 9401 15379 9459 15385
rect 9674 15376 9680 15388
rect 9732 15376 9738 15428
rect 6914 15348 6920 15360
rect 6875 15320 6920 15348
rect 6914 15308 6920 15320
rect 6972 15308 6978 15360
rect 8938 15348 8944 15360
rect 8899 15320 8944 15348
rect 8938 15308 8944 15320
rect 8996 15308 9002 15360
rect 11330 15308 11336 15360
rect 11388 15348 11394 15360
rect 12342 15348 12348 15360
rect 11388 15320 12348 15348
rect 11388 15308 11394 15320
rect 12342 15308 12348 15320
rect 12400 15348 12406 15360
rect 13173 15351 13231 15357
rect 13173 15348 13185 15351
rect 12400 15320 13185 15348
rect 12400 15308 12406 15320
rect 13173 15317 13185 15320
rect 13219 15317 13231 15351
rect 14366 15348 14372 15360
rect 14327 15320 14372 15348
rect 13173 15311 13231 15317
rect 14366 15308 14372 15320
rect 14424 15308 14430 15360
rect 14550 15308 14556 15360
rect 14608 15348 14614 15360
rect 15427 15351 15485 15357
rect 15427 15348 15439 15351
rect 14608 15320 15439 15348
rect 14608 15308 14614 15320
rect 15427 15317 15439 15320
rect 15473 15317 15485 15351
rect 15427 15311 15485 15317
rect 18690 15308 18696 15360
rect 18748 15348 18754 15360
rect 19429 15351 19487 15357
rect 19429 15348 19441 15351
rect 18748 15320 19441 15348
rect 18748 15308 18754 15320
rect 19429 15317 19441 15320
rect 19475 15317 19487 15351
rect 19429 15311 19487 15317
rect 1104 15258 20884 15280
rect 1104 15206 4648 15258
rect 4700 15206 4712 15258
rect 4764 15206 4776 15258
rect 4828 15206 4840 15258
rect 4892 15206 11982 15258
rect 12034 15206 12046 15258
rect 12098 15206 12110 15258
rect 12162 15206 12174 15258
rect 12226 15206 19315 15258
rect 19367 15206 19379 15258
rect 19431 15206 19443 15258
rect 19495 15206 19507 15258
rect 19559 15206 20884 15258
rect 1104 15184 20884 15206
rect 6270 15144 6276 15156
rect 6231 15116 6276 15144
rect 6270 15104 6276 15116
rect 6328 15104 6334 15156
rect 7926 15144 7932 15156
rect 7839 15116 7932 15144
rect 7926 15104 7932 15116
rect 7984 15144 7990 15156
rect 9861 15147 9919 15153
rect 9861 15144 9873 15147
rect 7984 15116 9873 15144
rect 7984 15104 7990 15116
rect 9861 15113 9873 15116
rect 9907 15144 9919 15147
rect 10226 15144 10232 15156
rect 9907 15116 10232 15144
rect 9907 15113 9919 15116
rect 9861 15107 9919 15113
rect 10226 15104 10232 15116
rect 10284 15104 10290 15156
rect 11698 15144 11704 15156
rect 11659 15116 11704 15144
rect 11698 15104 11704 15116
rect 11756 15104 11762 15156
rect 13357 15147 13415 15153
rect 13357 15113 13369 15147
rect 13403 15144 13415 15147
rect 13814 15144 13820 15156
rect 13403 15116 13820 15144
rect 13403 15113 13415 15116
rect 13357 15107 13415 15113
rect 13786 15104 13820 15116
rect 13872 15104 13878 15156
rect 16393 15147 16451 15153
rect 16393 15113 16405 15147
rect 16439 15144 16451 15147
rect 16574 15144 16580 15156
rect 16439 15116 16580 15144
rect 16439 15113 16451 15116
rect 16393 15107 16451 15113
rect 16574 15104 16580 15116
rect 16632 15104 16638 15156
rect 17034 15144 17040 15156
rect 16995 15116 17040 15144
rect 17034 15104 17040 15116
rect 17092 15104 17098 15156
rect 18506 15104 18512 15156
rect 18564 15144 18570 15156
rect 19429 15147 19487 15153
rect 19429 15144 19441 15147
rect 18564 15116 19441 15144
rect 18564 15104 18570 15116
rect 19429 15113 19441 15116
rect 19475 15113 19487 15147
rect 19429 15107 19487 15113
rect 13786 15076 13814 15104
rect 14737 15079 14795 15085
rect 14737 15076 14749 15079
rect 13786 15048 14749 15076
rect 7558 15008 7564 15020
rect 7471 14980 7564 15008
rect 7558 14968 7564 14980
rect 7616 15008 7622 15020
rect 8205 15011 8263 15017
rect 8205 15008 8217 15011
rect 7616 14980 8217 15008
rect 7616 14968 7622 14980
rect 8205 14977 8217 14980
rect 8251 14977 8263 15011
rect 8205 14971 8263 14977
rect 8573 15011 8631 15017
rect 8573 14977 8585 15011
rect 8619 15008 8631 15011
rect 9306 15008 9312 15020
rect 8619 14980 9312 15008
rect 8619 14977 8631 14980
rect 8573 14971 8631 14977
rect 9306 14968 9312 14980
rect 9364 14968 9370 15020
rect 10045 15011 10103 15017
rect 10045 14977 10057 15011
rect 10091 15008 10103 15011
rect 10134 15008 10140 15020
rect 10091 14980 10140 15008
rect 10091 14977 10103 14980
rect 10045 14971 10103 14977
rect 10134 14968 10140 14980
rect 10192 15008 10198 15020
rect 11241 15011 11299 15017
rect 11241 15008 11253 15011
rect 10192 14980 11253 15008
rect 10192 14968 10198 14980
rect 11241 14977 11253 14980
rect 11287 14977 11299 15011
rect 13446 15008 13452 15020
rect 13407 14980 13452 15008
rect 11241 14971 11299 14977
rect 13446 14968 13452 14980
rect 13504 14968 13510 15020
rect 2222 14900 2228 14952
rect 2280 14940 2286 14952
rect 5788 14943 5846 14949
rect 5788 14940 5800 14943
rect 2280 14912 5800 14940
rect 2280 14900 2286 14912
rect 5788 14909 5800 14912
rect 5834 14940 5846 14943
rect 6270 14940 6276 14952
rect 5834 14912 6276 14940
rect 5834 14909 5846 14912
rect 5788 14903 5846 14909
rect 6270 14900 6276 14912
rect 6328 14900 6334 14952
rect 6641 14943 6699 14949
rect 6641 14909 6653 14943
rect 6687 14940 6699 14943
rect 6733 14943 6791 14949
rect 6733 14940 6745 14943
rect 6687 14912 6745 14940
rect 6687 14909 6699 14912
rect 6641 14903 6699 14909
rect 6733 14909 6745 14912
rect 6779 14940 6791 14943
rect 6822 14940 6828 14952
rect 6779 14912 6828 14940
rect 6779 14909 6791 14912
rect 6733 14903 6791 14909
rect 6822 14900 6828 14912
rect 6880 14900 6886 14952
rect 6914 14900 6920 14952
rect 6972 14940 6978 14952
rect 7285 14943 7343 14949
rect 7285 14940 7297 14943
rect 6972 14912 7297 14940
rect 6972 14900 6978 14912
rect 7285 14909 7297 14912
rect 7331 14909 7343 14943
rect 7285 14903 7343 14909
rect 12345 14943 12403 14949
rect 12345 14909 12357 14943
rect 12391 14909 12403 14943
rect 12894 14940 12900 14952
rect 12855 14912 12900 14940
rect 12345 14903 12403 14909
rect 8665 14875 8723 14881
rect 8665 14841 8677 14875
rect 8711 14841 8723 14875
rect 9214 14872 9220 14884
rect 9175 14844 9220 14872
rect 8665 14835 8723 14841
rect 5859 14807 5917 14813
rect 5859 14773 5871 14807
rect 5905 14804 5917 14807
rect 6086 14804 6092 14816
rect 5905 14776 6092 14804
rect 5905 14773 5917 14776
rect 5859 14767 5917 14773
rect 6086 14764 6092 14776
rect 6144 14764 6150 14816
rect 8680 14804 8708 14835
rect 9214 14832 9220 14844
rect 9272 14832 9278 14884
rect 9324 14844 10088 14872
rect 8938 14804 8944 14816
rect 8680 14776 8944 14804
rect 8938 14764 8944 14776
rect 8996 14804 9002 14816
rect 9324 14804 9352 14844
rect 8996 14776 9352 14804
rect 10060 14804 10088 14844
rect 10226 14832 10232 14884
rect 10284 14872 10290 14884
rect 10366 14875 10424 14881
rect 10366 14872 10378 14875
rect 10284 14844 10378 14872
rect 10284 14832 10290 14844
rect 10366 14841 10378 14844
rect 10412 14841 10424 14875
rect 10366 14835 10424 14841
rect 11146 14832 11152 14884
rect 11204 14872 11210 14884
rect 11606 14872 11612 14884
rect 11204 14844 11612 14872
rect 11204 14832 11210 14844
rect 11606 14832 11612 14844
rect 11664 14872 11670 14884
rect 11977 14875 12035 14881
rect 11977 14872 11989 14875
rect 11664 14844 11989 14872
rect 11664 14832 11670 14844
rect 11977 14841 11989 14844
rect 12023 14841 12035 14875
rect 12360 14872 12388 14903
rect 12894 14900 12900 14912
rect 12952 14900 12958 14952
rect 12912 14872 12940 14900
rect 13826 14881 13854 15048
rect 14737 15045 14749 15048
rect 14783 15076 14795 15079
rect 16761 15079 16819 15085
rect 16761 15076 16773 15079
rect 14783 15048 16773 15076
rect 14783 15045 14795 15048
rect 14737 15039 14795 15045
rect 16761 15045 16773 15048
rect 16807 15076 16819 15079
rect 17218 15076 17224 15088
rect 16807 15048 17224 15076
rect 16807 15045 16819 15048
rect 16761 15039 16819 15045
rect 17218 15036 17224 15048
rect 17276 15076 17282 15088
rect 18325 15079 18383 15085
rect 18325 15076 18337 15079
rect 17276 15048 18337 15076
rect 17276 15036 17282 15048
rect 18325 15045 18337 15048
rect 18371 15076 18383 15079
rect 18782 15076 18788 15088
rect 18371 15048 18788 15076
rect 18371 15045 18383 15048
rect 18325 15039 18383 15045
rect 18782 15036 18788 15048
rect 18840 15036 18846 15088
rect 19058 15076 19064 15088
rect 19019 15048 19064 15076
rect 19058 15036 19064 15048
rect 19116 15076 19122 15088
rect 19242 15076 19248 15088
rect 19116 15048 19248 15076
rect 19116 15036 19122 15048
rect 19242 15036 19248 15048
rect 19300 15036 19306 15088
rect 15102 14968 15108 15020
rect 15160 15008 15166 15020
rect 15565 15011 15623 15017
rect 15565 15008 15577 15011
rect 15160 14980 15577 15008
rect 15160 14968 15166 14980
rect 15565 14977 15577 14980
rect 15611 14977 15623 15011
rect 15565 14971 15623 14977
rect 15930 14968 15936 15020
rect 15988 15008 15994 15020
rect 17034 15008 17040 15020
rect 15988 14980 17040 15008
rect 15988 14968 15994 14980
rect 17034 14968 17040 14980
rect 17092 14968 17098 15020
rect 18509 15011 18567 15017
rect 18509 14977 18521 15011
rect 18555 15008 18567 15011
rect 18966 15008 18972 15020
rect 18555 14980 18972 15008
rect 18555 14977 18567 14980
rect 18509 14971 18567 14977
rect 18966 14968 18972 14980
rect 19024 15008 19030 15020
rect 19797 15011 19855 15017
rect 19797 15008 19809 15011
rect 19024 14980 19809 15008
rect 19024 14968 19030 14980
rect 19797 14977 19809 14980
rect 19843 14977 19855 15011
rect 19797 14971 19855 14977
rect 14369 14943 14427 14949
rect 14369 14909 14381 14943
rect 14415 14940 14427 14943
rect 16850 14940 16856 14952
rect 14415 14912 15148 14940
rect 16811 14912 16856 14940
rect 14415 14909 14427 14912
rect 14369 14903 14427 14909
rect 12360 14844 12940 14872
rect 13811 14875 13869 14881
rect 11977 14835 12035 14841
rect 13811 14841 13823 14875
rect 13857 14841 13869 14875
rect 13811 14835 13869 14841
rect 10686 14804 10692 14816
rect 10060 14776 10692 14804
rect 8996 14764 9002 14776
rect 10686 14764 10692 14776
rect 10744 14764 10750 14816
rect 10962 14804 10968 14816
rect 10923 14776 10968 14804
rect 10962 14764 10968 14776
rect 11020 14764 11026 14816
rect 12575 14807 12633 14813
rect 12575 14773 12587 14807
rect 12621 14804 12633 14807
rect 12802 14804 12808 14816
rect 12621 14776 12808 14804
rect 12621 14773 12633 14776
rect 12575 14767 12633 14773
rect 12802 14764 12808 14776
rect 12860 14764 12866 14816
rect 14734 14764 14740 14816
rect 14792 14804 14798 14816
rect 15013 14807 15071 14813
rect 15013 14804 15025 14807
rect 14792 14776 15025 14804
rect 14792 14764 14798 14776
rect 15013 14773 15025 14776
rect 15059 14773 15071 14807
rect 15120 14804 15148 14912
rect 16850 14900 16856 14912
rect 16908 14940 16914 14952
rect 17405 14943 17463 14949
rect 17405 14940 17417 14943
rect 16908 14912 17417 14940
rect 16908 14900 16914 14912
rect 17405 14909 17417 14912
rect 17451 14909 17463 14943
rect 17405 14903 17463 14909
rect 15286 14872 15292 14884
rect 15247 14844 15292 14872
rect 15286 14832 15292 14844
rect 15344 14832 15350 14884
rect 15381 14875 15439 14881
rect 15381 14841 15393 14875
rect 15427 14841 15439 14875
rect 15381 14835 15439 14841
rect 17865 14875 17923 14881
rect 17865 14841 17877 14875
rect 17911 14872 17923 14875
rect 18601 14875 18659 14881
rect 17911 14844 18460 14872
rect 17911 14841 17923 14844
rect 17865 14835 17923 14841
rect 15396 14804 15424 14835
rect 15470 14804 15476 14816
rect 15120 14776 15476 14804
rect 15013 14767 15071 14773
rect 15470 14764 15476 14776
rect 15528 14764 15534 14816
rect 18432 14804 18460 14844
rect 18601 14841 18613 14875
rect 18647 14872 18659 14875
rect 18690 14872 18696 14884
rect 18647 14844 18696 14872
rect 18647 14841 18659 14844
rect 18601 14835 18659 14841
rect 18616 14804 18644 14835
rect 18690 14832 18696 14844
rect 18748 14832 18754 14884
rect 18432 14776 18644 14804
rect 1104 14714 20884 14736
rect 1104 14662 8315 14714
rect 8367 14662 8379 14714
rect 8431 14662 8443 14714
rect 8495 14662 8507 14714
rect 8559 14662 15648 14714
rect 15700 14662 15712 14714
rect 15764 14662 15776 14714
rect 15828 14662 15840 14714
rect 15892 14662 20884 14714
rect 1104 14640 20884 14662
rect 6362 14560 6368 14612
rect 6420 14600 6426 14612
rect 9217 14603 9275 14609
rect 6420 14572 9162 14600
rect 6420 14560 6426 14572
rect 6914 14532 6920 14544
rect 5644 14504 6920 14532
rect 2866 14424 2872 14476
rect 2924 14464 2930 14476
rect 4408 14467 4466 14473
rect 4408 14464 4420 14467
rect 2924 14436 4420 14464
rect 2924 14424 2930 14436
rect 4408 14433 4420 14436
rect 4454 14464 4466 14467
rect 4982 14464 4988 14476
rect 4454 14436 4988 14464
rect 4454 14433 4466 14436
rect 4408 14427 4466 14433
rect 4982 14424 4988 14436
rect 5040 14424 5046 14476
rect 5261 14467 5319 14473
rect 5261 14433 5273 14467
rect 5307 14464 5319 14467
rect 5442 14464 5448 14476
rect 5307 14436 5448 14464
rect 5307 14433 5319 14436
rect 5261 14427 5319 14433
rect 5442 14424 5448 14436
rect 5500 14464 5506 14476
rect 5644 14473 5672 14504
rect 6914 14492 6920 14504
rect 6972 14492 6978 14544
rect 7279 14535 7337 14541
rect 7279 14501 7291 14535
rect 7325 14532 7337 14535
rect 7926 14532 7932 14544
rect 7325 14504 7932 14532
rect 7325 14501 7337 14504
rect 7279 14495 7337 14501
rect 7926 14492 7932 14504
rect 7984 14492 7990 14544
rect 5629 14467 5687 14473
rect 5629 14464 5641 14467
rect 5500 14436 5641 14464
rect 5500 14424 5506 14436
rect 5629 14433 5641 14436
rect 5675 14433 5687 14467
rect 5902 14464 5908 14476
rect 5815 14436 5908 14464
rect 5629 14427 5687 14433
rect 5902 14424 5908 14436
rect 5960 14464 5966 14476
rect 9030 14464 9036 14476
rect 5960 14436 9036 14464
rect 5960 14424 5966 14436
rect 9030 14424 9036 14436
rect 9088 14424 9094 14476
rect 9134 14464 9162 14572
rect 9217 14569 9229 14603
rect 9263 14600 9275 14603
rect 9306 14600 9312 14612
rect 9263 14572 9312 14600
rect 9263 14569 9275 14572
rect 9217 14563 9275 14569
rect 9306 14560 9312 14572
rect 9364 14560 9370 14612
rect 9858 14600 9864 14612
rect 9819 14572 9864 14600
rect 9858 14560 9864 14572
rect 9916 14560 9922 14612
rect 10226 14560 10232 14612
rect 10284 14600 10290 14612
rect 10505 14603 10563 14609
rect 10505 14600 10517 14603
rect 10284 14572 10517 14600
rect 10284 14560 10290 14572
rect 10505 14569 10517 14572
rect 10551 14600 10563 14603
rect 10873 14603 10931 14609
rect 10873 14600 10885 14603
rect 10551 14572 10885 14600
rect 10551 14569 10563 14572
rect 10505 14563 10563 14569
rect 10873 14569 10885 14572
rect 10919 14569 10931 14603
rect 12526 14600 12532 14612
rect 12487 14572 12532 14600
rect 10873 14563 10931 14569
rect 12526 14560 12532 14572
rect 12584 14560 12590 14612
rect 13265 14603 13323 14609
rect 13265 14569 13277 14603
rect 13311 14600 13323 14603
rect 13354 14600 13360 14612
rect 13311 14572 13360 14600
rect 13311 14569 13323 14572
rect 13265 14563 13323 14569
rect 13354 14560 13360 14572
rect 13412 14560 13418 14612
rect 14826 14600 14832 14612
rect 14108 14572 14832 14600
rect 10962 14492 10968 14544
rect 11020 14532 11026 14544
rect 11241 14535 11299 14541
rect 11241 14532 11253 14535
rect 11020 14504 11253 14532
rect 11020 14492 11026 14504
rect 11241 14501 11253 14504
rect 11287 14532 11299 14535
rect 11514 14532 11520 14544
rect 11287 14504 11520 14532
rect 11287 14501 11299 14504
rect 11241 14495 11299 14501
rect 11514 14492 11520 14504
rect 11572 14492 11578 14544
rect 11793 14535 11851 14541
rect 11793 14501 11805 14535
rect 11839 14532 11851 14535
rect 11882 14532 11888 14544
rect 11839 14504 11888 14532
rect 11839 14501 11851 14504
rect 11793 14495 11851 14501
rect 11882 14492 11888 14504
rect 11940 14492 11946 14544
rect 13538 14532 13544 14544
rect 13499 14504 13544 14532
rect 13538 14492 13544 14504
rect 13596 14492 13602 14544
rect 14108 14541 14136 14572
rect 14826 14560 14832 14572
rect 14884 14600 14890 14612
rect 15105 14603 15163 14609
rect 15105 14600 15117 14603
rect 14884 14572 15117 14600
rect 14884 14560 14890 14572
rect 15105 14569 15117 14572
rect 15151 14600 15163 14603
rect 15286 14600 15292 14612
rect 15151 14572 15292 14600
rect 15151 14569 15163 14572
rect 15105 14563 15163 14569
rect 15286 14560 15292 14572
rect 15344 14560 15350 14612
rect 15470 14600 15476 14612
rect 15431 14572 15476 14600
rect 15470 14560 15476 14572
rect 15528 14560 15534 14612
rect 15841 14603 15899 14609
rect 15841 14569 15853 14603
rect 15887 14600 15899 14603
rect 15930 14600 15936 14612
rect 15887 14572 15936 14600
rect 15887 14569 15899 14572
rect 15841 14563 15899 14569
rect 15930 14560 15936 14572
rect 15988 14560 15994 14612
rect 17681 14603 17739 14609
rect 17681 14569 17693 14603
rect 17727 14600 17739 14603
rect 17727 14572 18736 14600
rect 17727 14569 17739 14572
rect 17681 14563 17739 14569
rect 14093 14535 14151 14541
rect 14093 14501 14105 14535
rect 14139 14501 14151 14535
rect 14093 14495 14151 14501
rect 17123 14535 17181 14541
rect 17123 14501 17135 14535
rect 17169 14532 17181 14535
rect 17218 14532 17224 14544
rect 17169 14504 17224 14532
rect 17169 14501 17181 14504
rect 17123 14495 17181 14501
rect 17218 14492 17224 14504
rect 17276 14492 17282 14544
rect 18598 14532 18604 14544
rect 18559 14504 18604 14532
rect 18598 14492 18604 14504
rect 18656 14492 18662 14544
rect 18708 14541 18736 14572
rect 18693 14535 18751 14541
rect 18693 14501 18705 14535
rect 18739 14532 18751 14535
rect 19058 14532 19064 14544
rect 18739 14504 19064 14532
rect 18739 14501 18751 14504
rect 18693 14495 18751 14501
rect 19058 14492 19064 14504
rect 19116 14492 19122 14544
rect 19242 14532 19248 14544
rect 19203 14504 19248 14532
rect 19242 14492 19248 14504
rect 19300 14492 19306 14544
rect 10112 14467 10170 14473
rect 10112 14464 10124 14467
rect 9134 14436 10124 14464
rect 10112 14433 10124 14436
rect 10158 14464 10170 14467
rect 10318 14464 10324 14476
rect 10158 14436 10324 14464
rect 10158 14433 10170 14436
rect 10112 14427 10170 14433
rect 10318 14424 10324 14436
rect 10376 14424 10382 14476
rect 15654 14464 15660 14476
rect 14451 14436 15660 14464
rect 6089 14399 6147 14405
rect 6089 14365 6101 14399
rect 6135 14396 6147 14399
rect 6917 14399 6975 14405
rect 6917 14396 6929 14399
rect 6135 14368 6929 14396
rect 6135 14365 6147 14368
rect 6089 14359 6147 14365
rect 6917 14365 6929 14368
rect 6963 14396 6975 14399
rect 8018 14396 8024 14408
rect 6963 14368 8024 14396
rect 6963 14365 6975 14368
rect 6917 14359 6975 14365
rect 8018 14356 8024 14368
rect 8076 14356 8082 14408
rect 9214 14356 9220 14408
rect 9272 14396 9278 14408
rect 11149 14399 11207 14405
rect 11149 14396 11161 14399
rect 9272 14368 11161 14396
rect 9272 14356 9278 14368
rect 11149 14365 11161 14368
rect 11195 14396 11207 14399
rect 11790 14396 11796 14408
rect 11195 14368 11796 14396
rect 11195 14365 11207 14368
rect 11149 14359 11207 14365
rect 11790 14356 11796 14368
rect 11848 14356 11854 14408
rect 13449 14399 13507 14405
rect 13449 14365 13461 14399
rect 13495 14396 13507 14399
rect 13722 14396 13728 14408
rect 13495 14368 13728 14396
rect 13495 14365 13507 14368
rect 13449 14359 13507 14365
rect 13722 14356 13728 14368
rect 13780 14356 13786 14408
rect 4479 14331 4537 14337
rect 4479 14297 4491 14331
rect 4525 14328 4537 14331
rect 6730 14328 6736 14340
rect 4525 14300 6736 14328
rect 4525 14297 4537 14300
rect 4479 14291 4537 14297
rect 6730 14288 6736 14300
rect 6788 14288 6794 14340
rect 6822 14288 6828 14340
rect 6880 14328 6886 14340
rect 9858 14328 9864 14340
rect 6880 14300 9864 14328
rect 6880 14288 6886 14300
rect 9858 14288 9864 14300
rect 9916 14328 9922 14340
rect 10594 14328 10600 14340
rect 9916 14300 10600 14328
rect 9916 14288 9922 14300
rect 10594 14288 10600 14300
rect 10652 14288 10658 14340
rect 12986 14288 12992 14340
rect 13044 14328 13050 14340
rect 14451 14328 14479 14436
rect 15654 14424 15660 14436
rect 15712 14464 15718 14476
rect 16390 14464 16396 14476
rect 15712 14436 16396 14464
rect 15712 14424 15718 14436
rect 16390 14424 16396 14436
rect 16448 14424 16454 14476
rect 16482 14424 16488 14476
rect 16540 14464 16546 14476
rect 16758 14464 16764 14476
rect 16540 14436 16764 14464
rect 16540 14424 16546 14436
rect 16758 14424 16764 14436
rect 16816 14424 16822 14476
rect 16206 14356 16212 14408
rect 16264 14396 16270 14408
rect 16301 14399 16359 14405
rect 16301 14396 16313 14399
rect 16264 14368 16313 14396
rect 16264 14356 16270 14368
rect 16301 14365 16313 14368
rect 16347 14396 16359 14399
rect 17862 14396 17868 14408
rect 16347 14368 17868 14396
rect 16347 14365 16359 14368
rect 16301 14359 16359 14365
rect 17862 14356 17868 14368
rect 17920 14356 17926 14408
rect 13044 14300 14479 14328
rect 13044 14288 13050 14300
rect 4246 14220 4252 14272
rect 4304 14260 4310 14272
rect 4801 14263 4859 14269
rect 4801 14260 4813 14263
rect 4304 14232 4813 14260
rect 4304 14220 4310 14232
rect 4801 14229 4813 14232
rect 4847 14260 4859 14263
rect 5626 14260 5632 14272
rect 4847 14232 5632 14260
rect 4847 14229 4859 14232
rect 4801 14223 4859 14229
rect 5626 14220 5632 14232
rect 5684 14220 5690 14272
rect 7834 14260 7840 14272
rect 7795 14232 7840 14260
rect 7834 14220 7840 14232
rect 7892 14220 7898 14272
rect 8754 14260 8760 14272
rect 8715 14232 8760 14260
rect 8754 14220 8760 14232
rect 8812 14220 8818 14272
rect 10183 14263 10241 14269
rect 10183 14229 10195 14263
rect 10229 14260 10241 14263
rect 10410 14260 10416 14272
rect 10229 14232 10416 14260
rect 10229 14229 10241 14232
rect 10183 14223 10241 14229
rect 10410 14220 10416 14232
rect 10468 14220 10474 14272
rect 12897 14263 12955 14269
rect 12897 14229 12909 14263
rect 12943 14260 12955 14263
rect 13446 14260 13452 14272
rect 12943 14232 13452 14260
rect 12943 14229 12955 14232
rect 12897 14223 12955 14229
rect 13446 14220 13452 14232
rect 13504 14220 13510 14272
rect 14182 14220 14188 14272
rect 14240 14260 14246 14272
rect 14369 14263 14427 14269
rect 14369 14260 14381 14263
rect 14240 14232 14381 14260
rect 14240 14220 14246 14232
rect 14369 14229 14381 14232
rect 14415 14229 14427 14263
rect 14369 14223 14427 14229
rect 1104 14170 20884 14192
rect 1104 14118 4648 14170
rect 4700 14118 4712 14170
rect 4764 14118 4776 14170
rect 4828 14118 4840 14170
rect 4892 14118 11982 14170
rect 12034 14118 12046 14170
rect 12098 14118 12110 14170
rect 12162 14118 12174 14170
rect 12226 14118 19315 14170
rect 19367 14118 19379 14170
rect 19431 14118 19443 14170
rect 19495 14118 19507 14170
rect 19559 14118 20884 14170
rect 1104 14096 20884 14118
rect 4709 14059 4767 14065
rect 4709 14025 4721 14059
rect 4755 14056 4767 14059
rect 4982 14056 4988 14068
rect 4755 14028 4988 14056
rect 4755 14025 4767 14028
rect 4709 14019 4767 14025
rect 4982 14016 4988 14028
rect 5040 14016 5046 14068
rect 5077 14059 5135 14065
rect 5077 14025 5089 14059
rect 5123 14056 5135 14059
rect 5166 14056 5172 14068
rect 5123 14028 5172 14056
rect 5123 14025 5135 14028
rect 5077 14019 5135 14025
rect 5092 13920 5120 14019
rect 5166 14016 5172 14028
rect 5224 14016 5230 14068
rect 8018 14056 8024 14068
rect 7979 14028 8024 14056
rect 8018 14016 8024 14028
rect 8076 14016 8082 14068
rect 13446 14016 13452 14068
rect 13504 14056 13510 14068
rect 13722 14056 13728 14068
rect 13504 14028 13728 14056
rect 13504 14016 13510 14028
rect 13722 14016 13728 14028
rect 13780 14016 13786 14068
rect 14185 14059 14243 14065
rect 14185 14025 14197 14059
rect 14231 14056 14243 14059
rect 14366 14056 14372 14068
rect 14231 14028 14372 14056
rect 14231 14025 14243 14028
rect 14185 14019 14243 14025
rect 14366 14016 14372 14028
rect 14424 14016 14430 14068
rect 15010 14016 15016 14068
rect 15068 14056 15074 14068
rect 15654 14056 15660 14068
rect 15068 14028 15240 14056
rect 15615 14028 15660 14056
rect 15068 14016 15074 14028
rect 6457 13991 6515 13997
rect 6457 13957 6469 13991
rect 6503 13988 6515 13991
rect 7190 13988 7196 14000
rect 6503 13960 7196 13988
rect 6503 13957 6515 13960
rect 6457 13951 6515 13957
rect 7190 13948 7196 13960
rect 7248 13948 7254 14000
rect 7742 13948 7748 14000
rect 7800 13988 7806 14000
rect 10226 13988 10232 14000
rect 7800 13960 10232 13988
rect 7800 13948 7806 13960
rect 10226 13948 10232 13960
rect 10284 13948 10290 14000
rect 5000 13892 5120 13920
rect 5905 13923 5963 13929
rect 4154 13812 4160 13864
rect 4212 13861 4218 13864
rect 4212 13855 4266 13861
rect 4212 13821 4220 13855
rect 4254 13852 4266 13855
rect 5000 13852 5028 13892
rect 5905 13889 5917 13923
rect 5951 13920 5963 13923
rect 8754 13920 8760 13932
rect 5951 13892 8760 13920
rect 5951 13889 5963 13892
rect 5905 13883 5963 13889
rect 8754 13880 8760 13892
rect 8812 13880 8818 13932
rect 9582 13920 9588 13932
rect 8864 13892 9588 13920
rect 4254 13824 5028 13852
rect 4254 13821 4266 13824
rect 4212 13815 4266 13821
rect 4212 13812 4218 13815
rect 5074 13812 5080 13864
rect 5132 13852 5138 13864
rect 5442 13852 5448 13864
rect 5132 13824 5448 13852
rect 5132 13812 5138 13824
rect 5442 13812 5448 13824
rect 5500 13812 5506 13864
rect 5626 13852 5632 13864
rect 5587 13824 5632 13852
rect 5626 13812 5632 13824
rect 5684 13812 5690 13864
rect 6825 13855 6883 13861
rect 6564 13824 6684 13852
rect 5534 13744 5540 13796
rect 5592 13784 5598 13796
rect 6564 13784 6592 13824
rect 6656 13814 6684 13824
rect 6825 13821 6837 13855
rect 6871 13852 6883 13855
rect 6914 13852 6920 13864
rect 6871 13824 6920 13852
rect 6871 13821 6883 13824
rect 6825 13815 6883 13821
rect 6656 13786 6776 13814
rect 6914 13812 6920 13824
rect 6972 13812 6978 13864
rect 8864 13852 8892 13892
rect 9582 13880 9588 13892
rect 9640 13920 9646 13932
rect 10134 13920 10140 13932
rect 9640 13892 10140 13920
rect 9640 13880 9646 13892
rect 10134 13880 10140 13892
rect 10192 13880 10198 13932
rect 10502 13920 10508 13932
rect 10463 13892 10508 13920
rect 10502 13880 10508 13892
rect 10560 13920 10566 13932
rect 11701 13923 11759 13929
rect 11701 13920 11713 13923
rect 10560 13892 11713 13920
rect 10560 13880 10566 13892
rect 11701 13889 11713 13892
rect 11747 13889 11759 13923
rect 11701 13883 11759 13889
rect 12437 13923 12495 13929
rect 12437 13889 12449 13923
rect 12483 13920 12495 13923
rect 12526 13920 12532 13932
rect 12483 13892 12532 13920
rect 12483 13889 12495 13892
rect 12437 13883 12495 13889
rect 12526 13880 12532 13892
rect 12584 13880 12590 13932
rect 15013 13923 15071 13929
rect 15013 13889 15025 13923
rect 15059 13920 15071 13923
rect 15102 13920 15108 13932
rect 15059 13892 15108 13920
rect 15059 13889 15071 13892
rect 15013 13883 15071 13889
rect 15102 13880 15108 13892
rect 15160 13880 15166 13932
rect 9674 13852 9680 13864
rect 7070 13824 8892 13852
rect 9635 13824 9680 13852
rect 5592 13756 6592 13784
rect 6748 13784 6776 13786
rect 7070 13784 7098 13824
rect 9674 13812 9680 13824
rect 9732 13812 9738 13864
rect 10045 13855 10103 13861
rect 10045 13821 10057 13855
rect 10091 13852 10103 13855
rect 10318 13852 10324 13864
rect 10091 13824 10324 13852
rect 10091 13821 10103 13824
rect 10045 13815 10103 13821
rect 10318 13812 10324 13824
rect 10376 13852 10382 13864
rect 15212 13852 15240 14028
rect 15654 14016 15660 14028
rect 15712 14016 15718 14068
rect 17129 14059 17187 14065
rect 17129 14025 17141 14059
rect 17175 14056 17187 14059
rect 17494 14056 17500 14068
rect 17175 14028 17500 14056
rect 17175 14025 17187 14028
rect 17129 14019 17187 14025
rect 17494 14016 17500 14028
rect 17552 14056 17558 14068
rect 17773 14059 17831 14065
rect 17773 14056 17785 14059
rect 17552 14028 17785 14056
rect 17552 14016 17558 14028
rect 17773 14025 17785 14028
rect 17819 14025 17831 14059
rect 19058 14056 19064 14068
rect 19019 14028 19064 14056
rect 17773 14019 17831 14025
rect 17218 13948 17224 14000
rect 17276 13988 17282 14000
rect 17405 13991 17463 13997
rect 17405 13988 17417 13991
rect 17276 13960 17417 13988
rect 17276 13948 17282 13960
rect 17405 13957 17417 13960
rect 17451 13957 17463 13991
rect 17405 13951 17463 13957
rect 16206 13920 16212 13932
rect 16167 13892 16212 13920
rect 16206 13880 16212 13892
rect 16264 13880 16270 13932
rect 10376 13824 13814 13852
rect 10376 13812 10382 13824
rect 8573 13787 8631 13793
rect 8573 13784 8585 13787
rect 6748 13756 7098 13784
rect 7208 13756 8585 13784
rect 5592 13744 5598 13756
rect 7208 13728 7236 13756
rect 8573 13753 8585 13756
rect 8619 13784 8631 13787
rect 9078 13787 9136 13793
rect 9078 13784 9090 13787
rect 8619 13756 9090 13784
rect 8619 13753 8631 13756
rect 8573 13747 8631 13753
rect 9078 13753 9090 13756
rect 9124 13784 9136 13787
rect 10867 13787 10925 13793
rect 9124 13756 9674 13784
rect 9124 13753 9136 13756
rect 9078 13747 9136 13753
rect 4295 13719 4353 13725
rect 4295 13685 4307 13719
rect 4341 13716 4353 13719
rect 5994 13716 6000 13728
rect 4341 13688 6000 13716
rect 4341 13685 4353 13688
rect 4295 13679 4353 13685
rect 5994 13676 6000 13688
rect 6052 13676 6058 13728
rect 6273 13719 6331 13725
rect 6273 13685 6285 13719
rect 6319 13716 6331 13719
rect 6457 13719 6515 13725
rect 6457 13716 6469 13719
rect 6319 13688 6469 13716
rect 6319 13685 6331 13688
rect 6273 13679 6331 13685
rect 6457 13685 6469 13688
rect 6503 13716 6515 13719
rect 6549 13719 6607 13725
rect 6549 13716 6561 13719
rect 6503 13688 6561 13716
rect 6503 13685 6515 13688
rect 6457 13679 6515 13685
rect 6549 13685 6561 13688
rect 6595 13685 6607 13719
rect 7190 13716 7196 13728
rect 7151 13688 7196 13716
rect 6549 13679 6607 13685
rect 7190 13676 7196 13688
rect 7248 13676 7254 13728
rect 7650 13676 7656 13728
rect 7708 13716 7714 13728
rect 7745 13719 7803 13725
rect 7745 13716 7757 13719
rect 7708 13688 7757 13716
rect 7708 13676 7714 13688
rect 7745 13685 7757 13688
rect 7791 13685 7803 13719
rect 9646 13716 9674 13756
rect 10867 13753 10879 13787
rect 10913 13784 10925 13787
rect 12758 13787 12816 13793
rect 12758 13784 12770 13787
rect 10913 13756 12296 13784
rect 10913 13753 10925 13756
rect 10867 13747 10925 13753
rect 10882 13716 10910 13747
rect 11422 13716 11428 13728
rect 9646 13688 10910 13716
rect 11383 13688 11428 13716
rect 7745 13679 7803 13685
rect 11422 13676 11428 13688
rect 11480 13676 11486 13728
rect 12268 13725 12296 13756
rect 12636 13756 12770 13784
rect 12636 13728 12664 13756
rect 12758 13753 12770 13756
rect 12804 13753 12816 13787
rect 12758 13747 12816 13753
rect 12253 13719 12311 13725
rect 12253 13685 12265 13719
rect 12299 13716 12311 13719
rect 12618 13716 12624 13728
rect 12299 13688 12624 13716
rect 12299 13685 12311 13688
rect 12253 13679 12311 13685
rect 12618 13676 12624 13688
rect 12676 13676 12682 13728
rect 13354 13716 13360 13728
rect 13315 13688 13360 13716
rect 13354 13676 13360 13688
rect 13412 13716 13418 13728
rect 13538 13716 13544 13728
rect 13412 13688 13544 13716
rect 13412 13676 13418 13688
rect 13538 13676 13544 13688
rect 13596 13716 13602 13728
rect 13633 13719 13691 13725
rect 13633 13716 13645 13719
rect 13596 13688 13645 13716
rect 13596 13676 13602 13688
rect 13633 13685 13645 13688
rect 13679 13685 13691 13719
rect 13786 13716 13814 13824
rect 15028 13824 15240 13852
rect 16117 13855 16175 13861
rect 15028 13796 15056 13824
rect 16117 13821 16129 13855
rect 16163 13852 16175 13855
rect 17236 13852 17264 13948
rect 16163 13824 17264 13852
rect 16163 13821 16175 13824
rect 16117 13815 16175 13821
rect 16592 13796 16620 13824
rect 14182 13744 14188 13796
rect 14240 13784 14246 13796
rect 14366 13784 14372 13796
rect 14240 13756 14372 13784
rect 14240 13744 14246 13756
rect 14366 13744 14372 13756
rect 14424 13744 14430 13796
rect 14458 13744 14464 13796
rect 14516 13784 14522 13796
rect 14516 13756 14561 13784
rect 14516 13744 14522 13756
rect 15010 13744 15016 13796
rect 15068 13744 15074 13796
rect 16574 13793 16580 13796
rect 16571 13747 16580 13793
rect 16632 13784 16638 13796
rect 17788 13784 17816 14019
rect 19058 14016 19064 14028
rect 19116 14016 19122 14068
rect 19886 14056 19892 14068
rect 19847 14028 19892 14056
rect 19886 14016 19892 14028
rect 19944 14016 19950 14068
rect 19610 13948 19616 14000
rect 19668 13988 19674 14000
rect 20073 13991 20131 13997
rect 20073 13988 20085 13991
rect 19668 13960 20085 13988
rect 19668 13948 19674 13960
rect 20073 13957 20085 13960
rect 20119 13957 20131 13991
rect 20073 13951 20131 13957
rect 18138 13920 18144 13932
rect 18099 13892 18144 13920
rect 18138 13880 18144 13892
rect 18196 13880 18202 13932
rect 19645 13852 19651 13864
rect 19606 13824 19651 13852
rect 19645 13812 19651 13824
rect 19703 13812 19709 13864
rect 18233 13787 18291 13793
rect 18233 13784 18245 13787
rect 16632 13756 16719 13784
rect 17788 13756 18245 13784
rect 16574 13744 16580 13747
rect 16632 13744 16638 13756
rect 18233 13753 18245 13756
rect 18279 13753 18291 13787
rect 18233 13747 18291 13753
rect 18785 13787 18843 13793
rect 18785 13753 18797 13787
rect 18831 13753 18843 13787
rect 18785 13747 18843 13753
rect 15470 13716 15476 13728
rect 13786 13688 15476 13716
rect 13633 13679 13691 13685
rect 15470 13676 15476 13688
rect 15528 13676 15534 13728
rect 18800 13716 18828 13747
rect 18874 13716 18880 13728
rect 18800 13688 18880 13716
rect 18874 13676 18880 13688
rect 18932 13676 18938 13728
rect 19426 13716 19432 13728
rect 19387 13688 19432 13716
rect 19426 13676 19432 13688
rect 19484 13676 19490 13728
rect 1104 13626 20884 13648
rect 1104 13574 8315 13626
rect 8367 13574 8379 13626
rect 8431 13574 8443 13626
rect 8495 13574 8507 13626
rect 8559 13574 15648 13626
rect 15700 13574 15712 13626
rect 15764 13574 15776 13626
rect 15828 13574 15840 13626
rect 15892 13574 20884 13626
rect 1104 13552 20884 13574
rect 2869 13515 2927 13521
rect 2869 13481 2881 13515
rect 2915 13512 2927 13515
rect 5534 13512 5540 13524
rect 2915 13484 5540 13512
rect 2915 13481 2927 13484
rect 2869 13475 2927 13481
rect 5534 13472 5540 13484
rect 5592 13472 5598 13524
rect 5718 13472 5724 13524
rect 5776 13512 5782 13524
rect 11330 13512 11336 13524
rect 5776 13484 11336 13512
rect 5776 13472 5782 13484
rect 11330 13472 11336 13484
rect 11388 13472 11394 13524
rect 11514 13512 11520 13524
rect 11475 13484 11520 13512
rect 11514 13472 11520 13484
rect 11572 13472 11578 13524
rect 13446 13512 13452 13524
rect 13407 13484 13452 13512
rect 13446 13472 13452 13484
rect 13504 13472 13510 13524
rect 16209 13515 16267 13521
rect 16209 13481 16221 13515
rect 16255 13512 16267 13515
rect 16298 13512 16304 13524
rect 16255 13484 16304 13512
rect 16255 13481 16267 13484
rect 16209 13475 16267 13481
rect 16298 13472 16304 13484
rect 16356 13472 16362 13524
rect 16758 13472 16764 13524
rect 16816 13512 16822 13524
rect 17497 13515 17555 13521
rect 17497 13512 17509 13515
rect 16816 13484 17509 13512
rect 16816 13472 16822 13484
rect 17497 13481 17509 13484
rect 17543 13481 17555 13515
rect 18138 13512 18144 13524
rect 18099 13484 18144 13512
rect 17497 13475 17555 13481
rect 18138 13472 18144 13484
rect 18196 13472 18202 13524
rect 3970 13404 3976 13456
rect 4028 13444 4034 13456
rect 6546 13444 6552 13456
rect 4028 13416 5396 13444
rect 6507 13416 6552 13444
rect 4028 13404 4034 13416
rect 5368 13388 5396 13416
rect 6546 13404 6552 13416
rect 6604 13404 6610 13456
rect 6822 13404 6828 13456
rect 6880 13444 6886 13456
rect 7377 13447 7435 13453
rect 7377 13444 7389 13447
rect 6880 13416 7389 13444
rect 6880 13404 6886 13416
rect 7377 13413 7389 13416
rect 7423 13413 7435 13447
rect 7377 13407 7435 13413
rect 7834 13404 7840 13456
rect 7892 13444 7898 13456
rect 8113 13447 8171 13453
rect 8113 13444 8125 13447
rect 7892 13416 8125 13444
rect 7892 13404 7898 13416
rect 8113 13413 8125 13416
rect 8159 13413 8171 13447
rect 10686 13444 10692 13456
rect 10599 13416 10692 13444
rect 8113 13407 8171 13413
rect 10686 13404 10692 13416
rect 10744 13444 10750 13456
rect 11422 13444 11428 13456
rect 10744 13416 11428 13444
rect 10744 13404 10750 13416
rect 11422 13404 11428 13416
rect 11480 13404 11486 13456
rect 11882 13404 11888 13456
rect 11940 13444 11946 13456
rect 12253 13447 12311 13453
rect 12253 13444 12265 13447
rect 11940 13416 12265 13444
rect 11940 13404 11946 13416
rect 12253 13413 12265 13416
rect 12299 13444 12311 13447
rect 13354 13444 13360 13456
rect 12299 13416 13360 13444
rect 12299 13413 12311 13416
rect 12253 13407 12311 13413
rect 13354 13404 13360 13416
rect 13412 13404 13418 13456
rect 13814 13404 13820 13456
rect 13872 13444 13878 13456
rect 13872 13416 13917 13444
rect 13872 13404 13878 13416
rect 16390 13404 16396 13456
rect 16448 13444 16454 13456
rect 16574 13444 16580 13456
rect 16448 13416 16580 13444
rect 16448 13404 16454 13416
rect 16574 13404 16580 13416
rect 16632 13453 16638 13456
rect 16632 13447 16680 13453
rect 16632 13413 16634 13447
rect 16668 13413 16680 13447
rect 18414 13444 18420 13456
rect 18375 13416 18420 13444
rect 16632 13407 16680 13413
rect 16632 13404 16638 13407
rect 18414 13404 18420 13416
rect 18472 13404 18478 13456
rect 5074 13376 5080 13388
rect 4987 13348 5080 13376
rect 5074 13336 5080 13348
rect 5132 13376 5138 13388
rect 5350 13376 5356 13388
rect 5132 13348 5212 13376
rect 5311 13348 5356 13376
rect 5132 13336 5138 13348
rect 2682 13268 2688 13320
rect 2740 13308 2746 13320
rect 2866 13308 2872 13320
rect 2740 13280 2872 13308
rect 2740 13268 2746 13280
rect 2866 13268 2872 13280
rect 2924 13268 2930 13320
rect 5184 13240 5212 13348
rect 5350 13336 5356 13348
rect 5408 13336 5414 13388
rect 5537 13379 5595 13385
rect 5537 13345 5549 13379
rect 5583 13376 5595 13379
rect 6270 13376 6276 13388
rect 5583 13348 6276 13376
rect 5583 13345 5595 13348
rect 5537 13339 5595 13345
rect 6270 13336 6276 13348
rect 6328 13336 6334 13388
rect 15356 13379 15414 13385
rect 15356 13345 15368 13379
rect 15402 13376 15414 13379
rect 15470 13376 15476 13388
rect 15402 13348 15476 13376
rect 15402 13345 15414 13348
rect 15356 13339 15414 13345
rect 15470 13336 15476 13348
rect 15528 13376 15534 13388
rect 17402 13376 17408 13388
rect 15528 13348 17408 13376
rect 15528 13336 15534 13348
rect 17402 13336 17408 13348
rect 17460 13336 17466 13388
rect 5994 13268 6000 13320
rect 6052 13308 6058 13320
rect 6457 13311 6515 13317
rect 6457 13308 6469 13311
rect 6052 13280 6469 13308
rect 6052 13268 6058 13280
rect 6457 13277 6469 13280
rect 6503 13277 6515 13311
rect 6457 13271 6515 13277
rect 7101 13311 7159 13317
rect 7101 13277 7113 13311
rect 7147 13308 7159 13311
rect 7558 13308 7564 13320
rect 7147 13280 7564 13308
rect 7147 13277 7159 13280
rect 7101 13271 7159 13277
rect 7558 13268 7564 13280
rect 7616 13268 7622 13320
rect 8021 13311 8079 13317
rect 8021 13308 8033 13311
rect 7760 13280 8033 13308
rect 5184 13212 5580 13240
rect 5552 13184 5580 13212
rect 7760 13184 7788 13280
rect 8021 13277 8033 13280
rect 8067 13277 8079 13311
rect 8662 13308 8668 13320
rect 8623 13280 8668 13308
rect 8021 13271 8079 13277
rect 8662 13268 8668 13280
rect 8720 13268 8726 13320
rect 9950 13268 9956 13320
rect 10008 13308 10014 13320
rect 10597 13311 10655 13317
rect 10597 13308 10609 13311
rect 10008 13280 10609 13308
rect 10008 13268 10014 13280
rect 10597 13277 10609 13280
rect 10643 13308 10655 13311
rect 10686 13308 10692 13320
rect 10643 13280 10692 13308
rect 10643 13277 10655 13280
rect 10597 13271 10655 13277
rect 10686 13268 10692 13280
rect 10744 13268 10750 13320
rect 12161 13311 12219 13317
rect 12161 13308 12173 13311
rect 10882 13280 12173 13308
rect 10410 13200 10416 13252
rect 10468 13240 10474 13252
rect 10882 13240 10910 13280
rect 12161 13277 12173 13280
rect 12207 13308 12219 13311
rect 12342 13308 12348 13320
rect 12207 13280 12348 13308
rect 12207 13277 12219 13280
rect 12161 13271 12219 13277
rect 12342 13268 12348 13280
rect 12400 13268 12406 13320
rect 12802 13268 12808 13320
rect 12860 13308 12866 13320
rect 13446 13308 13452 13320
rect 12860 13280 13452 13308
rect 12860 13268 12866 13280
rect 13446 13268 13452 13280
rect 13504 13308 13510 13320
rect 13725 13311 13783 13317
rect 13725 13308 13737 13311
rect 13504 13280 13737 13308
rect 13504 13268 13510 13280
rect 13725 13277 13737 13280
rect 13771 13277 13783 13311
rect 14366 13308 14372 13320
rect 14279 13280 14372 13308
rect 13725 13271 13783 13277
rect 14366 13268 14372 13280
rect 14424 13308 14430 13320
rect 16022 13308 16028 13320
rect 14424 13280 16028 13308
rect 14424 13268 14430 13280
rect 16022 13268 16028 13280
rect 16080 13268 16086 13320
rect 16114 13268 16120 13320
rect 16172 13308 16178 13320
rect 16301 13311 16359 13317
rect 16301 13308 16313 13311
rect 16172 13280 16313 13308
rect 16172 13268 16178 13280
rect 16301 13277 16313 13280
rect 16347 13308 16359 13311
rect 16666 13308 16672 13320
rect 16347 13280 16672 13308
rect 16347 13277 16359 13280
rect 16301 13271 16359 13277
rect 16666 13268 16672 13280
rect 16724 13268 16730 13320
rect 18322 13308 18328 13320
rect 18283 13280 18328 13308
rect 18322 13268 18328 13280
rect 18380 13268 18386 13320
rect 18598 13308 18604 13320
rect 18511 13280 18604 13308
rect 18598 13268 18604 13280
rect 18656 13308 18662 13320
rect 19426 13308 19432 13320
rect 18656 13280 19432 13308
rect 18656 13268 18662 13280
rect 19426 13268 19432 13280
rect 19484 13268 19490 13320
rect 11146 13240 11152 13252
rect 10468 13212 10910 13240
rect 11107 13212 11152 13240
rect 10468 13200 10474 13212
rect 11146 13200 11152 13212
rect 11204 13200 11210 13252
rect 12713 13243 12771 13249
rect 12713 13209 12725 13243
rect 12759 13240 12771 13243
rect 14384 13240 14412 13268
rect 12759 13212 14412 13240
rect 12759 13209 12771 13212
rect 12713 13203 12771 13209
rect 16206 13200 16212 13252
rect 16264 13240 16270 13252
rect 18616 13240 18644 13268
rect 16264 13212 18644 13240
rect 16264 13200 16270 13212
rect 2866 13172 2872 13184
rect 2827 13144 2872 13172
rect 2866 13132 2872 13144
rect 2924 13132 2930 13184
rect 3099 13175 3157 13181
rect 3099 13141 3111 13175
rect 3145 13172 3157 13175
rect 4982 13172 4988 13184
rect 3145 13144 4988 13172
rect 3145 13141 3157 13144
rect 3099 13135 3157 13141
rect 4982 13132 4988 13144
rect 5040 13132 5046 13184
rect 5534 13132 5540 13184
rect 5592 13172 5598 13184
rect 5813 13175 5871 13181
rect 5813 13172 5825 13175
rect 5592 13144 5825 13172
rect 5592 13132 5598 13144
rect 5813 13141 5825 13144
rect 5859 13141 5871 13175
rect 5813 13135 5871 13141
rect 5902 13132 5908 13184
rect 5960 13172 5966 13184
rect 6270 13172 6276 13184
rect 5960 13144 6276 13172
rect 5960 13132 5966 13144
rect 6270 13132 6276 13144
rect 6328 13132 6334 13184
rect 7742 13172 7748 13184
rect 7703 13144 7748 13172
rect 7742 13132 7748 13144
rect 7800 13132 7806 13184
rect 10318 13172 10324 13184
rect 10279 13144 10324 13172
rect 10318 13132 10324 13144
rect 10376 13132 10382 13184
rect 11514 13132 11520 13184
rect 11572 13172 11578 13184
rect 11790 13172 11796 13184
rect 11572 13144 11796 13172
rect 11572 13132 11578 13144
rect 11790 13132 11796 13144
rect 11848 13172 11854 13184
rect 11885 13175 11943 13181
rect 11885 13172 11897 13175
rect 11848 13144 11897 13172
rect 11848 13132 11854 13144
rect 11885 13141 11897 13144
rect 11931 13141 11943 13175
rect 11885 13135 11943 13141
rect 15427 13175 15485 13181
rect 15427 13141 15439 13175
rect 15473 13172 15485 13175
rect 16482 13172 16488 13184
rect 15473 13144 16488 13172
rect 15473 13141 15485 13144
rect 15427 13135 15485 13141
rect 16482 13132 16488 13144
rect 16540 13132 16546 13184
rect 16574 13132 16580 13184
rect 16632 13172 16638 13184
rect 17221 13175 17279 13181
rect 17221 13172 17233 13175
rect 16632 13144 17233 13172
rect 16632 13132 16638 13144
rect 17221 13141 17233 13144
rect 17267 13141 17279 13175
rect 17221 13135 17279 13141
rect 1104 13082 20884 13104
rect 1104 13030 4648 13082
rect 4700 13030 4712 13082
rect 4764 13030 4776 13082
rect 4828 13030 4840 13082
rect 4892 13030 11982 13082
rect 12034 13030 12046 13082
rect 12098 13030 12110 13082
rect 12162 13030 12174 13082
rect 12226 13030 19315 13082
rect 19367 13030 19379 13082
rect 19431 13030 19443 13082
rect 19495 13030 19507 13082
rect 19559 13030 20884 13082
rect 1104 13008 20884 13030
rect 2685 12971 2743 12977
rect 2685 12937 2697 12971
rect 2731 12968 2743 12971
rect 2774 12968 2780 12980
rect 2731 12940 2780 12968
rect 2731 12937 2743 12940
rect 2685 12931 2743 12937
rect 2200 12767 2258 12773
rect 2200 12733 2212 12767
rect 2246 12764 2258 12767
rect 2700 12764 2728 12931
rect 2774 12928 2780 12940
rect 2832 12928 2838 12980
rect 2866 12928 2872 12980
rect 2924 12968 2930 12980
rect 2961 12971 3019 12977
rect 2961 12968 2973 12971
rect 2924 12940 2973 12968
rect 2924 12928 2930 12940
rect 2961 12937 2973 12940
rect 3007 12937 3019 12971
rect 3970 12968 3976 12980
rect 3931 12940 3976 12968
rect 2961 12931 3019 12937
rect 3970 12928 3976 12940
rect 4028 12928 4034 12980
rect 4295 12971 4353 12977
rect 4295 12937 4307 12971
rect 4341 12968 4353 12971
rect 9766 12968 9772 12980
rect 4341 12940 9772 12968
rect 4341 12937 4353 12940
rect 4295 12931 4353 12937
rect 9766 12928 9772 12940
rect 9824 12928 9830 12980
rect 11422 12968 11428 12980
rect 11383 12940 11428 12968
rect 11422 12928 11428 12940
rect 11480 12928 11486 12980
rect 13633 12971 13691 12977
rect 13633 12937 13645 12971
rect 13679 12968 13691 12971
rect 13814 12968 13820 12980
rect 13679 12940 13820 12968
rect 13679 12937 13691 12940
rect 13633 12931 13691 12937
rect 13814 12928 13820 12940
rect 13872 12968 13878 12980
rect 13909 12971 13967 12977
rect 13909 12968 13921 12971
rect 13872 12940 13921 12968
rect 13872 12928 13878 12940
rect 13909 12937 13921 12940
rect 13955 12968 13967 12971
rect 14277 12971 14335 12977
rect 14277 12968 14289 12971
rect 13955 12940 14289 12968
rect 13955 12937 13967 12940
rect 13909 12931 13967 12937
rect 14277 12937 14289 12940
rect 14323 12937 14335 12971
rect 15470 12968 15476 12980
rect 15431 12940 15476 12968
rect 14277 12931 14335 12937
rect 4614 12860 4620 12912
rect 4672 12900 4678 12912
rect 10318 12900 10324 12912
rect 4672 12872 10324 12900
rect 4672 12860 4678 12872
rect 10318 12860 10324 12872
rect 10376 12900 10382 12912
rect 11882 12900 11888 12912
rect 10376 12872 10456 12900
rect 11843 12872 11888 12900
rect 10376 12860 10382 12872
rect 6086 12792 6092 12844
rect 6144 12832 6150 12844
rect 7101 12835 7159 12841
rect 7101 12832 7113 12835
rect 6144 12804 7113 12832
rect 6144 12792 6150 12804
rect 7101 12801 7113 12804
rect 7147 12832 7159 12835
rect 7374 12832 7380 12844
rect 7147 12804 7380 12832
rect 7147 12801 7159 12804
rect 7101 12795 7159 12801
rect 7374 12792 7380 12804
rect 7432 12792 7438 12844
rect 7558 12792 7564 12844
rect 7616 12832 7622 12844
rect 7616 12804 8248 12832
rect 7616 12792 7622 12804
rect 2246 12736 2728 12764
rect 2246 12733 2258 12736
rect 2200 12727 2258 12733
rect 2958 12724 2964 12776
rect 3016 12764 3022 12776
rect 3180 12767 3238 12773
rect 3180 12764 3192 12767
rect 3016 12736 3192 12764
rect 3016 12724 3022 12736
rect 3180 12733 3192 12736
rect 3226 12764 3238 12767
rect 3605 12767 3663 12773
rect 3605 12764 3617 12767
rect 3226 12736 3617 12764
rect 3226 12733 3238 12736
rect 3180 12727 3238 12733
rect 3605 12733 3617 12736
rect 3651 12764 3663 12767
rect 4224 12767 4282 12773
rect 4224 12764 4236 12767
rect 3651 12736 4236 12764
rect 3651 12733 3663 12736
rect 3605 12727 3663 12733
rect 4224 12733 4236 12736
rect 4270 12764 4282 12767
rect 5077 12767 5135 12773
rect 4270 12736 4752 12764
rect 4270 12733 4282 12736
rect 4224 12727 4282 12733
rect 2271 12631 2329 12637
rect 2271 12597 2283 12631
rect 2317 12628 2329 12631
rect 3050 12628 3056 12640
rect 2317 12600 3056 12628
rect 2317 12597 2329 12600
rect 2271 12591 2329 12597
rect 3050 12588 3056 12600
rect 3108 12588 3114 12640
rect 3283 12631 3341 12637
rect 3283 12597 3295 12631
rect 3329 12628 3341 12631
rect 3510 12628 3516 12640
rect 3329 12600 3516 12628
rect 3329 12597 3341 12600
rect 3283 12591 3341 12597
rect 3510 12588 3516 12600
rect 3568 12588 3574 12640
rect 4724 12637 4752 12736
rect 5077 12733 5089 12767
rect 5123 12764 5135 12767
rect 5445 12767 5503 12773
rect 5445 12764 5457 12767
rect 5123 12736 5457 12764
rect 5123 12733 5135 12736
rect 5077 12727 5135 12733
rect 5445 12733 5457 12736
rect 5491 12764 5503 12767
rect 5534 12764 5540 12776
rect 5491 12736 5540 12764
rect 5491 12733 5503 12736
rect 5445 12727 5503 12733
rect 5534 12724 5540 12736
rect 5592 12724 5598 12776
rect 5721 12767 5779 12773
rect 5721 12733 5733 12767
rect 5767 12733 5779 12767
rect 5721 12727 5779 12733
rect 5905 12767 5963 12773
rect 5905 12733 5917 12767
rect 5951 12764 5963 12767
rect 6178 12764 6184 12776
rect 5951 12736 6184 12764
rect 5951 12733 5963 12736
rect 5905 12727 5963 12733
rect 5626 12656 5632 12708
rect 5684 12696 5690 12708
rect 5736 12696 5764 12727
rect 6178 12724 6184 12736
rect 6236 12724 6242 12776
rect 8220 12764 8248 12804
rect 8662 12792 8668 12844
rect 8720 12832 8726 12844
rect 10428 12841 10456 12872
rect 11882 12860 11888 12872
rect 11940 12860 11946 12912
rect 9125 12835 9183 12841
rect 9125 12832 9137 12835
rect 8720 12804 9137 12832
rect 8720 12792 8726 12804
rect 9125 12801 9137 12804
rect 9171 12801 9183 12835
rect 9125 12795 9183 12801
rect 10413 12835 10471 12841
rect 10413 12801 10425 12835
rect 10459 12801 10471 12835
rect 10413 12795 10471 12801
rect 12253 12835 12311 12841
rect 12253 12801 12265 12835
rect 12299 12832 12311 12835
rect 12710 12832 12716 12844
rect 12299 12804 12716 12832
rect 12299 12801 12311 12804
rect 12253 12795 12311 12801
rect 12710 12792 12716 12804
rect 12768 12792 12774 12844
rect 8220 12736 8708 12764
rect 7193 12699 7251 12705
rect 5684 12668 6316 12696
rect 5684 12656 5690 12668
rect 4709 12631 4767 12637
rect 4709 12597 4721 12631
rect 4755 12628 4767 12631
rect 4982 12628 4988 12640
rect 4755 12600 4988 12628
rect 4755 12597 4767 12600
rect 4709 12591 4767 12597
rect 4982 12588 4988 12600
rect 5040 12588 5046 12640
rect 6288 12637 6316 12668
rect 7193 12665 7205 12699
rect 7239 12665 7251 12699
rect 7742 12696 7748 12708
rect 7655 12668 7748 12696
rect 7193 12659 7251 12665
rect 6273 12631 6331 12637
rect 6273 12597 6285 12631
rect 6319 12628 6331 12631
rect 6362 12628 6368 12640
rect 6319 12600 6368 12628
rect 6319 12597 6331 12600
rect 6273 12591 6331 12597
rect 6362 12588 6368 12600
rect 6420 12588 6426 12640
rect 6546 12588 6552 12640
rect 6604 12628 6610 12640
rect 6641 12631 6699 12637
rect 6641 12628 6653 12631
rect 6604 12600 6653 12628
rect 6604 12588 6610 12600
rect 6641 12597 6653 12600
rect 6687 12628 6699 12631
rect 7208 12628 7236 12659
rect 7742 12656 7748 12668
rect 7800 12696 7806 12708
rect 8202 12696 8208 12708
rect 7800 12668 8208 12696
rect 7800 12656 7806 12668
rect 8202 12656 8208 12668
rect 8260 12656 8266 12708
rect 8680 12696 8708 12736
rect 8846 12696 8852 12708
rect 8680 12668 8852 12696
rect 8846 12656 8852 12668
rect 8904 12656 8910 12708
rect 8941 12699 8999 12705
rect 8941 12665 8953 12699
rect 8987 12696 8999 12699
rect 9674 12696 9680 12708
rect 8987 12668 9680 12696
rect 8987 12665 8999 12668
rect 8941 12659 8999 12665
rect 7650 12628 7656 12640
rect 6687 12600 7656 12628
rect 6687 12597 6699 12600
rect 6641 12591 6699 12597
rect 7650 12588 7656 12600
rect 7708 12628 7714 12640
rect 8021 12631 8079 12637
rect 8021 12628 8033 12631
rect 7708 12600 8033 12628
rect 7708 12588 7714 12600
rect 8021 12597 8033 12600
rect 8067 12597 8079 12631
rect 8021 12591 8079 12597
rect 8665 12631 8723 12637
rect 8665 12597 8677 12631
rect 8711 12628 8723 12631
rect 8956 12628 8984 12659
rect 9674 12656 9680 12668
rect 9732 12656 9738 12708
rect 10502 12656 10508 12708
rect 10560 12696 10566 12708
rect 11057 12699 11115 12705
rect 10560 12668 10605 12696
rect 10560 12656 10566 12668
rect 11057 12665 11069 12699
rect 11103 12696 11115 12699
rect 11146 12696 11152 12708
rect 11103 12668 11152 12696
rect 11103 12665 11115 12668
rect 11057 12659 11115 12665
rect 11146 12656 11152 12668
rect 11204 12696 11210 12708
rect 11882 12696 11888 12708
rect 11204 12668 11888 12696
rect 11204 12656 11210 12668
rect 11882 12656 11888 12668
rect 11940 12656 11946 12708
rect 12710 12656 12716 12708
rect 12768 12696 12774 12708
rect 13034 12699 13092 12705
rect 13034 12696 13046 12699
rect 12768 12668 13046 12696
rect 12768 12656 12774 12668
rect 13034 12665 13046 12668
rect 13080 12665 13092 12699
rect 14292 12696 14320 12931
rect 15470 12928 15476 12940
rect 15528 12928 15534 12980
rect 18046 12968 18052 12980
rect 17925 12940 18052 12968
rect 14458 12860 14464 12912
rect 14516 12900 14522 12912
rect 17925 12900 17953 12940
rect 18046 12928 18052 12940
rect 18104 12968 18110 12980
rect 18690 12968 18696 12980
rect 18104 12940 18696 12968
rect 18104 12928 18110 12940
rect 18690 12928 18696 12940
rect 18748 12928 18754 12980
rect 18782 12900 18788 12912
rect 14516 12872 17953 12900
rect 18616 12872 18788 12900
rect 14516 12860 14522 12872
rect 14550 12832 14556 12844
rect 14511 12804 14556 12832
rect 14550 12792 14556 12804
rect 14608 12792 14614 12844
rect 14826 12832 14832 12844
rect 14787 12804 14832 12832
rect 14826 12792 14832 12804
rect 14884 12792 14890 12844
rect 16117 12835 16175 12841
rect 16117 12801 16129 12835
rect 16163 12832 16175 12835
rect 16298 12832 16304 12844
rect 16163 12804 16304 12832
rect 16163 12801 16175 12804
rect 16117 12795 16175 12801
rect 16298 12792 16304 12804
rect 16356 12792 16362 12844
rect 18616 12841 18644 12872
rect 18782 12860 18788 12872
rect 18840 12900 18846 12912
rect 19150 12900 19156 12912
rect 18840 12872 19156 12900
rect 18840 12860 18846 12872
rect 19150 12860 19156 12872
rect 19208 12860 19214 12912
rect 18601 12835 18659 12841
rect 18601 12801 18613 12835
rect 18647 12801 18659 12835
rect 18874 12832 18880 12844
rect 18835 12804 18880 12832
rect 18601 12795 18659 12801
rect 18874 12792 18880 12804
rect 18932 12792 18938 12844
rect 17037 12767 17095 12773
rect 17037 12733 17049 12767
rect 17083 12764 17095 12767
rect 17773 12767 17831 12773
rect 17773 12764 17785 12767
rect 17083 12736 17785 12764
rect 17083 12733 17095 12736
rect 17037 12727 17095 12733
rect 17773 12733 17785 12736
rect 17819 12764 17831 12767
rect 18325 12767 18383 12773
rect 18325 12764 18337 12767
rect 17819 12736 18337 12764
rect 17819 12733 17831 12736
rect 17773 12727 17831 12733
rect 18325 12733 18337 12736
rect 18371 12764 18383 12767
rect 18414 12764 18420 12776
rect 18371 12736 18420 12764
rect 18371 12733 18383 12736
rect 18325 12727 18383 12733
rect 14645 12699 14703 12705
rect 14645 12696 14657 12699
rect 14292 12668 14657 12696
rect 13034 12659 13092 12665
rect 14645 12665 14657 12668
rect 14691 12665 14703 12699
rect 16390 12696 16396 12708
rect 14645 12659 14703 12665
rect 15948 12668 16396 12696
rect 8711 12600 8984 12628
rect 10229 12631 10287 12637
rect 8711 12597 8723 12600
rect 8665 12591 8723 12597
rect 10229 12597 10241 12631
rect 10275 12628 10287 12631
rect 10520 12628 10548 12656
rect 15948 12640 15976 12668
rect 16390 12656 16396 12668
rect 16448 12705 16454 12708
rect 16448 12699 16496 12705
rect 16448 12665 16450 12699
rect 16484 12665 16496 12699
rect 16448 12659 16496 12665
rect 16448 12656 16454 12659
rect 15930 12628 15936 12640
rect 10275 12600 10548 12628
rect 15891 12600 15936 12628
rect 10275 12597 10287 12600
rect 10229 12591 10287 12597
rect 15930 12588 15936 12600
rect 15988 12588 15994 12640
rect 18340 12628 18368 12727
rect 18414 12724 18420 12736
rect 18472 12724 18478 12776
rect 18693 12699 18751 12705
rect 18693 12665 18705 12699
rect 18739 12665 18751 12699
rect 18693 12659 18751 12665
rect 18708 12628 18736 12659
rect 18340 12600 18736 12628
rect 1104 12538 20884 12560
rect 1104 12486 8315 12538
rect 8367 12486 8379 12538
rect 8431 12486 8443 12538
rect 8495 12486 8507 12538
rect 8559 12486 15648 12538
rect 15700 12486 15712 12538
rect 15764 12486 15776 12538
rect 15828 12486 15840 12538
rect 15892 12486 20884 12538
rect 1104 12464 20884 12486
rect 3099 12427 3157 12433
rect 3099 12393 3111 12427
rect 3145 12424 3157 12427
rect 4614 12424 4620 12436
rect 3145 12396 4620 12424
rect 3145 12393 3157 12396
rect 3099 12387 3157 12393
rect 4614 12384 4620 12396
rect 4672 12384 4678 12436
rect 5994 12424 6000 12436
rect 5955 12396 6000 12424
rect 5994 12384 6000 12396
rect 6052 12384 6058 12436
rect 7374 12424 7380 12436
rect 7335 12396 7380 12424
rect 7374 12384 7380 12396
rect 7432 12384 7438 12436
rect 7834 12424 7840 12436
rect 7795 12396 7840 12424
rect 7834 12384 7840 12396
rect 7892 12384 7898 12436
rect 8846 12384 8852 12436
rect 8904 12424 8910 12436
rect 8941 12427 8999 12433
rect 8941 12424 8953 12427
rect 8904 12396 8953 12424
rect 8904 12384 8910 12396
rect 8941 12393 8953 12396
rect 8987 12424 8999 12427
rect 10686 12424 10692 12436
rect 8987 12396 10456 12424
rect 10647 12396 10692 12424
rect 8987 12393 8999 12396
rect 8941 12387 8999 12393
rect 5534 12356 5540 12368
rect 4908 12328 5540 12356
rect 1949 12291 2007 12297
rect 1949 12257 1961 12291
rect 1995 12288 2007 12291
rect 2038 12288 2044 12300
rect 1995 12260 2044 12288
rect 1995 12257 2007 12260
rect 1949 12251 2007 12257
rect 2038 12248 2044 12260
rect 2096 12248 2102 12300
rect 2774 12248 2780 12300
rect 2832 12288 2838 12300
rect 4908 12297 4936 12328
rect 5534 12316 5540 12328
rect 5592 12316 5598 12368
rect 6454 12356 6460 12368
rect 6415 12328 6460 12356
rect 6454 12316 6460 12328
rect 6512 12316 6518 12368
rect 8113 12359 8171 12365
rect 8113 12356 8125 12359
rect 7116 12328 8125 12356
rect 2996 12291 3054 12297
rect 2996 12288 3008 12291
rect 2832 12260 3008 12288
rect 2832 12248 2838 12260
rect 2996 12257 3008 12260
rect 3042 12257 3054 12291
rect 2996 12251 3054 12257
rect 4893 12291 4951 12297
rect 4893 12257 4905 12291
rect 4939 12257 4951 12291
rect 4893 12251 4951 12257
rect 5169 12291 5227 12297
rect 5169 12257 5181 12291
rect 5215 12288 5227 12291
rect 5258 12288 5264 12300
rect 5215 12260 5264 12288
rect 5215 12257 5227 12260
rect 5169 12251 5227 12257
rect 3697 12223 3755 12229
rect 3697 12189 3709 12223
rect 3743 12220 3755 12223
rect 3878 12220 3884 12232
rect 3743 12192 3884 12220
rect 3743 12189 3755 12192
rect 3697 12183 3755 12189
rect 3878 12180 3884 12192
rect 3936 12220 3942 12232
rect 5184 12220 5212 12251
rect 5258 12248 5264 12260
rect 5316 12248 5322 12300
rect 7116 12297 7144 12328
rect 8113 12325 8125 12328
rect 8159 12356 8171 12359
rect 9030 12356 9036 12368
rect 8159 12328 9036 12356
rect 8159 12325 8171 12328
rect 8113 12319 8171 12325
rect 9030 12316 9036 12328
rect 9088 12356 9094 12368
rect 10428 12365 10456 12396
rect 10686 12384 10692 12396
rect 10744 12384 10750 12436
rect 12342 12424 12348 12436
rect 12303 12396 12348 12424
rect 12342 12384 12348 12396
rect 12400 12384 12406 12436
rect 13446 12424 13452 12436
rect 13407 12396 13452 12424
rect 13446 12384 13452 12396
rect 13504 12384 13510 12436
rect 14550 12384 14556 12436
rect 14608 12424 14614 12436
rect 14645 12427 14703 12433
rect 14645 12424 14657 12427
rect 14608 12396 14657 12424
rect 14608 12384 14614 12396
rect 14645 12393 14657 12396
rect 14691 12393 14703 12427
rect 16666 12424 16672 12436
rect 16627 12396 16672 12424
rect 14645 12387 14703 12393
rect 16666 12384 16672 12396
rect 16724 12384 16730 12436
rect 17402 12384 17408 12436
rect 17460 12424 17466 12436
rect 17497 12427 17555 12433
rect 17497 12424 17509 12427
rect 17460 12396 17509 12424
rect 17460 12384 17466 12396
rect 17497 12393 17509 12396
rect 17543 12393 17555 12427
rect 18322 12424 18328 12436
rect 18283 12396 18328 12424
rect 17497 12387 17555 12393
rect 18322 12384 18328 12396
rect 18380 12384 18386 12436
rect 18782 12424 18788 12436
rect 18743 12396 18788 12424
rect 18782 12384 18788 12396
rect 18840 12384 18846 12436
rect 9861 12359 9919 12365
rect 9861 12356 9873 12359
rect 9088 12328 9873 12356
rect 9088 12316 9094 12328
rect 9861 12325 9873 12328
rect 9907 12325 9919 12359
rect 9861 12319 9919 12325
rect 10413 12359 10471 12365
rect 10413 12325 10425 12359
rect 10459 12325 10471 12359
rect 10413 12319 10471 12325
rect 11425 12359 11483 12365
rect 11425 12325 11437 12359
rect 11471 12356 11483 12359
rect 11606 12356 11612 12368
rect 11471 12328 11612 12356
rect 11471 12325 11483 12328
rect 11425 12319 11483 12325
rect 11606 12316 11612 12328
rect 11664 12316 11670 12368
rect 13814 12316 13820 12368
rect 13872 12356 13878 12368
rect 14369 12359 14427 12365
rect 13872 12328 13917 12356
rect 13872 12316 13878 12328
rect 14369 12325 14381 12359
rect 14415 12356 14427 12359
rect 14826 12356 14832 12368
rect 14415 12328 14832 12356
rect 14415 12325 14427 12328
rect 14369 12319 14427 12325
rect 14826 12316 14832 12328
rect 14884 12316 14890 12368
rect 15470 12356 15476 12368
rect 15431 12328 15476 12356
rect 15470 12316 15476 12328
rect 15528 12316 15534 12368
rect 16022 12356 16028 12368
rect 15983 12328 16028 12356
rect 16022 12316 16028 12328
rect 16080 12316 16086 12368
rect 19058 12356 19064 12368
rect 19019 12328 19064 12356
rect 19058 12316 19064 12328
rect 19116 12316 19122 12368
rect 7101 12291 7159 12297
rect 7101 12257 7113 12291
rect 7147 12257 7159 12291
rect 7101 12251 7159 12257
rect 16758 12248 16764 12300
rect 16816 12288 16822 12300
rect 17129 12291 17187 12297
rect 17129 12288 17141 12291
rect 16816 12260 17141 12288
rect 16816 12248 16822 12260
rect 17129 12257 17141 12260
rect 17175 12288 17187 12291
rect 17770 12288 17776 12300
rect 17175 12260 17776 12288
rect 17175 12257 17187 12260
rect 17129 12251 17187 12257
rect 17770 12248 17776 12260
rect 17828 12248 17834 12300
rect 5350 12220 5356 12232
rect 3936 12192 5212 12220
rect 5311 12192 5356 12220
rect 3936 12180 3942 12192
rect 5350 12180 5356 12192
rect 5408 12180 5414 12232
rect 6178 12220 6184 12232
rect 6139 12192 6184 12220
rect 6178 12180 6184 12192
rect 6236 12180 6242 12232
rect 8021 12223 8079 12229
rect 8021 12189 8033 12223
rect 8067 12189 8079 12223
rect 8021 12183 8079 12189
rect 1854 12112 1860 12164
rect 1912 12152 1918 12164
rect 8036 12152 8064 12183
rect 8202 12180 8208 12232
rect 8260 12220 8266 12232
rect 8297 12223 8355 12229
rect 8297 12220 8309 12223
rect 8260 12192 8309 12220
rect 8260 12180 8266 12192
rect 8297 12189 8309 12192
rect 8343 12189 8355 12223
rect 9766 12220 9772 12232
rect 9727 12192 9772 12220
rect 8297 12183 8355 12189
rect 9766 12180 9772 12192
rect 9824 12180 9830 12232
rect 11333 12223 11391 12229
rect 11333 12189 11345 12223
rect 11379 12189 11391 12223
rect 11333 12183 11391 12189
rect 8662 12152 8668 12164
rect 1912 12124 8668 12152
rect 1912 12112 1918 12124
rect 8662 12112 8668 12124
rect 8720 12112 8726 12164
rect 11238 12112 11244 12164
rect 11296 12152 11302 12164
rect 11348 12152 11376 12183
rect 11514 12180 11520 12232
rect 11572 12220 11578 12232
rect 11609 12223 11667 12229
rect 11609 12220 11621 12223
rect 11572 12192 11621 12220
rect 11572 12180 11578 12192
rect 11609 12189 11621 12192
rect 11655 12189 11667 12223
rect 11609 12183 11667 12189
rect 13725 12223 13783 12229
rect 13725 12189 13737 12223
rect 13771 12220 13783 12223
rect 14182 12220 14188 12232
rect 13771 12192 14188 12220
rect 13771 12189 13783 12192
rect 13725 12183 13783 12189
rect 14182 12180 14188 12192
rect 14240 12180 14246 12232
rect 15381 12223 15439 12229
rect 15381 12220 15393 12223
rect 15028 12192 15393 12220
rect 11296 12124 11376 12152
rect 11296 12112 11302 12124
rect 2087 12087 2145 12093
rect 2087 12053 2099 12087
rect 2133 12084 2145 12087
rect 3142 12084 3148 12096
rect 2133 12056 3148 12084
rect 2133 12053 2145 12056
rect 2087 12047 2145 12053
rect 3142 12044 3148 12056
rect 3200 12044 3206 12096
rect 5534 12044 5540 12096
rect 5592 12084 5598 12096
rect 5721 12087 5779 12093
rect 5721 12084 5733 12087
rect 5592 12056 5733 12084
rect 5592 12044 5598 12056
rect 5721 12053 5733 12056
rect 5767 12084 5779 12087
rect 7190 12084 7196 12096
rect 5767 12056 7196 12084
rect 5767 12053 5779 12056
rect 5721 12047 5779 12053
rect 7190 12044 7196 12056
rect 7248 12044 7254 12096
rect 7466 12044 7472 12096
rect 7524 12084 7530 12096
rect 9122 12084 9128 12096
rect 7524 12056 9128 12084
rect 7524 12044 7530 12056
rect 9122 12044 9128 12056
rect 9180 12044 9186 12096
rect 9858 12044 9864 12096
rect 9916 12084 9922 12096
rect 11054 12084 11060 12096
rect 9916 12056 11060 12084
rect 9916 12044 9922 12056
rect 11054 12044 11060 12056
rect 11112 12044 11118 12096
rect 12710 12084 12716 12096
rect 12671 12056 12716 12084
rect 12710 12044 12716 12056
rect 12768 12044 12774 12096
rect 12802 12044 12808 12096
rect 12860 12084 12866 12096
rect 15028 12093 15056 12192
rect 15381 12189 15393 12192
rect 15427 12189 15439 12223
rect 15381 12183 15439 12189
rect 16482 12180 16488 12232
rect 16540 12220 16546 12232
rect 18966 12220 18972 12232
rect 16540 12192 18972 12220
rect 16540 12180 16546 12192
rect 18966 12180 18972 12192
rect 19024 12180 19030 12232
rect 19150 12180 19156 12232
rect 19208 12220 19214 12232
rect 19245 12223 19303 12229
rect 19245 12220 19257 12223
rect 19208 12192 19257 12220
rect 19208 12180 19214 12192
rect 19245 12189 19257 12192
rect 19291 12189 19303 12223
rect 19245 12183 19303 12189
rect 18049 12155 18107 12161
rect 18049 12121 18061 12155
rect 18095 12152 18107 12155
rect 18782 12152 18788 12164
rect 18095 12124 18788 12152
rect 18095 12121 18107 12124
rect 18049 12115 18107 12121
rect 18782 12112 18788 12124
rect 18840 12112 18846 12164
rect 15013 12087 15071 12093
rect 15013 12084 15025 12087
rect 12860 12056 15025 12084
rect 12860 12044 12866 12056
rect 15013 12053 15025 12056
rect 15059 12053 15071 12087
rect 15013 12047 15071 12053
rect 16022 12044 16028 12096
rect 16080 12084 16086 12096
rect 16301 12087 16359 12093
rect 16301 12084 16313 12087
rect 16080 12056 16313 12084
rect 16080 12044 16086 12056
rect 16301 12053 16313 12056
rect 16347 12053 16359 12087
rect 16301 12047 16359 12053
rect 1104 11994 20884 12016
rect 1104 11942 4648 11994
rect 4700 11942 4712 11994
rect 4764 11942 4776 11994
rect 4828 11942 4840 11994
rect 4892 11942 11982 11994
rect 12034 11942 12046 11994
rect 12098 11942 12110 11994
rect 12162 11942 12174 11994
rect 12226 11942 19315 11994
rect 19367 11942 19379 11994
rect 19431 11942 19443 11994
rect 19495 11942 19507 11994
rect 19559 11942 20884 11994
rect 1104 11920 20884 11942
rect 2774 11840 2780 11892
rect 2832 11880 2838 11892
rect 3053 11883 3111 11889
rect 3053 11880 3065 11883
rect 2832 11852 3065 11880
rect 2832 11840 2838 11852
rect 3053 11849 3065 11852
rect 3099 11849 3111 11883
rect 3053 11843 3111 11849
rect 4709 11883 4767 11889
rect 4709 11849 4721 11883
rect 4755 11880 4767 11883
rect 5534 11880 5540 11892
rect 4755 11852 5540 11880
rect 4755 11849 4767 11852
rect 4709 11843 4767 11849
rect 5534 11840 5540 11852
rect 5592 11840 5598 11892
rect 8018 11880 8024 11892
rect 5803 11852 8024 11880
rect 2869 11815 2927 11821
rect 2869 11781 2881 11815
rect 2915 11812 2927 11815
rect 5803 11812 5831 11852
rect 8018 11840 8024 11852
rect 8076 11840 8082 11892
rect 8113 11883 8171 11889
rect 8113 11849 8125 11883
rect 8159 11880 8171 11883
rect 9030 11880 9036 11892
rect 8159 11852 9036 11880
rect 8159 11849 8171 11852
rect 8113 11843 8171 11849
rect 9030 11840 9036 11852
rect 9088 11840 9094 11892
rect 9766 11840 9772 11892
rect 9824 11880 9830 11892
rect 10689 11883 10747 11889
rect 10689 11880 10701 11883
rect 9824 11852 10701 11880
rect 9824 11840 9830 11852
rect 10689 11849 10701 11852
rect 10735 11849 10747 11883
rect 10689 11843 10747 11849
rect 13814 11840 13820 11892
rect 13872 11880 13878 11892
rect 14185 11883 14243 11889
rect 14185 11880 14197 11883
rect 13872 11852 14197 11880
rect 13872 11840 13878 11852
rect 14185 11849 14197 11852
rect 14231 11880 14243 11883
rect 15470 11880 15476 11892
rect 14231 11852 15476 11880
rect 14231 11849 14243 11852
rect 14185 11843 14243 11849
rect 15470 11840 15476 11852
rect 15528 11880 15534 11892
rect 15841 11883 15899 11889
rect 15841 11880 15853 11883
rect 15528 11852 15853 11880
rect 15528 11840 15534 11852
rect 15841 11849 15853 11852
rect 15887 11849 15899 11883
rect 17770 11880 17776 11892
rect 17731 11852 17776 11880
rect 15841 11843 15899 11849
rect 17770 11840 17776 11852
rect 17828 11840 17834 11892
rect 19058 11840 19064 11892
rect 19116 11880 19122 11892
rect 19613 11883 19671 11889
rect 19613 11880 19625 11883
rect 19116 11852 19625 11880
rect 19116 11840 19122 11852
rect 19613 11849 19625 11852
rect 19659 11849 19671 11883
rect 19613 11843 19671 11849
rect 2915 11784 5831 11812
rect 5997 11815 6055 11821
rect 2915 11781 2927 11784
rect 2869 11775 2927 11781
rect 5997 11781 6009 11815
rect 6043 11812 6055 11815
rect 11701 11815 11759 11821
rect 11701 11812 11713 11815
rect 6043 11784 11713 11812
rect 6043 11781 6055 11784
rect 5997 11775 6055 11781
rect 11701 11781 11713 11784
rect 11747 11781 11759 11815
rect 11701 11775 11759 11781
rect 11790 11772 11796 11824
rect 11848 11812 11854 11824
rect 13909 11815 13967 11821
rect 13909 11812 13921 11815
rect 11848 11784 13921 11812
rect 11848 11772 11854 11784
rect 13909 11781 13921 11784
rect 13955 11781 13967 11815
rect 13909 11775 13967 11781
rect 13998 11772 14004 11824
rect 14056 11812 14062 11824
rect 18506 11812 18512 11824
rect 14056 11784 18512 11812
rect 14056 11772 14062 11784
rect 18506 11772 18512 11784
rect 18564 11772 18570 11824
rect 18966 11772 18972 11824
rect 19024 11812 19030 11824
rect 19981 11815 20039 11821
rect 19981 11812 19993 11815
rect 19024 11784 19993 11812
rect 19024 11772 19030 11784
rect 19981 11781 19993 11784
rect 20027 11781 20039 11815
rect 19981 11775 20039 11781
rect 5077 11747 5135 11753
rect 5077 11713 5089 11747
rect 5123 11744 5135 11747
rect 5123 11716 5304 11744
rect 5123 11713 5135 11716
rect 5077 11707 5135 11713
rect 1632 11679 1690 11685
rect 1632 11645 1644 11679
rect 1678 11676 1690 11679
rect 2660 11679 2718 11685
rect 1678 11648 2544 11676
rect 1678 11645 1690 11648
rect 1632 11639 1690 11645
rect 1719 11611 1777 11617
rect 1719 11577 1731 11611
rect 1765 11608 1777 11611
rect 1854 11608 1860 11620
rect 1765 11580 1860 11608
rect 1765 11577 1777 11580
rect 1719 11571 1777 11577
rect 1854 11568 1860 11580
rect 1912 11568 1918 11620
rect 2038 11540 2044 11552
rect 1999 11512 2044 11540
rect 2038 11500 2044 11512
rect 2096 11500 2102 11552
rect 2516 11549 2544 11648
rect 2660 11645 2672 11679
rect 2706 11676 2718 11679
rect 3421 11679 3479 11685
rect 3421 11676 3433 11679
rect 2706 11648 3433 11676
rect 2706 11645 2718 11648
rect 2660 11639 2718 11645
rect 3421 11645 3433 11648
rect 3467 11645 3479 11679
rect 3878 11676 3884 11688
rect 3839 11648 3884 11676
rect 3421 11639 3479 11645
rect 3436 11608 3464 11639
rect 3878 11636 3884 11648
rect 3936 11636 3942 11688
rect 4157 11679 4215 11685
rect 4157 11645 4169 11679
rect 4203 11676 4215 11679
rect 4982 11676 4988 11688
rect 4203 11648 4988 11676
rect 4203 11645 4215 11648
rect 4157 11639 4215 11645
rect 4982 11636 4988 11648
rect 5040 11636 5046 11688
rect 5166 11676 5172 11688
rect 5127 11648 5172 11676
rect 5166 11636 5172 11648
rect 5224 11636 5230 11688
rect 5276 11676 5304 11716
rect 5350 11704 5356 11756
rect 5408 11744 5414 11756
rect 6825 11747 6883 11753
rect 6825 11744 6837 11747
rect 5408 11716 6837 11744
rect 5408 11704 5414 11716
rect 6825 11713 6837 11716
rect 6871 11744 6883 11747
rect 7098 11744 7104 11756
rect 6871 11716 7104 11744
rect 6871 11713 6883 11716
rect 6825 11707 6883 11713
rect 7098 11704 7104 11716
rect 7156 11704 7162 11756
rect 8110 11704 8116 11756
rect 8168 11744 8174 11756
rect 11471 11747 11529 11753
rect 8168 11716 11411 11744
rect 8168 11704 8174 11716
rect 5718 11676 5724 11688
rect 5276 11648 5724 11676
rect 5718 11636 5724 11648
rect 5776 11636 5782 11688
rect 8573 11679 8631 11685
rect 8573 11676 8585 11679
rect 6885 11648 8585 11676
rect 4341 11611 4399 11617
rect 3436 11580 4154 11608
rect 2501 11543 2559 11549
rect 2501 11509 2513 11543
rect 2547 11540 2559 11543
rect 2590 11540 2596 11552
rect 2547 11512 2596 11540
rect 2547 11509 2559 11512
rect 2501 11503 2559 11509
rect 2590 11500 2596 11512
rect 2648 11500 2654 11552
rect 4126 11540 4154 11580
rect 4341 11577 4353 11611
rect 4387 11608 4399 11611
rect 6885 11608 6913 11648
rect 8573 11645 8585 11648
rect 8619 11676 8631 11679
rect 9493 11679 9551 11685
rect 9493 11676 9505 11679
rect 8619 11648 9505 11676
rect 8619 11645 8631 11648
rect 8573 11639 8631 11645
rect 9493 11645 9505 11648
rect 9539 11645 9551 11679
rect 9493 11639 9551 11645
rect 10413 11679 10471 11685
rect 10413 11645 10425 11679
rect 10459 11676 10471 11679
rect 10502 11676 10508 11688
rect 10459 11648 10508 11676
rect 10459 11645 10471 11648
rect 10413 11639 10471 11645
rect 10502 11636 10508 11648
rect 10560 11676 10566 11688
rect 10870 11676 10876 11688
rect 10560 11648 10876 11676
rect 10560 11636 10566 11648
rect 10870 11636 10876 11648
rect 10928 11636 10934 11688
rect 11383 11685 11411 11716
rect 11471 11713 11483 11747
rect 11517 11744 11529 11747
rect 14734 11744 14740 11756
rect 11517 11716 14740 11744
rect 11517 11713 11529 11716
rect 11471 11707 11529 11713
rect 14734 11704 14740 11716
rect 14792 11704 14798 11756
rect 14921 11747 14979 11753
rect 14921 11713 14933 11747
rect 14967 11744 14979 11747
rect 15194 11744 15200 11756
rect 14967 11716 15200 11744
rect 14967 11713 14979 11716
rect 14921 11707 14979 11713
rect 15194 11704 15200 11716
rect 15252 11704 15258 11756
rect 15565 11747 15623 11753
rect 15565 11713 15577 11747
rect 15611 11744 15623 11747
rect 16206 11744 16212 11756
rect 15611 11716 16212 11744
rect 15611 11713 15623 11716
rect 15565 11707 15623 11713
rect 16206 11704 16212 11716
rect 16264 11704 16270 11756
rect 16485 11747 16543 11753
rect 16485 11713 16497 11747
rect 16531 11744 16543 11747
rect 16850 11744 16856 11756
rect 16531 11716 16856 11744
rect 16531 11713 16543 11716
rect 16485 11707 16543 11713
rect 16850 11704 16856 11716
rect 16908 11704 16914 11756
rect 17129 11747 17187 11753
rect 17129 11713 17141 11747
rect 17175 11744 17187 11747
rect 18874 11744 18880 11756
rect 17175 11716 18880 11744
rect 17175 11713 17187 11716
rect 17129 11707 17187 11713
rect 18874 11704 18880 11716
rect 18932 11704 18938 11756
rect 19337 11747 19395 11753
rect 19337 11713 19349 11747
rect 19383 11744 19395 11747
rect 19610 11744 19616 11756
rect 19383 11716 19616 11744
rect 19383 11713 19395 11716
rect 19337 11707 19395 11713
rect 19610 11704 19616 11716
rect 19668 11704 19674 11756
rect 11368 11679 11426 11685
rect 11368 11645 11380 11679
rect 11414 11645 11426 11679
rect 11368 11639 11426 11645
rect 11701 11679 11759 11685
rect 11701 11645 11713 11679
rect 11747 11676 11759 11679
rect 12894 11676 12900 11688
rect 11747 11648 12900 11676
rect 11747 11645 11759 11648
rect 11701 11639 11759 11645
rect 4387 11580 6913 11608
rect 7187 11611 7245 11617
rect 4387 11577 4399 11580
rect 4341 11571 4399 11577
rect 7187 11577 7199 11611
rect 7233 11608 7245 11611
rect 9855 11611 9913 11617
rect 7233 11580 9444 11608
rect 7233 11577 7245 11580
rect 7187 11571 7245 11577
rect 6086 11540 6092 11552
rect 4126 11512 6092 11540
rect 6086 11500 6092 11512
rect 6144 11500 6150 11552
rect 6273 11543 6331 11549
rect 6273 11509 6285 11543
rect 6319 11540 6331 11543
rect 6454 11540 6460 11552
rect 6319 11512 6460 11540
rect 6319 11509 6331 11512
rect 6273 11503 6331 11509
rect 6454 11500 6460 11512
rect 6512 11540 6518 11552
rect 6641 11543 6699 11549
rect 6641 11540 6653 11543
rect 6512 11512 6653 11540
rect 6512 11500 6518 11512
rect 6641 11509 6653 11512
rect 6687 11540 6699 11543
rect 7202 11540 7230 11571
rect 6687 11512 7230 11540
rect 6687 11509 6699 11512
rect 6641 11503 6699 11509
rect 7466 11500 7472 11552
rect 7524 11540 7530 11552
rect 9416 11549 9444 11580
rect 9855 11577 9867 11611
rect 9901 11577 9913 11611
rect 11383 11608 11411 11639
rect 12894 11636 12900 11648
rect 12952 11636 12958 11688
rect 13909 11679 13967 11685
rect 13909 11645 13921 11679
rect 13955 11676 13967 11679
rect 14458 11676 14464 11688
rect 13955 11648 14464 11676
rect 13955 11645 13967 11648
rect 13909 11639 13967 11645
rect 14458 11636 14464 11648
rect 14516 11636 14522 11688
rect 11790 11608 11796 11620
rect 11383 11580 11796 11608
rect 9855 11571 9913 11577
rect 7745 11543 7803 11549
rect 7745 11540 7757 11543
rect 7524 11512 7757 11540
rect 7524 11500 7530 11512
rect 7745 11509 7757 11512
rect 7791 11509 7803 11543
rect 7745 11503 7803 11509
rect 9401 11543 9459 11549
rect 9401 11509 9413 11543
rect 9447 11540 9459 11543
rect 9876 11540 9904 11571
rect 11790 11568 11796 11580
rect 11848 11568 11854 11620
rect 13259 11611 13317 11617
rect 13259 11577 13271 11611
rect 13305 11608 13317 11611
rect 14550 11608 14556 11620
rect 13305 11580 14556 11608
rect 13305 11577 13317 11580
rect 13259 11571 13317 11577
rect 10410 11540 10416 11552
rect 9447 11512 10416 11540
rect 9447 11509 9459 11512
rect 9401 11503 9459 11509
rect 10410 11500 10416 11512
rect 10468 11500 10474 11552
rect 11241 11543 11299 11549
rect 11241 11509 11253 11543
rect 11287 11540 11299 11543
rect 11606 11540 11612 11552
rect 11287 11512 11612 11540
rect 11287 11509 11299 11512
rect 11241 11503 11299 11509
rect 11606 11500 11612 11512
rect 11664 11500 11670 11552
rect 12710 11500 12716 11552
rect 12768 11540 12774 11552
rect 12805 11543 12863 11549
rect 12805 11540 12817 11543
rect 12768 11512 12817 11540
rect 12768 11500 12774 11512
rect 12805 11509 12817 11512
rect 12851 11540 12863 11543
rect 13274 11540 13302 11571
rect 14550 11568 14556 11580
rect 14608 11568 14614 11620
rect 14737 11611 14795 11617
rect 14737 11577 14749 11611
rect 14783 11608 14795 11611
rect 15013 11611 15071 11617
rect 15013 11608 15025 11611
rect 14783 11580 15025 11608
rect 14783 11577 14795 11580
rect 14737 11571 14795 11577
rect 15013 11577 15025 11580
rect 15059 11577 15071 11611
rect 15013 11571 15071 11577
rect 16301 11611 16359 11617
rect 16301 11577 16313 11611
rect 16347 11608 16359 11611
rect 16574 11608 16580 11620
rect 16347 11580 16580 11608
rect 16347 11577 16359 11580
rect 16301 11571 16359 11577
rect 13354 11540 13360 11552
rect 12851 11512 13360 11540
rect 12851 11509 12863 11512
rect 12805 11503 12863 11509
rect 13354 11500 13360 11512
rect 13412 11500 13418 11552
rect 15028 11540 15056 11571
rect 16316 11540 16344 11571
rect 16574 11568 16580 11580
rect 16632 11568 16638 11620
rect 18509 11611 18567 11617
rect 18509 11577 18521 11611
rect 18555 11608 18567 11611
rect 18690 11608 18696 11620
rect 18555 11580 18696 11608
rect 18555 11577 18567 11580
rect 18509 11571 18567 11577
rect 18690 11568 18696 11580
rect 18748 11568 18754 11620
rect 18782 11568 18788 11620
rect 18840 11608 18846 11620
rect 18840 11580 18885 11608
rect 18840 11568 18846 11580
rect 17402 11540 17408 11552
rect 15028 11512 16344 11540
rect 17363 11512 17408 11540
rect 17402 11500 17408 11512
rect 17460 11500 17466 11552
rect 1104 11450 20884 11472
rect 1104 11398 8315 11450
rect 8367 11398 8379 11450
rect 8431 11398 8443 11450
rect 8495 11398 8507 11450
rect 8559 11398 15648 11450
rect 15700 11398 15712 11450
rect 15764 11398 15776 11450
rect 15828 11398 15840 11450
rect 15892 11398 20884 11450
rect 1104 11376 20884 11398
rect 1578 11336 1584 11348
rect 1539 11308 1584 11336
rect 1578 11296 1584 11308
rect 1636 11296 1642 11348
rect 5166 11336 5172 11348
rect 5127 11308 5172 11336
rect 5166 11296 5172 11308
rect 5224 11336 5230 11348
rect 5350 11336 5356 11348
rect 5224 11308 5356 11336
rect 5224 11296 5230 11308
rect 5350 11296 5356 11308
rect 5408 11336 5414 11348
rect 5537 11339 5595 11345
rect 5537 11336 5549 11339
rect 5408 11308 5549 11336
rect 5408 11296 5414 11308
rect 5537 11305 5549 11308
rect 5583 11305 5595 11339
rect 5537 11299 5595 11305
rect 6178 11296 6184 11348
rect 6236 11336 6242 11348
rect 6733 11339 6791 11345
rect 6733 11336 6745 11339
rect 6236 11308 6745 11336
rect 6236 11296 6242 11308
rect 6733 11305 6745 11308
rect 6779 11305 6791 11339
rect 7098 11336 7104 11348
rect 7059 11308 7104 11336
rect 6733 11299 6791 11305
rect 7098 11296 7104 11308
rect 7156 11296 7162 11348
rect 10689 11339 10747 11345
rect 7253 11308 9812 11336
rect 4430 11268 4436 11280
rect 4172 11240 4436 11268
rect 1397 11203 1455 11209
rect 1397 11169 1409 11203
rect 1443 11200 1455 11203
rect 2222 11200 2228 11212
rect 1443 11172 2228 11200
rect 1443 11169 1455 11172
rect 1397 11163 1455 11169
rect 2222 11160 2228 11172
rect 2280 11160 2286 11212
rect 2590 11160 2596 11212
rect 2648 11200 2654 11212
rect 3028 11203 3086 11209
rect 3028 11200 3040 11203
rect 2648 11172 3040 11200
rect 2648 11160 2654 11172
rect 3028 11169 3040 11172
rect 3074 11200 3086 11203
rect 3418 11200 3424 11212
rect 3074 11172 3424 11200
rect 3074 11169 3086 11172
rect 3028 11163 3086 11169
rect 3418 11160 3424 11172
rect 3476 11160 3482 11212
rect 4172 11209 4200 11240
rect 4430 11228 4436 11240
rect 4488 11228 4494 11280
rect 4893 11271 4951 11277
rect 4893 11237 4905 11271
rect 4939 11268 4951 11271
rect 7253 11268 7281 11308
rect 7466 11268 7472 11280
rect 4939 11240 7281 11268
rect 7427 11240 7472 11268
rect 4939 11237 4951 11240
rect 4893 11231 4951 11237
rect 7466 11228 7472 11240
rect 7524 11228 7530 11280
rect 8021 11271 8079 11277
rect 8021 11237 8033 11271
rect 8067 11268 8079 11271
rect 8202 11268 8208 11280
rect 8067 11240 8208 11268
rect 8067 11237 8079 11240
rect 8021 11231 8079 11237
rect 8202 11228 8208 11240
rect 8260 11228 8266 11280
rect 8662 11268 8668 11280
rect 8623 11240 8668 11268
rect 8662 11228 8668 11240
rect 8720 11228 8726 11280
rect 4157 11203 4215 11209
rect 4157 11169 4169 11203
rect 4203 11169 4215 11203
rect 4709 11203 4767 11209
rect 4709 11200 4721 11203
rect 4157 11163 4215 11169
rect 4264 11172 4721 11200
rect 3697 11135 3755 11141
rect 3697 11101 3709 11135
rect 3743 11132 3755 11135
rect 4264 11132 4292 11172
rect 4709 11169 4721 11172
rect 4755 11200 4767 11203
rect 5074 11200 5080 11212
rect 4755 11172 5080 11200
rect 4755 11169 4767 11172
rect 4709 11163 4767 11169
rect 5074 11160 5080 11172
rect 5132 11160 5138 11212
rect 5442 11160 5448 11212
rect 5500 11200 5506 11212
rect 5721 11203 5779 11209
rect 5721 11200 5733 11203
rect 5500 11172 5733 11200
rect 5500 11160 5506 11172
rect 5721 11169 5733 11172
rect 5767 11169 5779 11203
rect 6178 11200 6184 11212
rect 6139 11172 6184 11200
rect 5721 11163 5779 11169
rect 6178 11160 6184 11172
rect 6236 11160 6242 11212
rect 9784 11209 9812 11308
rect 10689 11305 10701 11339
rect 10735 11305 10747 11339
rect 11238 11336 11244 11348
rect 11199 11308 11244 11336
rect 10689 11299 10747 11305
rect 10131 11271 10189 11277
rect 10131 11237 10143 11271
rect 10177 11268 10189 11271
rect 10410 11268 10416 11280
rect 10177 11240 10416 11268
rect 10177 11237 10189 11240
rect 10131 11231 10189 11237
rect 10410 11228 10416 11240
rect 10468 11228 10474 11280
rect 10704 11268 10732 11299
rect 11238 11296 11244 11308
rect 11296 11296 11302 11348
rect 12894 11336 12900 11348
rect 12855 11308 12900 11336
rect 12894 11296 12900 11308
rect 12952 11296 12958 11348
rect 14921 11339 14979 11345
rect 14921 11305 14933 11339
rect 14967 11336 14979 11339
rect 15194 11336 15200 11348
rect 14967 11308 15200 11336
rect 14967 11305 14979 11308
rect 14921 11299 14979 11305
rect 15194 11296 15200 11308
rect 15252 11296 15258 11348
rect 16850 11336 16856 11348
rect 16811 11308 16856 11336
rect 16850 11296 16856 11308
rect 16908 11296 16914 11348
rect 18693 11339 18751 11345
rect 18693 11305 18705 11339
rect 18739 11336 18751 11339
rect 18782 11336 18788 11348
rect 18739 11308 18788 11336
rect 18739 11305 18751 11308
rect 18693 11299 18751 11305
rect 18782 11296 18788 11308
rect 18840 11296 18846 11348
rect 11606 11268 11612 11280
rect 10704 11240 11612 11268
rect 11606 11228 11612 11240
rect 11664 11268 11670 11280
rect 11701 11271 11759 11277
rect 11701 11268 11713 11271
rect 11664 11240 11713 11268
rect 11664 11228 11670 11240
rect 11701 11237 11713 11240
rect 11747 11237 11759 11271
rect 11701 11231 11759 11237
rect 13449 11271 13507 11277
rect 13449 11237 13461 11271
rect 13495 11268 13507 11271
rect 13538 11268 13544 11280
rect 13495 11240 13544 11268
rect 13495 11237 13507 11240
rect 13449 11231 13507 11237
rect 13538 11228 13544 11240
rect 13596 11228 13602 11280
rect 14550 11228 14556 11280
rect 14608 11268 14614 11280
rect 15927 11271 15985 11277
rect 15927 11268 15939 11271
rect 14608 11240 15939 11268
rect 14608 11228 14614 11240
rect 15927 11237 15939 11240
rect 15973 11268 15985 11271
rect 16022 11268 16028 11280
rect 15973 11240 16028 11268
rect 15973 11237 15985 11240
rect 15927 11231 15985 11237
rect 16022 11228 16028 11240
rect 16080 11268 16086 11280
rect 17402 11268 17408 11280
rect 16080 11240 17408 11268
rect 16080 11228 16086 11240
rect 17402 11228 17408 11240
rect 17460 11268 17466 11280
rect 17634 11271 17692 11277
rect 17634 11268 17646 11271
rect 17460 11240 17646 11268
rect 17460 11228 17466 11240
rect 17634 11237 17646 11240
rect 17680 11237 17692 11271
rect 19245 11271 19303 11277
rect 19245 11268 19257 11271
rect 17634 11231 17692 11237
rect 18661 11240 19257 11268
rect 9769 11203 9827 11209
rect 9769 11169 9781 11203
rect 9815 11200 9827 11203
rect 9858 11200 9864 11212
rect 9815 11172 9864 11200
rect 9815 11169 9827 11172
rect 9769 11163 9827 11169
rect 9858 11160 9864 11172
rect 9916 11160 9922 11212
rect 15378 11160 15384 11212
rect 15436 11200 15442 11212
rect 15565 11203 15623 11209
rect 15565 11200 15577 11203
rect 15436 11172 15577 11200
rect 15436 11160 15442 11172
rect 15565 11169 15577 11172
rect 15611 11169 15623 11203
rect 15565 11163 15623 11169
rect 18233 11203 18291 11209
rect 18233 11169 18245 11203
rect 18279 11200 18291 11203
rect 18661 11200 18689 11240
rect 19245 11237 19257 11240
rect 19291 11268 19303 11271
rect 19610 11268 19616 11280
rect 19291 11240 19616 11268
rect 19291 11237 19303 11240
rect 19245 11231 19303 11237
rect 19610 11228 19616 11240
rect 19668 11228 19674 11280
rect 18279 11172 18689 11200
rect 18279 11169 18291 11172
rect 18233 11163 18291 11169
rect 3743 11104 4292 11132
rect 3743 11101 3755 11104
rect 3697 11095 3755 11101
rect 4522 11092 4528 11144
rect 4580 11132 4586 11144
rect 5460 11132 5488 11160
rect 6454 11132 6460 11144
rect 4580 11104 5488 11132
rect 6415 11104 6460 11132
rect 4580 11092 4586 11104
rect 6454 11092 6460 11104
rect 6512 11092 6518 11144
rect 7374 11132 7380 11144
rect 7335 11104 7380 11132
rect 7374 11092 7380 11104
rect 7432 11092 7438 11144
rect 8205 11135 8263 11141
rect 8205 11101 8217 11135
rect 8251 11132 8263 11135
rect 11422 11132 11428 11144
rect 8251 11104 11428 11132
rect 8251 11101 8263 11104
rect 8205 11095 8263 11101
rect 11422 11092 11428 11104
rect 11480 11132 11486 11144
rect 11609 11135 11667 11141
rect 11609 11132 11621 11135
rect 11480 11104 11621 11132
rect 11480 11092 11486 11104
rect 11609 11101 11621 11104
rect 11655 11101 11667 11135
rect 11882 11132 11888 11144
rect 11843 11104 11888 11132
rect 11609 11095 11667 11101
rect 11882 11092 11888 11104
rect 11940 11092 11946 11144
rect 12434 11092 12440 11144
rect 12492 11132 12498 11144
rect 13357 11135 13415 11141
rect 13357 11132 13369 11135
rect 12492 11104 13369 11132
rect 12492 11092 12498 11104
rect 13357 11101 13369 11104
rect 13403 11101 13415 11135
rect 13998 11132 14004 11144
rect 13959 11104 14004 11132
rect 13357 11095 13415 11101
rect 13998 11092 14004 11104
rect 14056 11092 14062 11144
rect 14734 11092 14740 11144
rect 14792 11132 14798 11144
rect 16482 11132 16488 11144
rect 14792 11104 16488 11132
rect 14792 11092 14798 11104
rect 16482 11092 16488 11104
rect 16540 11132 16546 11144
rect 17129 11135 17187 11141
rect 17129 11132 17141 11135
rect 16540 11104 17141 11132
rect 16540 11092 16546 11104
rect 17129 11101 17141 11104
rect 17175 11101 17187 11135
rect 17129 11095 17187 11101
rect 17313 11135 17371 11141
rect 17313 11101 17325 11135
rect 17359 11132 17371 11135
rect 17678 11132 17684 11144
rect 17359 11104 17684 11132
rect 17359 11101 17371 11104
rect 17313 11095 17371 11101
rect 17678 11092 17684 11104
rect 17736 11092 17742 11144
rect 18782 11092 18788 11144
rect 18840 11132 18846 11144
rect 19150 11132 19156 11144
rect 18840 11104 19156 11132
rect 18840 11092 18846 11104
rect 19150 11092 19156 11104
rect 19208 11092 19214 11144
rect 19518 11132 19524 11144
rect 19479 11104 19524 11132
rect 19518 11092 19524 11104
rect 19576 11092 19582 11144
rect 3099 11067 3157 11073
rect 3099 11033 3111 11067
rect 3145 11064 3157 11067
rect 3145 11036 5764 11064
rect 3145 11033 3157 11036
rect 3099 11027 3157 11033
rect 5736 10996 5764 11036
rect 5810 11024 5816 11076
rect 5868 11064 5874 11076
rect 12526 11064 12532 11076
rect 5868 11036 12532 11064
rect 5868 11024 5874 11036
rect 12526 11024 12532 11036
rect 12584 11024 12590 11076
rect 19536 11064 19564 11092
rect 19702 11064 19708 11076
rect 19536 11036 19708 11064
rect 19702 11024 19708 11036
rect 19760 11024 19766 11076
rect 8205 10999 8263 11005
rect 8205 10996 8217 10999
rect 5736 10968 8217 10996
rect 8205 10965 8217 10968
rect 8251 10965 8263 10999
rect 8386 10996 8392 11008
rect 8347 10968 8392 10996
rect 8205 10959 8263 10965
rect 8386 10956 8392 10968
rect 8444 10956 8450 11008
rect 14274 10996 14280 11008
rect 14235 10968 14280 10996
rect 14274 10956 14280 10968
rect 14332 10956 14338 11008
rect 16298 10956 16304 11008
rect 16356 10996 16362 11008
rect 16485 10999 16543 11005
rect 16485 10996 16497 10999
rect 16356 10968 16497 10996
rect 16356 10956 16362 10968
rect 16485 10965 16497 10968
rect 16531 10996 16543 10999
rect 19058 10996 19064 11008
rect 16531 10968 19064 10996
rect 16531 10965 16543 10968
rect 16485 10959 16543 10965
rect 19058 10956 19064 10968
rect 19116 10956 19122 11008
rect 1104 10906 20884 10928
rect 1104 10854 4648 10906
rect 4700 10854 4712 10906
rect 4764 10854 4776 10906
rect 4828 10854 4840 10906
rect 4892 10854 11982 10906
rect 12034 10854 12046 10906
rect 12098 10854 12110 10906
rect 12162 10854 12174 10906
rect 12226 10854 19315 10906
rect 19367 10854 19379 10906
rect 19431 10854 19443 10906
rect 19495 10854 19507 10906
rect 19559 10854 20884 10906
rect 1104 10832 20884 10854
rect 2133 10795 2191 10801
rect 2133 10761 2145 10795
rect 2179 10792 2191 10795
rect 2222 10792 2228 10804
rect 2179 10764 2228 10792
rect 2179 10761 2191 10764
rect 2133 10755 2191 10761
rect 1670 10597 1676 10600
rect 1648 10591 1676 10597
rect 1648 10588 1660 10591
rect 1583 10560 1660 10588
rect 1648 10557 1660 10560
rect 1728 10588 1734 10600
rect 2148 10588 2176 10755
rect 2222 10752 2228 10764
rect 2280 10752 2286 10804
rect 3050 10752 3056 10804
rect 3108 10792 3114 10804
rect 4154 10792 4160 10804
rect 3108 10764 4160 10792
rect 3108 10752 3114 10764
rect 4154 10752 4160 10764
rect 4212 10752 4218 10804
rect 4709 10795 4767 10801
rect 4709 10761 4721 10795
rect 4755 10792 4767 10795
rect 5074 10792 5080 10804
rect 4755 10764 5080 10792
rect 4755 10761 4767 10764
rect 4709 10755 4767 10761
rect 5074 10752 5080 10764
rect 5132 10752 5138 10804
rect 5442 10752 5448 10804
rect 5500 10792 5506 10804
rect 6549 10795 6607 10801
rect 6549 10792 6561 10795
rect 5500 10764 6561 10792
rect 5500 10752 5506 10764
rect 6549 10761 6561 10764
rect 6595 10761 6607 10795
rect 8386 10792 8392 10804
rect 6549 10755 6607 10761
rect 7852 10764 8392 10792
rect 2501 10727 2559 10733
rect 2501 10693 2513 10727
rect 2547 10724 2559 10727
rect 3878 10724 3884 10736
rect 2547 10696 3884 10724
rect 2547 10693 2559 10696
rect 2501 10687 2559 10693
rect 3878 10684 3884 10696
rect 3936 10684 3942 10736
rect 7852 10665 7880 10764
rect 8386 10752 8392 10764
rect 8444 10792 8450 10804
rect 9447 10795 9505 10801
rect 9447 10792 9459 10795
rect 8444 10764 9459 10792
rect 8444 10752 8450 10764
rect 9447 10761 9459 10764
rect 9493 10761 9505 10795
rect 11606 10792 11612 10804
rect 11567 10764 11612 10792
rect 9447 10755 9505 10761
rect 11606 10752 11612 10764
rect 11664 10752 11670 10804
rect 16298 10792 16304 10804
rect 16259 10764 16304 10792
rect 16298 10752 16304 10764
rect 16356 10752 16362 10804
rect 19610 10792 19616 10804
rect 19571 10764 19616 10792
rect 19610 10752 19616 10764
rect 19668 10752 19674 10804
rect 9140 10696 10640 10724
rect 7837 10659 7895 10665
rect 7837 10625 7849 10659
rect 7883 10625 7895 10659
rect 7837 10619 7895 10625
rect 8481 10659 8539 10665
rect 8481 10625 8493 10659
rect 8527 10656 8539 10659
rect 8846 10656 8852 10668
rect 8527 10628 8852 10656
rect 8527 10625 8539 10628
rect 8481 10619 8539 10625
rect 8846 10616 8852 10628
rect 8904 10616 8910 10668
rect 1728 10560 2176 10588
rect 2660 10591 2718 10597
rect 1648 10551 1676 10557
rect 1670 10548 1676 10551
rect 1728 10548 1734 10560
rect 2660 10557 2672 10591
rect 2706 10588 2718 10591
rect 3878 10588 3884 10600
rect 2706 10560 3096 10588
rect 3839 10560 3884 10588
rect 2706 10557 2718 10560
rect 2660 10551 2718 10557
rect 3068 10464 3096 10560
rect 3878 10548 3884 10560
rect 3936 10548 3942 10600
rect 4062 10588 4068 10600
rect 4023 10560 4068 10588
rect 4062 10548 4068 10560
rect 4120 10548 4126 10600
rect 4430 10548 4436 10600
rect 4488 10588 4494 10600
rect 5442 10588 5448 10600
rect 4488 10560 5448 10588
rect 4488 10548 4494 10560
rect 5442 10548 5448 10560
rect 5500 10588 5506 10600
rect 5626 10588 5632 10600
rect 5500 10560 5632 10588
rect 5500 10548 5506 10560
rect 5626 10548 5632 10560
rect 5684 10548 5690 10600
rect 5721 10591 5779 10597
rect 5721 10557 5733 10591
rect 5767 10557 5779 10591
rect 5721 10551 5779 10557
rect 5905 10591 5963 10597
rect 5905 10557 5917 10591
rect 5951 10588 5963 10591
rect 7558 10588 7564 10600
rect 5951 10560 7564 10588
rect 5951 10557 5963 10560
rect 5905 10551 5963 10557
rect 1719 10455 1777 10461
rect 1719 10421 1731 10455
rect 1765 10452 1777 10455
rect 1946 10452 1952 10464
rect 1765 10424 1952 10452
rect 1765 10421 1777 10424
rect 1719 10415 1777 10421
rect 1946 10412 1952 10424
rect 2004 10412 2010 10464
rect 2731 10455 2789 10461
rect 2731 10421 2743 10455
rect 2777 10452 2789 10455
rect 2958 10452 2964 10464
rect 2777 10424 2964 10452
rect 2777 10421 2789 10424
rect 2731 10415 2789 10421
rect 2958 10412 2964 10424
rect 3016 10412 3022 10464
rect 3050 10412 3056 10464
rect 3108 10452 3114 10464
rect 3418 10452 3424 10464
rect 3108 10424 3153 10452
rect 3379 10424 3424 10452
rect 3108 10412 3114 10424
rect 3418 10412 3424 10424
rect 3476 10412 3482 10464
rect 3881 10455 3939 10461
rect 3881 10421 3893 10455
rect 3927 10452 3939 10455
rect 3970 10452 3976 10464
rect 3927 10424 3976 10452
rect 3927 10421 3939 10424
rect 3881 10415 3939 10421
rect 3970 10412 3976 10424
rect 4028 10412 4034 10464
rect 5077 10455 5135 10461
rect 5077 10421 5089 10455
rect 5123 10452 5135 10455
rect 5626 10452 5632 10464
rect 5123 10424 5632 10452
rect 5123 10421 5135 10424
rect 5077 10415 5135 10421
rect 5626 10412 5632 10424
rect 5684 10452 5690 10464
rect 5736 10452 5764 10551
rect 7558 10548 7564 10560
rect 7616 10548 7622 10600
rect 7377 10523 7435 10529
rect 7377 10489 7389 10523
rect 7423 10520 7435 10523
rect 7466 10520 7472 10532
rect 7423 10492 7472 10520
rect 7423 10489 7435 10492
rect 7377 10483 7435 10489
rect 7466 10480 7472 10492
rect 7524 10520 7530 10532
rect 7929 10523 7987 10529
rect 7929 10520 7941 10523
rect 7524 10492 7941 10520
rect 7524 10480 7530 10492
rect 7929 10489 7941 10492
rect 7975 10489 7987 10523
rect 7929 10483 7987 10489
rect 6178 10452 6184 10464
rect 5684 10424 6184 10452
rect 5684 10412 5690 10424
rect 6178 10412 6184 10424
rect 6236 10412 6242 10464
rect 7944 10452 7972 10483
rect 8018 10480 8024 10532
rect 8076 10520 8082 10532
rect 9140 10529 9168 10696
rect 10612 10665 10640 10696
rect 10597 10659 10655 10665
rect 10597 10625 10609 10659
rect 10643 10625 10655 10659
rect 10597 10619 10655 10625
rect 11241 10659 11299 10665
rect 11241 10625 11253 10659
rect 11287 10656 11299 10659
rect 11514 10656 11520 10668
rect 11287 10628 11520 10656
rect 11287 10625 11299 10628
rect 11241 10619 11299 10625
rect 11514 10616 11520 10628
rect 11572 10616 11578 10668
rect 12526 10616 12532 10668
rect 12584 10656 12590 10668
rect 12805 10659 12863 10665
rect 12805 10656 12817 10659
rect 12584 10628 12817 10656
rect 12584 10616 12590 10628
rect 12805 10625 12817 10628
rect 12851 10625 12863 10659
rect 12805 10619 12863 10625
rect 13998 10616 14004 10668
rect 14056 10656 14062 10668
rect 14369 10659 14427 10665
rect 14369 10656 14381 10659
rect 14056 10628 14381 10656
rect 14056 10616 14062 10628
rect 14369 10625 14381 10628
rect 14415 10625 14427 10659
rect 14642 10656 14648 10668
rect 14603 10628 14648 10656
rect 14369 10619 14427 10625
rect 14642 10616 14648 10628
rect 14700 10616 14706 10668
rect 16482 10656 16488 10668
rect 16443 10628 16488 10656
rect 16482 10616 16488 10628
rect 16540 10616 16546 10668
rect 19245 10659 19303 10665
rect 19245 10625 19257 10659
rect 19291 10656 19303 10659
rect 19702 10656 19708 10668
rect 19291 10628 19708 10656
rect 19291 10625 19303 10628
rect 19245 10619 19303 10625
rect 19702 10616 19708 10628
rect 19760 10616 19766 10668
rect 9376 10591 9434 10597
rect 9376 10557 9388 10591
rect 9422 10588 9434 10591
rect 9766 10588 9772 10600
rect 9422 10560 9772 10588
rect 9422 10557 9434 10560
rect 9376 10551 9434 10557
rect 9766 10548 9772 10560
rect 9824 10548 9830 10600
rect 9125 10523 9183 10529
rect 9125 10520 9137 10523
rect 8076 10492 9137 10520
rect 8076 10480 8082 10492
rect 9125 10489 9137 10492
rect 9171 10489 9183 10523
rect 9784 10520 9812 10548
rect 10689 10523 10747 10529
rect 9784 10492 10640 10520
rect 9125 10483 9183 10489
rect 8757 10455 8815 10461
rect 8757 10452 8769 10455
rect 7944 10424 8769 10452
rect 8757 10421 8769 10424
rect 8803 10421 8815 10455
rect 8757 10415 8815 10421
rect 10229 10455 10287 10461
rect 10229 10421 10241 10455
rect 10275 10452 10287 10455
rect 10410 10452 10416 10464
rect 10275 10424 10416 10452
rect 10275 10421 10287 10424
rect 10229 10415 10287 10421
rect 10410 10412 10416 10424
rect 10468 10412 10474 10464
rect 10612 10452 10640 10492
rect 10689 10489 10701 10523
rect 10735 10520 10747 10523
rect 10870 10520 10876 10532
rect 10735 10492 10876 10520
rect 10735 10489 10747 10492
rect 10689 10483 10747 10489
rect 10870 10480 10876 10492
rect 10928 10480 10934 10532
rect 12897 10523 12955 10529
rect 12897 10489 12909 10523
rect 12943 10489 12955 10523
rect 13446 10520 13452 10532
rect 13407 10492 13452 10520
rect 12897 10483 12955 10489
rect 11514 10452 11520 10464
rect 10612 10424 11520 10452
rect 11514 10412 11520 10424
rect 11572 10412 11578 10464
rect 12253 10455 12311 10461
rect 12253 10421 12265 10455
rect 12299 10452 12311 10455
rect 12912 10452 12940 10483
rect 13446 10480 13452 10492
rect 13504 10480 13510 10532
rect 14458 10480 14464 10532
rect 14516 10520 14522 10532
rect 14516 10492 14561 10520
rect 14516 10480 14522 10492
rect 16298 10480 16304 10532
rect 16356 10520 16362 10532
rect 16577 10523 16635 10529
rect 16577 10520 16589 10523
rect 16356 10492 16589 10520
rect 16356 10480 16362 10492
rect 16577 10489 16589 10492
rect 16623 10489 16635 10523
rect 17126 10520 17132 10532
rect 17087 10492 17132 10520
rect 16577 10483 16635 10489
rect 17126 10480 17132 10492
rect 17184 10520 17190 10532
rect 18598 10520 18604 10532
rect 17184 10492 18604 10520
rect 17184 10480 17190 10492
rect 18598 10480 18604 10492
rect 18656 10480 18662 10532
rect 18693 10523 18751 10529
rect 18693 10489 18705 10523
rect 18739 10489 18751 10523
rect 18693 10483 18751 10489
rect 13538 10452 13544 10464
rect 12299 10424 13544 10452
rect 12299 10421 12311 10424
rect 12253 10415 12311 10421
rect 13538 10412 13544 10424
rect 13596 10452 13602 10464
rect 13725 10455 13783 10461
rect 13725 10452 13737 10455
rect 13596 10424 13737 10452
rect 13596 10412 13602 10424
rect 13725 10421 13737 10424
rect 13771 10421 13783 10455
rect 13725 10415 13783 10421
rect 14185 10455 14243 10461
rect 14185 10421 14197 10455
rect 14231 10452 14243 10455
rect 14476 10452 14504 10480
rect 14231 10424 14504 10452
rect 15657 10455 15715 10461
rect 14231 10421 14243 10424
rect 14185 10415 14243 10421
rect 15657 10421 15669 10455
rect 15703 10452 15715 10455
rect 16022 10452 16028 10464
rect 15703 10424 16028 10452
rect 15703 10421 15715 10424
rect 15657 10415 15715 10421
rect 16022 10412 16028 10424
rect 16080 10452 16086 10464
rect 16942 10452 16948 10464
rect 16080 10424 16948 10452
rect 16080 10412 16086 10424
rect 16942 10412 16948 10424
rect 17000 10452 17006 10464
rect 17405 10455 17463 10461
rect 17405 10452 17417 10455
rect 17000 10424 17417 10452
rect 17000 10412 17006 10424
rect 17405 10421 17417 10424
rect 17451 10421 17463 10455
rect 17405 10415 17463 10421
rect 17678 10412 17684 10464
rect 17736 10452 17742 10464
rect 17773 10455 17831 10461
rect 17773 10452 17785 10455
rect 17736 10424 17785 10452
rect 17736 10412 17742 10424
rect 17773 10421 17785 10424
rect 17819 10421 17831 10455
rect 18322 10452 18328 10464
rect 18283 10424 18328 10452
rect 17773 10415 17831 10421
rect 18322 10412 18328 10424
rect 18380 10452 18386 10464
rect 18708 10452 18736 10483
rect 18380 10424 18736 10452
rect 18380 10412 18386 10424
rect 18782 10412 18788 10464
rect 18840 10452 18846 10464
rect 19889 10455 19947 10461
rect 19889 10452 19901 10455
rect 18840 10424 19901 10452
rect 18840 10412 18846 10424
rect 19889 10421 19901 10424
rect 19935 10421 19947 10455
rect 19889 10415 19947 10421
rect 1104 10362 20884 10384
rect 1104 10310 8315 10362
rect 8367 10310 8379 10362
rect 8431 10310 8443 10362
rect 8495 10310 8507 10362
rect 8559 10310 15648 10362
rect 15700 10310 15712 10362
rect 15764 10310 15776 10362
rect 15828 10310 15840 10362
rect 15892 10310 20884 10362
rect 1104 10288 20884 10310
rect 1670 10248 1676 10260
rect 1631 10220 1676 10248
rect 1670 10208 1676 10220
rect 1728 10208 1734 10260
rect 5442 10248 5448 10260
rect 5403 10220 5448 10248
rect 5442 10208 5448 10220
rect 5500 10248 5506 10260
rect 5813 10251 5871 10257
rect 5813 10248 5825 10251
rect 5500 10220 5825 10248
rect 5500 10208 5506 10220
rect 5813 10217 5825 10220
rect 5859 10217 5871 10251
rect 7374 10248 7380 10260
rect 7335 10220 7380 10248
rect 5813 10211 5871 10217
rect 7374 10208 7380 10220
rect 7432 10208 7438 10260
rect 7558 10208 7564 10260
rect 7616 10248 7622 10260
rect 9582 10248 9588 10260
rect 7616 10220 9588 10248
rect 7616 10208 7622 10220
rect 9582 10208 9588 10220
rect 9640 10208 9646 10260
rect 9858 10248 9864 10260
rect 9819 10220 9864 10248
rect 9858 10208 9864 10220
rect 9916 10208 9922 10260
rect 10870 10248 10876 10260
rect 10831 10220 10876 10248
rect 10870 10208 10876 10220
rect 10928 10208 10934 10260
rect 12802 10248 12808 10260
rect 10980 10220 12808 10248
rect 1688 10112 1716 10208
rect 2087 10183 2145 10189
rect 2087 10149 2099 10183
rect 2133 10180 2145 10183
rect 5718 10180 5724 10192
rect 2133 10152 5724 10180
rect 2133 10149 2145 10152
rect 2087 10143 2145 10149
rect 5718 10140 5724 10152
rect 5776 10140 5782 10192
rect 6086 10180 6092 10192
rect 6047 10152 6092 10180
rect 6086 10140 6092 10152
rect 6144 10140 6150 10192
rect 7650 10180 7656 10192
rect 7611 10152 7656 10180
rect 7650 10140 7656 10152
rect 7708 10140 7714 10192
rect 10183 10183 10241 10189
rect 10183 10149 10195 10183
rect 10229 10180 10241 10183
rect 10980 10180 11008 10220
rect 12802 10208 12808 10220
rect 12860 10208 12866 10260
rect 13538 10248 13544 10260
rect 13499 10220 13544 10248
rect 13538 10208 13544 10220
rect 13596 10208 13602 10260
rect 13998 10208 14004 10260
rect 14056 10248 14062 10260
rect 14277 10251 14335 10257
rect 14277 10248 14289 10251
rect 14056 10220 14289 10248
rect 14056 10208 14062 10220
rect 14277 10217 14289 10220
rect 14323 10217 14335 10251
rect 14277 10211 14335 10217
rect 15378 10208 15384 10260
rect 15436 10248 15442 10260
rect 15841 10251 15899 10257
rect 15841 10248 15853 10251
rect 15436 10220 15853 10248
rect 15436 10208 15442 10220
rect 15841 10217 15853 10220
rect 15887 10217 15899 10251
rect 15841 10211 15899 10217
rect 17313 10251 17371 10257
rect 17313 10217 17325 10251
rect 17359 10248 17371 10251
rect 18322 10248 18328 10260
rect 17359 10220 18328 10248
rect 17359 10217 17371 10220
rect 17313 10211 17371 10217
rect 18322 10208 18328 10220
rect 18380 10208 18386 10260
rect 18598 10208 18604 10260
rect 18656 10248 18662 10260
rect 19337 10251 19395 10257
rect 19337 10248 19349 10251
rect 18656 10220 19349 10248
rect 18656 10208 18662 10220
rect 19337 10217 19349 10220
rect 19383 10217 19395 10251
rect 19337 10211 19395 10217
rect 11238 10180 11244 10192
rect 10229 10152 11008 10180
rect 11199 10152 11244 10180
rect 10229 10149 10241 10152
rect 10183 10143 10241 10149
rect 11238 10140 11244 10152
rect 11296 10140 11302 10192
rect 11422 10140 11428 10192
rect 11480 10180 11486 10192
rect 12069 10183 12127 10189
rect 12069 10180 12081 10183
rect 11480 10152 12081 10180
rect 11480 10140 11486 10152
rect 12069 10149 12081 10152
rect 12115 10149 12127 10183
rect 12069 10143 12127 10149
rect 12983 10183 13041 10189
rect 12983 10149 12995 10183
rect 13029 10180 13041 10183
rect 13354 10180 13360 10192
rect 13029 10152 13360 10180
rect 13029 10149 13041 10152
rect 12983 10143 13041 10149
rect 13354 10140 13360 10152
rect 13412 10140 13418 10192
rect 16755 10183 16813 10189
rect 16755 10149 16767 10183
rect 16801 10180 16813 10183
rect 16942 10180 16948 10192
rect 16801 10152 16948 10180
rect 16801 10149 16813 10152
rect 16755 10143 16813 10149
rect 16942 10140 16948 10152
rect 17000 10140 17006 10192
rect 17770 10140 17776 10192
rect 17828 10180 17834 10192
rect 18509 10183 18567 10189
rect 18509 10180 18521 10183
rect 17828 10152 18521 10180
rect 17828 10140 17834 10152
rect 18509 10149 18521 10152
rect 18555 10149 18567 10183
rect 18509 10143 18567 10149
rect 1984 10115 2042 10121
rect 1984 10112 1996 10115
rect 1688 10084 1996 10112
rect 1984 10081 1996 10084
rect 2030 10112 2042 10115
rect 2314 10112 2320 10124
rect 2030 10084 2320 10112
rect 2030 10081 2042 10084
rect 1984 10075 2042 10081
rect 2314 10072 2320 10084
rect 2372 10072 2378 10124
rect 2961 10115 3019 10121
rect 2961 10081 2973 10115
rect 3007 10112 3019 10115
rect 3050 10112 3056 10124
rect 3007 10084 3056 10112
rect 3007 10081 3019 10084
rect 2961 10075 3019 10081
rect 3050 10072 3056 10084
rect 3108 10072 3114 10124
rect 4522 10112 4528 10124
rect 4483 10084 4528 10112
rect 4522 10072 4528 10084
rect 4580 10072 4586 10124
rect 4801 10115 4859 10121
rect 4801 10112 4813 10115
rect 4632 10084 4813 10112
rect 3510 10004 3516 10056
rect 3568 10044 3574 10056
rect 4062 10044 4068 10056
rect 3568 10016 4068 10044
rect 3568 10004 3574 10016
rect 4062 10004 4068 10016
rect 4120 10044 4126 10056
rect 4632 10044 4660 10084
rect 4801 10081 4813 10084
rect 4847 10081 4859 10115
rect 4801 10075 4859 10081
rect 9950 10072 9956 10124
rect 10008 10112 10014 10124
rect 10080 10115 10138 10121
rect 10080 10112 10092 10115
rect 10008 10084 10092 10112
rect 10008 10072 10014 10084
rect 10080 10081 10092 10084
rect 10126 10081 10138 10115
rect 12434 10112 12440 10124
rect 12395 10084 12440 10112
rect 10080 10075 10138 10081
rect 12434 10072 12440 10084
rect 12492 10072 12498 10124
rect 12618 10112 12624 10124
rect 12579 10084 12624 10112
rect 12618 10072 12624 10084
rect 12676 10072 12682 10124
rect 15102 10072 15108 10124
rect 15160 10112 15166 10124
rect 15289 10115 15347 10121
rect 15289 10112 15301 10115
rect 15160 10084 15301 10112
rect 15160 10072 15166 10084
rect 15289 10081 15301 10084
rect 15335 10081 15347 10115
rect 15289 10075 15347 10081
rect 4120 10016 4660 10044
rect 5077 10047 5135 10053
rect 4120 10004 4126 10016
rect 5077 10013 5089 10047
rect 5123 10044 5135 10047
rect 5123 10016 5948 10044
rect 5123 10013 5135 10016
rect 5077 10007 5135 10013
rect 3099 9979 3157 9985
rect 3099 9945 3111 9979
rect 3145 9976 3157 9979
rect 5810 9976 5816 9988
rect 3145 9948 5816 9976
rect 3145 9945 3157 9948
rect 3099 9939 3157 9945
rect 5810 9936 5816 9948
rect 5868 9936 5874 9988
rect 3510 9868 3516 9920
rect 3568 9908 3574 9920
rect 3605 9911 3663 9917
rect 3605 9908 3617 9911
rect 3568 9880 3617 9908
rect 3568 9868 3574 9880
rect 3605 9877 3617 9880
rect 3651 9877 3663 9911
rect 5920 9908 5948 10016
rect 5994 10004 6000 10056
rect 6052 10044 6058 10056
rect 7558 10044 7564 10056
rect 6052 10016 6097 10044
rect 7519 10016 7564 10044
rect 6052 10004 6058 10016
rect 7558 10004 7564 10016
rect 7616 10004 7622 10056
rect 7837 10047 7895 10053
rect 7837 10013 7849 10047
rect 7883 10013 7895 10047
rect 11146 10044 11152 10056
rect 11107 10016 11152 10044
rect 7837 10007 7895 10013
rect 6549 9979 6607 9985
rect 6549 9945 6561 9979
rect 6595 9976 6607 9979
rect 7852 9976 7880 10007
rect 11146 10004 11152 10016
rect 11204 10004 11210 10056
rect 16298 10004 16304 10056
rect 16356 10044 16362 10056
rect 16393 10047 16451 10053
rect 16393 10044 16405 10047
rect 16356 10016 16405 10044
rect 16356 10004 16362 10016
rect 16393 10013 16405 10016
rect 16439 10013 16451 10047
rect 16393 10007 16451 10013
rect 18417 10047 18475 10053
rect 18417 10013 18429 10047
rect 18463 10013 18475 10047
rect 18782 10044 18788 10056
rect 18743 10016 18788 10044
rect 18417 10007 18475 10013
rect 8846 9976 8852 9988
rect 6595 9948 8852 9976
rect 6595 9945 6607 9948
rect 6549 9939 6607 9945
rect 8846 9936 8852 9948
rect 8904 9936 8910 9988
rect 9858 9936 9864 9988
rect 9916 9976 9922 9988
rect 10134 9976 10140 9988
rect 9916 9948 10140 9976
rect 9916 9936 9922 9948
rect 10134 9936 10140 9948
rect 10192 9936 10198 9988
rect 11701 9979 11759 9985
rect 11701 9945 11713 9979
rect 11747 9976 11759 9979
rect 13078 9976 13084 9988
rect 11747 9948 13084 9976
rect 11747 9945 11759 9948
rect 11701 9939 11759 9945
rect 13078 9936 13084 9948
rect 13136 9976 13142 9988
rect 13998 9976 14004 9988
rect 13136 9948 14004 9976
rect 13136 9936 13142 9948
rect 13998 9936 14004 9948
rect 14056 9936 14062 9988
rect 15473 9979 15531 9985
rect 15473 9945 15485 9979
rect 15519 9976 15531 9979
rect 15930 9976 15936 9988
rect 15519 9948 15936 9976
rect 15519 9945 15531 9948
rect 15473 9939 15531 9945
rect 15930 9936 15936 9948
rect 15988 9936 15994 9988
rect 18432 9976 18460 10007
rect 18782 10004 18788 10016
rect 18840 10004 18846 10056
rect 19610 9976 19616 9988
rect 18432 9948 19616 9976
rect 19610 9936 19616 9948
rect 19668 9936 19674 9988
rect 6822 9908 6828 9920
rect 5920 9880 6828 9908
rect 3605 9871 3663 9877
rect 6822 9868 6828 9880
rect 6880 9908 6886 9920
rect 6917 9911 6975 9917
rect 6917 9908 6929 9911
rect 6880 9880 6929 9908
rect 6880 9868 6886 9880
rect 6917 9877 6929 9880
rect 6963 9877 6975 9911
rect 8662 9908 8668 9920
rect 8623 9880 8668 9908
rect 6917 9871 6975 9877
rect 8662 9868 8668 9880
rect 8720 9868 8726 9920
rect 10410 9868 10416 9920
rect 10468 9908 10474 9920
rect 10597 9911 10655 9917
rect 10597 9908 10609 9911
rect 10468 9880 10609 9908
rect 10468 9868 10474 9880
rect 10597 9877 10609 9880
rect 10643 9908 10655 9911
rect 10686 9908 10692 9920
rect 10643 9880 10692 9908
rect 10643 9877 10655 9880
rect 10597 9871 10655 9877
rect 10686 9868 10692 9880
rect 10744 9868 10750 9920
rect 13722 9868 13728 9920
rect 13780 9908 13786 9920
rect 13817 9911 13875 9917
rect 13817 9908 13829 9911
rect 13780 9880 13829 9908
rect 13780 9868 13786 9880
rect 13817 9877 13829 9880
rect 13863 9877 13875 9911
rect 13817 9871 13875 9877
rect 16301 9911 16359 9917
rect 16301 9877 16313 9911
rect 16347 9908 16359 9911
rect 16482 9908 16488 9920
rect 16347 9880 16488 9908
rect 16347 9877 16359 9880
rect 16301 9871 16359 9877
rect 16482 9868 16488 9880
rect 16540 9868 16546 9920
rect 1104 9818 20884 9840
rect 1104 9766 4648 9818
rect 4700 9766 4712 9818
rect 4764 9766 4776 9818
rect 4828 9766 4840 9818
rect 4892 9766 11982 9818
rect 12034 9766 12046 9818
rect 12098 9766 12110 9818
rect 12162 9766 12174 9818
rect 12226 9766 19315 9818
rect 19367 9766 19379 9818
rect 19431 9766 19443 9818
rect 19495 9766 19507 9818
rect 19559 9766 20884 9818
rect 1104 9744 20884 9766
rect 2314 9704 2320 9716
rect 2275 9676 2320 9704
rect 2314 9664 2320 9676
rect 2372 9664 2378 9716
rect 4246 9664 4252 9716
rect 4304 9704 4310 9716
rect 4430 9704 4436 9716
rect 4304 9676 4436 9704
rect 4304 9664 4310 9676
rect 4430 9664 4436 9676
rect 4488 9664 4494 9716
rect 4893 9707 4951 9713
rect 4893 9673 4905 9707
rect 4939 9704 4951 9707
rect 5077 9707 5135 9713
rect 5077 9704 5089 9707
rect 4939 9676 5089 9704
rect 4939 9673 4951 9676
rect 4893 9667 4951 9673
rect 5077 9673 5089 9676
rect 5123 9704 5135 9707
rect 5902 9704 5908 9716
rect 5123 9676 5908 9704
rect 5123 9673 5135 9676
rect 5077 9667 5135 9673
rect 5902 9664 5908 9676
rect 5960 9664 5966 9716
rect 6086 9664 6092 9716
rect 6144 9704 6150 9716
rect 6181 9707 6239 9713
rect 6181 9704 6193 9707
rect 6144 9676 6193 9704
rect 6144 9664 6150 9676
rect 6181 9673 6193 9676
rect 6227 9673 6239 9707
rect 6181 9667 6239 9673
rect 6638 9664 6644 9716
rect 6696 9704 6702 9716
rect 12802 9704 12808 9716
rect 6696 9676 11278 9704
rect 12763 9676 12808 9704
rect 6696 9664 6702 9676
rect 1578 9636 1584 9648
rect 1539 9608 1584 9636
rect 1578 9596 1584 9608
rect 1636 9596 1642 9648
rect 2731 9639 2789 9645
rect 2731 9605 2743 9639
rect 2777 9636 2789 9639
rect 9677 9639 9735 9645
rect 9677 9636 9689 9639
rect 2777 9608 9689 9636
rect 2777 9605 2789 9608
rect 2731 9599 2789 9605
rect 9677 9605 9689 9608
rect 9723 9636 9735 9639
rect 11146 9636 11152 9648
rect 9723 9608 11152 9636
rect 9723 9605 9735 9608
rect 9677 9599 9735 9605
rect 11146 9596 11152 9608
rect 11204 9596 11210 9648
rect 4893 9571 4951 9577
rect 4893 9568 4905 9571
rect 3620 9540 4905 9568
rect 3620 9512 3648 9540
rect 4893 9537 4905 9540
rect 4939 9537 4951 9571
rect 6822 9568 6828 9580
rect 6783 9540 6828 9568
rect 4893 9531 4951 9537
rect 6822 9528 6828 9540
rect 6880 9528 6886 9580
rect 6914 9528 6920 9580
rect 6972 9568 6978 9580
rect 8662 9568 8668 9580
rect 6972 9540 8668 9568
rect 6972 9528 6978 9540
rect 8662 9528 8668 9540
rect 8720 9528 8726 9580
rect 8938 9568 8944 9580
rect 8899 9540 8944 9568
rect 8938 9528 8944 9540
rect 8996 9528 9002 9580
rect 9582 9528 9588 9580
rect 9640 9568 9646 9580
rect 10505 9571 10563 9577
rect 10505 9568 10517 9571
rect 9640 9540 10517 9568
rect 9640 9528 9646 9540
rect 10505 9537 10517 9540
rect 10551 9568 10563 9571
rect 10594 9568 10600 9580
rect 10551 9540 10600 9568
rect 10551 9537 10563 9540
rect 10505 9531 10563 9537
rect 10594 9528 10600 9540
rect 10652 9528 10658 9580
rect 11250 9568 11278 9676
rect 12802 9664 12808 9676
rect 12860 9664 12866 9716
rect 14458 9664 14464 9716
rect 14516 9704 14522 9716
rect 14645 9707 14703 9713
rect 14645 9704 14657 9707
rect 14516 9676 14657 9704
rect 14516 9664 14522 9676
rect 14645 9673 14657 9676
rect 14691 9673 14703 9707
rect 14645 9667 14703 9673
rect 15102 9664 15108 9716
rect 15160 9704 15166 9716
rect 15289 9707 15347 9713
rect 15289 9704 15301 9707
rect 15160 9676 15301 9704
rect 15160 9664 15166 9676
rect 15289 9673 15301 9676
rect 15335 9704 15347 9707
rect 16022 9704 16028 9716
rect 15335 9676 16028 9704
rect 15335 9673 15347 9676
rect 15289 9667 15347 9673
rect 16022 9664 16028 9676
rect 16080 9664 16086 9716
rect 16298 9664 16304 9716
rect 16356 9704 16362 9716
rect 17405 9707 17463 9713
rect 17405 9704 17417 9707
rect 16356 9676 17417 9704
rect 16356 9664 16362 9676
rect 17405 9673 17417 9676
rect 17451 9673 17463 9707
rect 17405 9667 17463 9673
rect 17770 9664 17776 9716
rect 17828 9704 17834 9716
rect 19058 9704 19064 9716
rect 17828 9676 19064 9704
rect 17828 9664 17834 9676
rect 19058 9664 19064 9676
rect 19116 9664 19122 9716
rect 15933 9639 15991 9645
rect 15933 9605 15945 9639
rect 15979 9636 15991 9639
rect 16574 9636 16580 9648
rect 15979 9608 16580 9636
rect 15979 9605 15991 9608
rect 15933 9599 15991 9605
rect 16574 9596 16580 9608
rect 16632 9596 16638 9648
rect 17144 9608 18460 9636
rect 17144 9580 17172 9608
rect 13722 9568 13728 9580
rect 11250 9540 13728 9568
rect 13722 9528 13728 9540
rect 13780 9528 13786 9580
rect 16301 9571 16359 9577
rect 16301 9537 16313 9571
rect 16347 9568 16359 9571
rect 16942 9568 16948 9580
rect 16347 9540 16948 9568
rect 16347 9537 16359 9540
rect 16301 9531 16359 9537
rect 16942 9528 16948 9540
rect 17000 9528 17006 9580
rect 17126 9568 17132 9580
rect 17087 9540 17132 9568
rect 17126 9528 17132 9540
rect 17184 9528 17190 9580
rect 17586 9528 17592 9580
rect 17644 9568 17650 9580
rect 18138 9568 18144 9580
rect 17644 9540 18144 9568
rect 17644 9528 17650 9540
rect 18138 9528 18144 9540
rect 18196 9528 18202 9580
rect 18432 9577 18460 9608
rect 18690 9596 18696 9648
rect 18748 9596 18754 9648
rect 18417 9571 18475 9577
rect 18417 9537 18429 9571
rect 18463 9537 18475 9571
rect 18708 9568 18736 9596
rect 19613 9571 19671 9577
rect 19613 9568 19625 9571
rect 18708 9540 19625 9568
rect 18417 9531 18475 9537
rect 19613 9537 19625 9540
rect 19659 9537 19671 9571
rect 19613 9531 19671 9537
rect 1302 9460 1308 9512
rect 1360 9500 1366 9512
rect 1397 9503 1455 9509
rect 1397 9500 1409 9503
rect 1360 9472 1409 9500
rect 1360 9460 1366 9472
rect 1397 9469 1409 9472
rect 1443 9500 1455 9503
rect 1949 9503 2007 9509
rect 1949 9500 1961 9503
rect 1443 9472 1961 9500
rect 1443 9469 1455 9472
rect 1397 9463 1455 9469
rect 1949 9469 1961 9472
rect 1995 9469 2007 9503
rect 1949 9463 2007 9469
rect 2222 9460 2228 9512
rect 2280 9500 2286 9512
rect 2628 9503 2686 9509
rect 2628 9500 2640 9503
rect 2280 9472 2640 9500
rect 2280 9460 2286 9472
rect 2628 9469 2640 9472
rect 2674 9500 2686 9503
rect 3418 9500 3424 9512
rect 2674 9472 3424 9500
rect 2674 9469 2686 9472
rect 2628 9463 2686 9469
rect 3418 9460 3424 9472
rect 3476 9460 3482 9512
rect 3602 9500 3608 9512
rect 3563 9472 3608 9500
rect 3602 9460 3608 9472
rect 3660 9460 3666 9512
rect 3694 9460 3700 9512
rect 3752 9500 3758 9512
rect 4065 9503 4123 9509
rect 4065 9500 4077 9503
rect 3752 9472 4077 9500
rect 3752 9460 3758 9472
rect 4065 9469 4077 9472
rect 4111 9500 4123 9503
rect 4617 9503 4675 9509
rect 4617 9500 4629 9503
rect 4111 9472 4629 9500
rect 4111 9469 4123 9472
rect 4065 9463 4123 9469
rect 4617 9469 4629 9472
rect 4663 9469 4675 9503
rect 7650 9500 7656 9512
rect 4617 9463 4675 9469
rect 6472 9472 7656 9500
rect 2958 9392 2964 9444
rect 3016 9432 3022 9444
rect 5258 9432 5264 9444
rect 3016 9404 5264 9432
rect 3016 9392 3022 9404
rect 5258 9392 5264 9404
rect 5316 9392 5322 9444
rect 5353 9435 5411 9441
rect 5353 9401 5365 9435
rect 5399 9401 5411 9435
rect 5353 9395 5411 9401
rect 5905 9435 5963 9441
rect 5905 9401 5917 9435
rect 5951 9432 5963 9435
rect 6362 9432 6368 9444
rect 5951 9404 6368 9432
rect 5951 9401 5963 9404
rect 5905 9395 5963 9401
rect 3050 9364 3056 9376
rect 3011 9336 3056 9364
rect 3050 9324 3056 9336
rect 3108 9324 3114 9376
rect 3878 9364 3884 9376
rect 3839 9336 3884 9364
rect 3878 9324 3884 9336
rect 3936 9324 3942 9376
rect 5074 9324 5080 9376
rect 5132 9364 5138 9376
rect 5368 9364 5396 9395
rect 6362 9392 6368 9404
rect 6420 9392 6426 9444
rect 6472 9364 6500 9472
rect 7650 9460 7656 9472
rect 7708 9500 7714 9512
rect 7745 9503 7803 9509
rect 7745 9500 7757 9503
rect 7708 9472 7757 9500
rect 7708 9460 7714 9472
rect 7745 9469 7757 9472
rect 7791 9500 7803 9503
rect 8021 9503 8079 9509
rect 8021 9500 8033 9503
rect 7791 9472 8033 9500
rect 7791 9469 7803 9472
rect 7745 9463 7803 9469
rect 8021 9469 8033 9472
rect 8067 9469 8079 9503
rect 8021 9463 8079 9469
rect 12621 9503 12679 9509
rect 12621 9469 12633 9503
rect 12667 9500 12679 9503
rect 12989 9503 13047 9509
rect 12989 9500 13001 9503
rect 12667 9472 13001 9500
rect 12667 9469 12679 9472
rect 12621 9463 12679 9469
rect 12989 9469 13001 9472
rect 13035 9469 13047 9503
rect 12989 9463 13047 9469
rect 13556 9472 13768 9500
rect 7146 9435 7204 9441
rect 7146 9432 7158 9435
rect 6564 9404 7158 9432
rect 6564 9376 6592 9404
rect 7146 9401 7158 9404
rect 7192 9401 7204 9435
rect 7146 9395 7204 9401
rect 8757 9435 8815 9441
rect 8757 9401 8769 9435
rect 8803 9401 8815 9435
rect 8757 9395 8815 9401
rect 5132 9336 6500 9364
rect 5132 9324 5138 9336
rect 6546 9324 6552 9376
rect 6604 9364 6610 9376
rect 6604 9336 6649 9364
rect 6604 9324 6610 9336
rect 8202 9324 8208 9376
rect 8260 9364 8266 9376
rect 8389 9367 8447 9373
rect 8389 9364 8401 9367
rect 8260 9336 8401 9364
rect 8260 9324 8266 9336
rect 8389 9333 8401 9336
rect 8435 9364 8447 9367
rect 8772 9364 8800 9395
rect 10686 9392 10692 9444
rect 10744 9432 10750 9444
rect 10867 9435 10925 9441
rect 10867 9432 10879 9435
rect 10744 9404 10879 9432
rect 10744 9392 10750 9404
rect 10867 9401 10879 9404
rect 10913 9432 10925 9435
rect 11330 9432 11336 9444
rect 10913 9404 11336 9432
rect 10913 9401 10925 9404
rect 10867 9395 10925 9401
rect 11330 9392 11336 9404
rect 11388 9432 11394 9444
rect 12161 9435 12219 9441
rect 12161 9432 12173 9435
rect 11388 9404 12173 9432
rect 11388 9392 11394 9404
rect 12161 9401 12173 9404
rect 12207 9432 12219 9435
rect 13354 9432 13360 9444
rect 12207 9404 13360 9432
rect 12207 9401 12219 9404
rect 12161 9395 12219 9401
rect 13354 9392 13360 9404
rect 13412 9432 13418 9444
rect 13556 9441 13584 9472
rect 13541 9435 13599 9441
rect 13541 9432 13553 9435
rect 13412 9404 13553 9432
rect 13412 9392 13418 9404
rect 13541 9401 13553 9404
rect 13587 9401 13599 9435
rect 13740 9432 13768 9472
rect 14046 9435 14104 9441
rect 14046 9432 14058 9435
rect 13740 9404 14058 9432
rect 13541 9395 13599 9401
rect 14046 9401 14058 9404
rect 14092 9401 14104 9435
rect 16482 9432 16488 9444
rect 16443 9404 16488 9432
rect 14046 9395 14104 9401
rect 16482 9392 16488 9404
rect 16540 9392 16546 9444
rect 16574 9392 16580 9444
rect 16632 9432 16638 9444
rect 17770 9432 17776 9444
rect 16632 9404 17776 9432
rect 16632 9392 16638 9404
rect 17770 9392 17776 9404
rect 17828 9392 17834 9444
rect 18233 9435 18291 9441
rect 18233 9401 18245 9435
rect 18279 9401 18291 9435
rect 18233 9395 18291 9401
rect 8435 9336 8800 9364
rect 8435 9333 8447 9336
rect 8389 9327 8447 9333
rect 9950 9324 9956 9376
rect 10008 9364 10014 9376
rect 10045 9367 10103 9373
rect 10045 9364 10057 9367
rect 10008 9336 10057 9364
rect 10008 9324 10014 9336
rect 10045 9333 10057 9336
rect 10091 9333 10103 9367
rect 10045 9327 10103 9333
rect 11238 9324 11244 9376
rect 11296 9364 11302 9376
rect 11425 9367 11483 9373
rect 11425 9364 11437 9367
rect 11296 9336 11437 9364
rect 11296 9324 11302 9336
rect 11425 9333 11437 9336
rect 11471 9364 11483 9367
rect 11793 9367 11851 9373
rect 11793 9364 11805 9367
rect 11471 9336 11805 9364
rect 11471 9333 11483 9336
rect 11425 9327 11483 9333
rect 11793 9333 11805 9336
rect 11839 9364 11851 9367
rect 11882 9364 11888 9376
rect 11839 9336 11888 9364
rect 11839 9333 11851 9336
rect 11793 9327 11851 9333
rect 11882 9324 11888 9336
rect 11940 9324 11946 9376
rect 12989 9367 13047 9373
rect 12989 9333 13001 9367
rect 13035 9364 13047 9367
rect 13265 9367 13323 9373
rect 13265 9364 13277 9367
rect 13035 9336 13277 9364
rect 13035 9333 13047 9336
rect 12989 9327 13047 9333
rect 13265 9333 13277 9336
rect 13311 9364 13323 9367
rect 13814 9364 13820 9376
rect 13311 9336 13820 9364
rect 13311 9333 13323 9336
rect 13265 9327 13323 9333
rect 13814 9324 13820 9336
rect 13872 9364 13878 9376
rect 14182 9364 14188 9376
rect 13872 9336 14188 9364
rect 13872 9324 13878 9336
rect 14182 9324 14188 9336
rect 14240 9324 14246 9376
rect 17494 9324 17500 9376
rect 17552 9364 17558 9376
rect 17865 9367 17923 9373
rect 17865 9364 17877 9367
rect 17552 9336 17877 9364
rect 17552 9324 17558 9336
rect 17865 9333 17877 9336
rect 17911 9364 17923 9367
rect 18248 9364 18276 9395
rect 17911 9336 18276 9364
rect 19521 9367 19579 9373
rect 17911 9333 17923 9336
rect 17865 9327 17923 9333
rect 19521 9333 19533 9367
rect 19567 9364 19579 9367
rect 19610 9364 19616 9376
rect 19567 9336 19616 9364
rect 19567 9333 19579 9336
rect 19521 9327 19579 9333
rect 19610 9324 19616 9336
rect 19668 9324 19674 9376
rect 1104 9274 20884 9296
rect 1104 9222 8315 9274
rect 8367 9222 8379 9274
rect 8431 9222 8443 9274
rect 8495 9222 8507 9274
rect 8559 9222 15648 9274
rect 15700 9222 15712 9274
rect 15764 9222 15776 9274
rect 15828 9222 15840 9274
rect 15892 9222 20884 9274
rect 1104 9200 20884 9222
rect 2498 9120 2504 9172
rect 2556 9160 2562 9172
rect 3099 9163 3157 9169
rect 3099 9160 3111 9163
rect 2556 9132 3111 9160
rect 2556 9120 2562 9132
rect 3099 9129 3111 9132
rect 3145 9129 3157 9163
rect 3099 9123 3157 9129
rect 3789 9163 3847 9169
rect 3789 9129 3801 9163
rect 3835 9160 3847 9163
rect 4522 9160 4528 9172
rect 3835 9132 4528 9160
rect 3835 9129 3847 9132
rect 3789 9123 3847 9129
rect 4522 9120 4528 9132
rect 4580 9160 4586 9172
rect 4617 9163 4675 9169
rect 4617 9160 4629 9163
rect 4580 9132 4629 9160
rect 4580 9120 4586 9132
rect 4617 9129 4629 9132
rect 4663 9129 4675 9163
rect 5074 9160 5080 9172
rect 5035 9132 5080 9160
rect 4617 9123 4675 9129
rect 5074 9120 5080 9132
rect 5132 9120 5138 9172
rect 5258 9120 5264 9172
rect 5316 9160 5322 9172
rect 6181 9163 6239 9169
rect 6181 9160 6193 9163
rect 5316 9132 6193 9160
rect 5316 9120 5322 9132
rect 6181 9129 6193 9132
rect 6227 9129 6239 9163
rect 6181 9123 6239 9129
rect 6362 9120 6368 9172
rect 6420 9160 6426 9172
rect 7742 9160 7748 9172
rect 6420 9132 7748 9160
rect 6420 9120 6426 9132
rect 7742 9120 7748 9132
rect 7800 9160 7806 9172
rect 8297 9163 8355 9169
rect 8297 9160 8309 9163
rect 7800 9132 8309 9160
rect 7800 9120 7806 9132
rect 8297 9129 8309 9132
rect 8343 9160 8355 9163
rect 8938 9160 8944 9172
rect 8343 9132 8944 9160
rect 8343 9129 8355 9132
rect 8297 9123 8355 9129
rect 8938 9120 8944 9132
rect 8996 9120 9002 9172
rect 10594 9160 10600 9172
rect 10555 9132 10600 9160
rect 10594 9120 10600 9132
rect 10652 9120 10658 9172
rect 12618 9160 12624 9172
rect 12579 9132 12624 9160
rect 12618 9120 12624 9132
rect 12676 9120 12682 9172
rect 15010 9120 15016 9172
rect 15068 9160 15074 9172
rect 16025 9163 16083 9169
rect 16025 9160 16037 9163
rect 15068 9132 16037 9160
rect 15068 9120 15074 9132
rect 16025 9129 16037 9132
rect 16071 9160 16083 9163
rect 16390 9160 16396 9172
rect 16071 9132 16396 9160
rect 16071 9129 16083 9132
rect 16025 9123 16083 9129
rect 16390 9120 16396 9132
rect 16448 9120 16454 9172
rect 16942 9160 16948 9172
rect 16903 9132 16948 9160
rect 16942 9120 16948 9132
rect 17000 9120 17006 9172
rect 17494 9160 17500 9172
rect 17455 9132 17500 9160
rect 17494 9120 17500 9132
rect 17552 9120 17558 9172
rect 18138 9160 18144 9172
rect 18099 9132 18144 9160
rect 18138 9120 18144 9132
rect 18196 9120 18202 9172
rect 19058 9120 19064 9172
rect 19116 9160 19122 9172
rect 19245 9163 19303 9169
rect 19245 9160 19257 9163
rect 19116 9132 19257 9160
rect 19116 9120 19122 9132
rect 19245 9129 19257 9132
rect 19291 9129 19303 9163
rect 19245 9123 19303 9129
rect 2087 9095 2145 9101
rect 2087 9061 2099 9095
rect 2133 9092 2145 9095
rect 6914 9092 6920 9104
rect 2133 9064 6920 9092
rect 2133 9061 2145 9064
rect 2087 9055 2145 9061
rect 6914 9052 6920 9064
rect 6972 9052 6978 9104
rect 7095 9095 7153 9101
rect 7095 9061 7107 9095
rect 7141 9092 7153 9095
rect 7466 9092 7472 9104
rect 7141 9064 7472 9092
rect 7141 9061 7153 9064
rect 7095 9055 7153 9061
rect 7466 9052 7472 9064
rect 7524 9052 7530 9104
rect 7558 9052 7564 9104
rect 7616 9092 7622 9104
rect 7929 9095 7987 9101
rect 7929 9092 7941 9095
rect 7616 9064 7941 9092
rect 7616 9052 7622 9064
rect 7929 9061 7941 9064
rect 7975 9061 7987 9095
rect 8754 9092 8760 9104
rect 8715 9064 8760 9092
rect 7929 9055 7987 9061
rect 8754 9052 8760 9064
rect 8812 9052 8818 9104
rect 11333 9095 11391 9101
rect 11333 9061 11345 9095
rect 11379 9092 11391 9095
rect 11882 9092 11888 9104
rect 11379 9064 11888 9092
rect 11379 9061 11391 9064
rect 11333 9055 11391 9061
rect 11882 9052 11888 9064
rect 11940 9052 11946 9104
rect 13722 9052 13728 9104
rect 13780 9092 13786 9104
rect 13817 9095 13875 9101
rect 13817 9092 13829 9095
rect 13780 9064 13829 9092
rect 13780 9052 13786 9064
rect 13817 9061 13829 9064
rect 13863 9061 13875 9095
rect 13817 9055 13875 9061
rect 14369 9095 14427 9101
rect 14369 9061 14381 9095
rect 14415 9092 14427 9095
rect 14642 9092 14648 9104
rect 14415 9064 14648 9092
rect 14415 9061 14427 9064
rect 14369 9055 14427 9061
rect 14642 9052 14648 9064
rect 14700 9052 14706 9104
rect 16960 9092 16988 9120
rect 18646 9095 18704 9101
rect 18646 9092 18658 9095
rect 16960 9064 18658 9092
rect 18646 9061 18658 9064
rect 18692 9092 18704 9095
rect 19150 9092 19156 9104
rect 18692 9064 19156 9092
rect 18692 9061 18704 9064
rect 18646 9055 18704 9061
rect 19150 9052 19156 9064
rect 19208 9052 19214 9104
rect 1946 9024 1952 9036
rect 1907 8996 1952 9024
rect 1946 8984 1952 8996
rect 2004 8984 2010 9036
rect 2869 9027 2927 9033
rect 2869 8993 2881 9027
rect 2915 9024 2927 9027
rect 3028 9027 3086 9033
rect 3028 9024 3040 9027
rect 2915 8996 3040 9024
rect 2915 8993 2927 8996
rect 2869 8987 2927 8993
rect 3028 8993 3040 8996
rect 3074 9024 3086 9027
rect 5074 9024 5080 9036
rect 3074 8996 5080 9024
rect 3074 8993 3086 8996
rect 3028 8987 3086 8993
rect 5074 8984 5080 8996
rect 5132 8984 5138 9036
rect 5353 9027 5411 9033
rect 5353 8993 5365 9027
rect 5399 8993 5411 9027
rect 5626 9024 5632 9036
rect 5587 8996 5632 9024
rect 5353 8987 5411 8993
rect 4154 8916 4160 8968
rect 4212 8956 4218 8968
rect 5368 8956 5396 8987
rect 5626 8984 5632 8996
rect 5684 8984 5690 9036
rect 6086 8984 6092 9036
rect 6144 9024 6150 9036
rect 7653 9027 7711 9033
rect 7653 9024 7665 9027
rect 6144 8996 7665 9024
rect 6144 8984 6150 8996
rect 7653 8993 7665 8996
rect 7699 9024 7711 9027
rect 8202 9024 8208 9036
rect 7699 8996 8208 9024
rect 7699 8993 7711 8996
rect 7653 8987 7711 8993
rect 8202 8984 8208 8996
rect 8260 8984 8266 9036
rect 8481 9027 8539 9033
rect 8481 8993 8493 9027
rect 8527 9024 8539 9027
rect 8662 9024 8668 9036
rect 8527 8996 8668 9024
rect 8527 8993 8539 8996
rect 8481 8987 8539 8993
rect 8662 8984 8668 8996
rect 8720 8984 8726 9036
rect 10045 9027 10103 9033
rect 10045 8993 10057 9027
rect 10091 8993 10103 9027
rect 15470 9024 15476 9036
rect 15431 8996 15476 9024
rect 10045 8987 10103 8993
rect 5442 8956 5448 8968
rect 4212 8928 4257 8956
rect 5368 8928 5448 8956
rect 4212 8916 4218 8928
rect 5442 8916 5448 8928
rect 5500 8916 5506 8968
rect 5905 8959 5963 8965
rect 5905 8925 5917 8959
rect 5951 8956 5963 8959
rect 6638 8956 6644 8968
rect 5951 8928 6644 8956
rect 5951 8925 5963 8928
rect 5905 8919 5963 8925
rect 6638 8916 6644 8928
rect 6696 8916 6702 8968
rect 6733 8959 6791 8965
rect 6733 8925 6745 8959
rect 6779 8925 6791 8959
rect 6733 8919 6791 8925
rect 2498 8848 2504 8900
rect 2556 8888 2562 8900
rect 3789 8891 3847 8897
rect 3789 8888 3801 8891
rect 2556 8860 3801 8888
rect 2556 8848 2562 8860
rect 3789 8857 3801 8860
rect 3835 8857 3847 8891
rect 3789 8851 3847 8857
rect 3970 8848 3976 8900
rect 4028 8888 4034 8900
rect 6748 8888 6776 8919
rect 8110 8916 8116 8968
rect 8168 8956 8174 8968
rect 9306 8956 9312 8968
rect 8168 8928 9312 8956
rect 8168 8916 8174 8928
rect 9306 8916 9312 8928
rect 9364 8956 9370 8968
rect 10060 8956 10088 8987
rect 15470 8984 15476 8996
rect 15528 8984 15534 9036
rect 16482 8984 16488 9036
rect 16540 9024 16546 9036
rect 17586 9024 17592 9036
rect 16540 8996 17592 9024
rect 16540 8984 16546 8996
rect 17586 8984 17592 8996
rect 17644 8984 17650 9036
rect 10410 8956 10416 8968
rect 9364 8928 10416 8956
rect 9364 8916 9370 8928
rect 10410 8916 10416 8928
rect 10468 8916 10474 8968
rect 10962 8916 10968 8968
rect 11020 8956 11026 8968
rect 11241 8959 11299 8965
rect 11241 8956 11253 8959
rect 11020 8928 11253 8956
rect 11020 8916 11026 8928
rect 11241 8925 11253 8928
rect 11287 8925 11299 8959
rect 11241 8919 11299 8925
rect 11885 8959 11943 8965
rect 11885 8925 11897 8959
rect 11931 8956 11943 8959
rect 12342 8956 12348 8968
rect 11931 8928 12348 8956
rect 11931 8925 11943 8928
rect 11885 8919 11943 8925
rect 12342 8916 12348 8928
rect 12400 8956 12406 8968
rect 13446 8956 13452 8968
rect 12400 8928 13452 8956
rect 12400 8916 12406 8928
rect 13446 8916 13452 8928
rect 13504 8956 13510 8968
rect 13725 8959 13783 8965
rect 13725 8956 13737 8959
rect 13504 8928 13737 8956
rect 13504 8916 13510 8928
rect 13725 8925 13737 8928
rect 13771 8925 13783 8959
rect 13725 8919 13783 8925
rect 16577 8959 16635 8965
rect 16577 8925 16589 8959
rect 16623 8956 16635 8959
rect 17402 8956 17408 8968
rect 16623 8928 17408 8956
rect 16623 8925 16635 8928
rect 16577 8919 16635 8925
rect 17402 8916 17408 8928
rect 17460 8916 17466 8968
rect 18230 8916 18236 8968
rect 18288 8956 18294 8968
rect 18325 8959 18383 8965
rect 18325 8956 18337 8959
rect 18288 8928 18337 8956
rect 18288 8916 18294 8928
rect 18325 8925 18337 8928
rect 18371 8925 18383 8959
rect 18325 8919 18383 8925
rect 7374 8888 7380 8900
rect 4028 8860 7380 8888
rect 4028 8848 4034 8860
rect 7374 8848 7380 8860
rect 7432 8848 7438 8900
rect 10229 8891 10287 8897
rect 10229 8857 10241 8891
rect 10275 8888 10287 8891
rect 11698 8888 11704 8900
rect 10275 8860 11704 8888
rect 10275 8857 10287 8860
rect 10229 8851 10287 8857
rect 11698 8848 11704 8860
rect 11756 8848 11762 8900
rect 15657 8891 15715 8897
rect 15657 8857 15669 8891
rect 15703 8888 15715 8891
rect 21542 8888 21548 8900
rect 15703 8860 21548 8888
rect 15703 8857 15715 8860
rect 15657 8851 15715 8857
rect 21542 8848 21548 8860
rect 21600 8848 21606 8900
rect 3694 8820 3700 8832
rect 3655 8792 3700 8820
rect 3694 8780 3700 8792
rect 3752 8780 3758 8832
rect 5350 8780 5356 8832
rect 5408 8820 5414 8832
rect 5994 8820 6000 8832
rect 5408 8792 6000 8820
rect 5408 8780 5414 8792
rect 5994 8780 6000 8792
rect 6052 8820 6058 8832
rect 6549 8823 6607 8829
rect 6549 8820 6561 8823
rect 6052 8792 6561 8820
rect 6052 8780 6058 8792
rect 6549 8789 6561 8792
rect 6595 8789 6607 8823
rect 6549 8783 6607 8789
rect 7190 8780 7196 8832
rect 7248 8820 7254 8832
rect 10502 8820 10508 8832
rect 7248 8792 10508 8820
rect 7248 8780 7254 8792
rect 10502 8780 10508 8792
rect 10560 8780 10566 8832
rect 10962 8820 10968 8832
rect 10923 8792 10968 8820
rect 10962 8780 10968 8792
rect 11020 8780 11026 8832
rect 16206 8780 16212 8832
rect 16264 8820 16270 8832
rect 16393 8823 16451 8829
rect 16393 8820 16405 8823
rect 16264 8792 16405 8820
rect 16264 8780 16270 8792
rect 16393 8789 16405 8792
rect 16439 8789 16451 8823
rect 16393 8783 16451 8789
rect 1104 8730 20884 8752
rect 1104 8678 4648 8730
rect 4700 8678 4712 8730
rect 4764 8678 4776 8730
rect 4828 8678 4840 8730
rect 4892 8678 11982 8730
rect 12034 8678 12046 8730
rect 12098 8678 12110 8730
rect 12162 8678 12174 8730
rect 12226 8678 19315 8730
rect 19367 8678 19379 8730
rect 19431 8678 19443 8730
rect 19495 8678 19507 8730
rect 19559 8678 20884 8730
rect 1104 8656 20884 8678
rect 1946 8616 1952 8628
rect 1907 8588 1952 8616
rect 1946 8576 1952 8588
rect 2004 8576 2010 8628
rect 5442 8576 5448 8628
rect 5500 8616 5506 8628
rect 6270 8616 6276 8628
rect 5500 8588 6276 8616
rect 5500 8576 5506 8588
rect 6270 8576 6276 8588
rect 6328 8576 6334 8628
rect 7374 8616 7380 8628
rect 7335 8588 7380 8616
rect 7374 8576 7380 8588
rect 7432 8576 7438 8628
rect 7466 8576 7472 8628
rect 7524 8616 7530 8628
rect 9033 8619 9091 8625
rect 9033 8616 9045 8619
rect 7524 8588 9045 8616
rect 7524 8576 7530 8588
rect 9033 8585 9045 8588
rect 9079 8616 9091 8619
rect 9490 8616 9496 8628
rect 9079 8588 9496 8616
rect 9079 8585 9091 8588
rect 9033 8579 9091 8585
rect 9490 8576 9496 8588
rect 9548 8576 9554 8628
rect 10410 8616 10416 8628
rect 10371 8588 10416 8616
rect 10410 8576 10416 8588
rect 10468 8576 10474 8628
rect 11241 8619 11299 8625
rect 11241 8616 11253 8619
rect 10520 8588 11253 8616
rect 2958 8508 2964 8560
rect 3016 8548 3022 8560
rect 3694 8548 3700 8560
rect 3016 8520 3700 8548
rect 3016 8508 3022 8520
rect 2038 8412 2044 8424
rect 1997 8384 2044 8412
rect 2038 8372 2044 8384
rect 2096 8421 2102 8424
rect 2096 8415 2145 8421
rect 2096 8381 2099 8415
rect 2133 8381 2145 8415
rect 3326 8412 3332 8424
rect 3287 8384 3332 8412
rect 2096 8375 2145 8381
rect 2096 8372 2130 8375
rect 3326 8372 3332 8384
rect 3384 8372 3390 8424
rect 3620 8421 3648 8520
rect 3694 8508 3700 8520
rect 3752 8508 3758 8560
rect 3878 8508 3884 8560
rect 3936 8548 3942 8560
rect 4065 8551 4123 8557
rect 4065 8548 4077 8551
rect 3936 8520 4077 8548
rect 3936 8508 3942 8520
rect 4065 8517 4077 8520
rect 4111 8517 4123 8551
rect 4065 8511 4123 8517
rect 4525 8551 4583 8557
rect 4525 8517 4537 8551
rect 4571 8548 4583 8551
rect 5166 8548 5172 8560
rect 4571 8520 5172 8548
rect 4571 8517 4583 8520
rect 4525 8511 4583 8517
rect 4080 8480 4108 8511
rect 5166 8508 5172 8520
rect 5224 8548 5230 8560
rect 6454 8548 6460 8560
rect 5224 8520 6460 8548
rect 5224 8508 5230 8520
rect 6454 8508 6460 8520
rect 6512 8548 6518 8560
rect 7009 8551 7067 8557
rect 7009 8548 7021 8551
rect 6512 8520 7021 8548
rect 6512 8508 6518 8520
rect 7009 8517 7021 8520
rect 7055 8548 7067 8551
rect 7484 8548 7512 8576
rect 7055 8520 7512 8548
rect 7576 8520 9260 8548
rect 7055 8517 7067 8520
rect 7009 8511 7067 8517
rect 4617 8483 4675 8489
rect 4617 8480 4629 8483
rect 4080 8452 4629 8480
rect 4617 8449 4629 8452
rect 4663 8449 4675 8483
rect 4617 8443 4675 8449
rect 3605 8415 3663 8421
rect 3605 8381 3617 8415
rect 3651 8381 3663 8415
rect 3605 8375 3663 8381
rect 3789 8415 3847 8421
rect 3789 8381 3801 8415
rect 3835 8412 3847 8415
rect 7576 8412 7604 8520
rect 9232 8492 9260 8520
rect 10226 8508 10232 8560
rect 10284 8548 10290 8560
rect 10520 8548 10548 8588
rect 11241 8585 11253 8588
rect 11287 8585 11299 8619
rect 13722 8616 13728 8628
rect 13683 8588 13728 8616
rect 11241 8579 11299 8585
rect 13722 8576 13728 8588
rect 13780 8576 13786 8628
rect 15470 8616 15476 8628
rect 15431 8588 15476 8616
rect 15470 8576 15476 8588
rect 15528 8576 15534 8628
rect 17494 8576 17500 8628
rect 17552 8616 17558 8628
rect 17773 8619 17831 8625
rect 17773 8616 17785 8619
rect 17552 8588 17785 8616
rect 17552 8576 17558 8588
rect 17773 8585 17785 8588
rect 17819 8616 17831 8619
rect 18322 8616 18328 8628
rect 17819 8588 18328 8616
rect 17819 8585 17831 8588
rect 17773 8579 17831 8585
rect 18322 8576 18328 8588
rect 18380 8576 18386 8628
rect 19150 8616 19156 8628
rect 19111 8588 19156 8616
rect 19150 8576 19156 8588
rect 19208 8576 19214 8628
rect 10284 8520 10548 8548
rect 10284 8508 10290 8520
rect 11882 8508 11888 8560
rect 11940 8548 11946 8560
rect 12161 8551 12219 8557
rect 12161 8548 12173 8551
rect 11940 8520 12173 8548
rect 11940 8508 11946 8520
rect 12161 8517 12173 8520
rect 12207 8517 12219 8551
rect 13078 8548 13084 8560
rect 13039 8520 13084 8548
rect 12161 8511 12219 8517
rect 13078 8508 13084 8520
rect 13136 8508 13142 8560
rect 18782 8548 18788 8560
rect 18743 8520 18788 8548
rect 18782 8508 18788 8520
rect 18840 8508 18846 8560
rect 7742 8480 7748 8492
rect 7703 8452 7748 8480
rect 7742 8440 7748 8452
rect 7800 8440 7806 8492
rect 7926 8440 7932 8492
rect 7984 8480 7990 8492
rect 8021 8483 8079 8489
rect 8021 8480 8033 8483
rect 7984 8452 8033 8480
rect 7984 8440 7990 8452
rect 8021 8449 8033 8452
rect 8067 8449 8079 8483
rect 9214 8480 9220 8492
rect 9127 8452 9220 8480
rect 8021 8443 8079 8449
rect 9214 8440 9220 8452
rect 9272 8440 9278 8492
rect 12529 8483 12587 8489
rect 12529 8449 12541 8483
rect 12575 8480 12587 8483
rect 12710 8480 12716 8492
rect 12575 8452 12716 8480
rect 12575 8449 12587 8452
rect 12529 8443 12587 8449
rect 12710 8440 12716 8452
rect 12768 8440 12774 8492
rect 14642 8440 14648 8492
rect 14700 8480 14706 8492
rect 14737 8483 14795 8489
rect 14737 8480 14749 8483
rect 14700 8452 14749 8480
rect 14700 8440 14706 8452
rect 14737 8449 14749 8452
rect 14783 8449 14795 8483
rect 14737 8443 14795 8449
rect 14918 8440 14924 8492
rect 14976 8480 14982 8492
rect 16669 8483 16727 8489
rect 14976 8452 15332 8480
rect 14976 8440 14982 8452
rect 15304 8424 15332 8452
rect 16669 8449 16681 8483
rect 16715 8480 16727 8483
rect 17678 8480 17684 8492
rect 16715 8452 17684 8480
rect 16715 8449 16727 8452
rect 16669 8443 16727 8449
rect 17678 8440 17684 8452
rect 17736 8440 17742 8492
rect 18233 8483 18291 8489
rect 18233 8449 18245 8483
rect 18279 8480 18291 8483
rect 18279 8452 19656 8480
rect 18279 8449 18291 8452
rect 18233 8443 18291 8449
rect 11149 8415 11207 8421
rect 11149 8412 11161 8415
rect 3835 8384 7604 8412
rect 8496 8384 11161 8412
rect 3835 8381 3847 8384
rect 3789 8375 3847 8381
rect 2102 8276 2130 8372
rect 2179 8347 2237 8353
rect 2179 8313 2191 8347
rect 2225 8344 2237 8347
rect 4979 8347 5037 8353
rect 2225 8316 4844 8344
rect 2225 8313 2237 8316
rect 2179 8307 2237 8313
rect 2590 8276 2596 8288
rect 2102 8248 2596 8276
rect 2590 8236 2596 8248
rect 2648 8236 2654 8288
rect 2958 8276 2964 8288
rect 2919 8248 2964 8276
rect 2958 8236 2964 8248
rect 3016 8236 3022 8288
rect 3050 8236 3056 8288
rect 3108 8276 3114 8288
rect 4062 8276 4068 8288
rect 3108 8248 4068 8276
rect 3108 8236 3114 8248
rect 4062 8236 4068 8248
rect 4120 8236 4126 8288
rect 4816 8276 4844 8316
rect 4979 8313 4991 8347
rect 5025 8344 5037 8347
rect 5166 8344 5172 8356
rect 5025 8316 5172 8344
rect 5025 8313 5037 8316
rect 4979 8307 5037 8313
rect 5166 8304 5172 8316
rect 5224 8304 5230 8356
rect 7846 8347 7904 8353
rect 7846 8313 7858 8347
rect 7892 8344 7904 8347
rect 7892 8316 7972 8344
rect 7892 8313 7904 8316
rect 7846 8307 7904 8313
rect 5350 8276 5356 8288
rect 4816 8248 5356 8276
rect 5350 8236 5356 8248
rect 5408 8236 5414 8288
rect 5534 8276 5540 8288
rect 5495 8248 5540 8276
rect 5534 8236 5540 8248
rect 5592 8236 5598 8288
rect 5626 8236 5632 8288
rect 5684 8276 5690 8288
rect 5813 8279 5871 8285
rect 5813 8276 5825 8279
rect 5684 8248 5825 8276
rect 5684 8236 5690 8248
rect 5813 8245 5825 8248
rect 5859 8245 5871 8279
rect 7944 8276 7972 8316
rect 8018 8304 8024 8356
rect 8076 8344 8082 8356
rect 8496 8344 8524 8384
rect 11149 8381 11161 8384
rect 11195 8412 11207 8415
rect 11793 8415 11851 8421
rect 11793 8412 11805 8415
rect 11195 8384 11805 8412
rect 11195 8381 11207 8384
rect 11149 8375 11207 8381
rect 11793 8381 11805 8384
rect 11839 8381 11851 8415
rect 11793 8375 11851 8381
rect 9490 8344 9496 8356
rect 8076 8316 8524 8344
rect 8588 8316 9168 8344
rect 9451 8316 9496 8344
rect 8076 8304 8082 8316
rect 8110 8276 8116 8288
rect 7944 8248 8116 8276
rect 5813 8239 5871 8245
rect 8110 8236 8116 8248
rect 8168 8276 8174 8288
rect 8588 8276 8616 8316
rect 8168 8248 8616 8276
rect 8168 8236 8174 8248
rect 8662 8236 8668 8288
rect 8720 8276 8726 8288
rect 9140 8276 9168 8316
rect 9490 8304 9496 8316
rect 9548 8304 9554 8356
rect 10318 8304 10324 8356
rect 10376 8344 10382 8356
rect 10873 8347 10931 8353
rect 10873 8344 10885 8347
rect 10376 8316 10885 8344
rect 10376 8304 10382 8316
rect 10873 8313 10885 8316
rect 10919 8344 10931 8347
rect 10965 8347 11023 8353
rect 10965 8344 10977 8347
rect 10919 8316 10977 8344
rect 10919 8313 10931 8316
rect 10873 8307 10931 8313
rect 10965 8313 10977 8316
rect 11011 8313 11023 8347
rect 11808 8344 11836 8375
rect 15286 8372 15292 8424
rect 15344 8412 15350 8424
rect 15933 8415 15991 8421
rect 15933 8412 15945 8415
rect 15344 8384 15945 8412
rect 15344 8372 15350 8384
rect 15933 8381 15945 8384
rect 15979 8412 15991 8415
rect 16206 8412 16212 8424
rect 15979 8384 16212 8412
rect 15979 8381 15991 8384
rect 15933 8375 15991 8381
rect 16206 8372 16212 8384
rect 16264 8372 16270 8424
rect 16390 8412 16396 8424
rect 16351 8384 16396 8412
rect 16390 8372 16396 8384
rect 16448 8372 16454 8424
rect 12526 8344 12532 8356
rect 11808 8316 12532 8344
rect 10965 8307 11023 8313
rect 12526 8304 12532 8316
rect 12584 8304 12590 8356
rect 12618 8304 12624 8356
rect 12676 8344 12682 8356
rect 12676 8316 12721 8344
rect 12676 8304 12682 8316
rect 13262 8304 13268 8356
rect 13320 8344 13326 8356
rect 14185 8347 14243 8353
rect 14185 8344 14197 8347
rect 13320 8316 14197 8344
rect 13320 8304 13326 8316
rect 14185 8313 14197 8316
rect 14231 8344 14243 8347
rect 14461 8347 14519 8353
rect 14461 8344 14473 8347
rect 14231 8316 14473 8344
rect 14231 8313 14243 8316
rect 14185 8307 14243 8313
rect 14461 8313 14473 8316
rect 14507 8313 14519 8347
rect 14461 8307 14519 8313
rect 14553 8347 14611 8353
rect 14553 8313 14565 8347
rect 14599 8344 14611 8347
rect 14642 8344 14648 8356
rect 14599 8316 14648 8344
rect 14599 8313 14611 8316
rect 14553 8307 14611 8313
rect 14642 8304 14648 8316
rect 14700 8304 14706 8356
rect 18322 8304 18328 8356
rect 18380 8344 18386 8356
rect 18380 8316 18425 8344
rect 18380 8304 18386 8316
rect 10137 8279 10195 8285
rect 10137 8276 10149 8279
rect 8720 8248 8765 8276
rect 9140 8248 10149 8276
rect 8720 8236 8726 8248
rect 10137 8245 10149 8248
rect 10183 8245 10195 8279
rect 16942 8276 16948 8288
rect 16903 8248 16948 8276
rect 10137 8239 10195 8245
rect 16942 8236 16948 8248
rect 17000 8236 17006 8288
rect 17402 8276 17408 8288
rect 17315 8248 17408 8276
rect 17402 8236 17408 8248
rect 17460 8276 17466 8288
rect 18966 8276 18972 8288
rect 17460 8248 18972 8276
rect 17460 8236 17466 8248
rect 18966 8236 18972 8248
rect 19024 8236 19030 8288
rect 19628 8285 19656 8452
rect 19613 8279 19671 8285
rect 19613 8245 19625 8279
rect 19659 8276 19671 8279
rect 19886 8276 19892 8288
rect 19659 8248 19892 8276
rect 19659 8245 19671 8248
rect 19613 8239 19671 8245
rect 19886 8236 19892 8248
rect 19944 8236 19950 8288
rect 1104 8186 20884 8208
rect 1104 8134 8315 8186
rect 8367 8134 8379 8186
rect 8431 8134 8443 8186
rect 8495 8134 8507 8186
rect 8559 8134 15648 8186
rect 15700 8134 15712 8186
rect 15764 8134 15776 8186
rect 15828 8134 15840 8186
rect 15892 8134 20884 8186
rect 1104 8112 20884 8134
rect 2498 8072 2504 8084
rect 2459 8044 2504 8072
rect 2498 8032 2504 8044
rect 2556 8032 2562 8084
rect 2869 8075 2927 8081
rect 2869 8041 2881 8075
rect 2915 8072 2927 8075
rect 3050 8072 3056 8084
rect 2915 8044 3056 8072
rect 2915 8041 2927 8044
rect 2869 8035 2927 8041
rect 3050 8032 3056 8044
rect 3108 8032 3114 8084
rect 3326 8032 3332 8084
rect 3384 8072 3390 8084
rect 3421 8075 3479 8081
rect 3421 8072 3433 8075
rect 3384 8044 3433 8072
rect 3384 8032 3390 8044
rect 3421 8041 3433 8044
rect 3467 8041 3479 8075
rect 3421 8035 3479 8041
rect 1946 7936 1952 7948
rect 1910 7908 1952 7936
rect 1946 7896 1952 7908
rect 2004 7945 2010 7948
rect 2004 7939 2058 7945
rect 2004 7905 2012 7939
rect 2046 7936 2058 7939
rect 2406 7936 2412 7948
rect 2046 7908 2412 7936
rect 2046 7905 2058 7908
rect 2004 7899 2058 7905
rect 2004 7896 2010 7899
rect 2406 7896 2412 7908
rect 2464 7896 2470 7948
rect 3028 7939 3086 7945
rect 3028 7905 3040 7939
rect 3074 7936 3086 7939
rect 3234 7936 3240 7948
rect 3074 7908 3240 7936
rect 3074 7905 3086 7908
rect 3028 7899 3086 7905
rect 3234 7896 3240 7908
rect 3292 7896 3298 7948
rect 3436 7936 3464 8035
rect 4154 8032 4160 8084
rect 4212 8072 4218 8084
rect 4709 8075 4767 8081
rect 4709 8072 4721 8075
rect 4212 8044 4721 8072
rect 4212 8032 4218 8044
rect 4709 8041 4721 8044
rect 4755 8041 4767 8075
rect 5534 8072 5540 8084
rect 4709 8035 4767 8041
rect 5092 8044 5540 8072
rect 3605 8007 3663 8013
rect 3605 7973 3617 8007
rect 3651 8004 3663 8007
rect 4249 8007 4307 8013
rect 4249 8004 4261 8007
rect 3651 7976 4261 8004
rect 3651 7973 3663 7976
rect 3605 7967 3663 7973
rect 4249 7973 4261 7976
rect 4295 7973 4307 8007
rect 4724 8004 4752 8035
rect 5092 8013 5120 8044
rect 5534 8032 5540 8044
rect 5592 8072 5598 8084
rect 5905 8075 5963 8081
rect 5905 8072 5917 8075
rect 5592 8044 5917 8072
rect 5592 8032 5598 8044
rect 5905 8041 5917 8044
rect 5951 8041 5963 8075
rect 8846 8072 8852 8084
rect 5905 8035 5963 8041
rect 7944 8044 8754 8072
rect 8807 8044 8852 8072
rect 7944 8016 7972 8044
rect 4985 8007 5043 8013
rect 4985 8004 4997 8007
rect 4724 7976 4997 8004
rect 4249 7967 4307 7973
rect 4985 7973 4997 7976
rect 5031 7973 5043 8007
rect 4985 7967 5043 7973
rect 5077 8007 5135 8013
rect 5077 7973 5089 8007
rect 5123 7973 5135 8007
rect 5077 7967 5135 7973
rect 5721 8007 5779 8013
rect 5721 7973 5733 8007
rect 5767 8004 5779 8007
rect 7926 8004 7932 8016
rect 5767 7976 7932 8004
rect 5767 7973 5779 7976
rect 5721 7967 5779 7973
rect 7926 7964 7932 7976
rect 7984 7964 7990 8016
rect 8021 8007 8079 8013
rect 8021 7973 8033 8007
rect 8067 8004 8079 8007
rect 8110 8004 8116 8016
rect 8067 7976 8116 8004
rect 8067 7973 8079 7976
rect 8021 7967 8079 7973
rect 8110 7964 8116 7976
rect 8168 7964 8174 8016
rect 8726 8004 8754 8044
rect 8846 8032 8852 8044
rect 8904 8032 8910 8084
rect 9214 8072 9220 8084
rect 9175 8044 9220 8072
rect 9214 8032 9220 8044
rect 9272 8032 9278 8084
rect 9861 8075 9919 8081
rect 9861 8041 9873 8075
rect 9907 8072 9919 8075
rect 13262 8072 13268 8084
rect 9907 8044 13268 8072
rect 9907 8041 9919 8044
rect 9861 8035 9919 8041
rect 13262 8032 13268 8044
rect 13320 8032 13326 8084
rect 13538 8032 13544 8084
rect 13596 8072 13602 8084
rect 13633 8075 13691 8081
rect 13633 8072 13645 8075
rect 13596 8044 13645 8072
rect 13596 8032 13602 8044
rect 13633 8041 13645 8044
rect 13679 8041 13691 8075
rect 13633 8035 13691 8041
rect 13722 8032 13728 8084
rect 13780 8072 13786 8084
rect 14185 8075 14243 8081
rect 14185 8072 14197 8075
rect 13780 8044 14197 8072
rect 13780 8032 13786 8044
rect 14185 8041 14197 8044
rect 14231 8041 14243 8075
rect 14185 8035 14243 8041
rect 15378 8032 15384 8084
rect 15436 8072 15442 8084
rect 18969 8075 19027 8081
rect 18969 8072 18981 8075
rect 15436 8044 18981 8072
rect 15436 8032 15442 8044
rect 18969 8041 18981 8044
rect 19015 8041 19027 8075
rect 18969 8035 19027 8041
rect 9398 8004 9404 8016
rect 8726 7976 9404 8004
rect 9398 7964 9404 7976
rect 9456 7964 9462 8016
rect 11235 8007 11293 8013
rect 11235 7973 11247 8007
rect 11281 8004 11293 8007
rect 11330 8004 11336 8016
rect 11281 7976 11336 8004
rect 11281 7973 11293 7976
rect 11235 7967 11293 7973
rect 11330 7964 11336 7976
rect 11388 7964 11394 8016
rect 16574 7964 16580 8016
rect 16632 8004 16638 8016
rect 16853 8007 16911 8013
rect 16853 8004 16865 8007
rect 16632 7976 16865 8004
rect 16632 7964 16638 7976
rect 16853 7973 16865 7976
rect 16899 8004 16911 8007
rect 17494 8004 17500 8016
rect 16899 7976 17500 8004
rect 16899 7973 16911 7976
rect 16853 7967 16911 7973
rect 17494 7964 17500 7976
rect 17552 7964 17558 8016
rect 18138 7964 18144 8016
rect 18196 8004 18202 8016
rect 18506 8004 18512 8016
rect 18196 7976 18512 8004
rect 18196 7964 18202 7976
rect 18506 7964 18512 7976
rect 18564 8004 18570 8016
rect 18693 8007 18751 8013
rect 18693 8004 18705 8007
rect 18564 7976 18705 8004
rect 18564 7964 18570 7976
rect 18693 7973 18705 7976
rect 18739 7973 18751 8007
rect 18693 7967 18751 7973
rect 4430 7936 4436 7948
rect 3436 7908 4436 7936
rect 4430 7896 4436 7908
rect 4488 7896 4494 7948
rect 6892 7939 6950 7945
rect 6892 7905 6904 7939
rect 6938 7936 6950 7939
rect 7098 7936 7104 7948
rect 6938 7908 7104 7936
rect 6938 7905 6950 7908
rect 6892 7899 6950 7905
rect 7098 7896 7104 7908
rect 7156 7896 7162 7948
rect 7650 7936 7656 7948
rect 7611 7908 7656 7936
rect 7650 7896 7656 7908
rect 7708 7896 7714 7948
rect 9766 7896 9772 7948
rect 9824 7936 9830 7948
rect 13265 7939 13323 7945
rect 13265 7936 13277 7939
rect 9824 7908 13277 7936
rect 9824 7896 9830 7908
rect 13265 7905 13277 7908
rect 13311 7936 13323 7939
rect 13446 7936 13452 7948
rect 13311 7908 13452 7936
rect 13311 7905 13323 7908
rect 13265 7899 13323 7905
rect 13446 7896 13452 7908
rect 13504 7896 13510 7948
rect 13906 7896 13912 7948
rect 13964 7936 13970 7948
rect 15749 7939 15807 7945
rect 15749 7936 15761 7939
rect 13964 7908 15761 7936
rect 13964 7896 13970 7908
rect 15749 7905 15761 7908
rect 15795 7936 15807 7939
rect 16114 7936 16120 7948
rect 15795 7908 16120 7936
rect 15795 7905 15807 7908
rect 15749 7899 15807 7905
rect 16114 7896 16120 7908
rect 16172 7896 16178 7948
rect 16301 7939 16359 7945
rect 16301 7905 16313 7939
rect 16347 7936 16359 7939
rect 16390 7936 16396 7948
rect 16347 7908 16396 7936
rect 16347 7905 16359 7908
rect 16301 7899 16359 7905
rect 16390 7896 16396 7908
rect 16448 7896 16454 7948
rect 18874 7936 18880 7948
rect 18835 7908 18880 7936
rect 18874 7896 18880 7908
rect 18932 7896 18938 7948
rect 19058 7896 19064 7948
rect 19116 7936 19122 7948
rect 19337 7939 19395 7945
rect 19337 7936 19349 7939
rect 19116 7908 19349 7936
rect 19116 7896 19122 7908
rect 19337 7905 19349 7908
rect 19383 7905 19395 7939
rect 19337 7899 19395 7905
rect 2087 7871 2145 7877
rect 2087 7837 2099 7871
rect 2133 7868 2145 7871
rect 7926 7868 7932 7880
rect 2133 7840 7932 7868
rect 2133 7837 2145 7840
rect 2087 7831 2145 7837
rect 7926 7828 7932 7840
rect 7984 7828 7990 7880
rect 8205 7871 8263 7877
rect 8205 7837 8217 7871
rect 8251 7837 8263 7871
rect 8205 7831 8263 7837
rect 1857 7803 1915 7809
rect 1857 7769 1869 7803
rect 1903 7800 1915 7803
rect 2866 7800 2872 7812
rect 1903 7772 2872 7800
rect 1903 7769 1915 7772
rect 1857 7763 1915 7769
rect 2866 7760 2872 7772
rect 2924 7760 2930 7812
rect 3099 7803 3157 7809
rect 3099 7769 3111 7803
rect 3145 7800 3157 7803
rect 3145 7772 5022 7800
rect 3145 7769 3157 7772
rect 3099 7763 3157 7769
rect 2884 7732 2912 7760
rect 3605 7735 3663 7741
rect 3605 7732 3617 7735
rect 2884 7704 3617 7732
rect 3605 7701 3617 7704
rect 3651 7701 3663 7735
rect 3605 7695 3663 7701
rect 3881 7735 3939 7741
rect 3881 7701 3893 7735
rect 3927 7732 3939 7735
rect 4430 7732 4436 7744
rect 3927 7704 4436 7732
rect 3927 7701 3939 7704
rect 3881 7695 3939 7701
rect 4430 7692 4436 7704
rect 4488 7692 4494 7744
rect 4994 7732 5022 7772
rect 5074 7760 5080 7812
rect 5132 7800 5138 7812
rect 5537 7803 5595 7809
rect 5537 7800 5549 7803
rect 5132 7772 5549 7800
rect 5132 7760 5138 7772
rect 5537 7769 5549 7772
rect 5583 7800 5595 7803
rect 5721 7803 5779 7809
rect 5721 7800 5733 7803
rect 5583 7772 5733 7800
rect 5583 7769 5595 7772
rect 5537 7763 5595 7769
rect 5721 7769 5733 7772
rect 5767 7769 5779 7803
rect 5721 7763 5779 7769
rect 6963 7803 7021 7809
rect 6963 7769 6975 7803
rect 7009 7800 7021 7803
rect 7009 7772 7465 7800
rect 7009 7769 7021 7772
rect 6963 7763 7021 7769
rect 5810 7732 5816 7744
rect 4994 7704 5816 7732
rect 5810 7692 5816 7704
rect 5868 7692 5874 7744
rect 7282 7732 7288 7744
rect 7243 7704 7288 7732
rect 7282 7692 7288 7704
rect 7340 7692 7346 7744
rect 7437 7732 7465 7772
rect 7742 7760 7748 7812
rect 7800 7800 7806 7812
rect 8220 7800 8248 7831
rect 8294 7828 8300 7880
rect 8352 7868 8358 7880
rect 10873 7871 10931 7877
rect 10873 7868 10885 7871
rect 8352 7840 10885 7868
rect 8352 7828 8358 7840
rect 10873 7837 10885 7840
rect 10919 7868 10931 7871
rect 11606 7868 11612 7880
rect 10919 7840 11612 7868
rect 10919 7837 10931 7840
rect 10873 7831 10931 7837
rect 11606 7828 11612 7840
rect 11664 7828 11670 7880
rect 16485 7871 16543 7877
rect 16485 7837 16497 7871
rect 16531 7868 16543 7871
rect 16531 7840 16941 7868
rect 16531 7837 16543 7840
rect 16485 7831 16543 7837
rect 11422 7800 11428 7812
rect 7800 7772 8248 7800
rect 8772 7772 11428 7800
rect 7800 7760 7806 7772
rect 8772 7732 8800 7772
rect 11422 7760 11428 7772
rect 11480 7760 11486 7812
rect 16913 7800 16941 7840
rect 17126 7828 17132 7880
rect 17184 7868 17190 7880
rect 17405 7871 17463 7877
rect 17405 7868 17417 7871
rect 17184 7840 17417 7868
rect 17184 7828 17190 7840
rect 17405 7837 17417 7840
rect 17451 7837 17463 7871
rect 18230 7868 18236 7880
rect 17405 7831 17463 7837
rect 17696 7840 18236 7868
rect 17696 7800 17724 7840
rect 18230 7828 18236 7840
rect 18288 7868 18294 7880
rect 18325 7871 18383 7877
rect 18325 7868 18337 7871
rect 18288 7840 18337 7868
rect 18288 7828 18294 7840
rect 18325 7837 18337 7840
rect 18371 7837 18383 7871
rect 18325 7831 18383 7837
rect 16913 7772 17724 7800
rect 17957 7803 18015 7809
rect 17957 7769 17969 7803
rect 18003 7800 18015 7803
rect 18414 7800 18420 7812
rect 18003 7772 18420 7800
rect 18003 7769 18015 7772
rect 17957 7763 18015 7769
rect 18414 7760 18420 7772
rect 18472 7760 18478 7812
rect 7437 7704 8800 7732
rect 9858 7692 9864 7744
rect 9916 7732 9922 7744
rect 10686 7732 10692 7744
rect 9916 7704 10692 7732
rect 9916 7692 9922 7704
rect 10686 7692 10692 7704
rect 10744 7692 10750 7744
rect 11790 7732 11796 7744
rect 11751 7704 11796 7732
rect 11790 7692 11796 7704
rect 11848 7732 11854 7744
rect 12437 7735 12495 7741
rect 12437 7732 12449 7735
rect 11848 7704 12449 7732
rect 11848 7692 11854 7704
rect 12437 7701 12449 7704
rect 12483 7732 12495 7735
rect 12618 7732 12624 7744
rect 12483 7704 12624 7732
rect 12483 7701 12495 7704
rect 12437 7695 12495 7701
rect 12618 7692 12624 7704
rect 12676 7692 12682 7744
rect 12710 7692 12716 7744
rect 12768 7732 12774 7744
rect 12805 7735 12863 7741
rect 12805 7732 12817 7735
rect 12768 7704 12817 7732
rect 12768 7692 12774 7704
rect 12805 7701 12817 7704
rect 12851 7701 12863 7735
rect 12805 7695 12863 7701
rect 14553 7735 14611 7741
rect 14553 7701 14565 7735
rect 14599 7732 14611 7735
rect 14642 7732 14648 7744
rect 14599 7704 14648 7732
rect 14599 7701 14611 7704
rect 14553 7695 14611 7701
rect 14642 7692 14648 7704
rect 14700 7692 14706 7744
rect 17126 7732 17132 7744
rect 17087 7704 17132 7732
rect 17126 7692 17132 7704
rect 17184 7692 17190 7744
rect 1104 7642 20884 7664
rect 1104 7590 4648 7642
rect 4700 7590 4712 7642
rect 4764 7590 4776 7642
rect 4828 7590 4840 7642
rect 4892 7590 11982 7642
rect 12034 7590 12046 7642
rect 12098 7590 12110 7642
rect 12162 7590 12174 7642
rect 12226 7590 19315 7642
rect 19367 7590 19379 7642
rect 19431 7590 19443 7642
rect 19495 7590 19507 7642
rect 19559 7590 20884 7642
rect 1104 7568 20884 7590
rect 106 7488 112 7540
rect 164 7528 170 7540
rect 1946 7528 1952 7540
rect 164 7500 1952 7528
rect 164 7488 170 7500
rect 1946 7488 1952 7500
rect 2004 7488 2010 7540
rect 3145 7531 3203 7537
rect 3145 7497 3157 7531
rect 3191 7528 3203 7531
rect 3234 7528 3240 7540
rect 3191 7500 3240 7528
rect 3191 7497 3203 7500
rect 3145 7491 3203 7497
rect 3234 7488 3240 7500
rect 3292 7488 3298 7540
rect 4522 7488 4528 7540
rect 4580 7528 4586 7540
rect 4617 7531 4675 7537
rect 4617 7528 4629 7531
rect 4580 7500 4629 7528
rect 4580 7488 4586 7500
rect 4617 7497 4629 7500
rect 4663 7497 4675 7531
rect 4617 7491 4675 7497
rect 6641 7531 6699 7537
rect 6641 7497 6653 7531
rect 6687 7528 6699 7531
rect 7098 7528 7104 7540
rect 6687 7500 7104 7528
rect 6687 7497 6699 7500
rect 6641 7491 6699 7497
rect 7098 7488 7104 7500
rect 7156 7488 7162 7540
rect 8846 7488 8852 7540
rect 8904 7528 8910 7540
rect 9674 7528 9680 7540
rect 8904 7500 9680 7528
rect 8904 7488 8910 7500
rect 9674 7488 9680 7500
rect 9732 7488 9738 7540
rect 9861 7531 9919 7537
rect 9861 7497 9873 7531
rect 9907 7528 9919 7531
rect 9907 7500 10364 7528
rect 9907 7497 9919 7500
rect 9861 7491 9919 7497
rect 3513 7463 3571 7469
rect 3513 7429 3525 7463
rect 3559 7460 3571 7463
rect 5534 7460 5540 7472
rect 3559 7432 5540 7460
rect 3559 7429 3571 7432
rect 3513 7423 3571 7429
rect 3050 7392 3056 7404
rect 2240 7364 3056 7392
rect 2240 7333 2268 7364
rect 3050 7352 3056 7364
rect 3108 7352 3114 7404
rect 2225 7327 2283 7333
rect 2225 7293 2237 7327
rect 2271 7293 2283 7327
rect 2225 7287 2283 7293
rect 2314 7284 2320 7336
rect 2372 7324 2378 7336
rect 2593 7327 2651 7333
rect 2593 7324 2605 7327
rect 2372 7296 2605 7324
rect 2372 7284 2378 7296
rect 2593 7293 2605 7296
rect 2639 7324 2651 7327
rect 2958 7324 2964 7336
rect 2639 7296 2964 7324
rect 2639 7293 2651 7296
rect 2593 7287 2651 7293
rect 2958 7284 2964 7296
rect 3016 7324 3022 7336
rect 3528 7324 3556 7423
rect 3786 7324 3792 7336
rect 3016 7296 3556 7324
rect 3747 7296 3792 7324
rect 3016 7284 3022 7296
rect 3786 7284 3792 7296
rect 3844 7284 3850 7336
rect 4080 7333 4108 7432
rect 5534 7420 5540 7432
rect 5592 7420 5598 7472
rect 9766 7460 9772 7472
rect 7713 7432 9772 7460
rect 4341 7395 4399 7401
rect 4341 7361 4353 7395
rect 4387 7392 4399 7395
rect 6917 7395 6975 7401
rect 6917 7392 6929 7395
rect 4387 7364 6929 7392
rect 4387 7361 4399 7364
rect 4341 7355 4399 7361
rect 6917 7361 6929 7364
rect 6963 7392 6975 7395
rect 7282 7392 7288 7404
rect 6963 7364 7288 7392
rect 6963 7361 6975 7364
rect 6917 7355 6975 7361
rect 7282 7352 7288 7364
rect 7340 7352 7346 7404
rect 4065 7327 4123 7333
rect 4065 7293 4077 7327
rect 4111 7293 4123 7327
rect 4065 7287 4123 7293
rect 4522 7284 4528 7336
rect 4580 7324 4586 7336
rect 4982 7324 4988 7336
rect 4580 7296 4988 7324
rect 4580 7284 4586 7296
rect 4982 7284 4988 7296
rect 5040 7324 5046 7336
rect 5169 7327 5227 7333
rect 5169 7324 5181 7327
rect 5040 7296 5181 7324
rect 5040 7284 5046 7296
rect 5169 7293 5181 7296
rect 5215 7293 5227 7327
rect 5626 7324 5632 7336
rect 5587 7296 5632 7324
rect 5169 7287 5227 7293
rect 5626 7284 5632 7296
rect 5684 7284 5690 7336
rect 5905 7327 5963 7333
rect 5905 7293 5917 7327
rect 5951 7324 5963 7327
rect 7713 7324 7741 7432
rect 9766 7420 9772 7432
rect 9824 7420 9830 7472
rect 10045 7463 10103 7469
rect 10045 7460 10057 7463
rect 9968 7432 10057 7460
rect 8110 7352 8116 7404
rect 8168 7392 8174 7404
rect 9968 7392 9996 7432
rect 10045 7429 10057 7432
rect 10091 7429 10103 7463
rect 10045 7423 10103 7429
rect 10336 7401 10364 7500
rect 10594 7488 10600 7540
rect 10652 7488 10658 7540
rect 11606 7528 11612 7540
rect 11567 7500 11612 7528
rect 11606 7488 11612 7500
rect 11664 7488 11670 7540
rect 14642 7528 14648 7540
rect 14603 7500 14648 7528
rect 14642 7488 14648 7500
rect 14700 7488 14706 7540
rect 15378 7528 15384 7540
rect 15339 7500 15384 7528
rect 15378 7488 15384 7500
rect 15436 7488 15442 7540
rect 16114 7528 16120 7540
rect 16075 7500 16120 7528
rect 16114 7488 16120 7500
rect 16172 7488 16178 7540
rect 17494 7528 17500 7540
rect 17455 7500 17500 7528
rect 17494 7488 17500 7500
rect 17552 7488 17558 7540
rect 17586 7488 17592 7540
rect 17644 7528 17650 7540
rect 19751 7531 19809 7537
rect 19751 7528 19763 7531
rect 17644 7500 19763 7528
rect 17644 7488 17650 7500
rect 19751 7497 19763 7500
rect 19797 7497 19809 7531
rect 19751 7491 19809 7497
rect 10612 7401 10640 7488
rect 13446 7420 13452 7472
rect 13504 7460 13510 7472
rect 14921 7463 14979 7469
rect 14921 7460 14933 7463
rect 13504 7432 14933 7460
rect 13504 7420 13510 7432
rect 14921 7429 14933 7432
rect 14967 7429 14979 7463
rect 14921 7423 14979 7429
rect 8168 7364 9996 7392
rect 8168 7352 8174 7364
rect 5951 7296 7741 7324
rect 7837 7327 7895 7333
rect 5951 7293 5963 7296
rect 5905 7287 5963 7293
rect 7837 7293 7849 7327
rect 7883 7324 7895 7327
rect 8481 7327 8539 7333
rect 8481 7324 8493 7327
rect 7883 7296 8493 7324
rect 7883 7293 7895 7296
rect 7837 7287 7895 7293
rect 8481 7293 8493 7296
rect 8527 7293 8539 7327
rect 8481 7287 8539 7293
rect 2777 7259 2835 7265
rect 2777 7225 2789 7259
rect 2823 7256 2835 7259
rect 3878 7256 3884 7268
rect 2823 7228 3884 7256
rect 2823 7225 2835 7228
rect 2777 7219 2835 7225
rect 3878 7216 3884 7228
rect 3936 7216 3942 7268
rect 7238 7259 7296 7265
rect 7238 7256 7250 7259
rect 6472 7228 7250 7256
rect 6472 7200 6500 7228
rect 7238 7225 7250 7228
rect 7284 7225 7296 7259
rect 7238 7219 7296 7225
rect 4614 7148 4620 7200
rect 4672 7188 4678 7200
rect 5077 7191 5135 7197
rect 5077 7188 5089 7191
rect 4672 7160 5089 7188
rect 4672 7148 4678 7160
rect 5077 7157 5089 7160
rect 5123 7188 5135 7191
rect 5626 7188 5632 7200
rect 5123 7160 5632 7188
rect 5123 7157 5135 7160
rect 5077 7151 5135 7157
rect 5626 7148 5632 7160
rect 5684 7148 5690 7200
rect 6273 7191 6331 7197
rect 6273 7157 6285 7191
rect 6319 7188 6331 7191
rect 6454 7188 6460 7200
rect 6319 7160 6460 7188
rect 6319 7157 6331 7160
rect 6273 7151 6331 7157
rect 6454 7148 6460 7160
rect 6512 7148 6518 7200
rect 8110 7188 8116 7200
rect 8071 7160 8116 7188
rect 8110 7148 8116 7160
rect 8168 7148 8174 7200
rect 8496 7188 8524 7287
rect 9398 7284 9404 7336
rect 9456 7324 9462 7336
rect 9769 7327 9827 7333
rect 9769 7324 9781 7327
rect 9456 7296 9501 7324
rect 9646 7296 9781 7324
rect 9456 7284 9462 7296
rect 8754 7256 8760 7268
rect 8715 7228 8760 7256
rect 8754 7216 8760 7228
rect 8812 7216 8818 7268
rect 8849 7259 8907 7265
rect 8849 7225 8861 7259
rect 8895 7225 8907 7259
rect 8849 7219 8907 7225
rect 8864 7188 8892 7219
rect 8496 7160 8892 7188
rect 9490 7148 9496 7200
rect 9548 7188 9554 7200
rect 9646 7188 9674 7296
rect 9769 7293 9781 7296
rect 9815 7324 9827 7327
rect 9861 7327 9919 7333
rect 9861 7324 9873 7327
rect 9815 7296 9873 7324
rect 9815 7293 9827 7296
rect 9769 7287 9827 7293
rect 9861 7293 9873 7296
rect 9907 7293 9919 7327
rect 9861 7287 9919 7293
rect 9548 7160 9674 7188
rect 9968 7188 9996 7364
rect 10321 7395 10379 7401
rect 10321 7361 10333 7395
rect 10367 7361 10379 7395
rect 10321 7355 10379 7361
rect 10597 7395 10655 7401
rect 10597 7361 10609 7395
rect 10643 7361 10655 7395
rect 10597 7355 10655 7361
rect 13725 7395 13783 7401
rect 13725 7361 13737 7395
rect 13771 7392 13783 7395
rect 15396 7392 15424 7488
rect 15470 7420 15476 7472
rect 15528 7460 15534 7472
rect 15841 7463 15899 7469
rect 15841 7460 15853 7463
rect 15528 7432 15853 7460
rect 15528 7420 15534 7432
rect 15841 7429 15853 7432
rect 15887 7460 15899 7463
rect 16390 7460 16396 7472
rect 15887 7432 16396 7460
rect 15887 7429 15899 7432
rect 15841 7423 15899 7429
rect 16390 7420 16396 7432
rect 16448 7420 16454 7472
rect 16666 7420 16672 7472
rect 16724 7460 16730 7472
rect 17037 7463 17095 7469
rect 17037 7460 17049 7463
rect 16724 7432 17049 7460
rect 16724 7420 16730 7432
rect 17037 7429 17049 7432
rect 17083 7460 17095 7463
rect 18693 7463 18751 7469
rect 18693 7460 18705 7463
rect 17083 7432 18705 7460
rect 17083 7429 17095 7432
rect 17037 7423 17095 7429
rect 18693 7429 18705 7432
rect 18739 7429 18751 7463
rect 18693 7423 18751 7429
rect 13771 7364 15424 7392
rect 13771 7361 13783 7364
rect 13725 7355 13783 7361
rect 16482 7352 16488 7404
rect 16540 7392 16546 7404
rect 18874 7392 18880 7404
rect 16540 7364 18880 7392
rect 16540 7352 16546 7364
rect 18874 7352 18880 7364
rect 18932 7392 18938 7404
rect 19429 7395 19487 7401
rect 19429 7392 19441 7395
rect 18932 7364 19441 7392
rect 18932 7352 18938 7364
rect 19429 7361 19441 7364
rect 19475 7361 19487 7395
rect 19429 7355 19487 7361
rect 11514 7284 11520 7336
rect 11572 7324 11578 7336
rect 12621 7327 12679 7333
rect 12621 7324 12633 7327
rect 11572 7296 12633 7324
rect 11572 7284 11578 7296
rect 12621 7293 12633 7296
rect 12667 7324 12679 7327
rect 13173 7327 13231 7333
rect 13173 7324 13185 7327
rect 12667 7296 13185 7324
rect 12667 7293 12679 7296
rect 12621 7287 12679 7293
rect 13173 7293 13185 7296
rect 13219 7293 13231 7327
rect 13173 7287 13231 7293
rect 19680 7327 19738 7333
rect 19680 7293 19692 7327
rect 19726 7293 19738 7327
rect 19680 7287 19738 7293
rect 10413 7259 10471 7265
rect 10413 7225 10425 7259
rect 10459 7225 10471 7259
rect 11330 7256 11336 7268
rect 11243 7228 11336 7256
rect 10413 7219 10471 7225
rect 10428 7188 10456 7219
rect 11330 7216 11336 7228
rect 11388 7256 11394 7268
rect 14046 7259 14104 7265
rect 14046 7256 14058 7259
rect 11388 7228 14058 7256
rect 11388 7216 11394 7228
rect 13556 7200 13584 7228
rect 14046 7225 14058 7228
rect 14092 7225 14104 7259
rect 14046 7219 14104 7225
rect 14366 7216 14372 7268
rect 14424 7256 14430 7268
rect 16485 7259 16543 7265
rect 16485 7256 16497 7259
rect 14424 7228 16497 7256
rect 14424 7216 14430 7228
rect 16485 7225 16497 7228
rect 16531 7225 16543 7259
rect 16485 7219 16543 7225
rect 12802 7188 12808 7200
rect 9968 7160 10456 7188
rect 12763 7160 12808 7188
rect 9548 7148 9554 7160
rect 12802 7148 12808 7160
rect 12860 7148 12866 7200
rect 13538 7188 13544 7200
rect 13499 7160 13544 7188
rect 13538 7148 13544 7160
rect 13596 7148 13602 7200
rect 16500 7188 16528 7219
rect 16574 7216 16580 7268
rect 16632 7256 16638 7268
rect 18138 7256 18144 7268
rect 16632 7228 16677 7256
rect 18099 7228 18144 7256
rect 16632 7216 16638 7228
rect 18138 7216 18144 7228
rect 18196 7216 18202 7268
rect 18233 7259 18291 7265
rect 18233 7225 18245 7259
rect 18279 7225 18291 7259
rect 18233 7219 18291 7225
rect 17034 7188 17040 7200
rect 16500 7160 17040 7188
rect 17034 7148 17040 7160
rect 17092 7148 17098 7200
rect 17865 7191 17923 7197
rect 17865 7157 17877 7191
rect 17911 7188 17923 7191
rect 18248 7188 18276 7219
rect 18322 7216 18328 7268
rect 18380 7256 18386 7268
rect 18380 7228 19334 7256
rect 18380 7216 18386 7228
rect 18506 7188 18512 7200
rect 17911 7160 18512 7188
rect 17911 7157 17923 7160
rect 17865 7151 17923 7157
rect 18506 7148 18512 7160
rect 18564 7148 18570 7200
rect 19058 7188 19064 7200
rect 19019 7160 19064 7188
rect 19058 7148 19064 7160
rect 19116 7148 19122 7200
rect 19306 7188 19334 7228
rect 19695 7200 19723 7287
rect 19695 7188 19708 7200
rect 19306 7160 19708 7188
rect 19702 7148 19708 7160
rect 19760 7188 19766 7200
rect 20073 7191 20131 7197
rect 20073 7188 20085 7191
rect 19760 7160 20085 7188
rect 19760 7148 19766 7160
rect 20073 7157 20085 7160
rect 20119 7157 20131 7191
rect 20073 7151 20131 7157
rect 1104 7098 20884 7120
rect 1104 7046 8315 7098
rect 8367 7046 8379 7098
rect 8431 7046 8443 7098
rect 8495 7046 8507 7098
rect 8559 7046 15648 7098
rect 15700 7046 15712 7098
rect 15764 7046 15776 7098
rect 15828 7046 15840 7098
rect 15892 7046 20884 7098
rect 1104 7024 20884 7046
rect 1535 6987 1593 6993
rect 1535 6953 1547 6987
rect 1581 6984 1593 6987
rect 7469 6987 7527 6993
rect 1581 6956 7420 6984
rect 1581 6953 1593 6956
rect 1535 6947 1593 6953
rect 2314 6916 2320 6928
rect 2275 6888 2320 6916
rect 2314 6876 2320 6888
rect 2372 6876 2378 6928
rect 3697 6919 3755 6925
rect 3697 6885 3709 6919
rect 3743 6916 3755 6919
rect 3786 6916 3792 6928
rect 3743 6888 3792 6916
rect 3743 6885 3755 6888
rect 3697 6879 3755 6885
rect 3786 6876 3792 6888
rect 3844 6876 3850 6928
rect 4062 6876 4068 6928
rect 4120 6916 4126 6928
rect 5997 6919 6055 6925
rect 5997 6916 6009 6919
rect 4120 6888 6009 6916
rect 4120 6876 4126 6888
rect 5997 6885 6009 6888
rect 6043 6885 6055 6919
rect 5997 6879 6055 6885
rect 6454 6876 6460 6928
rect 6512 6916 6518 6928
rect 6870 6919 6928 6925
rect 6870 6916 6882 6919
rect 6512 6888 6882 6916
rect 6512 6876 6518 6888
rect 6870 6885 6882 6888
rect 6916 6885 6928 6919
rect 7392 6916 7420 6956
rect 7469 6953 7481 6987
rect 7515 6984 7527 6987
rect 8110 6984 8116 6996
rect 7515 6956 8116 6984
rect 7515 6953 7527 6956
rect 7469 6947 7527 6953
rect 8110 6944 8116 6956
rect 8168 6944 8174 6996
rect 8711 6987 8769 6993
rect 8711 6953 8723 6987
rect 8757 6984 8769 6987
rect 10962 6984 10968 6996
rect 8757 6956 10968 6984
rect 8757 6953 8769 6956
rect 8711 6947 8769 6953
rect 10962 6944 10968 6956
rect 11020 6944 11026 6996
rect 11054 6944 11060 6996
rect 11112 6984 11118 6996
rect 11330 6984 11336 6996
rect 11112 6956 11336 6984
rect 11112 6944 11118 6956
rect 11330 6944 11336 6956
rect 11388 6984 11394 6996
rect 16482 6984 16488 6996
rect 11388 6956 16488 6984
rect 11388 6944 11394 6956
rect 16482 6944 16488 6956
rect 16540 6944 16546 6996
rect 16574 6944 16580 6996
rect 16632 6984 16638 6996
rect 16761 6987 16819 6993
rect 16761 6984 16773 6987
rect 16632 6956 16773 6984
rect 16632 6944 16638 6956
rect 16761 6953 16773 6956
rect 16807 6953 16819 6987
rect 17034 6984 17040 6996
rect 16995 6956 17040 6984
rect 16761 6947 16819 6953
rect 17034 6944 17040 6956
rect 17092 6944 17098 6996
rect 19518 6984 19524 6996
rect 19479 6956 19524 6984
rect 19518 6944 19524 6956
rect 19576 6944 19582 6996
rect 8938 6916 8944 6928
rect 7392 6888 8944 6916
rect 6870 6879 6928 6885
rect 8938 6876 8944 6888
rect 8996 6916 9002 6928
rect 9033 6919 9091 6925
rect 9033 6916 9045 6919
rect 8996 6888 9045 6916
rect 8996 6876 9002 6888
rect 9033 6885 9045 6888
rect 9079 6885 9091 6919
rect 9033 6879 9091 6885
rect 11422 6876 11428 6928
rect 11480 6916 11486 6928
rect 11609 6919 11667 6925
rect 11609 6916 11621 6919
rect 11480 6888 11621 6916
rect 11480 6876 11486 6888
rect 11609 6885 11621 6888
rect 11655 6885 11667 6919
rect 11609 6879 11667 6885
rect 11701 6919 11759 6925
rect 11701 6885 11713 6919
rect 11747 6916 11759 6919
rect 11790 6916 11796 6928
rect 11747 6888 11796 6916
rect 11747 6885 11759 6888
rect 11701 6879 11759 6885
rect 11790 6876 11796 6888
rect 11848 6876 11854 6928
rect 12253 6919 12311 6925
rect 12253 6885 12265 6919
rect 12299 6916 12311 6919
rect 12342 6916 12348 6928
rect 12299 6888 12348 6916
rect 12299 6885 12311 6888
rect 12253 6879 12311 6885
rect 12342 6876 12348 6888
rect 12400 6876 12406 6928
rect 14369 6919 14427 6925
rect 14369 6885 14381 6919
rect 14415 6916 14427 6919
rect 15470 6916 15476 6928
rect 14415 6888 15476 6916
rect 14415 6885 14427 6888
rect 14369 6879 14427 6885
rect 15470 6876 15476 6888
rect 15528 6876 15534 6928
rect 16203 6919 16261 6925
rect 16203 6885 16215 6919
rect 16249 6885 16261 6919
rect 16203 6879 16261 6885
rect 17910 6919 17968 6925
rect 17910 6885 17922 6919
rect 17956 6885 17968 6919
rect 17910 6879 17968 6885
rect 1464 6851 1522 6857
rect 1464 6817 1476 6851
rect 1510 6848 1522 6851
rect 2498 6848 2504 6860
rect 1510 6820 1900 6848
rect 2459 6820 2504 6848
rect 1510 6817 1522 6820
rect 1464 6811 1522 6817
rect 1872 6653 1900 6820
rect 2498 6808 2504 6820
rect 2556 6808 2562 6860
rect 2866 6848 2872 6860
rect 2827 6820 2872 6848
rect 2866 6808 2872 6820
rect 2924 6808 2930 6860
rect 5258 6848 5264 6860
rect 5219 6820 5264 6848
rect 5258 6808 5264 6820
rect 5316 6808 5322 6860
rect 5537 6851 5595 6857
rect 5537 6817 5549 6851
rect 5583 6848 5595 6851
rect 5626 6848 5632 6860
rect 5583 6820 5632 6848
rect 5583 6817 5595 6820
rect 5537 6811 5595 6817
rect 5626 6808 5632 6820
rect 5684 6808 5690 6860
rect 5721 6851 5779 6857
rect 5721 6817 5733 6851
rect 5767 6848 5779 6851
rect 8202 6848 8208 6860
rect 5767 6820 8208 6848
rect 5767 6817 5779 6820
rect 5721 6811 5779 6817
rect 8202 6808 8208 6820
rect 8260 6808 8266 6860
rect 8640 6851 8698 6857
rect 8640 6817 8652 6851
rect 8686 6848 8698 6851
rect 8754 6848 8760 6860
rect 8686 6820 8760 6848
rect 8686 6817 8698 6820
rect 8640 6811 8698 6817
rect 8754 6808 8760 6820
rect 8812 6808 8818 6860
rect 9953 6851 10011 6857
rect 9953 6817 9965 6851
rect 9999 6817 10011 6851
rect 9953 6811 10011 6817
rect 3142 6780 3148 6792
rect 3103 6752 3148 6780
rect 3142 6740 3148 6752
rect 3200 6740 3206 6792
rect 3878 6740 3884 6792
rect 3936 6780 3942 6792
rect 6549 6783 6607 6789
rect 6549 6780 6561 6783
rect 3936 6752 6561 6780
rect 3936 6740 3942 6752
rect 6549 6749 6561 6752
rect 6595 6780 6607 6783
rect 7374 6780 7380 6792
rect 6595 6752 7380 6780
rect 6595 6749 6607 6752
rect 6549 6743 6607 6749
rect 7374 6740 7380 6752
rect 7432 6740 7438 6792
rect 7926 6780 7932 6792
rect 7887 6752 7932 6780
rect 7926 6740 7932 6752
rect 7984 6740 7990 6792
rect 1946 6672 1952 6724
rect 2004 6712 2010 6724
rect 9401 6715 9459 6721
rect 9401 6712 9413 6715
rect 2004 6684 9413 6712
rect 2004 6672 2010 6684
rect 9401 6681 9413 6684
rect 9447 6712 9459 6715
rect 9766 6712 9772 6724
rect 9447 6684 9772 6712
rect 9447 6681 9459 6684
rect 9401 6675 9459 6681
rect 9766 6672 9772 6684
rect 9824 6672 9830 6724
rect 9968 6656 9996 6811
rect 10134 6808 10140 6860
rect 10192 6848 10198 6860
rect 10229 6851 10287 6857
rect 10229 6848 10241 6851
rect 10192 6820 10241 6848
rect 10192 6808 10198 6820
rect 10229 6817 10241 6820
rect 10275 6817 10287 6851
rect 10229 6811 10287 6817
rect 12526 6808 12532 6860
rect 12584 6848 12590 6860
rect 13446 6848 13452 6860
rect 12584 6820 13452 6848
rect 12584 6808 12590 6820
rect 13446 6808 13452 6820
rect 13504 6848 13510 6860
rect 13633 6851 13691 6857
rect 13633 6848 13645 6851
rect 13504 6820 13645 6848
rect 13504 6808 13510 6820
rect 13633 6817 13645 6820
rect 13679 6817 13691 6851
rect 13633 6811 13691 6817
rect 13909 6851 13967 6857
rect 13909 6817 13921 6851
rect 13955 6817 13967 6851
rect 16218 6848 16246 6879
rect 16574 6848 16580 6860
rect 16218 6820 16580 6848
rect 13909 6811 13967 6817
rect 10502 6780 10508 6792
rect 10463 6752 10508 6780
rect 10502 6740 10508 6752
rect 10560 6740 10566 6792
rect 13170 6740 13176 6792
rect 13228 6780 13234 6792
rect 13924 6780 13952 6811
rect 16574 6808 16580 6820
rect 16632 6848 16638 6860
rect 16942 6848 16948 6860
rect 16632 6820 16948 6848
rect 16632 6808 16638 6820
rect 16942 6808 16948 6820
rect 17000 6848 17006 6860
rect 17925 6848 17953 6879
rect 17000 6820 17953 6848
rect 17000 6808 17006 6820
rect 18046 6808 18052 6860
rect 18104 6848 18110 6860
rect 19150 6848 19156 6860
rect 18104 6820 19156 6848
rect 18104 6808 18110 6820
rect 19150 6808 19156 6820
rect 19208 6848 19214 6860
rect 19337 6851 19395 6857
rect 19337 6848 19349 6851
rect 19208 6820 19349 6848
rect 19208 6808 19214 6820
rect 19337 6817 19349 6820
rect 19383 6817 19395 6851
rect 19337 6811 19395 6817
rect 13228 6752 13952 6780
rect 13228 6740 13234 6752
rect 15010 6740 15016 6792
rect 15068 6780 15074 6792
rect 15841 6783 15899 6789
rect 15841 6780 15853 6783
rect 15068 6752 15853 6780
rect 15068 6740 15074 6752
rect 15841 6749 15853 6752
rect 15887 6749 15899 6783
rect 17589 6783 17647 6789
rect 17589 6780 17601 6783
rect 15841 6743 15899 6749
rect 17420 6752 17601 6780
rect 10042 6672 10048 6724
rect 10100 6712 10106 6724
rect 13722 6712 13728 6724
rect 10100 6684 10145 6712
rect 13683 6684 13728 6712
rect 10100 6672 10106 6684
rect 13722 6672 13728 6684
rect 13780 6672 13786 6724
rect 1857 6647 1915 6653
rect 1857 6613 1869 6647
rect 1903 6644 1915 6647
rect 2038 6644 2044 6656
rect 1903 6616 2044 6644
rect 1903 6613 1915 6616
rect 1857 6607 1915 6613
rect 2038 6604 2044 6616
rect 2096 6604 2102 6656
rect 3970 6604 3976 6656
rect 4028 6644 4034 6656
rect 4249 6647 4307 6653
rect 4249 6644 4261 6647
rect 4028 6616 4261 6644
rect 4028 6604 4034 6616
rect 4249 6613 4261 6616
rect 4295 6613 4307 6647
rect 4249 6607 4307 6613
rect 4430 6604 4436 6656
rect 4488 6644 4494 6656
rect 4617 6647 4675 6653
rect 4617 6644 4629 6647
rect 4488 6616 4629 6644
rect 4488 6604 4494 6616
rect 4617 6613 4629 6616
rect 4663 6613 4675 6647
rect 4617 6607 4675 6613
rect 5166 6604 5172 6656
rect 5224 6644 5230 6656
rect 9950 6644 9956 6656
rect 5224 6616 9956 6644
rect 5224 6604 5230 6616
rect 9950 6604 9956 6616
rect 10008 6604 10014 6656
rect 10962 6644 10968 6656
rect 10923 6616 10968 6644
rect 10962 6604 10968 6616
rect 11020 6604 11026 6656
rect 13357 6647 13415 6653
rect 13357 6613 13369 6647
rect 13403 6644 13415 6647
rect 13538 6644 13544 6656
rect 13403 6616 13544 6644
rect 13403 6613 13415 6616
rect 13357 6607 13415 6613
rect 13538 6604 13544 6616
rect 13596 6604 13602 6656
rect 17310 6604 17316 6656
rect 17368 6644 17374 6656
rect 17420 6653 17448 6752
rect 17589 6749 17601 6752
rect 17635 6749 17647 6783
rect 17589 6743 17647 6749
rect 17405 6647 17463 6653
rect 17405 6644 17417 6647
rect 17368 6616 17417 6644
rect 17368 6604 17374 6616
rect 17405 6613 17417 6616
rect 17451 6613 17463 6647
rect 18506 6644 18512 6656
rect 18467 6616 18512 6644
rect 17405 6607 17463 6613
rect 18506 6604 18512 6616
rect 18564 6604 18570 6656
rect 1104 6554 20884 6576
rect 1104 6502 4648 6554
rect 4700 6502 4712 6554
rect 4764 6502 4776 6554
rect 4828 6502 4840 6554
rect 4892 6502 11982 6554
rect 12034 6502 12046 6554
rect 12098 6502 12110 6554
rect 12162 6502 12174 6554
rect 12226 6502 19315 6554
rect 19367 6502 19379 6554
rect 19431 6502 19443 6554
rect 19495 6502 19507 6554
rect 19559 6502 20884 6554
rect 1104 6480 20884 6502
rect 2869 6443 2927 6449
rect 2869 6409 2881 6443
rect 2915 6440 2927 6443
rect 3513 6443 3571 6449
rect 3513 6440 3525 6443
rect 2915 6412 3525 6440
rect 2915 6409 2927 6412
rect 2869 6403 2927 6409
rect 3513 6409 3525 6412
rect 3559 6440 3571 6443
rect 6270 6440 6276 6452
rect 3559 6412 6276 6440
rect 3559 6409 3571 6412
rect 3513 6403 3571 6409
rect 6270 6400 6276 6412
rect 6328 6400 6334 6452
rect 6730 6400 6736 6452
rect 6788 6440 6794 6452
rect 8021 6443 8079 6449
rect 8021 6440 8033 6443
rect 6788 6412 8033 6440
rect 6788 6400 6794 6412
rect 8021 6409 8033 6412
rect 8067 6440 8079 6443
rect 8110 6440 8116 6452
rect 8067 6412 8116 6440
rect 8067 6409 8079 6412
rect 8021 6403 8079 6409
rect 8110 6400 8116 6412
rect 8168 6400 8174 6452
rect 9950 6400 9956 6452
rect 10008 6440 10014 6452
rect 11517 6443 11575 6449
rect 11517 6440 11529 6443
rect 10008 6412 11529 6440
rect 10008 6400 10014 6412
rect 11517 6409 11529 6412
rect 11563 6440 11575 6443
rect 11606 6440 11612 6452
rect 11563 6412 11612 6440
rect 11563 6409 11575 6412
rect 11517 6403 11575 6409
rect 11606 6400 11612 6412
rect 11664 6400 11670 6452
rect 11790 6440 11796 6452
rect 11751 6412 11796 6440
rect 11790 6400 11796 6412
rect 11848 6400 11854 6452
rect 13446 6400 13452 6452
rect 13504 6440 13510 6452
rect 14369 6443 14427 6449
rect 14369 6440 14381 6443
rect 13504 6412 14381 6440
rect 13504 6400 13510 6412
rect 14369 6409 14381 6412
rect 14415 6409 14427 6443
rect 15470 6440 15476 6452
rect 15431 6412 15476 6440
rect 14369 6403 14427 6409
rect 15470 6400 15476 6412
rect 15528 6400 15534 6452
rect 19150 6400 19156 6452
rect 19208 6440 19214 6452
rect 19337 6443 19395 6449
rect 19337 6440 19349 6443
rect 19208 6412 19349 6440
rect 19208 6400 19214 6412
rect 19337 6409 19349 6412
rect 19383 6409 19395 6443
rect 19337 6403 19395 6409
rect 19610 6400 19616 6452
rect 19668 6440 19674 6452
rect 19751 6443 19809 6449
rect 19751 6440 19763 6443
rect 19668 6412 19763 6440
rect 19668 6400 19674 6412
rect 19751 6409 19763 6412
rect 19797 6409 19809 6443
rect 19751 6403 19809 6409
rect 1949 6375 2007 6381
rect 1949 6341 1961 6375
rect 1995 6372 2007 6375
rect 2133 6375 2191 6381
rect 2133 6372 2145 6375
rect 1995 6344 2145 6372
rect 1995 6341 2007 6344
rect 1949 6335 2007 6341
rect 2133 6341 2145 6344
rect 2179 6372 2191 6375
rect 4246 6372 4252 6384
rect 2179 6344 4252 6372
rect 2179 6341 2191 6344
rect 2133 6335 2191 6341
rect 4246 6332 4252 6344
rect 4304 6372 4310 6384
rect 10042 6372 10048 6384
rect 4304 6344 10048 6372
rect 4304 6332 4310 6344
rect 10042 6332 10048 6344
rect 10100 6332 10106 6384
rect 11422 6332 11428 6384
rect 11480 6372 11486 6384
rect 12161 6375 12219 6381
rect 12161 6372 12173 6375
rect 11480 6344 12173 6372
rect 11480 6332 11486 6344
rect 12161 6341 12173 6344
rect 12207 6341 12219 6375
rect 12161 6335 12219 6341
rect 2869 6307 2927 6313
rect 2869 6304 2881 6307
rect 2056 6276 2881 6304
rect 2056 6245 2084 6276
rect 2869 6273 2881 6276
rect 2915 6273 2927 6307
rect 2869 6267 2927 6273
rect 2958 6264 2964 6316
rect 3016 6304 3022 6316
rect 3970 6304 3976 6316
rect 3016 6276 3976 6304
rect 3016 6264 3022 6276
rect 3970 6264 3976 6276
rect 4028 6304 4034 6316
rect 4341 6307 4399 6313
rect 4028 6276 4108 6304
rect 4028 6264 4034 6276
rect 2041 6239 2099 6245
rect 2041 6205 2053 6239
rect 2087 6205 2099 6239
rect 2041 6199 2099 6205
rect 2317 6239 2375 6245
rect 2317 6205 2329 6239
rect 2363 6205 2375 6239
rect 2317 6199 2375 6205
rect 2332 6168 2360 6199
rect 3234 6196 3240 6248
rect 3292 6236 3298 6248
rect 3878 6236 3884 6248
rect 3292 6208 3884 6236
rect 3292 6196 3298 6208
rect 3878 6196 3884 6208
rect 3936 6196 3942 6248
rect 4080 6245 4108 6276
rect 4341 6273 4353 6307
rect 4387 6304 4399 6307
rect 9030 6304 9036 6316
rect 4387 6276 9036 6304
rect 4387 6273 4399 6276
rect 4341 6267 4399 6273
rect 9030 6264 9036 6276
rect 9088 6264 9094 6316
rect 9950 6264 9956 6316
rect 10008 6304 10014 6316
rect 10781 6307 10839 6313
rect 10781 6304 10793 6307
rect 10008 6276 10793 6304
rect 10008 6264 10014 6276
rect 10781 6273 10793 6276
rect 10827 6273 10839 6307
rect 15010 6304 15016 6316
rect 14971 6276 15016 6304
rect 10781 6267 10839 6273
rect 15010 6264 15016 6276
rect 15068 6264 15074 6316
rect 15488 6304 15516 6400
rect 16022 6332 16028 6384
rect 16080 6372 16086 6384
rect 20073 6375 20131 6381
rect 20073 6372 20085 6375
rect 16080 6344 20085 6372
rect 16080 6332 16086 6344
rect 16298 6304 16304 6316
rect 15488 6276 16068 6304
rect 16259 6276 16304 6304
rect 4065 6239 4123 6245
rect 4065 6205 4077 6239
rect 4111 6205 4123 6239
rect 4065 6199 4123 6205
rect 4525 6239 4583 6245
rect 4525 6205 4537 6239
rect 4571 6236 4583 6239
rect 5077 6239 5135 6245
rect 5077 6236 5089 6239
rect 4571 6208 5089 6236
rect 4571 6205 4583 6208
rect 4525 6199 4583 6205
rect 5077 6205 5089 6208
rect 5123 6236 5135 6239
rect 5813 6239 5871 6245
rect 5813 6236 5825 6239
rect 5123 6208 5825 6236
rect 5123 6205 5135 6208
rect 5077 6199 5135 6205
rect 5813 6205 5825 6208
rect 5859 6205 5871 6239
rect 6178 6236 6184 6248
rect 6139 6208 6184 6236
rect 5813 6199 5871 6205
rect 3145 6171 3203 6177
rect 3145 6168 3157 6171
rect 2332 6140 3157 6168
rect 3145 6137 3157 6140
rect 3191 6168 3203 6171
rect 5828 6168 5856 6199
rect 6178 6196 6184 6208
rect 6236 6236 6242 6248
rect 6825 6239 6883 6245
rect 6825 6236 6837 6239
rect 6236 6208 6837 6236
rect 6236 6196 6242 6208
rect 6825 6205 6837 6208
rect 6871 6205 6883 6239
rect 7282 6236 7288 6248
rect 7243 6208 7288 6236
rect 6825 6199 6883 6205
rect 7282 6196 7288 6208
rect 7340 6196 7346 6248
rect 10045 6239 10103 6245
rect 10045 6205 10057 6239
rect 10091 6236 10103 6239
rect 10134 6236 10140 6248
rect 10091 6208 10140 6236
rect 10091 6205 10103 6208
rect 10045 6199 10103 6205
rect 10134 6196 10140 6208
rect 10192 6196 10198 6248
rect 12342 6196 12348 6248
rect 12400 6236 12406 6248
rect 13265 6239 13323 6245
rect 13265 6236 13277 6239
rect 12400 6208 13277 6236
rect 12400 6196 12406 6208
rect 13265 6205 13277 6208
rect 13311 6236 13323 6239
rect 14001 6239 14059 6245
rect 14001 6236 14013 6239
rect 13311 6208 14013 6236
rect 13311 6205 13323 6208
rect 13265 6199 13323 6205
rect 14001 6205 14013 6208
rect 14047 6236 14059 6239
rect 15102 6236 15108 6248
rect 14047 6208 15108 6236
rect 14047 6205 14059 6208
rect 14001 6199 14059 6205
rect 15102 6196 15108 6208
rect 15160 6196 15166 6248
rect 15470 6196 15476 6248
rect 15528 6236 15534 6248
rect 16040 6245 16068 6276
rect 16298 6264 16304 6276
rect 16356 6264 16362 6316
rect 18414 6304 18420 6316
rect 18375 6276 18420 6304
rect 18414 6264 18420 6276
rect 18472 6264 18478 6316
rect 15565 6239 15623 6245
rect 15565 6236 15577 6239
rect 15528 6208 15577 6236
rect 15528 6196 15534 6208
rect 15565 6205 15577 6208
rect 15611 6205 15623 6239
rect 15565 6199 15623 6205
rect 16025 6239 16083 6245
rect 16025 6205 16037 6239
rect 16071 6236 16083 6239
rect 17494 6236 17500 6248
rect 16071 6208 17500 6236
rect 16071 6205 16083 6208
rect 16025 6199 16083 6205
rect 17494 6196 17500 6208
rect 17552 6196 17558 6248
rect 19679 6245 19707 6344
rect 20073 6341 20085 6344
rect 20119 6341 20131 6375
rect 20073 6335 20131 6341
rect 19664 6239 19722 6245
rect 19664 6205 19676 6239
rect 19710 6205 19722 6239
rect 19664 6199 19722 6205
rect 6362 6168 6368 6180
rect 3191 6140 5488 6168
rect 5828 6140 6368 6168
rect 3191 6137 3203 6140
rect 3145 6131 3203 6137
rect 5460 6112 5488 6140
rect 6362 6128 6368 6140
rect 6420 6128 6426 6180
rect 7466 6128 7472 6180
rect 7524 6168 7530 6180
rect 7561 6171 7619 6177
rect 7561 6168 7573 6171
rect 7524 6140 7573 6168
rect 7524 6128 7530 6140
rect 7561 6137 7573 6140
rect 7607 6137 7619 6171
rect 8938 6168 8944 6180
rect 8899 6140 8944 6168
rect 7561 6131 7619 6137
rect 8938 6128 8944 6140
rect 8996 6128 9002 6180
rect 9042 6171 9100 6177
rect 9042 6137 9054 6171
rect 9088 6168 9100 6171
rect 9582 6168 9588 6180
rect 9088 6140 9168 6168
rect 9543 6140 9588 6168
rect 9088 6137 9100 6140
rect 9042 6131 9100 6137
rect 2314 6060 2320 6112
rect 2372 6100 2378 6112
rect 2501 6103 2559 6109
rect 2501 6100 2513 6103
rect 2372 6072 2513 6100
rect 2372 6060 2378 6072
rect 2501 6069 2513 6072
rect 2547 6069 2559 6103
rect 2501 6063 2559 6069
rect 3326 6060 3332 6112
rect 3384 6100 3390 6112
rect 4525 6103 4583 6109
rect 4525 6100 4537 6103
rect 3384 6072 4537 6100
rect 3384 6060 3390 6072
rect 4525 6069 4537 6072
rect 4571 6069 4583 6103
rect 4525 6063 4583 6069
rect 4614 6060 4620 6112
rect 4672 6100 4678 6112
rect 5442 6100 5448 6112
rect 4672 6072 4717 6100
rect 5403 6072 5448 6100
rect 4672 6060 4678 6072
rect 5442 6060 5448 6072
rect 5500 6060 5506 6112
rect 6454 6060 6460 6112
rect 6512 6100 6518 6112
rect 6641 6103 6699 6109
rect 6641 6100 6653 6103
rect 6512 6072 6653 6100
rect 6512 6060 6518 6072
rect 6641 6069 6653 6072
rect 6687 6100 6699 6103
rect 7834 6100 7840 6112
rect 6687 6072 7840 6100
rect 6687 6069 6699 6072
rect 6641 6063 6699 6069
rect 7834 6060 7840 6072
rect 7892 6060 7898 6112
rect 8665 6103 8723 6109
rect 8665 6069 8677 6103
rect 8711 6100 8723 6103
rect 8754 6100 8760 6112
rect 8711 6072 8760 6100
rect 8711 6069 8723 6072
rect 8665 6063 8723 6069
rect 8754 6060 8760 6072
rect 8812 6060 8818 6112
rect 9140 6100 9168 6140
rect 9582 6128 9588 6140
rect 9640 6128 9646 6180
rect 10502 6168 10508 6180
rect 9692 6140 10088 6168
rect 10463 6140 10508 6168
rect 9398 6100 9404 6112
rect 9140 6072 9404 6100
rect 9398 6060 9404 6072
rect 9456 6100 9462 6112
rect 9692 6100 9720 6140
rect 9456 6072 9720 6100
rect 10060 6100 10088 6140
rect 10502 6128 10508 6140
rect 10560 6128 10566 6180
rect 10597 6171 10655 6177
rect 10597 6137 10609 6171
rect 10643 6168 10655 6171
rect 10962 6168 10968 6180
rect 10643 6140 10968 6168
rect 10643 6137 10655 6140
rect 10597 6131 10655 6137
rect 10612 6100 10640 6131
rect 10962 6128 10968 6140
rect 11020 6128 11026 6180
rect 12526 6128 12532 6180
rect 12584 6168 12590 6180
rect 13357 6171 13415 6177
rect 13357 6168 13369 6171
rect 12584 6140 13369 6168
rect 12584 6128 12590 6140
rect 13357 6137 13369 6140
rect 13403 6168 13415 6171
rect 13722 6168 13728 6180
rect 13403 6140 13728 6168
rect 13403 6137 13415 6140
rect 13357 6131 13415 6137
rect 13722 6128 13728 6140
rect 13780 6168 13786 6180
rect 14182 6168 14188 6180
rect 13780 6140 14188 6168
rect 13780 6128 13786 6140
rect 14182 6128 14188 6140
rect 14240 6128 14246 6180
rect 17313 6171 17371 6177
rect 17313 6137 17325 6171
rect 17359 6168 17371 6171
rect 18138 6168 18144 6180
rect 17359 6140 17953 6168
rect 18099 6140 18144 6168
rect 17359 6137 17371 6140
rect 17313 6131 17371 6137
rect 10060 6072 10640 6100
rect 12897 6103 12955 6109
rect 9456 6060 9462 6072
rect 12897 6069 12909 6103
rect 12943 6100 12955 6103
rect 13170 6100 13176 6112
rect 12943 6072 13176 6100
rect 12943 6069 12955 6072
rect 12897 6063 12955 6069
rect 13170 6060 13176 6072
rect 13228 6060 13234 6112
rect 16574 6100 16580 6112
rect 16535 6072 16580 6100
rect 16574 6060 16580 6072
rect 16632 6100 16638 6112
rect 17589 6103 17647 6109
rect 17589 6100 17601 6103
rect 16632 6072 17601 6100
rect 16632 6060 16638 6072
rect 17589 6069 17601 6072
rect 17635 6069 17647 6103
rect 17925 6100 17953 6140
rect 18138 6128 18144 6140
rect 18196 6128 18202 6180
rect 18233 6171 18291 6177
rect 18233 6137 18245 6171
rect 18279 6168 18291 6171
rect 18506 6168 18512 6180
rect 18279 6140 18512 6168
rect 18279 6137 18291 6140
rect 18233 6131 18291 6137
rect 18248 6100 18276 6131
rect 18506 6128 18512 6140
rect 18564 6128 18570 6180
rect 17925 6072 18276 6100
rect 17589 6063 17647 6069
rect 1104 6010 20884 6032
rect 1104 5958 8315 6010
rect 8367 5958 8379 6010
rect 8431 5958 8443 6010
rect 8495 5958 8507 6010
rect 8559 5958 15648 6010
rect 15700 5958 15712 6010
rect 15764 5958 15776 6010
rect 15828 5958 15840 6010
rect 15892 5958 20884 6010
rect 1104 5936 20884 5958
rect 4338 5856 4344 5908
rect 4396 5896 4402 5908
rect 4801 5899 4859 5905
rect 4801 5896 4813 5899
rect 4396 5868 4813 5896
rect 4396 5856 4402 5868
rect 4801 5865 4813 5868
rect 4847 5865 4859 5899
rect 4801 5859 4859 5865
rect 5258 5856 5264 5908
rect 5316 5896 5322 5908
rect 5721 5899 5779 5905
rect 5721 5896 5733 5899
rect 5316 5868 5733 5896
rect 5316 5856 5322 5868
rect 5721 5865 5733 5868
rect 5767 5865 5779 5899
rect 6546 5896 6552 5908
rect 6507 5868 6552 5896
rect 5721 5859 5779 5865
rect 6546 5856 6552 5868
rect 6604 5856 6610 5908
rect 7009 5899 7067 5905
rect 7009 5865 7021 5899
rect 7055 5896 7067 5899
rect 7282 5896 7288 5908
rect 7055 5868 7288 5896
rect 7055 5865 7067 5868
rect 7009 5859 7067 5865
rect 7282 5856 7288 5868
rect 7340 5856 7346 5908
rect 7374 5856 7380 5908
rect 7432 5896 7438 5908
rect 7834 5896 7840 5908
rect 7432 5868 7477 5896
rect 7795 5868 7840 5896
rect 7432 5856 7438 5868
rect 7834 5856 7840 5868
rect 7892 5856 7898 5908
rect 9122 5856 9128 5908
rect 9180 5896 9186 5908
rect 9217 5899 9275 5905
rect 9217 5896 9229 5899
rect 9180 5868 9229 5896
rect 9180 5856 9186 5868
rect 9217 5865 9229 5868
rect 9263 5865 9275 5899
rect 9217 5859 9275 5865
rect 10042 5856 10048 5908
rect 10100 5896 10106 5908
rect 10689 5899 10747 5905
rect 10689 5896 10701 5899
rect 10100 5868 10701 5896
rect 10100 5856 10106 5868
rect 10689 5865 10701 5868
rect 10735 5865 10747 5899
rect 14001 5899 14059 5905
rect 14001 5896 14013 5899
rect 10689 5859 10747 5865
rect 12084 5868 14013 5896
rect 1535 5831 1593 5837
rect 1535 5797 1547 5831
rect 1581 5828 1593 5831
rect 1581 5800 9260 5828
rect 1581 5797 1593 5800
rect 1535 5791 1593 5797
rect 1448 5763 1506 5769
rect 1448 5729 1460 5763
rect 1494 5760 1506 5763
rect 1857 5763 1915 5769
rect 1857 5760 1869 5763
rect 1494 5732 1869 5760
rect 1494 5729 1506 5732
rect 1448 5723 1506 5729
rect 1857 5729 1869 5732
rect 1903 5760 1915 5763
rect 2222 5760 2228 5772
rect 1903 5732 2228 5760
rect 1903 5729 1915 5732
rect 1857 5723 1915 5729
rect 2222 5720 2228 5732
rect 2280 5720 2286 5772
rect 2314 5720 2320 5772
rect 2372 5760 2378 5772
rect 2409 5763 2467 5769
rect 2409 5760 2421 5763
rect 2372 5732 2421 5760
rect 2372 5720 2378 5732
rect 2409 5729 2421 5732
rect 2455 5729 2467 5763
rect 2409 5723 2467 5729
rect 2685 5763 2743 5769
rect 2685 5729 2697 5763
rect 2731 5760 2743 5763
rect 3605 5763 3663 5769
rect 3605 5760 3617 5763
rect 2731 5732 3617 5760
rect 2731 5729 2743 5732
rect 2685 5723 2743 5729
rect 3605 5729 3617 5732
rect 3651 5760 3663 5763
rect 3878 5760 3884 5772
rect 3651 5732 3884 5760
rect 3651 5729 3663 5732
rect 3605 5723 3663 5729
rect 3878 5720 3884 5732
rect 3936 5760 3942 5772
rect 4338 5760 4344 5772
rect 3936 5732 4154 5760
rect 4299 5732 4344 5760
rect 3936 5720 3942 5732
rect 3142 5692 3148 5704
rect 3103 5664 3148 5692
rect 3142 5652 3148 5664
rect 3200 5652 3206 5704
rect 4126 5692 4154 5732
rect 4338 5720 4344 5732
rect 4396 5720 4402 5772
rect 4617 5763 4675 5769
rect 4617 5729 4629 5763
rect 4663 5729 4675 5763
rect 5902 5760 5908 5772
rect 5863 5732 5908 5760
rect 4617 5723 4675 5729
rect 4632 5692 4660 5723
rect 5902 5720 5908 5732
rect 5960 5720 5966 5772
rect 9232 5760 9260 5800
rect 9306 5788 9312 5840
rect 9364 5828 9370 5840
rect 9861 5831 9919 5837
rect 9861 5828 9873 5831
rect 9364 5800 9873 5828
rect 9364 5788 9370 5800
rect 9861 5797 9873 5800
rect 9907 5797 9919 5831
rect 9861 5791 9919 5797
rect 9490 5760 9496 5772
rect 9232 5732 9496 5760
rect 9490 5720 9496 5732
rect 9548 5720 9554 5772
rect 10704 5760 10732 5859
rect 12084 5837 12112 5868
rect 14001 5865 14013 5868
rect 14047 5865 14059 5899
rect 14182 5896 14188 5908
rect 14143 5868 14188 5896
rect 14001 5859 14059 5865
rect 14182 5856 14188 5868
rect 14240 5856 14246 5908
rect 17402 5856 17408 5908
rect 17460 5896 17466 5908
rect 19521 5899 19579 5905
rect 19521 5896 19533 5899
rect 17460 5868 19533 5896
rect 17460 5856 17466 5868
rect 19521 5865 19533 5868
rect 19567 5865 19579 5899
rect 19521 5859 19579 5865
rect 12069 5831 12127 5837
rect 12069 5797 12081 5831
rect 12115 5797 12127 5831
rect 13170 5828 13176 5840
rect 13131 5800 13176 5828
rect 12069 5791 12127 5797
rect 11425 5763 11483 5769
rect 11425 5760 11437 5763
rect 10704 5732 11437 5760
rect 11425 5729 11437 5732
rect 11471 5760 11483 5763
rect 11790 5760 11796 5772
rect 11471 5732 11796 5760
rect 11471 5729 11483 5732
rect 11425 5723 11483 5729
rect 11790 5720 11796 5732
rect 11848 5720 11854 5772
rect 4126 5664 4660 5692
rect 6273 5695 6331 5701
rect 6273 5661 6285 5695
rect 6319 5692 6331 5695
rect 6362 5692 6368 5704
rect 6319 5664 6368 5692
rect 6319 5661 6331 5664
rect 6273 5655 6331 5661
rect 6362 5652 6368 5664
rect 6420 5652 6426 5704
rect 7466 5692 7472 5704
rect 7427 5664 7472 5692
rect 7466 5652 7472 5664
rect 7524 5652 7530 5704
rect 8941 5695 8999 5701
rect 8941 5661 8953 5695
rect 8987 5692 8999 5695
rect 9033 5695 9091 5701
rect 9033 5692 9045 5695
rect 8987 5664 9045 5692
rect 8987 5661 8999 5664
rect 8941 5655 8999 5661
rect 9033 5661 9045 5664
rect 9079 5692 9091 5695
rect 9398 5692 9404 5704
rect 9079 5664 9404 5692
rect 9079 5661 9091 5664
rect 9033 5655 9091 5661
rect 9398 5652 9404 5664
rect 9456 5652 9462 5704
rect 9766 5692 9772 5704
rect 9727 5664 9772 5692
rect 9766 5652 9772 5664
rect 9824 5652 9830 5704
rect 10410 5692 10416 5704
rect 10371 5664 10416 5692
rect 10410 5652 10416 5664
rect 10468 5652 10474 5704
rect 10502 5652 10508 5704
rect 10560 5692 10566 5704
rect 11057 5695 11115 5701
rect 11057 5692 11069 5695
rect 10560 5664 11069 5692
rect 10560 5652 10566 5664
rect 11057 5661 11069 5664
rect 11103 5661 11115 5695
rect 11057 5655 11115 5661
rect 2498 5624 2504 5636
rect 2459 5596 2504 5624
rect 2498 5584 2504 5596
rect 2556 5584 2562 5636
rect 4430 5624 4436 5636
rect 4391 5596 4436 5624
rect 4430 5584 4436 5596
rect 4488 5584 4494 5636
rect 6178 5624 6184 5636
rect 6091 5596 6184 5624
rect 6178 5584 6184 5596
rect 6236 5624 6242 5636
rect 12084 5624 12112 5791
rect 13170 5788 13176 5800
rect 13228 5788 13234 5840
rect 16114 5828 16120 5840
rect 16075 5800 16120 5828
rect 16114 5788 16120 5800
rect 16172 5788 16178 5840
rect 16666 5828 16672 5840
rect 16627 5800 16672 5828
rect 16666 5788 16672 5800
rect 16724 5788 16730 5840
rect 17678 5828 17684 5840
rect 17639 5800 17684 5828
rect 17678 5788 17684 5800
rect 17736 5788 17742 5840
rect 18233 5831 18291 5837
rect 18233 5797 18245 5831
rect 18279 5828 18291 5831
rect 18414 5828 18420 5840
rect 18279 5800 18420 5828
rect 18279 5797 18291 5800
rect 18233 5791 18291 5797
rect 18414 5788 18420 5800
rect 18472 5788 18478 5840
rect 12529 5763 12587 5769
rect 12529 5729 12541 5763
rect 12575 5760 12587 5763
rect 13446 5760 13452 5772
rect 12575 5732 13452 5760
rect 12575 5729 12587 5732
rect 12529 5723 12587 5729
rect 13446 5720 13452 5732
rect 13504 5720 13510 5772
rect 19061 5763 19119 5769
rect 19061 5729 19073 5763
rect 19107 5729 19119 5763
rect 19061 5723 19119 5729
rect 13630 5652 13636 5704
rect 13688 5692 13694 5704
rect 16025 5695 16083 5701
rect 16025 5692 16037 5695
rect 13688 5664 16037 5692
rect 13688 5652 13694 5664
rect 16025 5661 16037 5664
rect 16071 5692 16083 5695
rect 16942 5692 16948 5704
rect 16071 5664 16948 5692
rect 16071 5661 16083 5664
rect 16025 5655 16083 5661
rect 16942 5652 16948 5664
rect 17000 5652 17006 5704
rect 17405 5695 17463 5701
rect 17405 5661 17417 5695
rect 17451 5692 17463 5695
rect 17586 5692 17592 5704
rect 17451 5664 17592 5692
rect 17451 5661 17463 5664
rect 17405 5655 17463 5661
rect 17586 5652 17592 5664
rect 17644 5652 17650 5704
rect 19076 5692 19104 5723
rect 19150 5720 19156 5772
rect 19208 5760 19214 5772
rect 19337 5763 19395 5769
rect 19337 5760 19349 5763
rect 19208 5732 19349 5760
rect 19208 5720 19214 5732
rect 19337 5729 19349 5732
rect 19383 5729 19395 5763
rect 19337 5723 19395 5729
rect 17696 5664 19472 5692
rect 15470 5624 15476 5636
rect 6236 5596 12112 5624
rect 12360 5596 15476 5624
rect 6236 5584 6242 5596
rect 2314 5556 2320 5568
rect 2275 5528 2320 5556
rect 2314 5516 2320 5528
rect 2372 5516 2378 5568
rect 5166 5516 5172 5568
rect 5224 5556 5230 5568
rect 5353 5559 5411 5565
rect 5353 5556 5365 5559
rect 5224 5528 5365 5556
rect 5224 5516 5230 5528
rect 5353 5525 5365 5528
rect 5399 5525 5411 5559
rect 5353 5519 5411 5525
rect 6070 5559 6128 5565
rect 6070 5525 6082 5559
rect 6116 5556 6128 5559
rect 6270 5556 6276 5568
rect 6116 5528 6276 5556
rect 6116 5525 6128 5528
rect 6070 5519 6128 5525
rect 6270 5516 6276 5528
rect 6328 5516 6334 5568
rect 8389 5559 8447 5565
rect 8389 5525 8401 5559
rect 8435 5556 8447 5559
rect 9033 5559 9091 5565
rect 9033 5556 9045 5559
rect 8435 5528 9045 5556
rect 8435 5525 8447 5528
rect 8389 5519 8447 5525
rect 9033 5525 9045 5528
rect 9079 5525 9091 5559
rect 9033 5519 9091 5525
rect 11238 5516 11244 5568
rect 11296 5556 11302 5568
rect 12360 5556 12388 5596
rect 15470 5584 15476 5596
rect 15528 5624 15534 5636
rect 15565 5627 15623 5633
rect 15565 5624 15577 5627
rect 15528 5596 15577 5624
rect 15528 5584 15534 5596
rect 15565 5593 15577 5596
rect 15611 5593 15623 5627
rect 15565 5587 15623 5593
rect 16758 5584 16764 5636
rect 16816 5624 16822 5636
rect 17696 5624 17724 5664
rect 19058 5624 19064 5636
rect 16816 5596 17724 5624
rect 17925 5596 19064 5624
rect 16816 5584 16822 5596
rect 11296 5528 12388 5556
rect 11296 5516 11302 5528
rect 12434 5516 12440 5568
rect 12492 5556 12498 5568
rect 12805 5559 12863 5565
rect 12805 5556 12817 5559
rect 12492 5528 12817 5556
rect 12492 5516 12498 5528
rect 12805 5525 12817 5528
rect 12851 5525 12863 5559
rect 12805 5519 12863 5525
rect 14001 5559 14059 5565
rect 14001 5525 14013 5559
rect 14047 5556 14059 5559
rect 17925 5556 17953 5596
rect 19058 5584 19064 5596
rect 19116 5624 19122 5636
rect 19153 5627 19211 5633
rect 19153 5624 19165 5627
rect 19116 5596 19165 5624
rect 19116 5584 19122 5596
rect 19153 5593 19165 5596
rect 19199 5593 19211 5627
rect 19444 5624 19472 5664
rect 19610 5624 19616 5636
rect 19444 5596 19616 5624
rect 19153 5587 19211 5593
rect 19610 5584 19616 5596
rect 19668 5584 19674 5636
rect 14047 5528 17953 5556
rect 14047 5525 14059 5528
rect 14001 5519 14059 5525
rect 18230 5516 18236 5568
rect 18288 5556 18294 5568
rect 18509 5559 18567 5565
rect 18509 5556 18521 5559
rect 18288 5528 18521 5556
rect 18288 5516 18294 5528
rect 18509 5525 18521 5528
rect 18555 5525 18567 5559
rect 18509 5519 18567 5525
rect 1104 5466 20884 5488
rect 1104 5414 4648 5466
rect 4700 5414 4712 5466
rect 4764 5414 4776 5466
rect 4828 5414 4840 5466
rect 4892 5414 11982 5466
rect 12034 5414 12046 5466
rect 12098 5414 12110 5466
rect 12162 5414 12174 5466
rect 12226 5414 19315 5466
rect 19367 5414 19379 5466
rect 19431 5414 19443 5466
rect 19495 5414 19507 5466
rect 19559 5414 20884 5466
rect 1104 5392 20884 5414
rect 1719 5355 1777 5361
rect 1719 5321 1731 5355
rect 1765 5352 1777 5355
rect 1946 5352 1952 5364
rect 1765 5324 1952 5352
rect 1765 5321 1777 5324
rect 1719 5315 1777 5321
rect 1946 5312 1952 5324
rect 2004 5312 2010 5364
rect 2682 5312 2688 5364
rect 2740 5352 2746 5364
rect 3053 5355 3111 5361
rect 3053 5352 3065 5355
rect 2740 5324 3065 5352
rect 2740 5312 2746 5324
rect 3053 5321 3065 5324
rect 3099 5321 3111 5355
rect 3053 5315 3111 5321
rect 4246 5312 4252 5364
rect 4304 5352 4310 5364
rect 4985 5355 5043 5361
rect 4985 5352 4997 5355
rect 4304 5324 4997 5352
rect 4304 5312 4310 5324
rect 4985 5321 4997 5324
rect 5031 5352 5043 5355
rect 5031 5324 5304 5352
rect 5031 5321 5043 5324
rect 4985 5315 5043 5321
rect 5276 5293 5304 5324
rect 7466 5312 7472 5364
rect 7524 5352 7530 5364
rect 8573 5355 8631 5361
rect 8573 5352 8585 5355
rect 7524 5324 8585 5352
rect 7524 5312 7530 5324
rect 8573 5321 8585 5324
rect 8619 5321 8631 5355
rect 10318 5352 10324 5364
rect 8573 5315 8631 5321
rect 8772 5324 10324 5352
rect 5261 5287 5319 5293
rect 5261 5253 5273 5287
rect 5307 5253 5319 5287
rect 5261 5247 5319 5253
rect 5902 5244 5908 5296
rect 5960 5284 5966 5296
rect 6641 5287 6699 5293
rect 6641 5284 6653 5287
rect 5960 5256 6653 5284
rect 5960 5244 5966 5256
rect 6641 5253 6653 5256
rect 6687 5284 6699 5287
rect 8772 5284 8800 5324
rect 10318 5312 10324 5324
rect 10376 5312 10382 5364
rect 11790 5352 11796 5364
rect 11751 5324 11796 5352
rect 11790 5312 11796 5324
rect 11848 5312 11854 5364
rect 13725 5355 13783 5361
rect 13725 5352 13737 5355
rect 11900 5324 13737 5352
rect 6687 5256 8800 5284
rect 6687 5253 6699 5256
rect 6641 5247 6699 5253
rect 9122 5244 9128 5296
rect 9180 5284 9186 5296
rect 11900 5284 11928 5324
rect 13725 5321 13737 5324
rect 13771 5352 13783 5355
rect 13817 5355 13875 5361
rect 13817 5352 13829 5355
rect 13771 5324 13829 5352
rect 13771 5321 13783 5324
rect 13725 5315 13783 5321
rect 13817 5321 13829 5324
rect 13863 5321 13875 5355
rect 13817 5315 13875 5321
rect 15289 5355 15347 5361
rect 15289 5321 15301 5355
rect 15335 5352 15347 5355
rect 16114 5352 16120 5364
rect 15335 5324 16120 5352
rect 15335 5321 15347 5324
rect 15289 5315 15347 5321
rect 16114 5312 16120 5324
rect 16172 5352 16178 5364
rect 16669 5355 16727 5361
rect 16669 5352 16681 5355
rect 16172 5324 16681 5352
rect 16172 5312 16178 5324
rect 16669 5321 16681 5324
rect 16715 5352 16727 5355
rect 17497 5355 17555 5361
rect 17497 5352 17509 5355
rect 16715 5324 17509 5352
rect 16715 5321 16727 5324
rect 16669 5315 16727 5321
rect 17497 5321 17509 5324
rect 17543 5352 17555 5355
rect 17678 5352 17684 5364
rect 17543 5324 17684 5352
rect 17543 5321 17555 5324
rect 17497 5315 17555 5321
rect 17678 5312 17684 5324
rect 17736 5312 17742 5364
rect 19058 5312 19064 5364
rect 19116 5352 19122 5364
rect 19429 5355 19487 5361
rect 19429 5352 19441 5355
rect 19116 5324 19441 5352
rect 19116 5312 19122 5324
rect 19429 5321 19441 5324
rect 19475 5321 19487 5355
rect 19429 5315 19487 5321
rect 19751 5355 19809 5361
rect 19751 5321 19763 5355
rect 19797 5352 19809 5355
rect 19886 5352 19892 5364
rect 19797 5324 19892 5352
rect 19797 5321 19809 5324
rect 19751 5315 19809 5321
rect 19886 5312 19892 5324
rect 19944 5312 19950 5364
rect 9180 5256 9260 5284
rect 9180 5244 9186 5256
rect 2498 5216 2504 5228
rect 2411 5188 2504 5216
rect 2498 5176 2504 5188
rect 2556 5216 2562 5228
rect 3513 5219 3571 5225
rect 3513 5216 3525 5219
rect 2556 5188 3525 5216
rect 2556 5176 2562 5188
rect 3513 5185 3525 5188
rect 3559 5216 3571 5219
rect 3559 5188 3740 5216
rect 3559 5185 3571 5188
rect 3513 5179 3571 5185
rect 3712 5160 3740 5188
rect 3970 5176 3976 5228
rect 4028 5216 4034 5228
rect 4065 5219 4123 5225
rect 4065 5216 4077 5219
rect 4028 5188 4077 5216
rect 4028 5176 4034 5188
rect 4065 5185 4077 5188
rect 4111 5216 4123 5219
rect 4154 5216 4160 5228
rect 4111 5188 4160 5216
rect 4111 5185 4123 5188
rect 4065 5179 4123 5185
rect 4154 5176 4160 5188
rect 4212 5216 4218 5228
rect 5350 5216 5356 5228
rect 4212 5188 5356 5216
rect 4212 5176 4218 5188
rect 5350 5176 5356 5188
rect 5408 5176 5414 5228
rect 5534 5176 5540 5228
rect 5592 5216 5598 5228
rect 5629 5219 5687 5225
rect 5629 5216 5641 5219
rect 5592 5188 5641 5216
rect 5592 5176 5598 5188
rect 5629 5185 5641 5188
rect 5675 5185 5687 5219
rect 5629 5179 5687 5185
rect 6273 5219 6331 5225
rect 6273 5185 6285 5219
rect 6319 5216 6331 5219
rect 6362 5216 6368 5228
rect 6319 5188 6368 5216
rect 6319 5185 6331 5188
rect 6273 5179 6331 5185
rect 6362 5176 6368 5188
rect 6420 5216 6426 5228
rect 8662 5216 8668 5228
rect 6420 5188 8668 5216
rect 6420 5176 6426 5188
rect 8662 5176 8668 5188
rect 8720 5176 8726 5228
rect 9232 5225 9260 5256
rect 10888 5256 11928 5284
rect 13265 5287 13323 5293
rect 9217 5219 9275 5225
rect 9217 5185 9229 5219
rect 9263 5185 9275 5219
rect 9217 5179 9275 5185
rect 9861 5219 9919 5225
rect 9861 5185 9873 5219
rect 9907 5216 9919 5219
rect 9950 5216 9956 5228
rect 9907 5188 9956 5216
rect 9907 5185 9919 5188
rect 9861 5179 9919 5185
rect 9950 5176 9956 5188
rect 10008 5176 10014 5228
rect 1648 5151 1706 5157
rect 1648 5117 1660 5151
rect 1694 5148 1706 5151
rect 2593 5151 2651 5157
rect 1694 5120 2176 5148
rect 1694 5117 1706 5120
rect 1648 5111 1706 5117
rect 2148 5024 2176 5120
rect 2593 5117 2605 5151
rect 2639 5148 2651 5151
rect 2682 5148 2688 5160
rect 2639 5120 2688 5148
rect 2639 5117 2651 5120
rect 2593 5111 2651 5117
rect 2682 5108 2688 5120
rect 2740 5108 2746 5160
rect 3605 5151 3663 5157
rect 3605 5117 3617 5151
rect 3651 5117 3663 5151
rect 3605 5111 3663 5117
rect 3620 5080 3648 5111
rect 3694 5108 3700 5160
rect 3752 5148 3758 5160
rect 3878 5148 3884 5160
rect 3752 5120 3797 5148
rect 3839 5120 3884 5148
rect 3752 5108 3758 5120
rect 3878 5108 3884 5120
rect 3936 5148 3942 5160
rect 4522 5148 4528 5160
rect 3936 5120 4528 5148
rect 3936 5108 3942 5120
rect 4522 5108 4528 5120
rect 4580 5108 4586 5160
rect 5166 5148 5172 5160
rect 5127 5120 5172 5148
rect 5166 5108 5172 5120
rect 5224 5108 5230 5160
rect 5442 5148 5448 5160
rect 5403 5120 5448 5148
rect 5442 5108 5448 5120
rect 5500 5108 5506 5160
rect 7374 5148 7380 5160
rect 7335 5120 7380 5148
rect 7374 5108 7380 5120
rect 7432 5108 7438 5160
rect 10321 5151 10379 5157
rect 10321 5117 10333 5151
rect 10367 5148 10379 5151
rect 10778 5148 10784 5160
rect 10367 5120 10784 5148
rect 10367 5117 10379 5120
rect 10321 5111 10379 5117
rect 10778 5108 10784 5120
rect 10836 5108 10842 5160
rect 10888 5157 10916 5256
rect 13265 5253 13277 5287
rect 13311 5284 13323 5287
rect 16758 5284 16764 5296
rect 13311 5256 16764 5284
rect 13311 5253 13323 5256
rect 13265 5247 13323 5253
rect 16758 5244 16764 5256
rect 16816 5244 16822 5296
rect 16942 5284 16948 5296
rect 16903 5256 16948 5284
rect 16942 5244 16948 5256
rect 17000 5244 17006 5296
rect 12253 5219 12311 5225
rect 12253 5185 12265 5219
rect 12299 5216 12311 5219
rect 12342 5216 12348 5228
rect 12299 5188 12348 5216
rect 12299 5185 12311 5188
rect 12253 5179 12311 5185
rect 12342 5176 12348 5188
rect 12400 5216 12406 5228
rect 12529 5219 12587 5225
rect 12529 5216 12541 5219
rect 12400 5188 12541 5216
rect 12400 5176 12406 5188
rect 12529 5185 12541 5188
rect 12575 5185 12587 5219
rect 12529 5179 12587 5185
rect 16666 5176 16672 5228
rect 16724 5216 16730 5228
rect 18141 5219 18199 5225
rect 18141 5216 18153 5219
rect 16724 5188 18153 5216
rect 16724 5176 16730 5188
rect 18141 5185 18153 5188
rect 18187 5216 18199 5219
rect 18322 5216 18328 5228
rect 18187 5188 18328 5216
rect 18187 5185 18199 5188
rect 18141 5179 18199 5185
rect 18322 5176 18328 5188
rect 18380 5176 18386 5228
rect 18506 5176 18512 5228
rect 18564 5216 18570 5228
rect 18564 5188 19707 5216
rect 18564 5176 18570 5188
rect 10873 5151 10931 5157
rect 10873 5117 10885 5151
rect 10919 5117 10931 5151
rect 11054 5148 11060 5160
rect 11015 5120 11060 5148
rect 10873 5111 10931 5117
rect 4338 5080 4344 5092
rect 3620 5052 4344 5080
rect 4338 5040 4344 5052
rect 4396 5040 4402 5092
rect 4709 5083 4767 5089
rect 4709 5049 4721 5083
rect 4755 5080 4767 5083
rect 5460 5080 5488 5108
rect 4755 5052 5488 5080
rect 7698 5083 7756 5089
rect 4755 5049 4767 5052
rect 4709 5043 4767 5049
rect 7698 5049 7710 5083
rect 7744 5080 7756 5083
rect 7834 5080 7840 5092
rect 7744 5052 7840 5080
rect 7744 5049 7756 5052
rect 7698 5043 7756 5049
rect 2130 5012 2136 5024
rect 2091 4984 2136 5012
rect 2130 4972 2136 4984
rect 2188 4972 2194 5024
rect 2731 5015 2789 5021
rect 2731 4981 2743 5015
rect 2777 5012 2789 5015
rect 2866 5012 2872 5024
rect 2777 4984 2872 5012
rect 2777 4981 2789 4984
rect 2731 4975 2789 4981
rect 2866 4972 2872 4984
rect 2924 4972 2930 5024
rect 7285 5015 7343 5021
rect 7285 4981 7297 5015
rect 7331 5012 7343 5015
rect 7466 5012 7472 5024
rect 7331 4984 7472 5012
rect 7331 4981 7343 4984
rect 7285 4975 7343 4981
rect 7466 4972 7472 4984
rect 7524 5012 7530 5024
rect 7713 5012 7741 5043
rect 7834 5040 7840 5052
rect 7892 5040 7898 5092
rect 9306 5040 9312 5092
rect 9364 5080 9370 5092
rect 10594 5080 10600 5092
rect 9364 5052 9409 5080
rect 10555 5052 10600 5080
rect 9364 5040 9370 5052
rect 10594 5040 10600 5052
rect 10652 5080 10658 5092
rect 10888 5080 10916 5111
rect 11054 5108 11060 5120
rect 11112 5108 11118 5160
rect 12434 5148 12440 5160
rect 12395 5120 12440 5148
rect 12434 5108 12440 5120
rect 12492 5108 12498 5160
rect 12713 5151 12771 5157
rect 12713 5117 12725 5151
rect 12759 5148 12771 5151
rect 13446 5148 13452 5160
rect 12759 5120 13452 5148
rect 12759 5117 12771 5120
rect 12713 5111 12771 5117
rect 13446 5108 13452 5120
rect 13504 5108 13510 5160
rect 13725 5151 13783 5157
rect 13725 5117 13737 5151
rect 13771 5148 13783 5151
rect 14093 5151 14151 5157
rect 14093 5148 14105 5151
rect 13771 5120 14105 5148
rect 13771 5117 13783 5120
rect 13725 5111 13783 5117
rect 14093 5117 14105 5120
rect 14139 5117 14151 5151
rect 14093 5111 14151 5117
rect 15470 5108 15476 5160
rect 15528 5148 15534 5160
rect 19679 5157 19707 5188
rect 15749 5151 15807 5157
rect 15749 5148 15761 5151
rect 15528 5120 15761 5148
rect 15528 5108 15534 5120
rect 15749 5117 15761 5120
rect 15795 5117 15807 5151
rect 15749 5111 15807 5117
rect 19664 5151 19722 5157
rect 19664 5117 19676 5151
rect 19710 5148 19722 5151
rect 20073 5151 20131 5157
rect 20073 5148 20085 5151
rect 19710 5120 20085 5148
rect 19710 5117 19722 5120
rect 19664 5111 19722 5117
rect 20073 5117 20085 5120
rect 20119 5117 20131 5151
rect 20073 5111 20131 5117
rect 10652 5052 10916 5080
rect 10652 5040 10658 5052
rect 11606 5040 11612 5092
rect 11664 5080 11670 5092
rect 11664 5052 12020 5080
rect 11664 5040 11670 5052
rect 7524 4984 7741 5012
rect 8297 5015 8355 5021
rect 7524 4972 7530 4984
rect 8297 4981 8309 5015
rect 8343 5012 8355 5015
rect 9033 5015 9091 5021
rect 9033 5012 9045 5015
rect 8343 4984 9045 5012
rect 8343 4981 8355 4984
rect 8297 4975 8355 4981
rect 9033 4981 9045 4984
rect 9079 5012 9091 5015
rect 9324 5012 9352 5040
rect 9079 4984 9352 5012
rect 9079 4981 9091 4984
rect 9033 4975 9091 4981
rect 10226 4972 10232 5024
rect 10284 5012 10290 5024
rect 11238 5012 11244 5024
rect 10284 4984 11244 5012
rect 10284 4972 10290 4984
rect 11238 4972 11244 4984
rect 11296 4972 11302 5024
rect 11992 5012 12020 5052
rect 12342 5040 12348 5092
rect 12400 5080 12406 5092
rect 14001 5083 14059 5089
rect 14001 5080 14013 5083
rect 12400 5052 14013 5080
rect 12400 5040 12406 5052
rect 14001 5049 14013 5052
rect 14047 5049 14059 5083
rect 14001 5043 14059 5049
rect 15657 5083 15715 5089
rect 15657 5049 15669 5083
rect 15703 5080 15715 5083
rect 16111 5083 16169 5089
rect 16111 5080 16123 5083
rect 15703 5052 16123 5080
rect 15703 5049 15715 5052
rect 15657 5043 15715 5049
rect 16111 5049 16123 5052
rect 16157 5080 16169 5083
rect 16574 5080 16580 5092
rect 16157 5052 16580 5080
rect 16157 5049 16169 5052
rect 16111 5043 16169 5049
rect 16574 5040 16580 5052
rect 16632 5080 16638 5092
rect 16758 5080 16764 5092
rect 16632 5052 16764 5080
rect 16632 5040 16638 5052
rect 16758 5040 16764 5052
rect 16816 5040 16822 5092
rect 18230 5040 18236 5092
rect 18288 5080 18294 5092
rect 18785 5083 18843 5089
rect 18288 5052 18333 5080
rect 18288 5040 18294 5052
rect 18785 5049 18797 5083
rect 18831 5080 18843 5083
rect 18966 5080 18972 5092
rect 18831 5052 18972 5080
rect 18831 5049 18843 5052
rect 18785 5043 18843 5049
rect 18966 5040 18972 5052
rect 19024 5040 19030 5092
rect 12897 5015 12955 5021
rect 12897 5012 12909 5015
rect 11992 4984 12909 5012
rect 12897 4981 12909 4984
rect 12943 5012 12955 5015
rect 13265 5015 13323 5021
rect 13265 5012 13277 5015
rect 12943 4984 13277 5012
rect 12943 4981 12955 4984
rect 12897 4975 12955 4981
rect 13265 4981 13277 4984
rect 13311 4981 13323 5015
rect 13446 5012 13452 5024
rect 13407 4984 13452 5012
rect 13265 4975 13323 4981
rect 13446 4972 13452 4984
rect 13504 4972 13510 5024
rect 17678 4972 17684 5024
rect 17736 5012 17742 5024
rect 19061 5015 19119 5021
rect 19061 5012 19073 5015
rect 17736 4984 19073 5012
rect 17736 4972 17742 4984
rect 19061 4981 19073 4984
rect 19107 5012 19119 5015
rect 19150 5012 19156 5024
rect 19107 4984 19156 5012
rect 19107 4981 19119 4984
rect 19061 4975 19119 4981
rect 19150 4972 19156 4984
rect 19208 4972 19214 5024
rect 1104 4922 20884 4944
rect 1104 4870 8315 4922
rect 8367 4870 8379 4922
rect 8431 4870 8443 4922
rect 8495 4870 8507 4922
rect 8559 4870 15648 4922
rect 15700 4870 15712 4922
rect 15764 4870 15776 4922
rect 15828 4870 15840 4922
rect 15892 4870 20884 4922
rect 1104 4848 20884 4870
rect 3513 4811 3571 4817
rect 3513 4777 3525 4811
rect 3559 4808 3571 4811
rect 4433 4811 4491 4817
rect 4433 4808 4445 4811
rect 3559 4780 4445 4808
rect 3559 4777 3571 4780
rect 3513 4771 3571 4777
rect 4433 4777 4445 4780
rect 4479 4808 4491 4811
rect 4522 4808 4528 4820
rect 4479 4780 4528 4808
rect 4479 4777 4491 4780
rect 4433 4771 4491 4777
rect 4522 4768 4528 4780
rect 4580 4768 4586 4820
rect 5997 4811 6055 4817
rect 5997 4777 6009 4811
rect 6043 4808 6055 4811
rect 6178 4808 6184 4820
rect 6043 4780 6184 4808
rect 6043 4777 6055 4780
rect 5997 4771 6055 4777
rect 6178 4768 6184 4780
rect 6236 4768 6242 4820
rect 6270 4768 6276 4820
rect 6328 4808 6334 4820
rect 9217 4811 9275 4817
rect 6328 4780 6373 4808
rect 6328 4768 6334 4780
rect 9217 4777 9229 4811
rect 9263 4808 9275 4811
rect 9306 4808 9312 4820
rect 9263 4780 9312 4808
rect 9263 4777 9275 4780
rect 9217 4771 9275 4777
rect 9306 4768 9312 4780
rect 9364 4768 9370 4820
rect 9582 4768 9588 4820
rect 9640 4808 9646 4820
rect 10410 4808 10416 4820
rect 9640 4780 10416 4808
rect 9640 4768 9646 4780
rect 10410 4768 10416 4780
rect 10468 4808 10474 4820
rect 12989 4811 13047 4817
rect 12989 4808 13001 4811
rect 10468 4780 13001 4808
rect 10468 4768 10474 4780
rect 12989 4777 13001 4780
rect 13035 4777 13047 4811
rect 17678 4808 17684 4820
rect 12989 4771 13047 4777
rect 13786 4780 17684 4808
rect 3145 4743 3203 4749
rect 3145 4709 3157 4743
rect 3191 4740 3203 4743
rect 3234 4740 3240 4752
rect 3191 4712 3240 4740
rect 3191 4709 3203 4712
rect 3145 4703 3203 4709
rect 3234 4700 3240 4712
rect 3292 4740 3298 4752
rect 6362 4740 6368 4752
rect 3292 4712 6368 4740
rect 3292 4700 3298 4712
rect 6362 4700 6368 4712
rect 6420 4700 6426 4752
rect 7193 4743 7251 4749
rect 7193 4709 7205 4743
rect 7239 4740 7251 4743
rect 7374 4740 7380 4752
rect 7239 4712 7380 4740
rect 7239 4709 7251 4712
rect 7193 4703 7251 4709
rect 7374 4700 7380 4712
rect 7432 4740 7438 4752
rect 7837 4743 7895 4749
rect 7837 4740 7849 4743
rect 7432 4712 7849 4740
rect 7432 4700 7438 4712
rect 7837 4709 7849 4712
rect 7883 4709 7895 4743
rect 8202 4740 8208 4752
rect 8163 4712 8208 4740
rect 7837 4703 7895 4709
rect 8202 4700 8208 4712
rect 8260 4700 8266 4752
rect 9858 4740 9864 4752
rect 9819 4712 9864 4740
rect 9858 4700 9864 4712
rect 9916 4700 9922 4752
rect 12434 4740 12440 4752
rect 11992 4712 12440 4740
rect 1302 4632 1308 4684
rect 1360 4672 1366 4684
rect 1432 4675 1490 4681
rect 1432 4672 1444 4675
rect 1360 4644 1444 4672
rect 1360 4632 1366 4644
rect 1432 4641 1444 4644
rect 1478 4672 1490 4675
rect 1854 4672 1860 4684
rect 1478 4644 1860 4672
rect 1478 4641 1490 4644
rect 1432 4635 1490 4641
rect 1854 4632 1860 4644
rect 1912 4632 1918 4684
rect 2406 4672 2412 4684
rect 2367 4644 2412 4672
rect 2406 4632 2412 4644
rect 2464 4632 2470 4684
rect 2685 4675 2743 4681
rect 2685 4641 2697 4675
rect 2731 4641 2743 4675
rect 3786 4672 3792 4684
rect 3747 4644 3792 4672
rect 2685 4635 2743 4641
rect 2314 4564 2320 4616
rect 2372 4604 2378 4616
rect 2700 4604 2728 4635
rect 3786 4632 3792 4644
rect 3844 4632 3850 4684
rect 4430 4632 4436 4684
rect 4488 4672 4494 4684
rect 4709 4675 4767 4681
rect 4709 4672 4721 4675
rect 4488 4644 4721 4672
rect 4488 4632 4494 4644
rect 4709 4641 4721 4644
rect 4755 4641 4767 4675
rect 5166 4672 5172 4684
rect 5127 4644 5172 4672
rect 4709 4635 4767 4641
rect 5166 4632 5172 4644
rect 5224 4632 5230 4684
rect 5350 4672 5356 4684
rect 5311 4644 5356 4672
rect 5350 4632 5356 4644
rect 5408 4632 5414 4684
rect 6457 4675 6515 4681
rect 6457 4672 6469 4675
rect 5460 4644 6469 4672
rect 2372 4576 2728 4604
rect 2372 4564 2378 4576
rect 2958 4564 2964 4616
rect 3016 4604 3022 4616
rect 5184 4604 5212 4632
rect 5460 4604 5488 4644
rect 6457 4641 6469 4644
rect 6503 4641 6515 4675
rect 7006 4672 7012 4684
rect 6919 4644 7012 4672
rect 6457 4635 6515 4641
rect 7006 4632 7012 4644
rect 7064 4672 7070 4684
rect 7282 4672 7288 4684
rect 7064 4644 7288 4672
rect 7064 4632 7070 4644
rect 7282 4632 7288 4644
rect 7340 4632 7346 4684
rect 11790 4672 11796 4684
rect 11751 4644 11796 4672
rect 11790 4632 11796 4644
rect 11848 4672 11854 4684
rect 11992 4681 12020 4712
rect 12434 4700 12440 4712
rect 12492 4700 12498 4752
rect 12618 4740 12624 4752
rect 12531 4712 12624 4740
rect 11977 4675 12035 4681
rect 11977 4672 11989 4675
rect 11848 4644 11989 4672
rect 11848 4632 11854 4644
rect 11977 4641 11989 4644
rect 12023 4641 12035 4675
rect 11977 4635 12035 4641
rect 12253 4675 12311 4681
rect 12253 4641 12265 4675
rect 12299 4672 12311 4675
rect 12544 4672 12572 4712
rect 12618 4700 12624 4712
rect 12676 4740 12682 4752
rect 13786 4740 13814 4780
rect 17678 4768 17684 4780
rect 17736 4768 17742 4820
rect 17773 4811 17831 4817
rect 17773 4777 17785 4811
rect 17819 4808 17831 4811
rect 18141 4811 18199 4817
rect 18141 4808 18153 4811
rect 17819 4780 18153 4808
rect 17819 4777 17831 4780
rect 17773 4771 17831 4777
rect 18141 4777 18153 4780
rect 18187 4808 18199 4811
rect 18230 4808 18236 4820
rect 18187 4780 18236 4808
rect 18187 4777 18199 4780
rect 18141 4771 18199 4777
rect 18230 4768 18236 4780
rect 18288 4768 18294 4820
rect 18322 4768 18328 4820
rect 18380 4808 18386 4820
rect 18417 4811 18475 4817
rect 18417 4808 18429 4811
rect 18380 4780 18429 4808
rect 18380 4768 18386 4780
rect 18417 4777 18429 4780
rect 18463 4777 18475 4811
rect 19610 4808 19616 4820
rect 19571 4780 19616 4808
rect 18417 4771 18475 4777
rect 19610 4768 19616 4780
rect 19668 4768 19674 4820
rect 15473 4743 15531 4749
rect 15473 4740 15485 4743
rect 12676 4712 13814 4740
rect 14844 4712 15485 4740
rect 12676 4700 12682 4712
rect 14844 4684 14872 4712
rect 15473 4709 15485 4712
rect 15519 4709 15531 4743
rect 15473 4703 15531 4709
rect 16758 4700 16764 4752
rect 16816 4740 16822 4752
rect 17174 4743 17232 4749
rect 17174 4740 17186 4743
rect 16816 4712 17186 4740
rect 16816 4700 16822 4712
rect 17174 4709 17186 4712
rect 17220 4709 17232 4743
rect 18782 4740 18788 4752
rect 18743 4712 18788 4740
rect 17174 4703 17232 4709
rect 18782 4700 18788 4712
rect 18840 4700 18846 4752
rect 12299 4644 12572 4672
rect 13541 4675 13599 4681
rect 12299 4641 12311 4644
rect 12253 4635 12311 4641
rect 13541 4641 13553 4675
rect 13587 4672 13599 4675
rect 13725 4675 13783 4681
rect 13725 4672 13737 4675
rect 13587 4644 13737 4672
rect 13587 4641 13599 4644
rect 13541 4635 13599 4641
rect 13725 4641 13737 4644
rect 13771 4672 13783 4675
rect 14826 4672 14832 4684
rect 13771 4644 14832 4672
rect 13771 4641 13783 4644
rect 13725 4635 13783 4641
rect 14826 4632 14832 4644
rect 14884 4632 14890 4684
rect 3016 4576 5488 4604
rect 5629 4607 5687 4613
rect 3016 4564 3022 4576
rect 5629 4573 5641 4607
rect 5675 4604 5687 4607
rect 7926 4604 7932 4616
rect 5675 4576 7932 4604
rect 5675 4573 5687 4576
rect 5629 4567 5687 4573
rect 7926 4564 7932 4576
rect 7984 4564 7990 4616
rect 8110 4604 8116 4616
rect 8071 4576 8116 4604
rect 8110 4564 8116 4576
rect 8168 4564 8174 4616
rect 8757 4607 8815 4613
rect 8757 4573 8769 4607
rect 8803 4604 8815 4607
rect 9769 4607 9827 4613
rect 9769 4604 9781 4607
rect 8803 4576 9781 4604
rect 8803 4573 8815 4576
rect 8757 4567 8815 4573
rect 9769 4573 9781 4576
rect 9815 4604 9827 4607
rect 9950 4604 9956 4616
rect 9815 4576 9956 4604
rect 9815 4573 9827 4576
rect 9769 4567 9827 4573
rect 9950 4564 9956 4576
rect 10008 4564 10014 4616
rect 10045 4607 10103 4613
rect 10045 4573 10057 4607
rect 10091 4573 10103 4607
rect 10045 4567 10103 4573
rect 2133 4539 2191 4545
rect 2133 4505 2145 4539
rect 2179 4536 2191 4539
rect 2222 4536 2228 4548
rect 2179 4508 2228 4536
rect 2179 4505 2191 4508
rect 2133 4499 2191 4505
rect 2222 4496 2228 4508
rect 2280 4536 2286 4548
rect 2501 4539 2559 4545
rect 2501 4536 2513 4539
rect 2280 4508 2513 4536
rect 2280 4496 2286 4508
rect 2501 4505 2513 4508
rect 2547 4505 2559 4539
rect 2501 4499 2559 4505
rect 9674 4496 9680 4548
rect 9732 4536 9738 4548
rect 10060 4536 10088 4567
rect 11514 4564 11520 4616
rect 11572 4604 11578 4616
rect 12434 4604 12440 4616
rect 11572 4576 12204 4604
rect 12395 4576 12440 4604
rect 11572 4564 11578 4576
rect 9732 4508 10088 4536
rect 9732 4496 9738 4508
rect 11882 4496 11888 4548
rect 11940 4536 11946 4548
rect 12069 4539 12127 4545
rect 12069 4536 12081 4539
rect 11940 4508 12081 4536
rect 11940 4496 11946 4508
rect 12069 4505 12081 4508
rect 12115 4505 12127 4539
rect 12176 4536 12204 4576
rect 12434 4564 12440 4576
rect 12492 4564 12498 4616
rect 14366 4604 14372 4616
rect 14327 4576 14372 4604
rect 14366 4564 14372 4576
rect 14424 4564 14430 4616
rect 15378 4604 15384 4616
rect 15339 4576 15384 4604
rect 15378 4564 15384 4576
rect 15436 4564 15442 4616
rect 16022 4604 16028 4616
rect 15983 4576 16028 4604
rect 16022 4564 16028 4576
rect 16080 4564 16086 4616
rect 16853 4607 16911 4613
rect 16853 4573 16865 4607
rect 16899 4604 16911 4607
rect 17126 4604 17132 4616
rect 16899 4576 17132 4604
rect 16899 4573 16911 4576
rect 16853 4567 16911 4573
rect 17126 4564 17132 4576
rect 17184 4564 17190 4616
rect 18414 4564 18420 4616
rect 18472 4604 18478 4616
rect 18693 4607 18751 4613
rect 18693 4604 18705 4607
rect 18472 4576 18705 4604
rect 18472 4564 18478 4576
rect 18693 4573 18705 4576
rect 18739 4573 18751 4607
rect 18966 4604 18972 4616
rect 18927 4576 18972 4604
rect 18693 4567 18751 4573
rect 18966 4564 18972 4576
rect 19024 4564 19030 4616
rect 15286 4536 15292 4548
rect 12176 4508 15292 4536
rect 12069 4499 12127 4505
rect 15286 4496 15292 4508
rect 15344 4496 15350 4548
rect 15470 4496 15476 4548
rect 15528 4536 15534 4548
rect 16301 4539 16359 4545
rect 16301 4536 16313 4539
rect 15528 4508 16313 4536
rect 15528 4496 15534 4508
rect 16301 4505 16313 4508
rect 16347 4505 16359 4539
rect 16301 4499 16359 4505
rect 1535 4471 1593 4477
rect 1535 4437 1547 4471
rect 1581 4468 1593 4471
rect 1946 4468 1952 4480
rect 1581 4440 1952 4468
rect 1581 4437 1593 4440
rect 1535 4431 1593 4437
rect 1946 4428 1952 4440
rect 2004 4428 2010 4480
rect 6638 4428 6644 4480
rect 6696 4468 6702 4480
rect 7466 4468 7472 4480
rect 6696 4440 7472 4468
rect 6696 4428 6702 4440
rect 7466 4428 7472 4440
rect 7524 4428 7530 4480
rect 7558 4428 7564 4480
rect 7616 4468 7622 4480
rect 10781 4471 10839 4477
rect 10781 4468 10793 4471
rect 7616 4440 10793 4468
rect 7616 4428 7622 4440
rect 10781 4437 10793 4440
rect 10827 4468 10839 4471
rect 11054 4468 11060 4480
rect 10827 4440 11060 4468
rect 10827 4437 10839 4440
rect 10781 4431 10839 4437
rect 11054 4428 11060 4440
rect 11112 4428 11118 4480
rect 11422 4468 11428 4480
rect 11383 4440 11428 4468
rect 11422 4428 11428 4440
rect 11480 4428 11486 4480
rect 1104 4378 20884 4400
rect 1104 4326 4648 4378
rect 4700 4326 4712 4378
rect 4764 4326 4776 4378
rect 4828 4326 4840 4378
rect 4892 4326 11982 4378
rect 12034 4326 12046 4378
rect 12098 4326 12110 4378
rect 12162 4326 12174 4378
rect 12226 4326 19315 4378
rect 19367 4326 19379 4378
rect 19431 4326 19443 4378
rect 19495 4326 19507 4378
rect 19559 4326 20884 4378
rect 1104 4304 20884 4326
rect 8662 4264 8668 4276
rect 4126 4236 8668 4264
rect 2133 4199 2191 4205
rect 2133 4165 2145 4199
rect 2179 4196 2191 4199
rect 2222 4196 2228 4208
rect 2179 4168 2228 4196
rect 2179 4165 2191 4168
rect 2133 4159 2191 4165
rect 2222 4156 2228 4168
rect 2280 4196 2286 4208
rect 2498 4196 2504 4208
rect 2280 4168 2504 4196
rect 2280 4156 2286 4168
rect 2498 4156 2504 4168
rect 2556 4156 2562 4208
rect 2866 4156 2872 4208
rect 2924 4196 2930 4208
rect 4126 4196 4154 4236
rect 8662 4224 8668 4236
rect 8720 4224 8726 4276
rect 9125 4267 9183 4273
rect 9125 4233 9137 4267
rect 9171 4264 9183 4267
rect 9858 4264 9864 4276
rect 9171 4236 9864 4264
rect 9171 4233 9183 4236
rect 9125 4227 9183 4233
rect 9858 4224 9864 4236
rect 9916 4264 9922 4276
rect 10505 4267 10563 4273
rect 10505 4264 10517 4267
rect 9916 4236 10517 4264
rect 9916 4224 9922 4236
rect 10505 4233 10517 4236
rect 10551 4233 10563 4267
rect 10505 4227 10563 4233
rect 11471 4267 11529 4273
rect 11471 4233 11483 4267
rect 11517 4264 11529 4267
rect 12710 4264 12716 4276
rect 11517 4236 12716 4264
rect 11517 4233 11529 4236
rect 11471 4227 11529 4233
rect 12710 4224 12716 4236
rect 12768 4224 12774 4276
rect 14366 4224 14372 4276
rect 14424 4264 14430 4276
rect 15473 4267 15531 4273
rect 15473 4264 15485 4267
rect 14424 4236 15485 4264
rect 14424 4224 14430 4236
rect 15473 4233 15485 4236
rect 15519 4264 15531 4267
rect 15838 4264 15844 4276
rect 15519 4236 15844 4264
rect 15519 4233 15531 4236
rect 15473 4227 15531 4233
rect 15838 4224 15844 4236
rect 15896 4224 15902 4276
rect 18782 4224 18788 4276
rect 18840 4264 18846 4276
rect 18969 4267 19027 4273
rect 18969 4264 18981 4267
rect 18840 4236 18981 4264
rect 18840 4224 18846 4236
rect 18969 4233 18981 4236
rect 19015 4264 19027 4267
rect 19245 4267 19303 4273
rect 19245 4264 19257 4267
rect 19015 4236 19257 4264
rect 19015 4233 19027 4236
rect 18969 4227 19027 4233
rect 19245 4233 19257 4236
rect 19291 4233 19303 4267
rect 19245 4227 19303 4233
rect 2924 4168 4154 4196
rect 4709 4199 4767 4205
rect 2924 4156 2930 4168
rect 4709 4165 4721 4199
rect 4755 4196 4767 4199
rect 4982 4196 4988 4208
rect 4755 4168 4988 4196
rect 4755 4165 4767 4168
rect 4709 4159 4767 4165
rect 4982 4156 4988 4168
rect 5040 4156 5046 4208
rect 6457 4199 6515 4205
rect 6457 4165 6469 4199
rect 6503 4196 6515 4199
rect 9674 4196 9680 4208
rect 6503 4168 9680 4196
rect 6503 4165 6515 4168
rect 6457 4159 6515 4165
rect 9674 4156 9680 4168
rect 9732 4156 9738 4208
rect 11241 4199 11299 4205
rect 11241 4165 11253 4199
rect 11287 4196 11299 4199
rect 11882 4196 11888 4208
rect 11287 4168 11888 4196
rect 11287 4165 11299 4168
rect 11241 4159 11299 4165
rect 11882 4156 11888 4168
rect 11940 4156 11946 4208
rect 12069 4199 12127 4205
rect 12069 4165 12081 4199
rect 12115 4196 12127 4199
rect 12618 4196 12624 4208
rect 12115 4168 12624 4196
rect 12115 4165 12127 4168
rect 12069 4159 12127 4165
rect 12618 4156 12624 4168
rect 12676 4156 12682 4208
rect 14826 4196 14832 4208
rect 14787 4168 14832 4196
rect 14826 4156 14832 4168
rect 14884 4196 14890 4208
rect 15105 4199 15163 4205
rect 15105 4196 15117 4199
rect 14884 4168 15117 4196
rect 14884 4156 14890 4168
rect 15105 4165 15117 4168
rect 15151 4165 15163 4199
rect 15105 4159 15163 4165
rect 1949 4131 2007 4137
rect 1949 4097 1961 4131
rect 1995 4128 2007 4131
rect 2777 4131 2835 4137
rect 1995 4100 2360 4128
rect 1995 4097 2007 4100
rect 1949 4091 2007 4097
rect 2332 4072 2360 4100
rect 2777 4097 2789 4131
rect 2823 4128 2835 4131
rect 2958 4128 2964 4140
rect 2823 4100 2964 4128
rect 2823 4097 2835 4100
rect 2777 4091 2835 4097
rect 2958 4088 2964 4100
rect 3016 4088 3022 4140
rect 3142 4088 3148 4140
rect 3200 4128 3206 4140
rect 5077 4131 5135 4137
rect 5077 4128 5089 4131
rect 3200 4100 5089 4128
rect 3200 4088 3206 4100
rect 5077 4097 5089 4100
rect 5123 4128 5135 4131
rect 5905 4131 5963 4137
rect 5123 4100 5672 4128
rect 5123 4097 5135 4100
rect 5077 4091 5135 4097
rect 2041 4063 2099 4069
rect 2041 4029 2053 4063
rect 2087 4029 2099 4063
rect 2314 4060 2320 4072
rect 2275 4032 2320 4060
rect 2041 4023 2099 4029
rect 2056 3992 2084 4023
rect 2314 4020 2320 4032
rect 2372 4020 2378 4072
rect 2498 4020 2504 4072
rect 2556 4060 2562 4072
rect 3421 4063 3479 4069
rect 3421 4060 3433 4063
rect 2556 4032 3433 4060
rect 2556 4020 2562 4032
rect 3421 4029 3433 4032
rect 3467 4060 3479 4063
rect 3602 4060 3608 4072
rect 3467 4032 3608 4060
rect 3467 4029 3479 4032
rect 3421 4023 3479 4029
rect 3602 4020 3608 4032
rect 3660 4020 3666 4072
rect 3878 4060 3884 4072
rect 3839 4032 3884 4060
rect 3878 4020 3884 4032
rect 3936 4020 3942 4072
rect 4154 4020 4160 4072
rect 4212 4060 4218 4072
rect 4341 4063 4399 4069
rect 4212 4032 4257 4060
rect 4212 4020 4218 4032
rect 4341 4029 4353 4063
rect 4387 4060 4399 4063
rect 4430 4060 4436 4072
rect 4387 4032 4436 4060
rect 4387 4029 4399 4032
rect 4341 4023 4399 4029
rect 4430 4020 4436 4032
rect 4488 4020 4494 4072
rect 4982 4020 4988 4072
rect 5040 4060 5046 4072
rect 5644 4069 5672 4100
rect 5905 4097 5917 4131
rect 5951 4128 5963 4131
rect 9585 4131 9643 4137
rect 9585 4128 9597 4131
rect 5951 4100 9597 4128
rect 5951 4097 5963 4100
rect 5905 4091 5963 4097
rect 9585 4097 9597 4100
rect 9631 4128 9643 4131
rect 10781 4131 10839 4137
rect 10781 4128 10793 4131
rect 9631 4100 10793 4128
rect 9631 4097 9643 4100
rect 9585 4091 9643 4097
rect 10781 4097 10793 4100
rect 10827 4097 10839 4131
rect 13538 4128 13544 4140
rect 10781 4091 10839 4097
rect 12360 4100 13544 4128
rect 5169 4063 5227 4069
rect 5169 4060 5181 4063
rect 5040 4032 5181 4060
rect 5040 4020 5046 4032
rect 5169 4029 5181 4032
rect 5215 4029 5227 4063
rect 5169 4023 5227 4029
rect 5629 4063 5687 4069
rect 5629 4029 5641 4063
rect 5675 4060 5687 4063
rect 6178 4060 6184 4072
rect 5675 4032 6184 4060
rect 5675 4029 5687 4032
rect 5629 4023 5687 4029
rect 6178 4020 6184 4032
rect 6236 4020 6242 4072
rect 7098 4060 7104 4072
rect 7059 4032 7104 4060
rect 7098 4020 7104 4032
rect 7156 4020 7162 4072
rect 8021 4063 8079 4069
rect 8021 4029 8033 4063
rect 8067 4060 8079 4063
rect 8202 4060 8208 4072
rect 8067 4032 8208 4060
rect 8067 4029 8079 4032
rect 8021 4023 8079 4029
rect 8202 4020 8208 4032
rect 8260 4060 8266 4072
rect 8260 4032 8524 4060
rect 8260 4020 8266 4032
rect 3510 3992 3516 4004
rect 2056 3964 3516 3992
rect 3510 3952 3516 3964
rect 3568 3952 3574 4004
rect 6457 3995 6515 4001
rect 6457 3992 6469 3995
rect 4448 3964 6469 3992
rect 2406 3884 2412 3936
rect 2464 3924 2470 3936
rect 3053 3927 3111 3933
rect 3053 3924 3065 3927
rect 2464 3896 3065 3924
rect 2464 3884 2470 3896
rect 3053 3893 3065 3896
rect 3099 3893 3111 3927
rect 3053 3887 3111 3893
rect 4062 3884 4068 3936
rect 4120 3924 4126 3936
rect 4448 3924 4476 3964
rect 6457 3961 6469 3964
rect 6503 3961 6515 3995
rect 6457 3955 6515 3961
rect 6638 3924 6644 3936
rect 4120 3896 4476 3924
rect 6599 3896 6644 3924
rect 4120 3884 4126 3896
rect 6638 3884 6644 3896
rect 6696 3884 6702 3936
rect 7466 3884 7472 3936
rect 7524 3924 7530 3936
rect 7524 3896 7569 3924
rect 7524 3884 7530 3896
rect 7650 3884 7656 3936
rect 7708 3924 7714 3936
rect 8297 3927 8355 3933
rect 8297 3924 8309 3927
rect 7708 3896 8309 3924
rect 7708 3884 7714 3896
rect 8297 3893 8309 3896
rect 8343 3893 8355 3927
rect 8496 3924 8524 4032
rect 8846 4020 8852 4072
rect 8904 4060 8910 4072
rect 11422 4069 11428 4072
rect 11368 4063 11428 4069
rect 11368 4060 11380 4063
rect 8904 4032 11380 4060
rect 8904 4020 8910 4032
rect 11368 4029 11380 4032
rect 11414 4029 11428 4063
rect 11368 4023 11428 4029
rect 11422 4020 11428 4023
rect 11480 4020 11486 4072
rect 9906 3995 9964 4001
rect 9906 3961 9918 3995
rect 9952 3992 9964 3995
rect 12360 3992 12388 4100
rect 13538 4088 13544 4100
rect 13596 4128 13602 4140
rect 13725 4131 13783 4137
rect 13725 4128 13737 4131
rect 13596 4100 13737 4128
rect 13596 4088 13602 4100
rect 13725 4097 13737 4100
rect 13771 4097 13783 4131
rect 13725 4091 13783 4097
rect 12713 4063 12771 4069
rect 12713 4029 12725 4063
rect 12759 4060 12771 4063
rect 13446 4060 13452 4072
rect 12759 4032 13452 4060
rect 12759 4029 12771 4032
rect 12713 4023 12771 4029
rect 13446 4020 13452 4032
rect 13504 4020 13510 4072
rect 12526 3992 12532 4004
rect 9952 3964 12388 3992
rect 12487 3964 12532 3992
rect 9952 3961 9964 3964
rect 9906 3955 9964 3961
rect 8754 3924 8760 3936
rect 8496 3896 8760 3924
rect 8297 3887 8355 3893
rect 8754 3884 8760 3896
rect 8812 3884 8818 3936
rect 8938 3884 8944 3936
rect 8996 3924 9002 3936
rect 9401 3927 9459 3933
rect 9401 3924 9413 3927
rect 8996 3896 9413 3924
rect 8996 3884 9002 3896
rect 9401 3893 9413 3896
rect 9447 3924 9459 3927
rect 9921 3924 9949 3955
rect 12526 3952 12532 3964
rect 12584 3952 12590 4004
rect 13740 3992 13768 4091
rect 13906 4060 13912 4072
rect 13867 4032 13912 4060
rect 13906 4020 13912 4032
rect 13964 4020 13970 4072
rect 18049 4063 18107 4069
rect 18049 4029 18061 4063
rect 18095 4060 18107 4063
rect 18230 4060 18236 4072
rect 18095 4032 18236 4060
rect 18095 4029 18107 4032
rect 18049 4023 18107 4029
rect 18230 4020 18236 4032
rect 18288 4020 18294 4072
rect 14230 3995 14288 4001
rect 14230 3992 14242 3995
rect 13740 3964 14242 3992
rect 14230 3961 14242 3964
rect 14276 3961 14288 3995
rect 14230 3955 14288 3961
rect 14918 3952 14924 4004
rect 14976 3992 14982 4004
rect 15749 3995 15807 4001
rect 15749 3992 15761 3995
rect 14976 3964 15761 3992
rect 14976 3952 14982 3964
rect 15749 3961 15761 3964
rect 15795 3961 15807 3995
rect 15749 3955 15807 3961
rect 15838 3952 15844 4004
rect 15896 3992 15902 4004
rect 15896 3964 15941 3992
rect 15896 3952 15902 3964
rect 16022 3952 16028 4004
rect 16080 3992 16086 4004
rect 16390 3992 16396 4004
rect 16080 3964 16396 3992
rect 16080 3952 16086 3964
rect 16390 3952 16396 3964
rect 16448 3952 16454 4004
rect 17773 3995 17831 4001
rect 17773 3992 17785 3995
rect 16960 3964 17785 3992
rect 16960 3936 16988 3964
rect 17773 3961 17785 3964
rect 17819 3992 17831 3995
rect 18370 3995 18428 4001
rect 18370 3992 18382 3995
rect 17819 3964 18382 3992
rect 17819 3961 17831 3964
rect 17773 3955 17831 3961
rect 18370 3961 18382 3964
rect 18416 3961 18428 3995
rect 18370 3955 18428 3961
rect 9447 3896 9949 3924
rect 9447 3893 9459 3896
rect 9401 3887 9459 3893
rect 10410 3884 10416 3936
rect 10468 3924 10474 3936
rect 12618 3924 12624 3936
rect 10468 3896 12624 3924
rect 10468 3884 10474 3896
rect 12618 3884 12624 3896
rect 12676 3924 12682 3936
rect 12805 3927 12863 3933
rect 12805 3924 12817 3927
rect 12676 3896 12817 3924
rect 12676 3884 12682 3896
rect 12805 3893 12817 3896
rect 12851 3893 12863 3927
rect 12805 3887 12863 3893
rect 16758 3884 16764 3936
rect 16816 3924 16822 3936
rect 16942 3924 16948 3936
rect 16816 3896 16948 3924
rect 16816 3884 16822 3896
rect 16942 3884 16948 3896
rect 17000 3884 17006 3936
rect 17126 3884 17132 3936
rect 17184 3924 17190 3936
rect 17221 3927 17279 3933
rect 17221 3924 17233 3927
rect 17184 3896 17233 3924
rect 17184 3884 17190 3896
rect 17221 3893 17233 3896
rect 17267 3893 17279 3927
rect 17221 3887 17279 3893
rect 1104 3834 20884 3856
rect 1104 3782 8315 3834
rect 8367 3782 8379 3834
rect 8431 3782 8443 3834
rect 8495 3782 8507 3834
rect 8559 3782 15648 3834
rect 15700 3782 15712 3834
rect 15764 3782 15776 3834
rect 15828 3782 15840 3834
rect 15892 3782 20884 3834
rect 1104 3760 20884 3782
rect 2774 3680 2780 3732
rect 2832 3720 2838 3732
rect 2869 3723 2927 3729
rect 2869 3720 2881 3723
rect 2832 3692 2881 3720
rect 2832 3680 2838 3692
rect 2869 3689 2881 3692
rect 2915 3689 2927 3723
rect 3510 3720 3516 3732
rect 3471 3692 3516 3720
rect 2869 3683 2927 3689
rect 3510 3680 3516 3692
rect 3568 3680 3574 3732
rect 3786 3720 3792 3732
rect 3747 3692 3792 3720
rect 3786 3680 3792 3692
rect 3844 3680 3850 3732
rect 3878 3680 3884 3732
rect 3936 3720 3942 3732
rect 4249 3723 4307 3729
rect 4249 3720 4261 3723
rect 3936 3692 4261 3720
rect 3936 3680 3942 3692
rect 4249 3689 4261 3692
rect 4295 3689 4307 3723
rect 4249 3683 4307 3689
rect 4982 3680 4988 3732
rect 5040 3720 5046 3732
rect 5905 3723 5963 3729
rect 5905 3720 5917 3723
rect 5040 3692 5917 3720
rect 5040 3680 5046 3692
rect 5905 3689 5917 3692
rect 5951 3689 5963 3723
rect 5905 3683 5963 3689
rect 6178 3680 6184 3732
rect 6236 3720 6242 3732
rect 7006 3720 7012 3732
rect 6236 3692 7012 3720
rect 6236 3680 6242 3692
rect 1397 3655 1455 3661
rect 1397 3621 1409 3655
rect 1443 3652 1455 3655
rect 4522 3652 4528 3664
rect 1443 3624 4528 3652
rect 1443 3621 1455 3624
rect 1397 3615 1455 3621
rect 4522 3612 4528 3624
rect 4580 3612 4586 3664
rect 4801 3655 4859 3661
rect 4801 3621 4813 3655
rect 4847 3652 4859 3655
rect 5258 3652 5264 3664
rect 4847 3624 5264 3652
rect 4847 3621 4859 3624
rect 4801 3615 4859 3621
rect 5258 3612 5264 3624
rect 5316 3652 5322 3664
rect 6273 3655 6331 3661
rect 6273 3652 6285 3655
rect 5316 3624 6285 3652
rect 5316 3612 5322 3624
rect 6273 3621 6285 3624
rect 6319 3621 6331 3655
rect 6273 3615 6331 3621
rect 2406 3584 2412 3596
rect 2367 3556 2412 3584
rect 2406 3544 2412 3556
rect 2464 3544 2470 3596
rect 2685 3587 2743 3593
rect 2685 3553 2697 3587
rect 2731 3584 2743 3587
rect 3418 3584 3424 3596
rect 2731 3556 3424 3584
rect 2731 3553 2743 3556
rect 2685 3547 2743 3553
rect 3418 3544 3424 3556
rect 3476 3584 3482 3596
rect 5534 3584 5540 3596
rect 3476 3556 4154 3584
rect 5495 3556 5540 3584
rect 3476 3544 3482 3556
rect 4126 3516 4154 3556
rect 5534 3544 5540 3556
rect 5592 3544 5598 3596
rect 6454 3584 6460 3596
rect 6415 3556 6460 3584
rect 6454 3544 6460 3556
rect 6512 3544 6518 3596
rect 6932 3593 6960 3692
rect 7006 3680 7012 3692
rect 7064 3680 7070 3732
rect 7282 3680 7288 3732
rect 7340 3720 7346 3732
rect 10134 3720 10140 3732
rect 7340 3692 10140 3720
rect 7340 3680 7346 3692
rect 7098 3612 7104 3664
rect 7156 3652 7162 3664
rect 8128 3661 8156 3692
rect 10134 3680 10140 3692
rect 10192 3680 10198 3732
rect 11238 3680 11244 3732
rect 11296 3720 11302 3732
rect 11885 3723 11943 3729
rect 11885 3720 11897 3723
rect 11296 3692 11897 3720
rect 11296 3680 11302 3692
rect 11885 3689 11897 3692
rect 11931 3689 11943 3723
rect 12526 3720 12532 3732
rect 12487 3692 12532 3720
rect 11885 3683 11943 3689
rect 12526 3680 12532 3692
rect 12584 3680 12590 3732
rect 13906 3680 13912 3732
rect 13964 3720 13970 3732
rect 14185 3723 14243 3729
rect 14185 3720 14197 3723
rect 13964 3692 14197 3720
rect 13964 3680 13970 3692
rect 14185 3689 14197 3692
rect 14231 3720 14243 3723
rect 14645 3723 14703 3729
rect 14645 3720 14657 3723
rect 14231 3692 14657 3720
rect 14231 3689 14243 3692
rect 14185 3683 14243 3689
rect 14645 3689 14657 3692
rect 14691 3689 14703 3723
rect 14645 3683 14703 3689
rect 15378 3680 15384 3732
rect 15436 3720 15442 3732
rect 15473 3723 15531 3729
rect 15473 3720 15485 3723
rect 15436 3692 15485 3720
rect 15436 3680 15442 3692
rect 15473 3689 15485 3692
rect 15519 3689 15531 3723
rect 16390 3720 16396 3732
rect 15473 3683 15531 3689
rect 15764 3692 16396 3720
rect 7193 3655 7251 3661
rect 7193 3652 7205 3655
rect 7156 3624 7205 3652
rect 7156 3612 7162 3624
rect 7193 3621 7205 3624
rect 7239 3652 7251 3655
rect 7837 3655 7895 3661
rect 7837 3652 7849 3655
rect 7239 3624 7849 3652
rect 7239 3621 7251 3624
rect 7193 3615 7251 3621
rect 7837 3621 7849 3624
rect 7883 3621 7895 3655
rect 7837 3615 7895 3621
rect 8113 3655 8171 3661
rect 8113 3621 8125 3655
rect 8159 3621 8171 3655
rect 8113 3615 8171 3621
rect 8205 3655 8263 3661
rect 8205 3621 8217 3655
rect 8251 3652 8263 3655
rect 8754 3652 8760 3664
rect 8251 3624 8760 3652
rect 8251 3621 8263 3624
rect 8205 3615 8263 3621
rect 8754 3612 8760 3624
rect 8812 3612 8818 3664
rect 9858 3652 9864 3664
rect 9819 3624 9864 3652
rect 9858 3612 9864 3624
rect 9916 3612 9922 3664
rect 9950 3612 9956 3664
rect 10008 3652 10014 3664
rect 15764 3661 15792 3692
rect 16390 3680 16396 3692
rect 16448 3720 16454 3732
rect 16669 3723 16727 3729
rect 16669 3720 16681 3723
rect 16448 3692 16681 3720
rect 16448 3680 16454 3692
rect 16669 3689 16681 3692
rect 16715 3689 16727 3723
rect 16669 3683 16727 3689
rect 18414 3680 18420 3732
rect 18472 3720 18478 3732
rect 18601 3723 18659 3729
rect 18601 3720 18613 3723
rect 18472 3692 18613 3720
rect 18472 3680 18478 3692
rect 18601 3689 18613 3692
rect 18647 3689 18659 3723
rect 19058 3720 19064 3732
rect 19019 3692 19064 3720
rect 18601 3683 18659 3689
rect 19058 3680 19064 3692
rect 19116 3680 19122 3732
rect 11149 3655 11207 3661
rect 11149 3652 11161 3655
rect 10008 3624 11161 3652
rect 10008 3612 10014 3624
rect 11149 3621 11161 3624
rect 11195 3621 11207 3655
rect 15749 3655 15807 3661
rect 11149 3615 11207 3621
rect 14108 3624 14412 3652
rect 6917 3587 6975 3593
rect 6917 3553 6929 3587
rect 6963 3553 6975 3587
rect 6917 3547 6975 3553
rect 7469 3587 7527 3593
rect 7469 3553 7481 3587
rect 7515 3584 7527 3587
rect 7650 3584 7656 3596
rect 7515 3556 7656 3584
rect 7515 3553 7527 3556
rect 7469 3547 7527 3553
rect 7650 3544 7656 3556
rect 7708 3544 7714 3596
rect 10778 3544 10784 3596
rect 10836 3584 10842 3596
rect 11238 3584 11244 3596
rect 10836 3556 11244 3584
rect 10836 3544 10842 3556
rect 11238 3544 11244 3556
rect 11296 3584 11302 3596
rect 11425 3587 11483 3593
rect 11425 3584 11437 3587
rect 11296 3556 11437 3584
rect 11296 3544 11302 3556
rect 11425 3553 11437 3556
rect 11471 3553 11483 3587
rect 11425 3547 11483 3553
rect 11701 3587 11759 3593
rect 11701 3553 11713 3587
rect 11747 3584 11759 3587
rect 11882 3584 11888 3596
rect 11747 3556 11888 3584
rect 11747 3553 11759 3556
rect 11701 3547 11759 3553
rect 11882 3544 11888 3556
rect 11940 3544 11946 3596
rect 12434 3544 12440 3596
rect 12492 3584 12498 3596
rect 13081 3587 13139 3593
rect 13081 3584 13093 3587
rect 12492 3556 13093 3584
rect 12492 3544 12498 3556
rect 13081 3553 13093 3556
rect 13127 3584 13139 3587
rect 13170 3584 13176 3596
rect 13127 3556 13176 3584
rect 13127 3553 13139 3556
rect 13081 3547 13139 3553
rect 13170 3544 13176 3556
rect 13228 3584 13234 3596
rect 13265 3587 13323 3593
rect 13265 3584 13277 3587
rect 13228 3556 13277 3584
rect 13228 3544 13234 3556
rect 13265 3553 13277 3556
rect 13311 3553 13323 3587
rect 13265 3547 13323 3553
rect 13354 3544 13360 3596
rect 13412 3584 13418 3596
rect 14108 3593 14136 3624
rect 14093 3587 14151 3593
rect 14093 3584 14105 3587
rect 13412 3556 14105 3584
rect 13412 3544 13418 3556
rect 14093 3553 14105 3556
rect 14139 3553 14151 3587
rect 14274 3584 14280 3596
rect 14235 3556 14280 3584
rect 14093 3547 14151 3553
rect 14274 3544 14280 3556
rect 14332 3544 14338 3596
rect 5629 3519 5687 3525
rect 5629 3516 5641 3519
rect 4126 3488 5641 3516
rect 5629 3485 5641 3488
rect 5675 3516 5687 3519
rect 7558 3516 7564 3528
rect 5675 3488 7564 3516
rect 5675 3485 5687 3488
rect 5629 3479 5687 3485
rect 7558 3476 7564 3488
rect 7616 3476 7622 3528
rect 8757 3519 8815 3525
rect 8757 3485 8769 3519
rect 8803 3516 8815 3519
rect 9582 3516 9588 3528
rect 8803 3488 9588 3516
rect 8803 3485 8815 3488
rect 8757 3479 8815 3485
rect 9582 3476 9588 3488
rect 9640 3516 9646 3528
rect 9769 3519 9827 3525
rect 9769 3516 9781 3519
rect 9640 3488 9781 3516
rect 9640 3476 9646 3488
rect 9769 3485 9781 3488
rect 9815 3485 9827 3519
rect 9769 3479 9827 3485
rect 12618 3476 12624 3528
rect 12676 3516 12682 3528
rect 13630 3516 13636 3528
rect 12676 3488 13636 3516
rect 12676 3476 12682 3488
rect 13630 3476 13636 3488
rect 13688 3516 13694 3528
rect 14292 3516 14320 3544
rect 13688 3488 14320 3516
rect 13688 3476 13694 3488
rect 1762 3408 1768 3460
rect 1820 3448 1826 3460
rect 2498 3448 2504 3460
rect 1820 3420 2504 3448
rect 1820 3408 1826 3420
rect 2498 3408 2504 3420
rect 2556 3408 2562 3460
rect 9674 3448 9680 3460
rect 9587 3420 9680 3448
rect 9674 3408 9680 3420
rect 9732 3448 9738 3460
rect 10318 3448 10324 3460
rect 9732 3420 10324 3448
rect 9732 3408 9738 3420
rect 10318 3408 10324 3420
rect 10376 3408 10382 3460
rect 10870 3448 10876 3460
rect 10783 3420 10876 3448
rect 10870 3408 10876 3420
rect 10928 3448 10934 3460
rect 11517 3451 11575 3457
rect 11517 3448 11529 3451
rect 10928 3420 11529 3448
rect 10928 3408 10934 3420
rect 11517 3417 11529 3420
rect 11563 3448 11575 3451
rect 12342 3448 12348 3460
rect 11563 3420 12348 3448
rect 11563 3417 11575 3420
rect 11517 3411 11575 3417
rect 12342 3408 12348 3420
rect 12400 3408 12406 3460
rect 14384 3448 14412 3624
rect 15749 3621 15761 3655
rect 15795 3621 15807 3655
rect 15749 3615 15807 3621
rect 15838 3612 15844 3664
rect 15896 3652 15902 3664
rect 17218 3652 17224 3664
rect 15896 3624 15941 3652
rect 16408 3624 17224 3652
rect 15896 3612 15902 3624
rect 16408 3596 16436 3624
rect 17218 3612 17224 3624
rect 17276 3612 17282 3664
rect 17402 3612 17408 3664
rect 17460 3652 17466 3664
rect 19150 3652 19156 3664
rect 17460 3624 19156 3652
rect 17460 3612 17466 3624
rect 19150 3612 19156 3624
rect 19208 3652 19214 3664
rect 19208 3624 19288 3652
rect 19208 3612 19214 3624
rect 16390 3544 16396 3596
rect 16448 3584 16454 3596
rect 17310 3584 17316 3596
rect 16448 3556 16541 3584
rect 17271 3556 17316 3584
rect 16448 3544 16454 3556
rect 17310 3544 17316 3556
rect 17368 3544 17374 3596
rect 18785 3587 18843 3593
rect 18785 3584 18797 3587
rect 18385 3556 18797 3584
rect 14550 3476 14556 3528
rect 14608 3516 14614 3528
rect 15838 3516 15844 3528
rect 14608 3488 15844 3516
rect 14608 3476 14614 3488
rect 15838 3476 15844 3488
rect 15896 3476 15902 3528
rect 16206 3476 16212 3528
rect 16264 3516 16270 3528
rect 17221 3519 17279 3525
rect 17221 3516 17233 3519
rect 16264 3488 17233 3516
rect 16264 3476 16270 3488
rect 17221 3485 17233 3488
rect 17267 3485 17279 3519
rect 17221 3479 17279 3485
rect 16758 3448 16764 3460
rect 14384 3420 16764 3448
rect 16758 3408 16764 3420
rect 16816 3408 16822 3460
rect 16850 3408 16856 3460
rect 16908 3448 16914 3460
rect 18385 3448 18413 3556
rect 18785 3553 18797 3556
rect 18831 3584 18843 3587
rect 19058 3584 19064 3596
rect 18831 3556 19064 3584
rect 18831 3553 18843 3556
rect 18785 3547 18843 3553
rect 19058 3544 19064 3556
rect 19116 3544 19122 3596
rect 19260 3593 19288 3624
rect 19245 3587 19303 3593
rect 19245 3553 19257 3587
rect 19291 3553 19303 3587
rect 19245 3547 19303 3553
rect 16908 3420 18413 3448
rect 16908 3408 16914 3420
rect 2133 3383 2191 3389
rect 2133 3349 2145 3383
rect 2179 3380 2191 3383
rect 2314 3380 2320 3392
rect 2179 3352 2320 3380
rect 2179 3349 2191 3352
rect 2133 3343 2191 3349
rect 2314 3340 2320 3352
rect 2372 3380 2378 3392
rect 5534 3380 5540 3392
rect 2372 3352 5540 3380
rect 2372 3340 2378 3352
rect 5534 3340 5540 3352
rect 5592 3340 5598 3392
rect 9030 3380 9036 3392
rect 8991 3352 9036 3380
rect 9030 3340 9036 3352
rect 9088 3340 9094 3392
rect 9306 3340 9312 3392
rect 9364 3380 9370 3392
rect 9401 3383 9459 3389
rect 9401 3380 9413 3383
rect 9364 3352 9413 3380
rect 9364 3340 9370 3352
rect 9401 3349 9413 3352
rect 9447 3349 9459 3383
rect 9401 3343 9459 3349
rect 14918 3340 14924 3392
rect 14976 3380 14982 3392
rect 15013 3383 15071 3389
rect 15013 3380 15025 3383
rect 14976 3352 15025 3380
rect 14976 3340 14982 3352
rect 15013 3349 15025 3352
rect 15059 3349 15071 3383
rect 18230 3380 18236 3392
rect 18191 3352 18236 3380
rect 15013 3343 15071 3349
rect 18230 3340 18236 3352
rect 18288 3340 18294 3392
rect 1104 3290 20884 3312
rect 1104 3238 4648 3290
rect 4700 3238 4712 3290
rect 4764 3238 4776 3290
rect 4828 3238 4840 3290
rect 4892 3238 11982 3290
rect 12034 3238 12046 3290
rect 12098 3238 12110 3290
rect 12162 3238 12174 3290
rect 12226 3238 19315 3290
rect 19367 3238 19379 3290
rect 19431 3238 19443 3290
rect 19495 3238 19507 3290
rect 19559 3238 20884 3290
rect 1104 3216 20884 3238
rect 2406 3136 2412 3188
rect 2464 3176 2470 3188
rect 3053 3179 3111 3185
rect 3053 3176 3065 3179
rect 2464 3148 3065 3176
rect 2464 3136 2470 3148
rect 3053 3145 3065 3148
rect 3099 3145 3111 3179
rect 3418 3176 3424 3188
rect 3379 3148 3424 3176
rect 3053 3139 3111 3145
rect 3068 3108 3096 3139
rect 3418 3136 3424 3148
rect 3476 3136 3482 3188
rect 4985 3179 5043 3185
rect 4985 3145 4997 3179
rect 5031 3176 5043 3179
rect 5534 3176 5540 3188
rect 5031 3148 5540 3176
rect 5031 3145 5043 3148
rect 4985 3139 5043 3145
rect 5534 3136 5540 3148
rect 5592 3136 5598 3188
rect 6178 3136 6184 3188
rect 6236 3176 6242 3188
rect 6457 3179 6515 3185
rect 6457 3176 6469 3179
rect 6236 3148 6469 3176
rect 6236 3136 6242 3148
rect 6457 3145 6469 3148
rect 6503 3145 6515 3179
rect 6457 3139 6515 3145
rect 7190 3136 7196 3188
rect 7248 3176 7254 3188
rect 8846 3176 8852 3188
rect 7248 3148 8852 3176
rect 7248 3136 7254 3148
rect 8846 3136 8852 3148
rect 8904 3136 8910 3188
rect 9125 3179 9183 3185
rect 9125 3145 9137 3179
rect 9171 3176 9183 3179
rect 9858 3176 9864 3188
rect 9171 3148 9864 3176
rect 9171 3145 9183 3148
rect 9125 3139 9183 3145
rect 9858 3136 9864 3148
rect 9916 3136 9922 3188
rect 10134 3176 10140 3188
rect 10095 3148 10140 3176
rect 10134 3136 10140 3148
rect 10192 3136 10198 3188
rect 11238 3136 11244 3188
rect 11296 3176 11302 3188
rect 11609 3179 11667 3185
rect 11609 3176 11621 3179
rect 11296 3148 11621 3176
rect 11296 3136 11302 3148
rect 11609 3145 11621 3148
rect 11655 3145 11667 3179
rect 11609 3139 11667 3145
rect 12253 3179 12311 3185
rect 12253 3145 12265 3179
rect 12299 3176 12311 3179
rect 12342 3176 12348 3188
rect 12299 3148 12348 3176
rect 12299 3145 12311 3148
rect 12253 3139 12311 3145
rect 12342 3136 12348 3148
rect 12400 3136 12406 3188
rect 12618 3176 12624 3188
rect 12579 3148 12624 3176
rect 12618 3136 12624 3148
rect 12676 3136 12682 3188
rect 14274 3136 14280 3188
rect 14332 3176 14338 3188
rect 14553 3179 14611 3185
rect 14553 3176 14565 3179
rect 14332 3148 14565 3176
rect 14332 3136 14338 3148
rect 14553 3145 14565 3148
rect 14599 3145 14611 3179
rect 14553 3139 14611 3145
rect 15838 3136 15844 3188
rect 15896 3176 15902 3188
rect 17037 3179 17095 3185
rect 17037 3176 17049 3179
rect 15896 3148 17049 3176
rect 15896 3136 15902 3148
rect 17037 3145 17049 3148
rect 17083 3176 17095 3179
rect 17310 3176 17316 3188
rect 17083 3148 17316 3176
rect 17083 3145 17095 3148
rect 17037 3139 17095 3145
rect 17310 3136 17316 3148
rect 17368 3176 17374 3188
rect 17405 3179 17463 3185
rect 17405 3176 17417 3179
rect 17368 3148 17417 3176
rect 17368 3136 17374 3148
rect 17405 3145 17417 3148
rect 17451 3145 17463 3179
rect 19150 3176 19156 3188
rect 19111 3148 19156 3176
rect 17405 3139 17463 3145
rect 19150 3136 19156 3148
rect 19208 3136 19214 3188
rect 7929 3111 7987 3117
rect 7929 3108 7941 3111
rect 3068 3080 7941 3108
rect 7929 3077 7941 3080
rect 7975 3077 7987 3111
rect 7929 3071 7987 3077
rect 8754 3068 8760 3120
rect 8812 3108 8818 3120
rect 9401 3111 9459 3117
rect 9401 3108 9413 3111
rect 8812 3080 9413 3108
rect 8812 3068 8818 3080
rect 9401 3077 9413 3080
rect 9447 3077 9459 3111
rect 10870 3108 10876 3120
rect 10831 3080 10876 3108
rect 9401 3071 9459 3077
rect 10870 3068 10876 3080
rect 10928 3068 10934 3120
rect 12989 3111 13047 3117
rect 12989 3108 13001 3111
rect 10980 3080 13001 3108
rect 2777 3043 2835 3049
rect 2777 3009 2789 3043
rect 2823 3040 2835 3043
rect 8205 3043 8263 3049
rect 8205 3040 8217 3043
rect 2823 3012 8217 3040
rect 2823 3009 2835 3012
rect 2777 3003 2835 3009
rect 8205 3009 8217 3012
rect 8251 3040 8263 3043
rect 9030 3040 9036 3052
rect 8251 3012 9036 3040
rect 8251 3009 8263 3012
rect 8205 3003 8263 3009
rect 9030 3000 9036 3012
rect 9088 3000 9094 3052
rect 10980 3040 11008 3080
rect 12989 3077 13001 3080
rect 13035 3108 13047 3111
rect 13354 3108 13360 3120
rect 13035 3080 13360 3108
rect 13035 3077 13047 3080
rect 12989 3071 13047 3077
rect 13354 3068 13360 3080
rect 13412 3068 13418 3120
rect 15013 3111 15071 3117
rect 15013 3077 15025 3111
rect 15059 3108 15071 3111
rect 15059 3080 16528 3108
rect 15059 3077 15071 3080
rect 15013 3071 15071 3077
rect 11514 3040 11520 3052
rect 10796 3012 11008 3040
rect 11475 3012 11520 3040
rect 10796 2984 10824 3012
rect 11514 3000 11520 3012
rect 11572 3000 11578 3052
rect 11609 3043 11667 3049
rect 11609 3009 11621 3043
rect 11655 3040 11667 3043
rect 11655 3012 14044 3040
rect 11655 3009 11667 3012
rect 11609 3003 11667 3009
rect 2317 2975 2375 2981
rect 2317 2941 2329 2975
rect 2363 2941 2375 2975
rect 2317 2935 2375 2941
rect 2593 2975 2651 2981
rect 2593 2941 2605 2975
rect 2639 2972 2651 2975
rect 3142 2972 3148 2984
rect 2639 2944 3148 2972
rect 2639 2941 2651 2944
rect 2593 2935 2651 2941
rect 2332 2904 2360 2935
rect 3142 2932 3148 2944
rect 3200 2932 3206 2984
rect 3786 2972 3792 2984
rect 3747 2944 3792 2972
rect 3786 2932 3792 2944
rect 3844 2932 3850 2984
rect 4154 2932 4160 2984
rect 4212 2972 4218 2984
rect 4212 2944 4257 2972
rect 4212 2932 4218 2944
rect 4982 2932 4988 2984
rect 5040 2972 5046 2984
rect 5169 2975 5227 2981
rect 5169 2972 5181 2975
rect 5040 2944 5181 2972
rect 5040 2932 5046 2944
rect 5169 2941 5181 2944
rect 5215 2941 5227 2975
rect 5718 2972 5724 2984
rect 5679 2944 5724 2972
rect 5169 2935 5227 2941
rect 5718 2932 5724 2944
rect 5776 2932 5782 2984
rect 5902 2972 5908 2984
rect 5863 2944 5908 2972
rect 5902 2932 5908 2944
rect 5960 2932 5966 2984
rect 6822 2932 6828 2984
rect 6880 2972 6886 2984
rect 7101 2975 7159 2981
rect 7101 2972 7113 2975
rect 6880 2944 7113 2972
rect 6880 2932 6886 2944
rect 7101 2941 7113 2944
rect 7147 2972 7159 2975
rect 7653 2975 7711 2981
rect 7653 2972 7665 2975
rect 7147 2944 7665 2972
rect 7147 2941 7159 2944
rect 7101 2935 7159 2941
rect 7653 2941 7665 2944
rect 7699 2941 7711 2975
rect 10778 2972 10784 2984
rect 7653 2935 7711 2941
rect 7760 2944 8708 2972
rect 10739 2944 10784 2972
rect 3878 2904 3884 2916
rect 2332 2876 3884 2904
rect 3878 2864 3884 2876
rect 3936 2864 3942 2916
rect 4338 2864 4344 2916
rect 4396 2904 4402 2916
rect 4396 2876 4441 2904
rect 4396 2864 4402 2876
rect 4522 2864 4528 2916
rect 4580 2904 4586 2916
rect 7760 2904 7788 2944
rect 8570 2913 8576 2916
rect 4580 2876 7788 2904
rect 7929 2907 7987 2913
rect 4580 2864 4586 2876
rect 7929 2873 7941 2907
rect 7975 2904 7987 2907
rect 8567 2904 8576 2913
rect 7975 2876 8293 2904
rect 8531 2876 8576 2904
rect 7975 2873 7987 2876
rect 7929 2867 7987 2873
rect 1762 2796 1768 2848
rect 1820 2836 1826 2848
rect 1857 2839 1915 2845
rect 1857 2836 1869 2839
rect 1820 2808 1869 2836
rect 1820 2796 1826 2808
rect 1857 2805 1869 2808
rect 1903 2805 1915 2839
rect 7282 2836 7288 2848
rect 7243 2808 7288 2836
rect 1857 2799 1915 2805
rect 7282 2796 7288 2808
rect 7340 2796 7346 2848
rect 7742 2796 7748 2848
rect 7800 2836 7806 2848
rect 8021 2839 8079 2845
rect 8021 2836 8033 2839
rect 7800 2808 8033 2836
rect 7800 2796 7806 2808
rect 8021 2805 8033 2808
rect 8067 2805 8079 2839
rect 8265 2836 8293 2876
rect 8567 2867 8576 2876
rect 8570 2864 8576 2867
rect 8628 2864 8634 2916
rect 8680 2904 8708 2944
rect 10778 2932 10784 2944
rect 10836 2932 10842 2984
rect 10870 2932 10876 2984
rect 10928 2972 10934 2984
rect 11057 2975 11115 2981
rect 11057 2972 11069 2975
rect 10928 2944 11069 2972
rect 10928 2932 10934 2944
rect 11057 2941 11069 2944
rect 11103 2972 11115 2975
rect 11882 2972 11888 2984
rect 11103 2944 11888 2972
rect 11103 2941 11115 2944
rect 11057 2935 11115 2941
rect 11882 2932 11888 2944
rect 11940 2932 11946 2984
rect 13170 2972 13176 2984
rect 13131 2944 13176 2972
rect 13170 2932 13176 2944
rect 13228 2932 13234 2984
rect 13630 2972 13636 2984
rect 13591 2944 13636 2972
rect 13630 2932 13636 2944
rect 13688 2932 13694 2984
rect 14016 2981 14044 3012
rect 14001 2975 14059 2981
rect 14001 2941 14013 2975
rect 14047 2972 14059 2975
rect 15028 2972 15056 3071
rect 16390 3040 16396 3052
rect 16351 3012 16396 3040
rect 16390 3000 16396 3012
rect 16448 3000 16454 3052
rect 16500 3040 16528 3080
rect 17586 3068 17592 3120
rect 17644 3108 17650 3120
rect 19751 3111 19809 3117
rect 19751 3108 19763 3111
rect 17644 3080 19763 3108
rect 17644 3068 17650 3080
rect 19751 3077 19763 3080
rect 19797 3077 19809 3111
rect 19751 3071 19809 3077
rect 18049 3043 18107 3049
rect 18049 3040 18061 3043
rect 16500 3012 18061 3040
rect 18049 3009 18061 3012
rect 18095 3009 18107 3043
rect 18049 3003 18107 3009
rect 19058 3000 19064 3052
rect 19116 3040 19122 3052
rect 19429 3043 19487 3049
rect 19429 3040 19441 3043
rect 19116 3012 19441 3040
rect 19116 3000 19122 3012
rect 19429 3009 19441 3012
rect 19475 3009 19487 3043
rect 19429 3003 19487 3009
rect 14047 2944 15056 2972
rect 14047 2941 14059 2944
rect 14001 2935 14059 2941
rect 16758 2932 16764 2984
rect 16816 2972 16822 2984
rect 17865 2975 17923 2981
rect 17865 2972 17877 2975
rect 16816 2944 17877 2972
rect 16816 2932 16822 2944
rect 17865 2941 17877 2944
rect 17911 2972 17923 2975
rect 18690 2972 18696 2984
rect 17911 2944 18696 2972
rect 17911 2941 17923 2944
rect 17865 2935 17923 2941
rect 18690 2932 18696 2944
rect 18748 2932 18754 2984
rect 19702 2981 19708 2984
rect 19680 2975 19708 2981
rect 19680 2941 19692 2975
rect 19760 2972 19766 2984
rect 20073 2975 20131 2981
rect 20073 2972 20085 2975
rect 19760 2944 20085 2972
rect 19680 2935 19708 2941
rect 19702 2932 19708 2935
rect 19760 2932 19766 2944
rect 20073 2941 20085 2944
rect 20119 2941 20131 2975
rect 20073 2935 20131 2941
rect 15473 2907 15531 2913
rect 15473 2904 15485 2907
rect 8680 2876 15485 2904
rect 15473 2873 15485 2876
rect 15519 2904 15531 2907
rect 16117 2907 16175 2913
rect 16117 2904 16129 2907
rect 15519 2876 16129 2904
rect 15519 2873 15531 2876
rect 15473 2867 15531 2873
rect 16117 2873 16129 2876
rect 16163 2873 16175 2907
rect 16117 2867 16175 2873
rect 16206 2864 16212 2916
rect 16264 2904 16270 2916
rect 16264 2876 16309 2904
rect 16264 2864 16270 2876
rect 10597 2839 10655 2845
rect 10597 2836 10609 2839
rect 8265 2808 10609 2836
rect 8021 2799 8079 2805
rect 10597 2805 10609 2808
rect 10643 2836 10655 2839
rect 10778 2836 10784 2848
rect 10643 2808 10784 2836
rect 10643 2805 10655 2808
rect 10597 2799 10655 2805
rect 10778 2796 10784 2808
rect 10836 2796 10842 2848
rect 11882 2836 11888 2848
rect 11843 2808 11888 2836
rect 11882 2796 11888 2808
rect 11940 2796 11946 2848
rect 14274 2836 14280 2848
rect 14235 2808 14280 2836
rect 14274 2796 14280 2808
rect 14332 2796 14338 2848
rect 15933 2839 15991 2845
rect 15933 2805 15945 2839
rect 15979 2836 15991 2839
rect 16224 2836 16252 2864
rect 15979 2808 16252 2836
rect 15979 2805 15991 2808
rect 15933 2799 15991 2805
rect 1104 2746 20884 2768
rect 1104 2694 8315 2746
rect 8367 2694 8379 2746
rect 8431 2694 8443 2746
rect 8495 2694 8507 2746
rect 8559 2694 15648 2746
rect 15700 2694 15712 2746
rect 15764 2694 15776 2746
rect 15828 2694 15840 2746
rect 15892 2694 20884 2746
rect 1104 2672 20884 2694
rect 1854 2632 1860 2644
rect 1815 2604 1860 2632
rect 1854 2592 1860 2604
rect 1912 2592 1918 2644
rect 2317 2635 2375 2641
rect 2317 2601 2329 2635
rect 2363 2632 2375 2635
rect 3142 2632 3148 2644
rect 2363 2604 3148 2632
rect 2363 2601 2375 2604
rect 2317 2595 2375 2601
rect 3142 2592 3148 2604
rect 3200 2632 3206 2644
rect 3421 2635 3479 2641
rect 3421 2632 3433 2635
rect 3200 2604 3433 2632
rect 3200 2592 3206 2604
rect 3421 2601 3433 2604
rect 3467 2601 3479 2635
rect 3786 2632 3792 2644
rect 3747 2604 3792 2632
rect 3421 2595 3479 2601
rect 3786 2592 3792 2604
rect 3844 2592 3850 2644
rect 4154 2592 4160 2644
rect 4212 2632 4218 2644
rect 4801 2635 4859 2641
rect 4801 2632 4813 2635
rect 4212 2604 4813 2632
rect 4212 2592 4218 2604
rect 4801 2601 4813 2604
rect 4847 2632 4859 2635
rect 5718 2632 5724 2644
rect 4847 2604 5724 2632
rect 4847 2601 4859 2604
rect 4801 2595 4859 2601
rect 5718 2592 5724 2604
rect 5776 2592 5782 2644
rect 6454 2632 6460 2644
rect 6415 2604 6460 2632
rect 6454 2592 6460 2604
rect 6512 2592 6518 2644
rect 6917 2635 6975 2641
rect 6917 2601 6929 2635
rect 6963 2632 6975 2635
rect 9401 2635 9459 2641
rect 9401 2632 9413 2635
rect 6963 2604 9413 2632
rect 6963 2601 6975 2604
rect 6917 2595 6975 2601
rect 9401 2601 9413 2604
rect 9447 2632 9459 2635
rect 9493 2635 9551 2641
rect 9493 2632 9505 2635
rect 9447 2604 9505 2632
rect 9447 2601 9459 2604
rect 9401 2595 9459 2601
rect 9493 2601 9505 2604
rect 9539 2601 9551 2635
rect 10870 2632 10876 2644
rect 10831 2604 10876 2632
rect 9493 2595 9551 2601
rect 10870 2592 10876 2604
rect 10928 2592 10934 2644
rect 11238 2632 11244 2644
rect 11199 2604 11244 2632
rect 11238 2592 11244 2604
rect 11296 2592 11302 2644
rect 13170 2632 13176 2644
rect 13131 2604 13176 2632
rect 13170 2592 13176 2604
rect 13228 2592 13234 2644
rect 13538 2632 13544 2644
rect 13499 2604 13544 2632
rect 13538 2592 13544 2604
rect 13596 2592 13602 2644
rect 14274 2632 14280 2644
rect 13648 2604 14280 2632
rect 3804 2564 3832 2592
rect 2700 2536 3832 2564
rect 4387 2567 4445 2573
rect 2700 2505 2728 2536
rect 4387 2533 4399 2567
rect 4433 2564 4445 2567
rect 5902 2564 5908 2576
rect 4433 2536 5908 2564
rect 4433 2533 4445 2536
rect 4387 2527 4445 2533
rect 5902 2524 5908 2536
rect 5960 2524 5966 2576
rect 5997 2567 6055 2573
rect 5997 2533 6009 2567
rect 6043 2564 6055 2567
rect 6362 2564 6368 2576
rect 6043 2536 6368 2564
rect 6043 2533 6055 2536
rect 5997 2527 6055 2533
rect 6362 2524 6368 2536
rect 6420 2524 6426 2576
rect 7469 2567 7527 2573
rect 7469 2533 7481 2567
rect 7515 2564 7527 2567
rect 7650 2564 7656 2576
rect 7515 2536 7656 2564
rect 7515 2533 7527 2536
rect 7469 2527 7527 2533
rect 2685 2499 2743 2505
rect 2685 2465 2697 2499
rect 2731 2465 2743 2499
rect 2685 2459 2743 2465
rect 2961 2499 3019 2505
rect 2961 2465 2973 2499
rect 3007 2496 3019 2499
rect 3050 2496 3056 2508
rect 3007 2468 3056 2496
rect 3007 2465 3019 2468
rect 2961 2459 3019 2465
rect 3050 2456 3056 2468
rect 3108 2456 3114 2508
rect 4062 2456 4068 2508
rect 4120 2496 4126 2508
rect 4157 2499 4215 2505
rect 4157 2496 4169 2499
rect 4120 2468 4169 2496
rect 4120 2456 4126 2468
rect 4157 2465 4169 2468
rect 4203 2465 4215 2499
rect 4157 2459 4215 2465
rect 5169 2499 5227 2505
rect 5169 2465 5181 2499
rect 5215 2496 5227 2499
rect 5353 2499 5411 2505
rect 5353 2496 5365 2499
rect 5215 2468 5365 2496
rect 5215 2465 5227 2468
rect 5169 2459 5227 2465
rect 5353 2465 5365 2468
rect 5399 2465 5411 2499
rect 5353 2459 5411 2465
rect 1394 2428 1400 2440
rect 1355 2400 1400 2428
rect 1394 2388 1400 2400
rect 1452 2388 1458 2440
rect 3145 2431 3203 2437
rect 3145 2397 3157 2431
rect 3191 2428 3203 2431
rect 4985 2431 5043 2437
rect 4985 2428 4997 2431
rect 3191 2400 4997 2428
rect 3191 2397 3203 2400
rect 3145 2391 3203 2397
rect 4985 2397 4997 2400
rect 5031 2397 5043 2431
rect 4985 2391 5043 2397
rect 3970 2320 3976 2372
rect 4028 2360 4034 2372
rect 5184 2360 5212 2459
rect 5718 2456 5724 2508
rect 5776 2496 5782 2508
rect 7484 2496 7512 2527
rect 7650 2524 7656 2536
rect 7708 2524 7714 2576
rect 7742 2524 7748 2576
rect 7800 2564 7806 2576
rect 8250 2567 8308 2573
rect 8250 2564 8262 2567
rect 7800 2536 8262 2564
rect 7800 2524 7806 2536
rect 8250 2533 8262 2536
rect 8296 2564 8308 2567
rect 8662 2564 8668 2576
rect 8296 2536 8668 2564
rect 8296 2533 8308 2536
rect 8250 2527 8308 2533
rect 8662 2524 8668 2536
rect 8720 2524 8726 2576
rect 9217 2567 9275 2573
rect 9217 2564 9229 2567
rect 8864 2536 9229 2564
rect 8864 2505 8892 2536
rect 9217 2533 9229 2536
rect 9263 2564 9275 2567
rect 9953 2567 10011 2573
rect 9953 2564 9965 2567
rect 9263 2536 9965 2564
rect 9263 2533 9275 2536
rect 9217 2527 9275 2533
rect 9953 2533 9965 2536
rect 9999 2533 10011 2567
rect 9953 2527 10011 2533
rect 5776 2468 7512 2496
rect 8849 2499 8907 2505
rect 5776 2456 5782 2468
rect 8849 2465 8861 2499
rect 8895 2465 8907 2499
rect 11422 2496 11428 2508
rect 11383 2468 11428 2496
rect 8849 2459 8907 2465
rect 11422 2456 11428 2468
rect 11480 2496 11486 2508
rect 11977 2499 12035 2505
rect 11977 2496 11989 2499
rect 11480 2468 11989 2496
rect 11480 2456 11486 2468
rect 11977 2465 11989 2468
rect 12023 2465 12035 2499
rect 12434 2496 12440 2508
rect 12395 2468 12440 2496
rect 11977 2459 12035 2465
rect 12434 2456 12440 2468
rect 12492 2496 12498 2508
rect 13648 2505 13676 2604
rect 14274 2592 14280 2604
rect 14332 2632 14338 2644
rect 14829 2635 14887 2641
rect 14829 2632 14841 2635
rect 14332 2604 14841 2632
rect 14332 2592 14338 2604
rect 14829 2601 14841 2604
rect 14875 2601 14887 2635
rect 14829 2595 14887 2601
rect 15611 2635 15669 2641
rect 15611 2601 15623 2635
rect 15657 2632 15669 2635
rect 18138 2632 18144 2644
rect 15657 2604 18144 2632
rect 15657 2601 15669 2604
rect 15611 2595 15669 2601
rect 18138 2592 18144 2604
rect 18196 2592 18202 2644
rect 13814 2524 13820 2576
rect 13872 2564 13878 2576
rect 13954 2567 14012 2573
rect 13954 2564 13966 2567
rect 13872 2536 13966 2564
rect 13872 2524 13878 2536
rect 13954 2533 13966 2536
rect 14000 2533 14012 2567
rect 16574 2564 16580 2576
rect 13954 2527 14012 2533
rect 15396 2536 16580 2564
rect 12656 2499 12714 2505
rect 12656 2496 12668 2499
rect 12492 2468 12668 2496
rect 12492 2456 12498 2468
rect 12656 2465 12668 2468
rect 12702 2465 12714 2499
rect 12656 2459 12714 2465
rect 13633 2499 13691 2505
rect 13633 2465 13645 2499
rect 13679 2465 13691 2499
rect 15396 2496 15424 2536
rect 16574 2524 16580 2536
rect 16632 2524 16638 2576
rect 16806 2567 16864 2573
rect 16806 2564 16818 2567
rect 16684 2536 16818 2564
rect 13633 2459 13691 2465
rect 13786 2468 15424 2496
rect 15540 2499 15598 2505
rect 7929 2431 7987 2437
rect 7929 2428 7941 2431
rect 4028 2332 5212 2360
rect 7116 2400 7941 2428
rect 4028 2320 4034 2332
rect 4985 2295 5043 2301
rect 4985 2261 4997 2295
rect 5031 2292 5043 2295
rect 7116 2292 7144 2400
rect 7929 2397 7941 2400
rect 7975 2428 7987 2431
rect 9306 2428 9312 2440
rect 7975 2400 9312 2428
rect 7975 2397 7987 2400
rect 7929 2391 7987 2397
rect 9306 2388 9312 2400
rect 9364 2388 9370 2440
rect 9401 2431 9459 2437
rect 9401 2397 9413 2431
rect 9447 2428 9459 2431
rect 9861 2431 9919 2437
rect 9861 2428 9873 2431
rect 9447 2400 9873 2428
rect 9447 2397 9459 2400
rect 9401 2391 9459 2397
rect 9861 2397 9873 2400
rect 9907 2397 9919 2431
rect 10318 2428 10324 2440
rect 10279 2400 10324 2428
rect 9861 2391 9919 2397
rect 10318 2388 10324 2400
rect 10376 2388 10382 2440
rect 12759 2431 12817 2437
rect 12759 2397 12771 2431
rect 12805 2428 12817 2431
rect 13786 2428 13814 2468
rect 15540 2465 15552 2499
rect 15586 2496 15598 2499
rect 15930 2496 15936 2508
rect 15586 2468 15936 2496
rect 15586 2465 15598 2468
rect 15540 2459 15598 2465
rect 15930 2456 15936 2468
rect 15988 2456 15994 2508
rect 16485 2431 16543 2437
rect 16485 2428 16497 2431
rect 12805 2400 13814 2428
rect 15212 2400 16497 2428
rect 12805 2397 12817 2400
rect 12759 2391 12817 2397
rect 11609 2363 11667 2369
rect 11609 2329 11621 2363
rect 11655 2360 11667 2363
rect 15010 2360 15016 2372
rect 11655 2332 15016 2360
rect 11655 2329 11667 2332
rect 11609 2323 11667 2329
rect 15010 2320 15016 2332
rect 15068 2320 15074 2372
rect 15212 2304 15240 2400
rect 16485 2397 16497 2400
rect 16531 2397 16543 2431
rect 16485 2391 16543 2397
rect 16301 2363 16359 2369
rect 16301 2329 16313 2363
rect 16347 2360 16359 2363
rect 16684 2360 16712 2536
rect 16806 2533 16818 2536
rect 16852 2564 16864 2567
rect 16942 2564 16948 2576
rect 16852 2536 16948 2564
rect 16852 2533 16864 2536
rect 16806 2527 16864 2533
rect 16942 2524 16948 2536
rect 17000 2524 17006 2576
rect 17773 2567 17831 2573
rect 17773 2533 17785 2567
rect 17819 2564 17831 2567
rect 18509 2567 18567 2573
rect 18509 2564 18521 2567
rect 17819 2536 18521 2564
rect 17819 2533 17831 2536
rect 17773 2527 17831 2533
rect 18509 2533 18521 2536
rect 18555 2533 18567 2567
rect 18509 2527 18567 2533
rect 17405 2499 17463 2505
rect 17405 2465 17417 2499
rect 17451 2496 17463 2499
rect 17788 2496 17816 2527
rect 17451 2468 17816 2496
rect 17451 2465 17463 2468
rect 17405 2459 17463 2465
rect 18417 2431 18475 2437
rect 18417 2397 18429 2431
rect 18463 2397 18475 2431
rect 18417 2391 18475 2397
rect 16347 2332 16712 2360
rect 16347 2329 16359 2332
rect 16301 2323 16359 2329
rect 7742 2292 7748 2304
rect 5031 2264 7144 2292
rect 7703 2264 7748 2292
rect 5031 2261 5043 2264
rect 4985 2255 5043 2261
rect 7742 2252 7748 2264
rect 7800 2252 7806 2304
rect 14550 2292 14556 2304
rect 14511 2264 14556 2292
rect 14550 2252 14556 2264
rect 14608 2252 14614 2304
rect 15194 2292 15200 2304
rect 15155 2264 15200 2292
rect 15194 2252 15200 2264
rect 15252 2252 15258 2304
rect 18046 2292 18052 2304
rect 18007 2264 18052 2292
rect 18046 2252 18052 2264
rect 18104 2292 18110 2304
rect 18432 2292 18460 2391
rect 18506 2388 18512 2440
rect 18564 2428 18570 2440
rect 18693 2431 18751 2437
rect 18693 2428 18705 2431
rect 18564 2400 18705 2428
rect 18564 2388 18570 2400
rect 18693 2397 18705 2400
rect 18739 2428 18751 2431
rect 18782 2428 18788 2440
rect 18739 2400 18788 2428
rect 18739 2397 18751 2400
rect 18693 2391 18751 2397
rect 18782 2388 18788 2400
rect 18840 2388 18846 2440
rect 18104 2264 18460 2292
rect 18104 2252 18110 2264
rect 1104 2202 20884 2224
rect 1104 2150 4648 2202
rect 4700 2150 4712 2202
rect 4764 2150 4776 2202
rect 4828 2150 4840 2202
rect 4892 2150 11982 2202
rect 12034 2150 12046 2202
rect 12098 2150 12110 2202
rect 12162 2150 12174 2202
rect 12226 2150 19315 2202
rect 19367 2150 19379 2202
rect 19431 2150 19443 2202
rect 19495 2150 19507 2202
rect 19559 2150 20884 2202
rect 1104 2128 20884 2150
rect 3142 2048 3148 2100
rect 3200 2088 3206 2100
rect 6638 2088 6644 2100
rect 3200 2060 6644 2088
rect 3200 2048 3206 2060
rect 6638 2048 6644 2060
rect 6696 2088 6702 2100
rect 7742 2088 7748 2100
rect 6696 2060 7748 2088
rect 6696 2048 6702 2060
rect 7742 2048 7748 2060
rect 7800 2048 7806 2100
rect 12434 2048 12440 2100
rect 12492 2088 12498 2100
rect 18506 2088 18512 2100
rect 12492 2060 18512 2088
rect 12492 2048 12498 2060
rect 18506 2048 18512 2060
rect 18564 2048 18570 2100
rect 934 76 940 128
rect 992 116 998 128
rect 3970 116 3976 128
rect 992 88 3976 116
rect 992 76 998 88
rect 3970 76 3976 88
rect 4028 76 4034 128
rect 7282 8 7288 60
rect 7340 48 7346 60
rect 12894 48 12900 60
rect 7340 20 12900 48
rect 7340 8 7346 20
rect 12894 8 12900 20
rect 12952 8 12958 60
<< via1 >>
rect 4648 19558 4700 19610
rect 4712 19558 4764 19610
rect 4776 19558 4828 19610
rect 4840 19558 4892 19610
rect 11982 19558 12034 19610
rect 12046 19558 12098 19610
rect 12110 19558 12162 19610
rect 12174 19558 12226 19610
rect 19315 19558 19367 19610
rect 19379 19558 19431 19610
rect 19443 19558 19495 19610
rect 19507 19558 19559 19610
rect 15752 19456 15804 19508
rect 13820 19252 13872 19304
rect 14004 19184 14056 19236
rect 15108 19252 15160 19304
rect 17868 19252 17920 19304
rect 17132 19184 17184 19236
rect 20628 19184 20680 19236
rect 14280 19116 14332 19168
rect 14832 19159 14884 19168
rect 14832 19125 14841 19159
rect 14841 19125 14875 19159
rect 14875 19125 14884 19159
rect 14832 19116 14884 19125
rect 17592 19116 17644 19168
rect 17868 19116 17920 19168
rect 18144 19116 18196 19168
rect 19800 19116 19852 19168
rect 8315 19014 8367 19066
rect 8379 19014 8431 19066
rect 8443 19014 8495 19066
rect 8507 19014 8559 19066
rect 15648 19014 15700 19066
rect 15712 19014 15764 19066
rect 15776 19014 15828 19066
rect 15840 19014 15892 19066
rect 14464 18912 14516 18964
rect 21640 18844 21692 18896
rect 11888 18776 11940 18828
rect 13452 18776 13504 18828
rect 14556 18776 14608 18828
rect 16028 18819 16080 18828
rect 16028 18785 16037 18819
rect 16037 18785 16071 18819
rect 16071 18785 16080 18819
rect 16028 18776 16080 18785
rect 16304 18819 16356 18828
rect 16304 18785 16313 18819
rect 16313 18785 16347 18819
rect 16347 18785 16356 18819
rect 16304 18776 16356 18785
rect 17500 18776 17552 18828
rect 18604 18819 18656 18828
rect 18604 18785 18613 18819
rect 18613 18785 18647 18819
rect 18647 18785 18656 18819
rect 18604 18776 18656 18785
rect 19984 18776 20036 18828
rect 16488 18751 16540 18760
rect 16488 18717 16497 18751
rect 16497 18717 16531 18751
rect 16531 18717 16540 18751
rect 16488 18708 16540 18717
rect 16948 18640 17000 18692
rect 12624 18615 12676 18624
rect 12624 18581 12633 18615
rect 12633 18581 12667 18615
rect 12667 18581 12676 18615
rect 12624 18572 12676 18581
rect 13636 18572 13688 18624
rect 15568 18615 15620 18624
rect 15568 18581 15577 18615
rect 15577 18581 15611 18615
rect 15611 18581 15620 18615
rect 15568 18572 15620 18581
rect 17960 18572 18012 18624
rect 21548 18572 21600 18624
rect 4648 18470 4700 18522
rect 4712 18470 4764 18522
rect 4776 18470 4828 18522
rect 4840 18470 4892 18522
rect 11982 18470 12034 18522
rect 12046 18470 12098 18522
rect 12110 18470 12162 18522
rect 12174 18470 12226 18522
rect 19315 18470 19367 18522
rect 19379 18470 19431 18522
rect 19443 18470 19495 18522
rect 19507 18470 19559 18522
rect 1584 18411 1636 18420
rect 1584 18377 1593 18411
rect 1593 18377 1627 18411
rect 1627 18377 1636 18411
rect 1584 18368 1636 18377
rect 2780 18368 2832 18420
rect 3332 18368 3384 18420
rect 8208 18368 8260 18420
rect 7380 18300 7432 18352
rect 13452 18368 13504 18420
rect 15936 18368 15988 18420
rect 18328 18368 18380 18420
rect 19984 18411 20036 18420
rect 19984 18377 19993 18411
rect 19993 18377 20027 18411
rect 20027 18377 20036 18411
rect 19984 18368 20036 18377
rect 10876 18300 10928 18352
rect 18604 18300 18656 18352
rect 9588 18096 9640 18148
rect 10600 18164 10652 18216
rect 12624 18164 12676 18216
rect 13176 18164 13228 18216
rect 14372 18207 14424 18216
rect 14372 18173 14381 18207
rect 14381 18173 14415 18207
rect 14415 18173 14424 18207
rect 14372 18164 14424 18173
rect 14832 18164 14884 18216
rect 15568 18164 15620 18216
rect 15936 18164 15988 18216
rect 13268 18139 13320 18148
rect 13268 18105 13277 18139
rect 13277 18105 13311 18139
rect 13311 18105 13320 18139
rect 13268 18096 13320 18105
rect 9312 18028 9364 18080
rect 10968 18071 11020 18080
rect 10968 18037 10977 18071
rect 10977 18037 11011 18071
rect 11011 18037 11020 18071
rect 10968 18028 11020 18037
rect 11888 18071 11940 18080
rect 11888 18037 11897 18071
rect 11897 18037 11931 18071
rect 11931 18037 11940 18071
rect 11888 18028 11940 18037
rect 12348 18028 12400 18080
rect 14556 18028 14608 18080
rect 15476 18028 15528 18080
rect 16120 18096 16172 18148
rect 16396 18096 16448 18148
rect 17500 18096 17552 18148
rect 16304 18028 16356 18080
rect 18420 18028 18472 18080
rect 19156 18028 19208 18080
rect 19616 18071 19668 18080
rect 19616 18037 19625 18071
rect 19625 18037 19659 18071
rect 19659 18037 19668 18071
rect 19616 18028 19668 18037
rect 8315 17926 8367 17978
rect 8379 17926 8431 17978
rect 8443 17926 8495 17978
rect 8507 17926 8559 17978
rect 15648 17926 15700 17978
rect 15712 17926 15764 17978
rect 15776 17926 15828 17978
rect 15840 17926 15892 17978
rect 15384 17867 15436 17876
rect 15384 17833 15393 17867
rect 15393 17833 15427 17867
rect 15427 17833 15436 17867
rect 15384 17824 15436 17833
rect 16304 17824 16356 17876
rect 18512 17867 18564 17876
rect 18512 17833 18521 17867
rect 18521 17833 18555 17867
rect 18555 17833 18564 17867
rect 18512 17824 18564 17833
rect 13544 17756 13596 17808
rect 14096 17756 14148 17808
rect 10692 17731 10744 17740
rect 10692 17697 10701 17731
rect 10701 17697 10735 17731
rect 10735 17697 10744 17731
rect 10692 17688 10744 17697
rect 12808 17731 12860 17740
rect 12808 17697 12817 17731
rect 12817 17697 12851 17731
rect 12851 17697 12860 17731
rect 12808 17688 12860 17697
rect 13176 17731 13228 17740
rect 13176 17697 13185 17731
rect 13185 17697 13219 17731
rect 13219 17697 13228 17731
rect 13176 17688 13228 17697
rect 14924 17688 14976 17740
rect 10600 17620 10652 17672
rect 10784 17663 10836 17672
rect 10784 17629 10793 17663
rect 10793 17629 10827 17663
rect 10827 17629 10836 17663
rect 10784 17620 10836 17629
rect 13360 17663 13412 17672
rect 13360 17629 13369 17663
rect 13369 17629 13403 17663
rect 13403 17629 13412 17663
rect 13360 17620 13412 17629
rect 15200 17620 15252 17672
rect 17224 17688 17276 17740
rect 17316 17731 17368 17740
rect 17316 17697 17325 17731
rect 17325 17697 17359 17731
rect 17359 17697 17368 17731
rect 18696 17731 18748 17740
rect 17316 17688 17368 17697
rect 18696 17697 18705 17731
rect 18705 17697 18739 17731
rect 18739 17697 18748 17731
rect 18696 17688 18748 17697
rect 18880 17731 18932 17740
rect 18880 17697 18889 17731
rect 18889 17697 18923 17731
rect 18923 17697 18932 17731
rect 18880 17688 18932 17697
rect 12808 17552 12860 17604
rect 16028 17552 16080 17604
rect 12716 17484 12768 17536
rect 13728 17484 13780 17536
rect 17776 17484 17828 17536
rect 4648 17382 4700 17434
rect 4712 17382 4764 17434
rect 4776 17382 4828 17434
rect 4840 17382 4892 17434
rect 11982 17382 12034 17434
rect 12046 17382 12098 17434
rect 12110 17382 12162 17434
rect 12174 17382 12226 17434
rect 19315 17382 19367 17434
rect 19379 17382 19431 17434
rect 19443 17382 19495 17434
rect 19507 17382 19559 17434
rect 15200 17280 15252 17332
rect 17224 17323 17276 17332
rect 12624 17212 12676 17264
rect 17224 17289 17233 17323
rect 17233 17289 17267 17323
rect 17267 17289 17276 17323
rect 17224 17280 17276 17289
rect 11060 17144 11112 17196
rect 12348 17144 12400 17196
rect 9496 17119 9548 17128
rect 9496 17085 9505 17119
rect 9505 17085 9539 17119
rect 9539 17085 9548 17119
rect 9496 17076 9548 17085
rect 12716 17119 12768 17128
rect 12716 17085 12725 17119
rect 12725 17085 12759 17119
rect 12759 17085 12768 17119
rect 12716 17076 12768 17085
rect 14464 17144 14516 17196
rect 13176 17076 13228 17128
rect 13544 17076 13596 17128
rect 17868 17144 17920 17196
rect 16212 17076 16264 17128
rect 10140 17051 10192 17060
rect 10140 17017 10149 17051
rect 10149 17017 10183 17051
rect 10183 17017 10192 17051
rect 10140 17008 10192 17017
rect 10600 17008 10652 17060
rect 14648 17008 14700 17060
rect 15108 17008 15160 17060
rect 16580 17051 16632 17060
rect 8668 16940 8720 16992
rect 9864 16940 9916 16992
rect 10692 16940 10744 16992
rect 11704 16940 11756 16992
rect 12348 16940 12400 16992
rect 12716 16983 12768 16992
rect 12716 16949 12725 16983
rect 12725 16949 12759 16983
rect 12759 16949 12768 16983
rect 12716 16940 12768 16949
rect 14096 16983 14148 16992
rect 14096 16949 14105 16983
rect 14105 16949 14139 16983
rect 14139 16949 14148 16983
rect 14096 16940 14148 16949
rect 15292 16983 15344 16992
rect 15292 16949 15301 16983
rect 15301 16949 15335 16983
rect 15335 16949 15344 16983
rect 15292 16940 15344 16949
rect 15476 16940 15528 16992
rect 16580 17017 16589 17051
rect 16589 17017 16623 17051
rect 16623 17017 16632 17051
rect 16580 17008 16632 17017
rect 17776 17076 17828 17128
rect 18880 17076 18932 17128
rect 17316 16940 17368 16992
rect 17868 16940 17920 16992
rect 8315 16838 8367 16890
rect 8379 16838 8431 16890
rect 8443 16838 8495 16890
rect 8507 16838 8559 16890
rect 15648 16838 15700 16890
rect 15712 16838 15764 16890
rect 15776 16838 15828 16890
rect 15840 16838 15892 16890
rect 10784 16779 10836 16788
rect 10784 16745 10793 16779
rect 10793 16745 10827 16779
rect 10827 16745 10836 16779
rect 10784 16736 10836 16745
rect 12532 16736 12584 16788
rect 13452 16736 13504 16788
rect 16212 16736 16264 16788
rect 17500 16736 17552 16788
rect 1492 16600 1544 16652
rect 2872 16600 2924 16652
rect 9036 16668 9088 16720
rect 11796 16711 11848 16720
rect 11796 16677 11805 16711
rect 11805 16677 11839 16711
rect 11839 16677 11848 16711
rect 11796 16668 11848 16677
rect 8484 16643 8536 16652
rect 8484 16609 8493 16643
rect 8493 16609 8527 16643
rect 8527 16609 8536 16643
rect 8484 16600 8536 16609
rect 9680 16643 9732 16652
rect 9680 16609 9689 16643
rect 9689 16609 9723 16643
rect 9723 16609 9732 16643
rect 9680 16600 9732 16609
rect 9864 16600 9916 16652
rect 12624 16600 12676 16652
rect 17776 16668 17828 16720
rect 17960 16711 18012 16720
rect 17960 16677 17969 16711
rect 17969 16677 18003 16711
rect 18003 16677 18012 16711
rect 17960 16668 18012 16677
rect 18696 16736 18748 16788
rect 21548 16736 21600 16788
rect 13544 16600 13596 16652
rect 15568 16643 15620 16652
rect 8760 16575 8812 16584
rect 8760 16541 8769 16575
rect 8769 16541 8803 16575
rect 8803 16541 8812 16575
rect 8760 16532 8812 16541
rect 10508 16532 10560 16584
rect 11704 16575 11756 16584
rect 11704 16541 11713 16575
rect 11713 16541 11747 16575
rect 11747 16541 11756 16575
rect 11704 16532 11756 16541
rect 11888 16532 11940 16584
rect 15568 16609 15577 16643
rect 15577 16609 15611 16643
rect 15611 16609 15620 16643
rect 15568 16600 15620 16609
rect 15752 16643 15804 16652
rect 15752 16609 15761 16643
rect 15761 16609 15795 16643
rect 15795 16609 15804 16643
rect 15752 16600 15804 16609
rect 19616 16600 19668 16652
rect 17776 16532 17828 16584
rect 18604 16575 18656 16584
rect 18604 16541 18613 16575
rect 18613 16541 18647 16575
rect 18647 16541 18656 16575
rect 18604 16532 18656 16541
rect 15568 16464 15620 16516
rect 18696 16464 18748 16516
rect 8116 16396 8168 16448
rect 9496 16439 9548 16448
rect 9496 16405 9505 16439
rect 9505 16405 9539 16439
rect 9539 16405 9548 16439
rect 9496 16396 9548 16405
rect 12808 16396 12860 16448
rect 14464 16396 14516 16448
rect 14648 16439 14700 16448
rect 14648 16405 14657 16439
rect 14657 16405 14691 16439
rect 14691 16405 14700 16439
rect 14648 16396 14700 16405
rect 14924 16396 14976 16448
rect 4648 16294 4700 16346
rect 4712 16294 4764 16346
rect 4776 16294 4828 16346
rect 4840 16294 4892 16346
rect 11982 16294 12034 16346
rect 12046 16294 12098 16346
rect 12110 16294 12162 16346
rect 12174 16294 12226 16346
rect 19315 16294 19367 16346
rect 19379 16294 19431 16346
rect 19443 16294 19495 16346
rect 19507 16294 19559 16346
rect 1584 16235 1636 16244
rect 1584 16201 1593 16235
rect 1593 16201 1627 16235
rect 1627 16201 1636 16235
rect 1584 16192 1636 16201
rect 11704 16192 11756 16244
rect 14648 16192 14700 16244
rect 14832 16235 14884 16244
rect 14832 16201 14841 16235
rect 14841 16201 14875 16235
rect 14875 16201 14884 16235
rect 14832 16192 14884 16201
rect 15568 16192 15620 16244
rect 17500 16235 17552 16244
rect 17500 16201 17509 16235
rect 17509 16201 17543 16235
rect 17543 16201 17552 16235
rect 17500 16192 17552 16201
rect 17776 16235 17828 16244
rect 17776 16201 17785 16235
rect 17785 16201 17819 16235
rect 17819 16201 17828 16235
rect 17776 16192 17828 16201
rect 9680 16124 9732 16176
rect 1308 16056 1360 16108
rect 10784 16056 10836 16108
rect 11796 16124 11848 16176
rect 12624 16099 12676 16108
rect 12624 16065 12633 16099
rect 12633 16065 12667 16099
rect 12667 16065 12676 16099
rect 12624 16056 12676 16065
rect 13268 16056 13320 16108
rect 14464 16056 14516 16108
rect 15752 16056 15804 16108
rect 17316 16056 17368 16108
rect 19064 16124 19116 16176
rect 19984 16124 20036 16176
rect 18328 16056 18380 16108
rect 7380 16031 7432 16040
rect 7380 15997 7389 16031
rect 7389 15997 7423 16031
rect 7423 15997 7432 16031
rect 7380 15988 7432 15997
rect 9588 16031 9640 16040
rect 9588 15997 9632 16031
rect 9632 15997 9640 16031
rect 9588 15988 9640 15997
rect 13912 15988 13964 16040
rect 16212 16031 16264 16040
rect 16212 15997 16221 16031
rect 16221 15997 16255 16031
rect 16255 15997 16264 16031
rect 16212 15988 16264 15997
rect 7472 15920 7524 15972
rect 8024 15963 8076 15972
rect 8024 15929 8033 15963
rect 8033 15929 8067 15963
rect 8067 15929 8076 15963
rect 8024 15920 8076 15929
rect 8116 15963 8168 15972
rect 8116 15929 8125 15963
rect 8125 15929 8159 15963
rect 8159 15929 8168 15963
rect 8116 15920 8168 15929
rect 8484 15920 8536 15972
rect 8668 15963 8720 15972
rect 8668 15929 8677 15963
rect 8677 15929 8711 15963
rect 8711 15929 8720 15963
rect 8668 15920 8720 15929
rect 2964 15852 3016 15904
rect 7748 15895 7800 15904
rect 7748 15861 7757 15895
rect 7757 15861 7791 15895
rect 7791 15861 7800 15895
rect 9864 15920 9916 15972
rect 10232 15920 10284 15972
rect 9036 15895 9088 15904
rect 7748 15852 7800 15861
rect 9036 15861 9045 15895
rect 9045 15861 9079 15895
rect 9079 15861 9088 15895
rect 9036 15852 9088 15861
rect 9956 15852 10008 15904
rect 17960 15988 18012 16040
rect 18880 15988 18932 16040
rect 16672 15963 16724 15972
rect 13820 15852 13872 15904
rect 15016 15852 15068 15904
rect 15292 15852 15344 15904
rect 16672 15929 16681 15963
rect 16681 15929 16715 15963
rect 16715 15929 16724 15963
rect 16672 15920 16724 15929
rect 18236 15963 18288 15972
rect 18236 15929 18245 15963
rect 18245 15929 18279 15963
rect 18279 15929 18288 15963
rect 18236 15920 18288 15929
rect 17408 15852 17460 15904
rect 19616 15852 19668 15904
rect 8315 15750 8367 15802
rect 8379 15750 8431 15802
rect 8443 15750 8495 15802
rect 8507 15750 8559 15802
rect 15648 15750 15700 15802
rect 15712 15750 15764 15802
rect 15776 15750 15828 15802
rect 15840 15750 15892 15802
rect 8024 15648 8076 15700
rect 8116 15648 8168 15700
rect 7932 15580 7984 15632
rect 13820 15691 13872 15700
rect 13820 15657 13829 15691
rect 13829 15657 13863 15691
rect 13863 15657 13872 15691
rect 13820 15648 13872 15657
rect 16212 15648 16264 15700
rect 18236 15648 18288 15700
rect 18788 15648 18840 15700
rect 10232 15580 10284 15632
rect 11704 15623 11756 15632
rect 11704 15589 11713 15623
rect 11713 15589 11747 15623
rect 11747 15589 11756 15623
rect 11704 15580 11756 15589
rect 8760 15512 8812 15564
rect 9864 15512 9916 15564
rect 13360 15512 13412 15564
rect 14740 15512 14792 15564
rect 16580 15512 16632 15564
rect 18512 15555 18564 15564
rect 18512 15521 18521 15555
rect 18521 15521 18555 15555
rect 18555 15521 18564 15555
rect 18512 15512 18564 15521
rect 7564 15444 7616 15496
rect 11612 15487 11664 15496
rect 11612 15453 11621 15487
rect 11621 15453 11655 15487
rect 11655 15453 11664 15487
rect 11612 15444 11664 15453
rect 11888 15487 11940 15496
rect 11888 15453 11897 15487
rect 11897 15453 11931 15487
rect 11931 15453 11940 15487
rect 11888 15444 11940 15453
rect 5356 15376 5408 15428
rect 9680 15376 9732 15428
rect 6920 15351 6972 15360
rect 6920 15317 6929 15351
rect 6929 15317 6963 15351
rect 6963 15317 6972 15351
rect 6920 15308 6972 15317
rect 8944 15351 8996 15360
rect 8944 15317 8953 15351
rect 8953 15317 8987 15351
rect 8987 15317 8996 15351
rect 8944 15308 8996 15317
rect 11336 15308 11388 15360
rect 12348 15308 12400 15360
rect 14372 15351 14424 15360
rect 14372 15317 14381 15351
rect 14381 15317 14415 15351
rect 14415 15317 14424 15351
rect 14372 15308 14424 15317
rect 14556 15308 14608 15360
rect 18696 15308 18748 15360
rect 4648 15206 4700 15258
rect 4712 15206 4764 15258
rect 4776 15206 4828 15258
rect 4840 15206 4892 15258
rect 11982 15206 12034 15258
rect 12046 15206 12098 15258
rect 12110 15206 12162 15258
rect 12174 15206 12226 15258
rect 19315 15206 19367 15258
rect 19379 15206 19431 15258
rect 19443 15206 19495 15258
rect 19507 15206 19559 15258
rect 6276 15147 6328 15156
rect 6276 15113 6285 15147
rect 6285 15113 6319 15147
rect 6319 15113 6328 15147
rect 6276 15104 6328 15113
rect 7932 15147 7984 15156
rect 7932 15113 7941 15147
rect 7941 15113 7975 15147
rect 7975 15113 7984 15147
rect 7932 15104 7984 15113
rect 10232 15104 10284 15156
rect 11704 15147 11756 15156
rect 11704 15113 11713 15147
rect 11713 15113 11747 15147
rect 11747 15113 11756 15147
rect 11704 15104 11756 15113
rect 13820 15104 13872 15156
rect 16580 15104 16632 15156
rect 17040 15147 17092 15156
rect 17040 15113 17049 15147
rect 17049 15113 17083 15147
rect 17083 15113 17092 15147
rect 17040 15104 17092 15113
rect 18512 15104 18564 15156
rect 7564 15011 7616 15020
rect 7564 14977 7573 15011
rect 7573 14977 7607 15011
rect 7607 14977 7616 15011
rect 7564 14968 7616 14977
rect 9312 14968 9364 15020
rect 10140 14968 10192 15020
rect 13452 15011 13504 15020
rect 13452 14977 13461 15011
rect 13461 14977 13495 15011
rect 13495 14977 13504 15011
rect 13452 14968 13504 14977
rect 2228 14900 2280 14952
rect 6276 14900 6328 14952
rect 6828 14900 6880 14952
rect 6920 14900 6972 14952
rect 12900 14943 12952 14952
rect 9220 14875 9272 14884
rect 6092 14764 6144 14816
rect 9220 14841 9229 14875
rect 9229 14841 9263 14875
rect 9263 14841 9272 14875
rect 9220 14832 9272 14841
rect 8944 14764 8996 14816
rect 10232 14832 10284 14884
rect 11152 14832 11204 14884
rect 11612 14832 11664 14884
rect 12900 14909 12909 14943
rect 12909 14909 12943 14943
rect 12943 14909 12952 14943
rect 12900 14900 12952 14909
rect 17224 15036 17276 15088
rect 18788 15036 18840 15088
rect 19064 15079 19116 15088
rect 19064 15045 19073 15079
rect 19073 15045 19107 15079
rect 19107 15045 19116 15079
rect 19064 15036 19116 15045
rect 19248 15036 19300 15088
rect 15108 14968 15160 15020
rect 15936 14968 15988 15020
rect 17040 14968 17092 15020
rect 18972 14968 19024 15020
rect 16856 14943 16908 14952
rect 10692 14764 10744 14816
rect 10968 14807 11020 14816
rect 10968 14773 10977 14807
rect 10977 14773 11011 14807
rect 11011 14773 11020 14807
rect 10968 14764 11020 14773
rect 12808 14764 12860 14816
rect 14740 14764 14792 14816
rect 16856 14909 16865 14943
rect 16865 14909 16899 14943
rect 16899 14909 16908 14943
rect 16856 14900 16908 14909
rect 15292 14875 15344 14884
rect 15292 14841 15301 14875
rect 15301 14841 15335 14875
rect 15335 14841 15344 14875
rect 15292 14832 15344 14841
rect 15476 14764 15528 14816
rect 18696 14832 18748 14884
rect 8315 14662 8367 14714
rect 8379 14662 8431 14714
rect 8443 14662 8495 14714
rect 8507 14662 8559 14714
rect 15648 14662 15700 14714
rect 15712 14662 15764 14714
rect 15776 14662 15828 14714
rect 15840 14662 15892 14714
rect 6368 14560 6420 14612
rect 2872 14424 2924 14476
rect 4988 14424 5040 14476
rect 5448 14424 5500 14476
rect 6920 14492 6972 14544
rect 7932 14492 7984 14544
rect 5908 14467 5960 14476
rect 5908 14433 5917 14467
rect 5917 14433 5951 14467
rect 5951 14433 5960 14467
rect 5908 14424 5960 14433
rect 9036 14424 9088 14476
rect 9312 14560 9364 14612
rect 9864 14603 9916 14612
rect 9864 14569 9873 14603
rect 9873 14569 9907 14603
rect 9907 14569 9916 14603
rect 9864 14560 9916 14569
rect 10232 14560 10284 14612
rect 12532 14603 12584 14612
rect 12532 14569 12541 14603
rect 12541 14569 12575 14603
rect 12575 14569 12584 14603
rect 12532 14560 12584 14569
rect 13360 14560 13412 14612
rect 10968 14492 11020 14544
rect 11520 14492 11572 14544
rect 11888 14492 11940 14544
rect 13544 14535 13596 14544
rect 13544 14501 13553 14535
rect 13553 14501 13587 14535
rect 13587 14501 13596 14535
rect 13544 14492 13596 14501
rect 14832 14560 14884 14612
rect 15292 14560 15344 14612
rect 15476 14603 15528 14612
rect 15476 14569 15485 14603
rect 15485 14569 15519 14603
rect 15519 14569 15528 14603
rect 15476 14560 15528 14569
rect 15936 14560 15988 14612
rect 17224 14492 17276 14544
rect 18604 14535 18656 14544
rect 18604 14501 18613 14535
rect 18613 14501 18647 14535
rect 18647 14501 18656 14535
rect 18604 14492 18656 14501
rect 19064 14492 19116 14544
rect 19248 14535 19300 14544
rect 19248 14501 19257 14535
rect 19257 14501 19291 14535
rect 19291 14501 19300 14535
rect 19248 14492 19300 14501
rect 10324 14424 10376 14476
rect 15660 14467 15712 14476
rect 8024 14356 8076 14408
rect 9220 14356 9272 14408
rect 11796 14356 11848 14408
rect 13728 14356 13780 14408
rect 6736 14288 6788 14340
rect 6828 14288 6880 14340
rect 9864 14288 9916 14340
rect 10600 14288 10652 14340
rect 12992 14288 13044 14340
rect 15660 14433 15669 14467
rect 15669 14433 15703 14467
rect 15703 14433 15712 14467
rect 15660 14424 15712 14433
rect 16396 14424 16448 14476
rect 16488 14424 16540 14476
rect 16764 14467 16816 14476
rect 16764 14433 16773 14467
rect 16773 14433 16807 14467
rect 16807 14433 16816 14467
rect 16764 14424 16816 14433
rect 16212 14356 16264 14408
rect 17868 14356 17920 14408
rect 4252 14220 4304 14272
rect 5632 14220 5684 14272
rect 7840 14263 7892 14272
rect 7840 14229 7849 14263
rect 7849 14229 7883 14263
rect 7883 14229 7892 14263
rect 7840 14220 7892 14229
rect 8760 14263 8812 14272
rect 8760 14229 8769 14263
rect 8769 14229 8803 14263
rect 8803 14229 8812 14263
rect 8760 14220 8812 14229
rect 10416 14220 10468 14272
rect 13452 14220 13504 14272
rect 14188 14220 14240 14272
rect 4648 14118 4700 14170
rect 4712 14118 4764 14170
rect 4776 14118 4828 14170
rect 4840 14118 4892 14170
rect 11982 14118 12034 14170
rect 12046 14118 12098 14170
rect 12110 14118 12162 14170
rect 12174 14118 12226 14170
rect 19315 14118 19367 14170
rect 19379 14118 19431 14170
rect 19443 14118 19495 14170
rect 19507 14118 19559 14170
rect 4988 14016 5040 14068
rect 5172 14016 5224 14068
rect 8024 14059 8076 14068
rect 8024 14025 8033 14059
rect 8033 14025 8067 14059
rect 8067 14025 8076 14059
rect 8024 14016 8076 14025
rect 13452 14016 13504 14068
rect 13728 14016 13780 14068
rect 14372 14016 14424 14068
rect 15016 14016 15068 14068
rect 15660 14059 15712 14068
rect 7196 13948 7248 14000
rect 7748 13948 7800 14000
rect 10232 13948 10284 14000
rect 4160 13812 4212 13864
rect 8760 13923 8812 13932
rect 8760 13889 8769 13923
rect 8769 13889 8803 13923
rect 8803 13889 8812 13923
rect 8760 13880 8812 13889
rect 5080 13812 5132 13864
rect 5448 13855 5500 13864
rect 5448 13821 5457 13855
rect 5457 13821 5491 13855
rect 5491 13821 5500 13855
rect 5448 13812 5500 13821
rect 5632 13855 5684 13864
rect 5632 13821 5641 13855
rect 5641 13821 5675 13855
rect 5675 13821 5684 13855
rect 5632 13812 5684 13821
rect 5540 13744 5592 13796
rect 6920 13812 6972 13864
rect 9588 13880 9640 13932
rect 10140 13880 10192 13932
rect 10508 13923 10560 13932
rect 10508 13889 10517 13923
rect 10517 13889 10551 13923
rect 10551 13889 10560 13923
rect 10508 13880 10560 13889
rect 12532 13880 12584 13932
rect 15108 13880 15160 13932
rect 9680 13855 9732 13864
rect 9680 13821 9689 13855
rect 9689 13821 9723 13855
rect 9723 13821 9732 13855
rect 9680 13812 9732 13821
rect 10324 13812 10376 13864
rect 15660 14025 15669 14059
rect 15669 14025 15703 14059
rect 15703 14025 15712 14059
rect 15660 14016 15712 14025
rect 17500 14016 17552 14068
rect 19064 14059 19116 14068
rect 17224 13948 17276 14000
rect 16212 13923 16264 13932
rect 16212 13889 16221 13923
rect 16221 13889 16255 13923
rect 16255 13889 16264 13923
rect 16212 13880 16264 13889
rect 6000 13676 6052 13728
rect 7196 13719 7248 13728
rect 7196 13685 7205 13719
rect 7205 13685 7239 13719
rect 7239 13685 7248 13719
rect 7196 13676 7248 13685
rect 7656 13676 7708 13728
rect 11428 13719 11480 13728
rect 11428 13685 11437 13719
rect 11437 13685 11471 13719
rect 11471 13685 11480 13719
rect 11428 13676 11480 13685
rect 12624 13676 12676 13728
rect 13360 13719 13412 13728
rect 13360 13685 13369 13719
rect 13369 13685 13403 13719
rect 13403 13685 13412 13719
rect 13360 13676 13412 13685
rect 13544 13676 13596 13728
rect 14188 13744 14240 13796
rect 14372 13787 14424 13796
rect 14372 13753 14381 13787
rect 14381 13753 14415 13787
rect 14415 13753 14424 13787
rect 14372 13744 14424 13753
rect 14464 13787 14516 13796
rect 14464 13753 14473 13787
rect 14473 13753 14507 13787
rect 14507 13753 14516 13787
rect 14464 13744 14516 13753
rect 15016 13744 15068 13796
rect 16580 13787 16632 13796
rect 16580 13753 16583 13787
rect 16583 13753 16617 13787
rect 16617 13753 16632 13787
rect 19064 14025 19073 14059
rect 19073 14025 19107 14059
rect 19107 14025 19116 14059
rect 19064 14016 19116 14025
rect 19892 14059 19944 14068
rect 19892 14025 19901 14059
rect 19901 14025 19935 14059
rect 19935 14025 19944 14059
rect 19892 14016 19944 14025
rect 19616 13948 19668 14000
rect 18144 13923 18196 13932
rect 18144 13889 18153 13923
rect 18153 13889 18187 13923
rect 18187 13889 18196 13923
rect 18144 13880 18196 13889
rect 19651 13855 19703 13864
rect 19651 13821 19660 13855
rect 19660 13821 19694 13855
rect 19694 13821 19703 13855
rect 19651 13812 19703 13821
rect 16580 13744 16632 13753
rect 15476 13676 15528 13728
rect 18880 13676 18932 13728
rect 19432 13719 19484 13728
rect 19432 13685 19441 13719
rect 19441 13685 19475 13719
rect 19475 13685 19484 13719
rect 19432 13676 19484 13685
rect 8315 13574 8367 13626
rect 8379 13574 8431 13626
rect 8443 13574 8495 13626
rect 8507 13574 8559 13626
rect 15648 13574 15700 13626
rect 15712 13574 15764 13626
rect 15776 13574 15828 13626
rect 15840 13574 15892 13626
rect 5540 13472 5592 13524
rect 5724 13472 5776 13524
rect 11336 13472 11388 13524
rect 11520 13515 11572 13524
rect 11520 13481 11529 13515
rect 11529 13481 11563 13515
rect 11563 13481 11572 13515
rect 11520 13472 11572 13481
rect 13452 13515 13504 13524
rect 13452 13481 13461 13515
rect 13461 13481 13495 13515
rect 13495 13481 13504 13515
rect 13452 13472 13504 13481
rect 16304 13472 16356 13524
rect 16764 13472 16816 13524
rect 18144 13515 18196 13524
rect 18144 13481 18153 13515
rect 18153 13481 18187 13515
rect 18187 13481 18196 13515
rect 18144 13472 18196 13481
rect 3976 13404 4028 13456
rect 6552 13447 6604 13456
rect 6552 13413 6561 13447
rect 6561 13413 6595 13447
rect 6595 13413 6604 13447
rect 6552 13404 6604 13413
rect 6828 13404 6880 13456
rect 7840 13404 7892 13456
rect 10692 13447 10744 13456
rect 10692 13413 10701 13447
rect 10701 13413 10735 13447
rect 10735 13413 10744 13447
rect 10692 13404 10744 13413
rect 11428 13404 11480 13456
rect 11888 13404 11940 13456
rect 13360 13404 13412 13456
rect 13820 13447 13872 13456
rect 13820 13413 13829 13447
rect 13829 13413 13863 13447
rect 13863 13413 13872 13447
rect 13820 13404 13872 13413
rect 16396 13404 16448 13456
rect 16580 13404 16632 13456
rect 18420 13447 18472 13456
rect 18420 13413 18429 13447
rect 18429 13413 18463 13447
rect 18463 13413 18472 13447
rect 18420 13404 18472 13413
rect 5080 13379 5132 13388
rect 5080 13345 5089 13379
rect 5089 13345 5123 13379
rect 5123 13345 5132 13379
rect 5356 13379 5408 13388
rect 5080 13336 5132 13345
rect 2688 13268 2740 13320
rect 2872 13268 2924 13320
rect 5356 13345 5365 13379
rect 5365 13345 5399 13379
rect 5399 13345 5408 13379
rect 5356 13336 5408 13345
rect 6276 13336 6328 13388
rect 15476 13336 15528 13388
rect 17408 13336 17460 13388
rect 6000 13268 6052 13320
rect 7564 13268 7616 13320
rect 8668 13311 8720 13320
rect 8668 13277 8677 13311
rect 8677 13277 8711 13311
rect 8711 13277 8720 13311
rect 8668 13268 8720 13277
rect 9956 13268 10008 13320
rect 10692 13268 10744 13320
rect 10416 13200 10468 13252
rect 12348 13268 12400 13320
rect 12808 13268 12860 13320
rect 13452 13268 13504 13320
rect 14372 13311 14424 13320
rect 14372 13277 14381 13311
rect 14381 13277 14415 13311
rect 14415 13277 14424 13311
rect 14372 13268 14424 13277
rect 16028 13268 16080 13320
rect 16120 13268 16172 13320
rect 16672 13268 16724 13320
rect 18328 13311 18380 13320
rect 18328 13277 18337 13311
rect 18337 13277 18371 13311
rect 18371 13277 18380 13311
rect 18328 13268 18380 13277
rect 18604 13311 18656 13320
rect 18604 13277 18613 13311
rect 18613 13277 18647 13311
rect 18647 13277 18656 13311
rect 18604 13268 18656 13277
rect 19432 13268 19484 13320
rect 11152 13243 11204 13252
rect 11152 13209 11161 13243
rect 11161 13209 11195 13243
rect 11195 13209 11204 13243
rect 11152 13200 11204 13209
rect 16212 13200 16264 13252
rect 2872 13175 2924 13184
rect 2872 13141 2881 13175
rect 2881 13141 2915 13175
rect 2915 13141 2924 13175
rect 2872 13132 2924 13141
rect 4988 13132 5040 13184
rect 5540 13132 5592 13184
rect 5908 13132 5960 13184
rect 6276 13175 6328 13184
rect 6276 13141 6285 13175
rect 6285 13141 6319 13175
rect 6319 13141 6328 13175
rect 6276 13132 6328 13141
rect 7748 13175 7800 13184
rect 7748 13141 7757 13175
rect 7757 13141 7791 13175
rect 7791 13141 7800 13175
rect 7748 13132 7800 13141
rect 10324 13175 10376 13184
rect 10324 13141 10333 13175
rect 10333 13141 10367 13175
rect 10367 13141 10376 13175
rect 10324 13132 10376 13141
rect 11520 13132 11572 13184
rect 11796 13132 11848 13184
rect 16488 13132 16540 13184
rect 16580 13132 16632 13184
rect 4648 13030 4700 13082
rect 4712 13030 4764 13082
rect 4776 13030 4828 13082
rect 4840 13030 4892 13082
rect 11982 13030 12034 13082
rect 12046 13030 12098 13082
rect 12110 13030 12162 13082
rect 12174 13030 12226 13082
rect 19315 13030 19367 13082
rect 19379 13030 19431 13082
rect 19443 13030 19495 13082
rect 19507 13030 19559 13082
rect 2780 12928 2832 12980
rect 2872 12928 2924 12980
rect 3976 12971 4028 12980
rect 3976 12937 3985 12971
rect 3985 12937 4019 12971
rect 4019 12937 4028 12971
rect 3976 12928 4028 12937
rect 9772 12928 9824 12980
rect 11428 12971 11480 12980
rect 11428 12937 11437 12971
rect 11437 12937 11471 12971
rect 11471 12937 11480 12971
rect 11428 12928 11480 12937
rect 13820 12928 13872 12980
rect 15476 12971 15528 12980
rect 4620 12860 4672 12912
rect 10324 12860 10376 12912
rect 11888 12903 11940 12912
rect 6092 12792 6144 12844
rect 7380 12792 7432 12844
rect 7564 12792 7616 12844
rect 2964 12724 3016 12776
rect 3056 12588 3108 12640
rect 3516 12588 3568 12640
rect 5540 12724 5592 12776
rect 5632 12656 5684 12708
rect 6184 12724 6236 12776
rect 8668 12792 8720 12844
rect 11888 12869 11897 12903
rect 11897 12869 11931 12903
rect 11931 12869 11940 12903
rect 11888 12860 11940 12869
rect 12716 12835 12768 12844
rect 12716 12801 12725 12835
rect 12725 12801 12759 12835
rect 12759 12801 12768 12835
rect 12716 12792 12768 12801
rect 4988 12588 5040 12640
rect 7748 12699 7800 12708
rect 6368 12588 6420 12640
rect 6552 12588 6604 12640
rect 7748 12665 7757 12699
rect 7757 12665 7791 12699
rect 7791 12665 7800 12699
rect 7748 12656 7800 12665
rect 8208 12656 8260 12708
rect 8852 12699 8904 12708
rect 8852 12665 8861 12699
rect 8861 12665 8895 12699
rect 8895 12665 8904 12699
rect 8852 12656 8904 12665
rect 7656 12588 7708 12640
rect 9680 12656 9732 12708
rect 10508 12699 10560 12708
rect 10508 12665 10517 12699
rect 10517 12665 10551 12699
rect 10551 12665 10560 12699
rect 10508 12656 10560 12665
rect 11152 12656 11204 12708
rect 11888 12656 11940 12708
rect 12716 12656 12768 12708
rect 15476 12937 15485 12971
rect 15485 12937 15519 12971
rect 15519 12937 15528 12971
rect 15476 12928 15528 12937
rect 14464 12860 14516 12912
rect 18052 12928 18104 12980
rect 18696 12928 18748 12980
rect 14556 12835 14608 12844
rect 14556 12801 14565 12835
rect 14565 12801 14599 12835
rect 14599 12801 14608 12835
rect 14556 12792 14608 12801
rect 14832 12835 14884 12844
rect 14832 12801 14841 12835
rect 14841 12801 14875 12835
rect 14875 12801 14884 12835
rect 14832 12792 14884 12801
rect 16304 12792 16356 12844
rect 18788 12860 18840 12912
rect 19156 12860 19208 12912
rect 18880 12835 18932 12844
rect 18880 12801 18889 12835
rect 18889 12801 18923 12835
rect 18923 12801 18932 12835
rect 18880 12792 18932 12801
rect 16396 12656 16448 12708
rect 15936 12631 15988 12640
rect 15936 12597 15945 12631
rect 15945 12597 15979 12631
rect 15979 12597 15988 12631
rect 15936 12588 15988 12597
rect 18420 12724 18472 12776
rect 8315 12486 8367 12538
rect 8379 12486 8431 12538
rect 8443 12486 8495 12538
rect 8507 12486 8559 12538
rect 15648 12486 15700 12538
rect 15712 12486 15764 12538
rect 15776 12486 15828 12538
rect 15840 12486 15892 12538
rect 4620 12384 4672 12436
rect 6000 12427 6052 12436
rect 6000 12393 6009 12427
rect 6009 12393 6043 12427
rect 6043 12393 6052 12427
rect 6000 12384 6052 12393
rect 7380 12427 7432 12436
rect 7380 12393 7389 12427
rect 7389 12393 7423 12427
rect 7423 12393 7432 12427
rect 7380 12384 7432 12393
rect 7840 12427 7892 12436
rect 7840 12393 7849 12427
rect 7849 12393 7883 12427
rect 7883 12393 7892 12427
rect 7840 12384 7892 12393
rect 8852 12384 8904 12436
rect 10692 12427 10744 12436
rect 2044 12248 2096 12300
rect 2780 12248 2832 12300
rect 5540 12316 5592 12368
rect 6460 12359 6512 12368
rect 6460 12325 6469 12359
rect 6469 12325 6503 12359
rect 6503 12325 6512 12359
rect 6460 12316 6512 12325
rect 3884 12180 3936 12232
rect 5264 12248 5316 12300
rect 9036 12316 9088 12368
rect 10692 12393 10701 12427
rect 10701 12393 10735 12427
rect 10735 12393 10744 12427
rect 10692 12384 10744 12393
rect 12348 12427 12400 12436
rect 12348 12393 12357 12427
rect 12357 12393 12391 12427
rect 12391 12393 12400 12427
rect 12348 12384 12400 12393
rect 13452 12427 13504 12436
rect 13452 12393 13461 12427
rect 13461 12393 13495 12427
rect 13495 12393 13504 12427
rect 13452 12384 13504 12393
rect 14556 12384 14608 12436
rect 16672 12427 16724 12436
rect 16672 12393 16681 12427
rect 16681 12393 16715 12427
rect 16715 12393 16724 12427
rect 16672 12384 16724 12393
rect 17408 12384 17460 12436
rect 18328 12427 18380 12436
rect 18328 12393 18337 12427
rect 18337 12393 18371 12427
rect 18371 12393 18380 12427
rect 18328 12384 18380 12393
rect 18788 12427 18840 12436
rect 18788 12393 18797 12427
rect 18797 12393 18831 12427
rect 18831 12393 18840 12427
rect 18788 12384 18840 12393
rect 11612 12316 11664 12368
rect 13820 12359 13872 12368
rect 13820 12325 13829 12359
rect 13829 12325 13863 12359
rect 13863 12325 13872 12359
rect 13820 12316 13872 12325
rect 14832 12316 14884 12368
rect 15476 12359 15528 12368
rect 15476 12325 15485 12359
rect 15485 12325 15519 12359
rect 15519 12325 15528 12359
rect 15476 12316 15528 12325
rect 16028 12359 16080 12368
rect 16028 12325 16037 12359
rect 16037 12325 16071 12359
rect 16071 12325 16080 12359
rect 16028 12316 16080 12325
rect 19064 12359 19116 12368
rect 19064 12325 19073 12359
rect 19073 12325 19107 12359
rect 19107 12325 19116 12359
rect 19064 12316 19116 12325
rect 16764 12248 16816 12300
rect 17776 12248 17828 12300
rect 5356 12223 5408 12232
rect 5356 12189 5365 12223
rect 5365 12189 5399 12223
rect 5399 12189 5408 12223
rect 5356 12180 5408 12189
rect 6184 12223 6236 12232
rect 6184 12189 6193 12223
rect 6193 12189 6227 12223
rect 6227 12189 6236 12223
rect 6184 12180 6236 12189
rect 1860 12112 1912 12164
rect 8208 12180 8260 12232
rect 9772 12223 9824 12232
rect 9772 12189 9781 12223
rect 9781 12189 9815 12223
rect 9815 12189 9824 12223
rect 9772 12180 9824 12189
rect 8668 12112 8720 12164
rect 11244 12112 11296 12164
rect 11520 12180 11572 12232
rect 14188 12180 14240 12232
rect 3148 12044 3200 12096
rect 5540 12044 5592 12096
rect 7196 12044 7248 12096
rect 7472 12044 7524 12096
rect 9128 12044 9180 12096
rect 9864 12044 9916 12096
rect 11060 12044 11112 12096
rect 12716 12087 12768 12096
rect 12716 12053 12725 12087
rect 12725 12053 12759 12087
rect 12759 12053 12768 12087
rect 12716 12044 12768 12053
rect 12808 12044 12860 12096
rect 16488 12180 16540 12232
rect 18972 12223 19024 12232
rect 18972 12189 18981 12223
rect 18981 12189 19015 12223
rect 19015 12189 19024 12223
rect 18972 12180 19024 12189
rect 19156 12180 19208 12232
rect 18788 12112 18840 12164
rect 16028 12044 16080 12096
rect 4648 11942 4700 11994
rect 4712 11942 4764 11994
rect 4776 11942 4828 11994
rect 4840 11942 4892 11994
rect 11982 11942 12034 11994
rect 12046 11942 12098 11994
rect 12110 11942 12162 11994
rect 12174 11942 12226 11994
rect 19315 11942 19367 11994
rect 19379 11942 19431 11994
rect 19443 11942 19495 11994
rect 19507 11942 19559 11994
rect 2780 11840 2832 11892
rect 5540 11840 5592 11892
rect 8024 11840 8076 11892
rect 9036 11883 9088 11892
rect 9036 11849 9045 11883
rect 9045 11849 9079 11883
rect 9079 11849 9088 11883
rect 9036 11840 9088 11849
rect 9772 11840 9824 11892
rect 13820 11883 13872 11892
rect 13820 11849 13829 11883
rect 13829 11849 13863 11883
rect 13863 11849 13872 11883
rect 13820 11840 13872 11849
rect 15476 11840 15528 11892
rect 17776 11883 17828 11892
rect 17776 11849 17785 11883
rect 17785 11849 17819 11883
rect 17819 11849 17828 11883
rect 17776 11840 17828 11849
rect 19064 11840 19116 11892
rect 11796 11772 11848 11824
rect 14004 11772 14056 11824
rect 18512 11772 18564 11824
rect 18972 11772 19024 11824
rect 1860 11568 1912 11620
rect 2044 11543 2096 11552
rect 2044 11509 2053 11543
rect 2053 11509 2087 11543
rect 2087 11509 2096 11543
rect 2044 11500 2096 11509
rect 3884 11679 3936 11688
rect 3884 11645 3893 11679
rect 3893 11645 3927 11679
rect 3927 11645 3936 11679
rect 3884 11636 3936 11645
rect 4988 11636 5040 11688
rect 5172 11679 5224 11688
rect 5172 11645 5181 11679
rect 5181 11645 5215 11679
rect 5215 11645 5224 11679
rect 5172 11636 5224 11645
rect 5356 11704 5408 11756
rect 7104 11704 7156 11756
rect 8116 11704 8168 11756
rect 5724 11679 5776 11688
rect 5724 11645 5733 11679
rect 5733 11645 5767 11679
rect 5767 11645 5776 11679
rect 5724 11636 5776 11645
rect 2596 11500 2648 11552
rect 10508 11636 10560 11688
rect 10876 11636 10928 11688
rect 14740 11704 14792 11756
rect 15200 11704 15252 11756
rect 16212 11704 16264 11756
rect 16856 11704 16908 11756
rect 18880 11704 18932 11756
rect 19616 11704 19668 11756
rect 12900 11679 12952 11688
rect 6092 11500 6144 11552
rect 6460 11500 6512 11552
rect 7472 11500 7524 11552
rect 12900 11645 12909 11679
rect 12909 11645 12943 11679
rect 12943 11645 12952 11679
rect 12900 11636 12952 11645
rect 14464 11636 14516 11688
rect 11796 11611 11848 11620
rect 11796 11577 11805 11611
rect 11805 11577 11839 11611
rect 11839 11577 11848 11611
rect 11796 11568 11848 11577
rect 10416 11500 10468 11552
rect 11612 11500 11664 11552
rect 12716 11500 12768 11552
rect 14556 11568 14608 11620
rect 16580 11611 16632 11620
rect 13360 11500 13412 11552
rect 16580 11577 16589 11611
rect 16589 11577 16623 11611
rect 16623 11577 16632 11611
rect 16580 11568 16632 11577
rect 18696 11611 18748 11620
rect 18696 11577 18705 11611
rect 18705 11577 18739 11611
rect 18739 11577 18748 11611
rect 18696 11568 18748 11577
rect 18788 11611 18840 11620
rect 18788 11577 18797 11611
rect 18797 11577 18831 11611
rect 18831 11577 18840 11611
rect 18788 11568 18840 11577
rect 17408 11543 17460 11552
rect 17408 11509 17417 11543
rect 17417 11509 17451 11543
rect 17451 11509 17460 11543
rect 17408 11500 17460 11509
rect 8315 11398 8367 11450
rect 8379 11398 8431 11450
rect 8443 11398 8495 11450
rect 8507 11398 8559 11450
rect 15648 11398 15700 11450
rect 15712 11398 15764 11450
rect 15776 11398 15828 11450
rect 15840 11398 15892 11450
rect 1584 11339 1636 11348
rect 1584 11305 1593 11339
rect 1593 11305 1627 11339
rect 1627 11305 1636 11339
rect 1584 11296 1636 11305
rect 5172 11339 5224 11348
rect 5172 11305 5181 11339
rect 5181 11305 5215 11339
rect 5215 11305 5224 11339
rect 5172 11296 5224 11305
rect 5356 11296 5408 11348
rect 6184 11296 6236 11348
rect 7104 11339 7156 11348
rect 7104 11305 7113 11339
rect 7113 11305 7147 11339
rect 7147 11305 7156 11339
rect 7104 11296 7156 11305
rect 2228 11160 2280 11212
rect 2596 11160 2648 11212
rect 3424 11160 3476 11212
rect 4436 11228 4488 11280
rect 7472 11271 7524 11280
rect 7472 11237 7481 11271
rect 7481 11237 7515 11271
rect 7515 11237 7524 11271
rect 7472 11228 7524 11237
rect 8208 11228 8260 11280
rect 8668 11271 8720 11280
rect 8668 11237 8677 11271
rect 8677 11237 8711 11271
rect 8711 11237 8720 11271
rect 8668 11228 8720 11237
rect 5080 11160 5132 11212
rect 5448 11160 5500 11212
rect 6184 11203 6236 11212
rect 6184 11169 6193 11203
rect 6193 11169 6227 11203
rect 6227 11169 6236 11203
rect 6184 11160 6236 11169
rect 11244 11339 11296 11348
rect 10416 11228 10468 11280
rect 11244 11305 11253 11339
rect 11253 11305 11287 11339
rect 11287 11305 11296 11339
rect 11244 11296 11296 11305
rect 12900 11339 12952 11348
rect 12900 11305 12909 11339
rect 12909 11305 12943 11339
rect 12943 11305 12952 11339
rect 12900 11296 12952 11305
rect 15200 11296 15252 11348
rect 16856 11339 16908 11348
rect 16856 11305 16865 11339
rect 16865 11305 16899 11339
rect 16899 11305 16908 11339
rect 16856 11296 16908 11305
rect 18788 11296 18840 11348
rect 11612 11228 11664 11280
rect 13544 11228 13596 11280
rect 14556 11228 14608 11280
rect 16028 11228 16080 11280
rect 17408 11228 17460 11280
rect 9864 11160 9916 11212
rect 15384 11160 15436 11212
rect 19616 11228 19668 11280
rect 4528 11092 4580 11144
rect 6460 11135 6512 11144
rect 6460 11101 6469 11135
rect 6469 11101 6503 11135
rect 6503 11101 6512 11135
rect 6460 11092 6512 11101
rect 7380 11135 7432 11144
rect 7380 11101 7389 11135
rect 7389 11101 7423 11135
rect 7423 11101 7432 11135
rect 7380 11092 7432 11101
rect 11428 11092 11480 11144
rect 11888 11135 11940 11144
rect 11888 11101 11897 11135
rect 11897 11101 11931 11135
rect 11931 11101 11940 11135
rect 11888 11092 11940 11101
rect 12440 11092 12492 11144
rect 14004 11135 14056 11144
rect 14004 11101 14013 11135
rect 14013 11101 14047 11135
rect 14047 11101 14056 11135
rect 14004 11092 14056 11101
rect 14740 11092 14792 11144
rect 16488 11092 16540 11144
rect 17684 11092 17736 11144
rect 18788 11092 18840 11144
rect 19156 11135 19208 11144
rect 19156 11101 19165 11135
rect 19165 11101 19199 11135
rect 19199 11101 19208 11135
rect 19156 11092 19208 11101
rect 19524 11135 19576 11144
rect 19524 11101 19533 11135
rect 19533 11101 19567 11135
rect 19567 11101 19576 11135
rect 19524 11092 19576 11101
rect 5816 11024 5868 11076
rect 12532 11067 12584 11076
rect 12532 11033 12541 11067
rect 12541 11033 12575 11067
rect 12575 11033 12584 11067
rect 12532 11024 12584 11033
rect 19708 11024 19760 11076
rect 8392 10999 8444 11008
rect 8392 10965 8401 10999
rect 8401 10965 8435 10999
rect 8435 10965 8444 10999
rect 8392 10956 8444 10965
rect 14280 10999 14332 11008
rect 14280 10965 14289 10999
rect 14289 10965 14323 10999
rect 14323 10965 14332 10999
rect 14280 10956 14332 10965
rect 16304 10956 16356 11008
rect 19064 10956 19116 11008
rect 4648 10854 4700 10906
rect 4712 10854 4764 10906
rect 4776 10854 4828 10906
rect 4840 10854 4892 10906
rect 11982 10854 12034 10906
rect 12046 10854 12098 10906
rect 12110 10854 12162 10906
rect 12174 10854 12226 10906
rect 19315 10854 19367 10906
rect 19379 10854 19431 10906
rect 19443 10854 19495 10906
rect 19507 10854 19559 10906
rect 1676 10591 1728 10600
rect 1676 10557 1694 10591
rect 1694 10557 1728 10591
rect 2228 10752 2280 10804
rect 3056 10752 3108 10804
rect 4160 10752 4212 10804
rect 5080 10752 5132 10804
rect 5448 10752 5500 10804
rect 3884 10684 3936 10736
rect 8392 10752 8444 10804
rect 11612 10795 11664 10804
rect 11612 10761 11621 10795
rect 11621 10761 11655 10795
rect 11655 10761 11664 10795
rect 11612 10752 11664 10761
rect 16304 10795 16356 10804
rect 16304 10761 16313 10795
rect 16313 10761 16347 10795
rect 16347 10761 16356 10795
rect 16304 10752 16356 10761
rect 19616 10795 19668 10804
rect 19616 10761 19625 10795
rect 19625 10761 19659 10795
rect 19659 10761 19668 10795
rect 19616 10752 19668 10761
rect 8852 10616 8904 10668
rect 1676 10548 1728 10557
rect 3884 10591 3936 10600
rect 3884 10557 3893 10591
rect 3893 10557 3927 10591
rect 3927 10557 3936 10591
rect 3884 10548 3936 10557
rect 4068 10591 4120 10600
rect 4068 10557 4077 10591
rect 4077 10557 4111 10591
rect 4111 10557 4120 10591
rect 4068 10548 4120 10557
rect 4436 10548 4488 10600
rect 5448 10591 5500 10600
rect 5448 10557 5457 10591
rect 5457 10557 5491 10591
rect 5491 10557 5500 10591
rect 5448 10548 5500 10557
rect 5632 10548 5684 10600
rect 1952 10412 2004 10464
rect 2964 10412 3016 10464
rect 3056 10455 3108 10464
rect 3056 10421 3065 10455
rect 3065 10421 3099 10455
rect 3099 10421 3108 10455
rect 3424 10455 3476 10464
rect 3056 10412 3108 10421
rect 3424 10421 3433 10455
rect 3433 10421 3467 10455
rect 3467 10421 3476 10455
rect 3424 10412 3476 10421
rect 3976 10412 4028 10464
rect 5632 10412 5684 10464
rect 7564 10548 7616 10600
rect 7472 10480 7524 10532
rect 6184 10455 6236 10464
rect 6184 10421 6193 10455
rect 6193 10421 6227 10455
rect 6227 10421 6236 10455
rect 6184 10412 6236 10421
rect 8024 10480 8076 10532
rect 11520 10616 11572 10668
rect 12532 10616 12584 10668
rect 14004 10616 14056 10668
rect 14648 10659 14700 10668
rect 14648 10625 14657 10659
rect 14657 10625 14691 10659
rect 14691 10625 14700 10659
rect 14648 10616 14700 10625
rect 16488 10659 16540 10668
rect 16488 10625 16497 10659
rect 16497 10625 16531 10659
rect 16531 10625 16540 10659
rect 16488 10616 16540 10625
rect 19708 10616 19760 10668
rect 9772 10591 9824 10600
rect 9772 10557 9781 10591
rect 9781 10557 9815 10591
rect 9815 10557 9824 10591
rect 9772 10548 9824 10557
rect 10416 10412 10468 10464
rect 10876 10480 10928 10532
rect 13452 10523 13504 10532
rect 11520 10412 11572 10464
rect 13452 10489 13461 10523
rect 13461 10489 13495 10523
rect 13495 10489 13504 10523
rect 13452 10480 13504 10489
rect 14464 10523 14516 10532
rect 14464 10489 14473 10523
rect 14473 10489 14507 10523
rect 14507 10489 14516 10523
rect 14464 10480 14516 10489
rect 16304 10480 16356 10532
rect 17132 10523 17184 10532
rect 17132 10489 17141 10523
rect 17141 10489 17175 10523
rect 17175 10489 17184 10523
rect 18604 10523 18656 10532
rect 17132 10480 17184 10489
rect 18604 10489 18613 10523
rect 18613 10489 18647 10523
rect 18647 10489 18656 10523
rect 18604 10480 18656 10489
rect 13544 10412 13596 10464
rect 16028 10412 16080 10464
rect 16948 10412 17000 10464
rect 17684 10412 17736 10464
rect 18328 10455 18380 10464
rect 18328 10421 18337 10455
rect 18337 10421 18371 10455
rect 18371 10421 18380 10455
rect 18328 10412 18380 10421
rect 18788 10412 18840 10464
rect 8315 10310 8367 10362
rect 8379 10310 8431 10362
rect 8443 10310 8495 10362
rect 8507 10310 8559 10362
rect 15648 10310 15700 10362
rect 15712 10310 15764 10362
rect 15776 10310 15828 10362
rect 15840 10310 15892 10362
rect 1676 10251 1728 10260
rect 1676 10217 1685 10251
rect 1685 10217 1719 10251
rect 1719 10217 1728 10251
rect 1676 10208 1728 10217
rect 5448 10251 5500 10260
rect 5448 10217 5457 10251
rect 5457 10217 5491 10251
rect 5491 10217 5500 10251
rect 5448 10208 5500 10217
rect 7380 10251 7432 10260
rect 7380 10217 7389 10251
rect 7389 10217 7423 10251
rect 7423 10217 7432 10251
rect 7380 10208 7432 10217
rect 7564 10208 7616 10260
rect 9588 10208 9640 10260
rect 9864 10251 9916 10260
rect 9864 10217 9873 10251
rect 9873 10217 9907 10251
rect 9907 10217 9916 10251
rect 9864 10208 9916 10217
rect 10876 10251 10928 10260
rect 10876 10217 10885 10251
rect 10885 10217 10919 10251
rect 10919 10217 10928 10251
rect 10876 10208 10928 10217
rect 5724 10140 5776 10192
rect 6092 10183 6144 10192
rect 6092 10149 6101 10183
rect 6101 10149 6135 10183
rect 6135 10149 6144 10183
rect 6092 10140 6144 10149
rect 7656 10183 7708 10192
rect 7656 10149 7665 10183
rect 7665 10149 7699 10183
rect 7699 10149 7708 10183
rect 7656 10140 7708 10149
rect 12808 10208 12860 10260
rect 13544 10251 13596 10260
rect 13544 10217 13553 10251
rect 13553 10217 13587 10251
rect 13587 10217 13596 10251
rect 13544 10208 13596 10217
rect 14004 10208 14056 10260
rect 15384 10208 15436 10260
rect 18328 10208 18380 10260
rect 18604 10208 18656 10260
rect 11244 10183 11296 10192
rect 11244 10149 11253 10183
rect 11253 10149 11287 10183
rect 11287 10149 11296 10183
rect 11244 10140 11296 10149
rect 11428 10140 11480 10192
rect 13360 10140 13412 10192
rect 16948 10140 17000 10192
rect 17776 10140 17828 10192
rect 2320 10072 2372 10124
rect 3056 10072 3108 10124
rect 4528 10115 4580 10124
rect 4528 10081 4537 10115
rect 4537 10081 4571 10115
rect 4571 10081 4580 10115
rect 4528 10072 4580 10081
rect 3516 10004 3568 10056
rect 4068 10004 4120 10056
rect 9956 10072 10008 10124
rect 12440 10115 12492 10124
rect 12440 10081 12449 10115
rect 12449 10081 12483 10115
rect 12483 10081 12492 10115
rect 12440 10072 12492 10081
rect 12624 10115 12676 10124
rect 12624 10081 12633 10115
rect 12633 10081 12667 10115
rect 12667 10081 12676 10115
rect 12624 10072 12676 10081
rect 15108 10072 15160 10124
rect 5816 9936 5868 9988
rect 3516 9868 3568 9920
rect 6000 10047 6052 10056
rect 6000 10013 6009 10047
rect 6009 10013 6043 10047
rect 6043 10013 6052 10047
rect 7564 10047 7616 10056
rect 6000 10004 6052 10013
rect 7564 10013 7573 10047
rect 7573 10013 7607 10047
rect 7607 10013 7616 10047
rect 7564 10004 7616 10013
rect 11152 10047 11204 10056
rect 11152 10013 11161 10047
rect 11161 10013 11195 10047
rect 11195 10013 11204 10047
rect 11152 10004 11204 10013
rect 16304 10004 16356 10056
rect 18788 10047 18840 10056
rect 8852 9936 8904 9988
rect 9864 9936 9916 9988
rect 10140 9936 10192 9988
rect 13084 9936 13136 9988
rect 14004 9936 14056 9988
rect 15936 9936 15988 9988
rect 18788 10013 18797 10047
rect 18797 10013 18831 10047
rect 18831 10013 18840 10047
rect 18788 10004 18840 10013
rect 19616 9936 19668 9988
rect 6828 9868 6880 9920
rect 8668 9911 8720 9920
rect 8668 9877 8677 9911
rect 8677 9877 8711 9911
rect 8711 9877 8720 9911
rect 8668 9868 8720 9877
rect 10416 9868 10468 9920
rect 10692 9868 10744 9920
rect 13728 9868 13780 9920
rect 16488 9868 16540 9920
rect 4648 9766 4700 9818
rect 4712 9766 4764 9818
rect 4776 9766 4828 9818
rect 4840 9766 4892 9818
rect 11982 9766 12034 9818
rect 12046 9766 12098 9818
rect 12110 9766 12162 9818
rect 12174 9766 12226 9818
rect 19315 9766 19367 9818
rect 19379 9766 19431 9818
rect 19443 9766 19495 9818
rect 19507 9766 19559 9818
rect 2320 9707 2372 9716
rect 2320 9673 2329 9707
rect 2329 9673 2363 9707
rect 2363 9673 2372 9707
rect 2320 9664 2372 9673
rect 4252 9664 4304 9716
rect 4436 9664 4488 9716
rect 5908 9664 5960 9716
rect 6092 9664 6144 9716
rect 6644 9664 6696 9716
rect 12808 9707 12860 9716
rect 1584 9639 1636 9648
rect 1584 9605 1593 9639
rect 1593 9605 1627 9639
rect 1627 9605 1636 9639
rect 1584 9596 1636 9605
rect 11152 9596 11204 9648
rect 6828 9571 6880 9580
rect 6828 9537 6837 9571
rect 6837 9537 6871 9571
rect 6871 9537 6880 9571
rect 6828 9528 6880 9537
rect 6920 9528 6972 9580
rect 8668 9571 8720 9580
rect 8668 9537 8677 9571
rect 8677 9537 8711 9571
rect 8711 9537 8720 9571
rect 8668 9528 8720 9537
rect 8944 9571 8996 9580
rect 8944 9537 8953 9571
rect 8953 9537 8987 9571
rect 8987 9537 8996 9571
rect 8944 9528 8996 9537
rect 9588 9528 9640 9580
rect 10600 9528 10652 9580
rect 12808 9673 12817 9707
rect 12817 9673 12851 9707
rect 12851 9673 12860 9707
rect 12808 9664 12860 9673
rect 14464 9664 14516 9716
rect 15108 9664 15160 9716
rect 16028 9664 16080 9716
rect 16304 9664 16356 9716
rect 17776 9664 17828 9716
rect 19064 9707 19116 9716
rect 19064 9673 19073 9707
rect 19073 9673 19107 9707
rect 19107 9673 19116 9707
rect 19064 9664 19116 9673
rect 16580 9596 16632 9648
rect 13728 9571 13780 9580
rect 13728 9537 13737 9571
rect 13737 9537 13771 9571
rect 13771 9537 13780 9571
rect 13728 9528 13780 9537
rect 16948 9528 17000 9580
rect 17132 9571 17184 9580
rect 17132 9537 17141 9571
rect 17141 9537 17175 9571
rect 17175 9537 17184 9571
rect 17132 9528 17184 9537
rect 17592 9528 17644 9580
rect 18144 9571 18196 9580
rect 18144 9537 18153 9571
rect 18153 9537 18187 9571
rect 18187 9537 18196 9571
rect 18144 9528 18196 9537
rect 18696 9596 18748 9648
rect 1308 9460 1360 9512
rect 2228 9460 2280 9512
rect 3424 9503 3476 9512
rect 3424 9469 3433 9503
rect 3433 9469 3467 9503
rect 3467 9469 3476 9503
rect 3424 9460 3476 9469
rect 3608 9503 3660 9512
rect 3608 9469 3617 9503
rect 3617 9469 3651 9503
rect 3651 9469 3660 9503
rect 3608 9460 3660 9469
rect 3700 9460 3752 9512
rect 2964 9392 3016 9444
rect 5264 9435 5316 9444
rect 5264 9401 5273 9435
rect 5273 9401 5307 9435
rect 5307 9401 5316 9435
rect 5264 9392 5316 9401
rect 3056 9367 3108 9376
rect 3056 9333 3065 9367
rect 3065 9333 3099 9367
rect 3099 9333 3108 9367
rect 3056 9324 3108 9333
rect 3884 9367 3936 9376
rect 3884 9333 3893 9367
rect 3893 9333 3927 9367
rect 3927 9333 3936 9367
rect 3884 9324 3936 9333
rect 5080 9324 5132 9376
rect 6368 9392 6420 9444
rect 7656 9460 7708 9512
rect 6552 9367 6604 9376
rect 6552 9333 6561 9367
rect 6561 9333 6595 9367
rect 6595 9333 6604 9367
rect 6552 9324 6604 9333
rect 8208 9324 8260 9376
rect 10692 9392 10744 9444
rect 11336 9392 11388 9444
rect 13360 9392 13412 9444
rect 16488 9435 16540 9444
rect 16488 9401 16497 9435
rect 16497 9401 16531 9435
rect 16531 9401 16540 9435
rect 16488 9392 16540 9401
rect 16580 9435 16632 9444
rect 16580 9401 16589 9435
rect 16589 9401 16623 9435
rect 16623 9401 16632 9435
rect 16580 9392 16632 9401
rect 17776 9392 17828 9444
rect 9956 9324 10008 9376
rect 11244 9324 11296 9376
rect 11888 9324 11940 9376
rect 13820 9324 13872 9376
rect 14188 9324 14240 9376
rect 17500 9324 17552 9376
rect 19616 9324 19668 9376
rect 8315 9222 8367 9274
rect 8379 9222 8431 9274
rect 8443 9222 8495 9274
rect 8507 9222 8559 9274
rect 15648 9222 15700 9274
rect 15712 9222 15764 9274
rect 15776 9222 15828 9274
rect 15840 9222 15892 9274
rect 2504 9120 2556 9172
rect 4528 9120 4580 9172
rect 5080 9163 5132 9172
rect 5080 9129 5089 9163
rect 5089 9129 5123 9163
rect 5123 9129 5132 9163
rect 5080 9120 5132 9129
rect 5264 9120 5316 9172
rect 6368 9120 6420 9172
rect 7748 9120 7800 9172
rect 8944 9120 8996 9172
rect 10600 9163 10652 9172
rect 10600 9129 10609 9163
rect 10609 9129 10643 9163
rect 10643 9129 10652 9163
rect 10600 9120 10652 9129
rect 12624 9163 12676 9172
rect 12624 9129 12633 9163
rect 12633 9129 12667 9163
rect 12667 9129 12676 9163
rect 12624 9120 12676 9129
rect 15016 9120 15068 9172
rect 16396 9120 16448 9172
rect 16948 9163 17000 9172
rect 16948 9129 16957 9163
rect 16957 9129 16991 9163
rect 16991 9129 17000 9163
rect 16948 9120 17000 9129
rect 17500 9163 17552 9172
rect 17500 9129 17509 9163
rect 17509 9129 17543 9163
rect 17543 9129 17552 9163
rect 17500 9120 17552 9129
rect 18144 9163 18196 9172
rect 18144 9129 18153 9163
rect 18153 9129 18187 9163
rect 18187 9129 18196 9163
rect 18144 9120 18196 9129
rect 19064 9120 19116 9172
rect 6920 9052 6972 9104
rect 7472 9052 7524 9104
rect 7564 9052 7616 9104
rect 8760 9095 8812 9104
rect 8760 9061 8769 9095
rect 8769 9061 8803 9095
rect 8803 9061 8812 9095
rect 8760 9052 8812 9061
rect 11888 9052 11940 9104
rect 13728 9052 13780 9104
rect 14648 9052 14700 9104
rect 19156 9052 19208 9104
rect 1952 9027 2004 9036
rect 1952 8993 1961 9027
rect 1961 8993 1995 9027
rect 1995 8993 2004 9027
rect 1952 8984 2004 8993
rect 5080 8984 5132 9036
rect 5632 9027 5684 9036
rect 4160 8959 4212 8968
rect 4160 8925 4169 8959
rect 4169 8925 4203 8959
rect 4203 8925 4212 8959
rect 5632 8993 5641 9027
rect 5641 8993 5675 9027
rect 5675 8993 5684 9027
rect 5632 8984 5684 8993
rect 6092 8984 6144 9036
rect 8208 8984 8260 9036
rect 8668 8984 8720 9036
rect 15476 9027 15528 9036
rect 4160 8916 4212 8925
rect 5448 8916 5500 8968
rect 6644 8916 6696 8968
rect 2504 8848 2556 8900
rect 3976 8848 4028 8900
rect 8116 8916 8168 8968
rect 9312 8916 9364 8968
rect 15476 8993 15485 9027
rect 15485 8993 15519 9027
rect 15519 8993 15528 9027
rect 15476 8984 15528 8993
rect 16488 8984 16540 9036
rect 17592 8984 17644 9036
rect 10416 8916 10468 8968
rect 10968 8916 11020 8968
rect 12348 8916 12400 8968
rect 13452 8959 13504 8968
rect 13452 8925 13461 8959
rect 13461 8925 13495 8959
rect 13495 8925 13504 8959
rect 13452 8916 13504 8925
rect 17408 8916 17460 8968
rect 18236 8916 18288 8968
rect 7380 8848 7432 8900
rect 11704 8848 11756 8900
rect 21548 8848 21600 8900
rect 3700 8823 3752 8832
rect 3700 8789 3709 8823
rect 3709 8789 3743 8823
rect 3743 8789 3752 8823
rect 3700 8780 3752 8789
rect 5356 8780 5408 8832
rect 6000 8780 6052 8832
rect 7196 8780 7248 8832
rect 10508 8780 10560 8832
rect 10968 8823 11020 8832
rect 10968 8789 10977 8823
rect 10977 8789 11011 8823
rect 11011 8789 11020 8823
rect 10968 8780 11020 8789
rect 16212 8780 16264 8832
rect 4648 8678 4700 8730
rect 4712 8678 4764 8730
rect 4776 8678 4828 8730
rect 4840 8678 4892 8730
rect 11982 8678 12034 8730
rect 12046 8678 12098 8730
rect 12110 8678 12162 8730
rect 12174 8678 12226 8730
rect 19315 8678 19367 8730
rect 19379 8678 19431 8730
rect 19443 8678 19495 8730
rect 19507 8678 19559 8730
rect 1952 8619 2004 8628
rect 1952 8585 1961 8619
rect 1961 8585 1995 8619
rect 1995 8585 2004 8619
rect 1952 8576 2004 8585
rect 5448 8576 5500 8628
rect 6276 8619 6328 8628
rect 6276 8585 6285 8619
rect 6285 8585 6319 8619
rect 6319 8585 6328 8619
rect 6276 8576 6328 8585
rect 7380 8619 7432 8628
rect 7380 8585 7389 8619
rect 7389 8585 7423 8619
rect 7423 8585 7432 8619
rect 7380 8576 7432 8585
rect 7472 8576 7524 8628
rect 9496 8576 9548 8628
rect 10416 8619 10468 8628
rect 10416 8585 10425 8619
rect 10425 8585 10459 8619
rect 10459 8585 10468 8619
rect 10416 8576 10468 8585
rect 2964 8508 3016 8560
rect 2044 8372 2096 8424
rect 3332 8415 3384 8424
rect 3332 8381 3341 8415
rect 3341 8381 3375 8415
rect 3375 8381 3384 8415
rect 3332 8372 3384 8381
rect 3700 8508 3752 8560
rect 3884 8508 3936 8560
rect 5172 8508 5224 8560
rect 6460 8508 6512 8560
rect 10232 8508 10284 8560
rect 13728 8619 13780 8628
rect 13728 8585 13737 8619
rect 13737 8585 13771 8619
rect 13771 8585 13780 8619
rect 13728 8576 13780 8585
rect 15476 8619 15528 8628
rect 15476 8585 15485 8619
rect 15485 8585 15519 8619
rect 15519 8585 15528 8619
rect 15476 8576 15528 8585
rect 17500 8576 17552 8628
rect 18328 8576 18380 8628
rect 19156 8619 19208 8628
rect 19156 8585 19165 8619
rect 19165 8585 19199 8619
rect 19199 8585 19208 8619
rect 19156 8576 19208 8585
rect 11888 8508 11940 8560
rect 13084 8551 13136 8560
rect 13084 8517 13093 8551
rect 13093 8517 13127 8551
rect 13127 8517 13136 8551
rect 13084 8508 13136 8517
rect 18788 8551 18840 8560
rect 18788 8517 18797 8551
rect 18797 8517 18831 8551
rect 18831 8517 18840 8551
rect 18788 8508 18840 8517
rect 7748 8483 7800 8492
rect 7748 8449 7757 8483
rect 7757 8449 7791 8483
rect 7791 8449 7800 8483
rect 7748 8440 7800 8449
rect 7932 8440 7984 8492
rect 9220 8483 9272 8492
rect 9220 8449 9229 8483
rect 9229 8449 9263 8483
rect 9263 8449 9272 8483
rect 9220 8440 9272 8449
rect 12716 8440 12768 8492
rect 14648 8440 14700 8492
rect 14924 8440 14976 8492
rect 17684 8440 17736 8492
rect 2596 8279 2648 8288
rect 2596 8245 2605 8279
rect 2605 8245 2639 8279
rect 2639 8245 2648 8279
rect 2596 8236 2648 8245
rect 2964 8279 3016 8288
rect 2964 8245 2973 8279
rect 2973 8245 3007 8279
rect 3007 8245 3016 8279
rect 2964 8236 3016 8245
rect 3056 8236 3108 8288
rect 4068 8236 4120 8288
rect 5172 8304 5224 8356
rect 5356 8236 5408 8288
rect 5540 8279 5592 8288
rect 5540 8245 5549 8279
rect 5549 8245 5583 8279
rect 5583 8245 5592 8279
rect 5540 8236 5592 8245
rect 5632 8236 5684 8288
rect 8024 8304 8076 8356
rect 9496 8347 9548 8356
rect 8116 8236 8168 8288
rect 8668 8279 8720 8288
rect 8668 8245 8677 8279
rect 8677 8245 8711 8279
rect 8711 8245 8720 8279
rect 9496 8313 9505 8347
rect 9505 8313 9539 8347
rect 9539 8313 9548 8347
rect 9496 8304 9548 8313
rect 10324 8304 10376 8356
rect 15292 8372 15344 8424
rect 16212 8372 16264 8424
rect 16396 8415 16448 8424
rect 16396 8381 16405 8415
rect 16405 8381 16439 8415
rect 16439 8381 16448 8415
rect 16396 8372 16448 8381
rect 12532 8304 12584 8356
rect 12624 8347 12676 8356
rect 12624 8313 12633 8347
rect 12633 8313 12667 8347
rect 12667 8313 12676 8347
rect 12624 8304 12676 8313
rect 13268 8304 13320 8356
rect 14648 8304 14700 8356
rect 18328 8347 18380 8356
rect 18328 8313 18337 8347
rect 18337 8313 18371 8347
rect 18371 8313 18380 8347
rect 18328 8304 18380 8313
rect 8668 8236 8720 8245
rect 16948 8279 17000 8288
rect 16948 8245 16957 8279
rect 16957 8245 16991 8279
rect 16991 8245 17000 8279
rect 16948 8236 17000 8245
rect 17408 8279 17460 8288
rect 17408 8245 17417 8279
rect 17417 8245 17451 8279
rect 17451 8245 17460 8279
rect 17408 8236 17460 8245
rect 18972 8236 19024 8288
rect 19892 8236 19944 8288
rect 8315 8134 8367 8186
rect 8379 8134 8431 8186
rect 8443 8134 8495 8186
rect 8507 8134 8559 8186
rect 15648 8134 15700 8186
rect 15712 8134 15764 8186
rect 15776 8134 15828 8186
rect 15840 8134 15892 8186
rect 2504 8075 2556 8084
rect 2504 8041 2513 8075
rect 2513 8041 2547 8075
rect 2547 8041 2556 8075
rect 2504 8032 2556 8041
rect 3056 8032 3108 8084
rect 3332 8032 3384 8084
rect 1952 7896 2004 7948
rect 2412 7896 2464 7948
rect 3240 7896 3292 7948
rect 4160 8032 4212 8084
rect 5540 8032 5592 8084
rect 8852 8075 8904 8084
rect 7932 7964 7984 8016
rect 8116 7964 8168 8016
rect 8852 8041 8861 8075
rect 8861 8041 8895 8075
rect 8895 8041 8904 8075
rect 8852 8032 8904 8041
rect 9220 8075 9272 8084
rect 9220 8041 9229 8075
rect 9229 8041 9263 8075
rect 9263 8041 9272 8075
rect 9220 8032 9272 8041
rect 13268 8032 13320 8084
rect 13544 8032 13596 8084
rect 13728 8032 13780 8084
rect 15384 8032 15436 8084
rect 9404 7964 9456 8016
rect 11336 7964 11388 8016
rect 16580 7964 16632 8016
rect 17500 8007 17552 8016
rect 17500 7973 17509 8007
rect 17509 7973 17543 8007
rect 17543 7973 17552 8007
rect 17500 7964 17552 7973
rect 18144 7964 18196 8016
rect 18512 7964 18564 8016
rect 4436 7896 4488 7948
rect 7104 7896 7156 7948
rect 7656 7939 7708 7948
rect 7656 7905 7665 7939
rect 7665 7905 7699 7939
rect 7699 7905 7708 7939
rect 7656 7896 7708 7905
rect 9772 7896 9824 7948
rect 13452 7896 13504 7948
rect 13912 7896 13964 7948
rect 16120 7896 16172 7948
rect 16396 7896 16448 7948
rect 18880 7939 18932 7948
rect 18880 7905 18889 7939
rect 18889 7905 18923 7939
rect 18923 7905 18932 7939
rect 18880 7896 18932 7905
rect 19064 7896 19116 7948
rect 7932 7871 7984 7880
rect 7932 7837 7941 7871
rect 7941 7837 7975 7871
rect 7975 7837 7984 7871
rect 7932 7828 7984 7837
rect 2872 7760 2924 7812
rect 4436 7692 4488 7744
rect 5080 7760 5132 7812
rect 5816 7692 5868 7744
rect 7288 7735 7340 7744
rect 7288 7701 7297 7735
rect 7297 7701 7331 7735
rect 7331 7701 7340 7735
rect 7288 7692 7340 7701
rect 7748 7760 7800 7812
rect 8300 7828 8352 7880
rect 11612 7828 11664 7880
rect 11428 7760 11480 7812
rect 17132 7828 17184 7880
rect 18236 7828 18288 7880
rect 18420 7760 18472 7812
rect 9864 7692 9916 7744
rect 10692 7692 10744 7744
rect 11796 7735 11848 7744
rect 11796 7701 11805 7735
rect 11805 7701 11839 7735
rect 11839 7701 11848 7735
rect 11796 7692 11848 7701
rect 12624 7692 12676 7744
rect 12716 7692 12768 7744
rect 14648 7692 14700 7744
rect 17132 7735 17184 7744
rect 17132 7701 17141 7735
rect 17141 7701 17175 7735
rect 17175 7701 17184 7735
rect 17132 7692 17184 7701
rect 4648 7590 4700 7642
rect 4712 7590 4764 7642
rect 4776 7590 4828 7642
rect 4840 7590 4892 7642
rect 11982 7590 12034 7642
rect 12046 7590 12098 7642
rect 12110 7590 12162 7642
rect 12174 7590 12226 7642
rect 19315 7590 19367 7642
rect 19379 7590 19431 7642
rect 19443 7590 19495 7642
rect 19507 7590 19559 7642
rect 112 7488 164 7540
rect 1952 7531 2004 7540
rect 1952 7497 1961 7531
rect 1961 7497 1995 7531
rect 1995 7497 2004 7531
rect 1952 7488 2004 7497
rect 3240 7488 3292 7540
rect 4528 7488 4580 7540
rect 7104 7488 7156 7540
rect 8852 7488 8904 7540
rect 9680 7488 9732 7540
rect 3056 7352 3108 7404
rect 2320 7284 2372 7336
rect 2964 7284 3016 7336
rect 3792 7327 3844 7336
rect 3792 7293 3801 7327
rect 3801 7293 3835 7327
rect 3835 7293 3844 7327
rect 3792 7284 3844 7293
rect 5540 7420 5592 7472
rect 7288 7352 7340 7404
rect 4528 7284 4580 7336
rect 4988 7284 5040 7336
rect 5632 7327 5684 7336
rect 5632 7293 5641 7327
rect 5641 7293 5675 7327
rect 5675 7293 5684 7327
rect 5632 7284 5684 7293
rect 9772 7420 9824 7472
rect 8116 7352 8168 7404
rect 10600 7488 10652 7540
rect 11612 7531 11664 7540
rect 11612 7497 11621 7531
rect 11621 7497 11655 7531
rect 11655 7497 11664 7531
rect 11612 7488 11664 7497
rect 14648 7531 14700 7540
rect 14648 7497 14657 7531
rect 14657 7497 14691 7531
rect 14691 7497 14700 7531
rect 14648 7488 14700 7497
rect 15384 7531 15436 7540
rect 15384 7497 15393 7531
rect 15393 7497 15427 7531
rect 15427 7497 15436 7531
rect 15384 7488 15436 7497
rect 16120 7531 16172 7540
rect 16120 7497 16129 7531
rect 16129 7497 16163 7531
rect 16163 7497 16172 7531
rect 16120 7488 16172 7497
rect 17500 7531 17552 7540
rect 17500 7497 17509 7531
rect 17509 7497 17543 7531
rect 17543 7497 17552 7531
rect 17500 7488 17552 7497
rect 17592 7488 17644 7540
rect 13452 7420 13504 7472
rect 3884 7216 3936 7268
rect 4620 7148 4672 7200
rect 5632 7148 5684 7200
rect 6460 7148 6512 7200
rect 8116 7191 8168 7200
rect 8116 7157 8125 7191
rect 8125 7157 8159 7191
rect 8159 7157 8168 7191
rect 8116 7148 8168 7157
rect 9404 7327 9456 7336
rect 9404 7293 9413 7327
rect 9413 7293 9447 7327
rect 9447 7293 9456 7327
rect 9404 7284 9456 7293
rect 8760 7259 8812 7268
rect 8760 7225 8769 7259
rect 8769 7225 8803 7259
rect 8803 7225 8812 7259
rect 8760 7216 8812 7225
rect 9496 7148 9548 7200
rect 15476 7420 15528 7472
rect 16396 7420 16448 7472
rect 16672 7420 16724 7472
rect 16488 7352 16540 7404
rect 18880 7352 18932 7404
rect 11520 7284 11572 7336
rect 11336 7259 11388 7268
rect 11336 7225 11345 7259
rect 11345 7225 11379 7259
rect 11379 7225 11388 7259
rect 11336 7216 11388 7225
rect 14372 7216 14424 7268
rect 12808 7191 12860 7200
rect 12808 7157 12817 7191
rect 12817 7157 12851 7191
rect 12851 7157 12860 7191
rect 12808 7148 12860 7157
rect 13544 7191 13596 7200
rect 13544 7157 13553 7191
rect 13553 7157 13587 7191
rect 13587 7157 13596 7191
rect 13544 7148 13596 7157
rect 16580 7259 16632 7268
rect 16580 7225 16589 7259
rect 16589 7225 16623 7259
rect 16623 7225 16632 7259
rect 18144 7259 18196 7268
rect 16580 7216 16632 7225
rect 18144 7225 18153 7259
rect 18153 7225 18187 7259
rect 18187 7225 18196 7259
rect 18144 7216 18196 7225
rect 17040 7148 17092 7200
rect 18328 7216 18380 7268
rect 18512 7148 18564 7200
rect 19064 7191 19116 7200
rect 19064 7157 19073 7191
rect 19073 7157 19107 7191
rect 19107 7157 19116 7191
rect 19064 7148 19116 7157
rect 19708 7148 19760 7200
rect 8315 7046 8367 7098
rect 8379 7046 8431 7098
rect 8443 7046 8495 7098
rect 8507 7046 8559 7098
rect 15648 7046 15700 7098
rect 15712 7046 15764 7098
rect 15776 7046 15828 7098
rect 15840 7046 15892 7098
rect 2320 6919 2372 6928
rect 2320 6885 2329 6919
rect 2329 6885 2363 6919
rect 2363 6885 2372 6919
rect 2320 6876 2372 6885
rect 3792 6876 3844 6928
rect 4068 6876 4120 6928
rect 6460 6876 6512 6928
rect 8116 6944 8168 6996
rect 10968 6944 11020 6996
rect 11060 6944 11112 6996
rect 11336 6944 11388 6996
rect 16488 6944 16540 6996
rect 16580 6944 16632 6996
rect 17040 6987 17092 6996
rect 17040 6953 17049 6987
rect 17049 6953 17083 6987
rect 17083 6953 17092 6987
rect 17040 6944 17092 6953
rect 19524 6987 19576 6996
rect 19524 6953 19533 6987
rect 19533 6953 19567 6987
rect 19567 6953 19576 6987
rect 19524 6944 19576 6953
rect 8944 6876 8996 6928
rect 11428 6876 11480 6928
rect 11796 6876 11848 6928
rect 12348 6876 12400 6928
rect 15476 6876 15528 6928
rect 2504 6851 2556 6860
rect 2504 6817 2513 6851
rect 2513 6817 2547 6851
rect 2547 6817 2556 6851
rect 2504 6808 2556 6817
rect 2872 6851 2924 6860
rect 2872 6817 2881 6851
rect 2881 6817 2915 6851
rect 2915 6817 2924 6851
rect 2872 6808 2924 6817
rect 5264 6851 5316 6860
rect 5264 6817 5273 6851
rect 5273 6817 5307 6851
rect 5307 6817 5316 6851
rect 5264 6808 5316 6817
rect 5632 6808 5684 6860
rect 8208 6808 8260 6860
rect 8760 6808 8812 6860
rect 3148 6783 3200 6792
rect 3148 6749 3157 6783
rect 3157 6749 3191 6783
rect 3191 6749 3200 6783
rect 3148 6740 3200 6749
rect 3884 6740 3936 6792
rect 7380 6740 7432 6792
rect 7932 6783 7984 6792
rect 7932 6749 7941 6783
rect 7941 6749 7975 6783
rect 7975 6749 7984 6783
rect 7932 6740 7984 6749
rect 1952 6672 2004 6724
rect 9772 6672 9824 6724
rect 10140 6808 10192 6860
rect 12532 6808 12584 6860
rect 13452 6808 13504 6860
rect 10508 6783 10560 6792
rect 10508 6749 10517 6783
rect 10517 6749 10551 6783
rect 10551 6749 10560 6783
rect 10508 6740 10560 6749
rect 13176 6740 13228 6792
rect 16580 6808 16632 6860
rect 16948 6808 17000 6860
rect 18052 6808 18104 6860
rect 19156 6808 19208 6860
rect 15016 6740 15068 6792
rect 10048 6715 10100 6724
rect 10048 6681 10057 6715
rect 10057 6681 10091 6715
rect 10091 6681 10100 6715
rect 13728 6715 13780 6724
rect 10048 6672 10100 6681
rect 13728 6681 13737 6715
rect 13737 6681 13771 6715
rect 13771 6681 13780 6715
rect 13728 6672 13780 6681
rect 2044 6604 2096 6656
rect 3976 6604 4028 6656
rect 4436 6604 4488 6656
rect 5172 6604 5224 6656
rect 9956 6604 10008 6656
rect 10968 6647 11020 6656
rect 10968 6613 10977 6647
rect 10977 6613 11011 6647
rect 11011 6613 11020 6647
rect 10968 6604 11020 6613
rect 13544 6604 13596 6656
rect 17316 6604 17368 6656
rect 18512 6647 18564 6656
rect 18512 6613 18521 6647
rect 18521 6613 18555 6647
rect 18555 6613 18564 6647
rect 18512 6604 18564 6613
rect 4648 6502 4700 6554
rect 4712 6502 4764 6554
rect 4776 6502 4828 6554
rect 4840 6502 4892 6554
rect 11982 6502 12034 6554
rect 12046 6502 12098 6554
rect 12110 6502 12162 6554
rect 12174 6502 12226 6554
rect 19315 6502 19367 6554
rect 19379 6502 19431 6554
rect 19443 6502 19495 6554
rect 19507 6502 19559 6554
rect 6276 6400 6328 6452
rect 6736 6400 6788 6452
rect 8116 6400 8168 6452
rect 9956 6400 10008 6452
rect 11612 6400 11664 6452
rect 11796 6443 11848 6452
rect 11796 6409 11805 6443
rect 11805 6409 11839 6443
rect 11839 6409 11848 6443
rect 11796 6400 11848 6409
rect 13452 6400 13504 6452
rect 15476 6443 15528 6452
rect 15476 6409 15485 6443
rect 15485 6409 15519 6443
rect 15519 6409 15528 6443
rect 15476 6400 15528 6409
rect 19156 6400 19208 6452
rect 19616 6400 19668 6452
rect 4252 6332 4304 6384
rect 10048 6332 10100 6384
rect 11428 6332 11480 6384
rect 2964 6264 3016 6316
rect 3976 6264 4028 6316
rect 3240 6196 3292 6248
rect 3884 6239 3936 6248
rect 3884 6205 3893 6239
rect 3893 6205 3927 6239
rect 3927 6205 3936 6239
rect 3884 6196 3936 6205
rect 9036 6264 9088 6316
rect 9956 6264 10008 6316
rect 15016 6307 15068 6316
rect 15016 6273 15025 6307
rect 15025 6273 15059 6307
rect 15059 6273 15068 6307
rect 15016 6264 15068 6273
rect 16028 6332 16080 6384
rect 16304 6307 16356 6316
rect 6184 6239 6236 6248
rect 6184 6205 6193 6239
rect 6193 6205 6227 6239
rect 6227 6205 6236 6239
rect 6184 6196 6236 6205
rect 7288 6239 7340 6248
rect 7288 6205 7297 6239
rect 7297 6205 7331 6239
rect 7331 6205 7340 6239
rect 7288 6196 7340 6205
rect 10140 6196 10192 6248
rect 12348 6196 12400 6248
rect 15108 6196 15160 6248
rect 15476 6196 15528 6248
rect 16304 6273 16313 6307
rect 16313 6273 16347 6307
rect 16347 6273 16356 6307
rect 16304 6264 16356 6273
rect 18420 6307 18472 6316
rect 18420 6273 18429 6307
rect 18429 6273 18463 6307
rect 18463 6273 18472 6307
rect 18420 6264 18472 6273
rect 17500 6196 17552 6248
rect 6368 6128 6420 6180
rect 7472 6128 7524 6180
rect 8944 6171 8996 6180
rect 8944 6137 8953 6171
rect 8953 6137 8987 6171
rect 8987 6137 8996 6171
rect 8944 6128 8996 6137
rect 9588 6171 9640 6180
rect 2320 6060 2372 6112
rect 3332 6060 3384 6112
rect 4620 6103 4672 6112
rect 4620 6069 4629 6103
rect 4629 6069 4663 6103
rect 4663 6069 4672 6103
rect 5448 6103 5500 6112
rect 4620 6060 4672 6069
rect 5448 6069 5457 6103
rect 5457 6069 5491 6103
rect 5491 6069 5500 6103
rect 5448 6060 5500 6069
rect 6460 6060 6512 6112
rect 7840 6060 7892 6112
rect 8760 6060 8812 6112
rect 9588 6137 9597 6171
rect 9597 6137 9631 6171
rect 9631 6137 9640 6171
rect 9588 6128 9640 6137
rect 10508 6171 10560 6180
rect 9404 6060 9456 6112
rect 10508 6137 10517 6171
rect 10517 6137 10551 6171
rect 10551 6137 10560 6171
rect 10508 6128 10560 6137
rect 10968 6128 11020 6180
rect 12532 6128 12584 6180
rect 13728 6128 13780 6180
rect 14188 6128 14240 6180
rect 18144 6171 18196 6180
rect 13176 6060 13228 6112
rect 16580 6103 16632 6112
rect 16580 6069 16589 6103
rect 16589 6069 16623 6103
rect 16623 6069 16632 6103
rect 16580 6060 16632 6069
rect 18144 6137 18153 6171
rect 18153 6137 18187 6171
rect 18187 6137 18196 6171
rect 18144 6128 18196 6137
rect 18512 6128 18564 6180
rect 8315 5958 8367 6010
rect 8379 5958 8431 6010
rect 8443 5958 8495 6010
rect 8507 5958 8559 6010
rect 15648 5958 15700 6010
rect 15712 5958 15764 6010
rect 15776 5958 15828 6010
rect 15840 5958 15892 6010
rect 4344 5856 4396 5908
rect 5264 5856 5316 5908
rect 6552 5899 6604 5908
rect 6552 5865 6561 5899
rect 6561 5865 6595 5899
rect 6595 5865 6604 5899
rect 6552 5856 6604 5865
rect 7288 5856 7340 5908
rect 7380 5899 7432 5908
rect 7380 5865 7389 5899
rect 7389 5865 7423 5899
rect 7423 5865 7432 5899
rect 7840 5899 7892 5908
rect 7380 5856 7432 5865
rect 7840 5865 7849 5899
rect 7849 5865 7883 5899
rect 7883 5865 7892 5899
rect 7840 5856 7892 5865
rect 9128 5856 9180 5908
rect 10048 5856 10100 5908
rect 2228 5720 2280 5772
rect 2320 5720 2372 5772
rect 3884 5720 3936 5772
rect 4344 5763 4396 5772
rect 3148 5695 3200 5704
rect 3148 5661 3157 5695
rect 3157 5661 3191 5695
rect 3191 5661 3200 5695
rect 3148 5652 3200 5661
rect 4344 5729 4353 5763
rect 4353 5729 4387 5763
rect 4387 5729 4396 5763
rect 4344 5720 4396 5729
rect 5908 5763 5960 5772
rect 5908 5729 5917 5763
rect 5917 5729 5951 5763
rect 5951 5729 5960 5763
rect 5908 5720 5960 5729
rect 9312 5788 9364 5840
rect 9496 5720 9548 5772
rect 14188 5899 14240 5908
rect 14188 5865 14197 5899
rect 14197 5865 14231 5899
rect 14231 5865 14240 5899
rect 14188 5856 14240 5865
rect 17408 5856 17460 5908
rect 13176 5831 13228 5840
rect 11796 5720 11848 5772
rect 6368 5652 6420 5704
rect 7472 5695 7524 5704
rect 7472 5661 7481 5695
rect 7481 5661 7515 5695
rect 7515 5661 7524 5695
rect 7472 5652 7524 5661
rect 9404 5652 9456 5704
rect 9772 5695 9824 5704
rect 9772 5661 9781 5695
rect 9781 5661 9815 5695
rect 9815 5661 9824 5695
rect 9772 5652 9824 5661
rect 10416 5695 10468 5704
rect 10416 5661 10425 5695
rect 10425 5661 10459 5695
rect 10459 5661 10468 5695
rect 10416 5652 10468 5661
rect 10508 5652 10560 5704
rect 2504 5627 2556 5636
rect 2504 5593 2513 5627
rect 2513 5593 2547 5627
rect 2547 5593 2556 5627
rect 2504 5584 2556 5593
rect 4436 5627 4488 5636
rect 4436 5593 4445 5627
rect 4445 5593 4479 5627
rect 4479 5593 4488 5627
rect 4436 5584 4488 5593
rect 6184 5627 6236 5636
rect 6184 5593 6193 5627
rect 6193 5593 6227 5627
rect 6227 5593 6236 5627
rect 13176 5797 13185 5831
rect 13185 5797 13219 5831
rect 13219 5797 13228 5831
rect 13176 5788 13228 5797
rect 16120 5831 16172 5840
rect 16120 5797 16129 5831
rect 16129 5797 16163 5831
rect 16163 5797 16172 5831
rect 16120 5788 16172 5797
rect 16672 5831 16724 5840
rect 16672 5797 16681 5831
rect 16681 5797 16715 5831
rect 16715 5797 16724 5831
rect 16672 5788 16724 5797
rect 17684 5831 17736 5840
rect 17684 5797 17693 5831
rect 17693 5797 17727 5831
rect 17727 5797 17736 5831
rect 17684 5788 17736 5797
rect 18420 5788 18472 5840
rect 13452 5763 13504 5772
rect 13452 5729 13461 5763
rect 13461 5729 13495 5763
rect 13495 5729 13504 5763
rect 13452 5720 13504 5729
rect 13636 5652 13688 5704
rect 16948 5652 17000 5704
rect 17592 5695 17644 5704
rect 17592 5661 17601 5695
rect 17601 5661 17635 5695
rect 17635 5661 17644 5695
rect 17592 5652 17644 5661
rect 19156 5720 19208 5772
rect 6184 5584 6236 5593
rect 2320 5559 2372 5568
rect 2320 5525 2329 5559
rect 2329 5525 2363 5559
rect 2363 5525 2372 5559
rect 2320 5516 2372 5525
rect 5172 5516 5224 5568
rect 6276 5516 6328 5568
rect 11244 5516 11296 5568
rect 15476 5584 15528 5636
rect 16764 5584 16816 5636
rect 12440 5516 12492 5568
rect 19064 5584 19116 5636
rect 19616 5584 19668 5636
rect 18236 5516 18288 5568
rect 4648 5414 4700 5466
rect 4712 5414 4764 5466
rect 4776 5414 4828 5466
rect 4840 5414 4892 5466
rect 11982 5414 12034 5466
rect 12046 5414 12098 5466
rect 12110 5414 12162 5466
rect 12174 5414 12226 5466
rect 19315 5414 19367 5466
rect 19379 5414 19431 5466
rect 19443 5414 19495 5466
rect 19507 5414 19559 5466
rect 1952 5312 2004 5364
rect 2688 5312 2740 5364
rect 4252 5312 4304 5364
rect 7472 5312 7524 5364
rect 5908 5244 5960 5296
rect 10324 5312 10376 5364
rect 11796 5355 11848 5364
rect 11796 5321 11805 5355
rect 11805 5321 11839 5355
rect 11839 5321 11848 5355
rect 11796 5312 11848 5321
rect 9128 5244 9180 5296
rect 16120 5312 16172 5364
rect 17684 5312 17736 5364
rect 19064 5312 19116 5364
rect 19892 5312 19944 5364
rect 2504 5219 2556 5228
rect 2504 5185 2513 5219
rect 2513 5185 2547 5219
rect 2547 5185 2556 5219
rect 2504 5176 2556 5185
rect 3976 5176 4028 5228
rect 4160 5176 4212 5228
rect 5356 5176 5408 5228
rect 5540 5176 5592 5228
rect 6368 5176 6420 5228
rect 8668 5176 8720 5228
rect 9956 5176 10008 5228
rect 2688 5108 2740 5160
rect 3700 5151 3752 5160
rect 3700 5117 3709 5151
rect 3709 5117 3743 5151
rect 3743 5117 3752 5151
rect 3884 5151 3936 5160
rect 3700 5108 3752 5117
rect 3884 5117 3893 5151
rect 3893 5117 3927 5151
rect 3927 5117 3936 5151
rect 3884 5108 3936 5117
rect 4528 5108 4580 5160
rect 5172 5151 5224 5160
rect 5172 5117 5181 5151
rect 5181 5117 5215 5151
rect 5215 5117 5224 5151
rect 5172 5108 5224 5117
rect 5448 5151 5500 5160
rect 5448 5117 5457 5151
rect 5457 5117 5491 5151
rect 5491 5117 5500 5151
rect 5448 5108 5500 5117
rect 7380 5151 7432 5160
rect 7380 5117 7389 5151
rect 7389 5117 7423 5151
rect 7423 5117 7432 5151
rect 7380 5108 7432 5117
rect 10784 5151 10836 5160
rect 10784 5117 10793 5151
rect 10793 5117 10827 5151
rect 10827 5117 10836 5151
rect 10784 5108 10836 5117
rect 16764 5244 16816 5296
rect 16948 5287 17000 5296
rect 16948 5253 16957 5287
rect 16957 5253 16991 5287
rect 16991 5253 17000 5287
rect 16948 5244 17000 5253
rect 12348 5176 12400 5228
rect 16672 5176 16724 5228
rect 18328 5176 18380 5228
rect 18512 5176 18564 5228
rect 11060 5151 11112 5160
rect 4344 5040 4396 5092
rect 2136 5015 2188 5024
rect 2136 4981 2145 5015
rect 2145 4981 2179 5015
rect 2179 4981 2188 5015
rect 2136 4972 2188 4981
rect 2872 4972 2924 5024
rect 7472 4972 7524 5024
rect 7840 5040 7892 5092
rect 9312 5083 9364 5092
rect 9312 5049 9321 5083
rect 9321 5049 9355 5083
rect 9355 5049 9364 5083
rect 10600 5083 10652 5092
rect 9312 5040 9364 5049
rect 10600 5049 10609 5083
rect 10609 5049 10643 5083
rect 10643 5049 10652 5083
rect 11060 5117 11069 5151
rect 11069 5117 11103 5151
rect 11103 5117 11112 5151
rect 11060 5108 11112 5117
rect 12440 5151 12492 5160
rect 12440 5117 12449 5151
rect 12449 5117 12483 5151
rect 12483 5117 12492 5151
rect 12440 5108 12492 5117
rect 13452 5108 13504 5160
rect 15476 5108 15528 5160
rect 10600 5040 10652 5049
rect 11612 5040 11664 5092
rect 10232 4972 10284 5024
rect 11244 5015 11296 5024
rect 11244 4981 11253 5015
rect 11253 4981 11287 5015
rect 11287 4981 11296 5015
rect 11244 4972 11296 4981
rect 12348 5040 12400 5092
rect 16580 5040 16632 5092
rect 16764 5040 16816 5092
rect 18236 5083 18288 5092
rect 18236 5049 18245 5083
rect 18245 5049 18279 5083
rect 18279 5049 18288 5083
rect 18236 5040 18288 5049
rect 18972 5040 19024 5092
rect 13452 5015 13504 5024
rect 13452 4981 13461 5015
rect 13461 4981 13495 5015
rect 13495 4981 13504 5015
rect 13452 4972 13504 4981
rect 17684 4972 17736 5024
rect 19156 4972 19208 5024
rect 8315 4870 8367 4922
rect 8379 4870 8431 4922
rect 8443 4870 8495 4922
rect 8507 4870 8559 4922
rect 15648 4870 15700 4922
rect 15712 4870 15764 4922
rect 15776 4870 15828 4922
rect 15840 4870 15892 4922
rect 4528 4768 4580 4820
rect 6184 4768 6236 4820
rect 6276 4811 6328 4820
rect 6276 4777 6285 4811
rect 6285 4777 6319 4811
rect 6319 4777 6328 4811
rect 6276 4768 6328 4777
rect 9312 4768 9364 4820
rect 9588 4768 9640 4820
rect 10416 4768 10468 4820
rect 3240 4700 3292 4752
rect 6368 4700 6420 4752
rect 7380 4700 7432 4752
rect 8208 4743 8260 4752
rect 8208 4709 8217 4743
rect 8217 4709 8251 4743
rect 8251 4709 8260 4743
rect 8208 4700 8260 4709
rect 9864 4743 9916 4752
rect 9864 4709 9873 4743
rect 9873 4709 9907 4743
rect 9907 4709 9916 4743
rect 9864 4700 9916 4709
rect 1308 4632 1360 4684
rect 1860 4632 1912 4684
rect 2412 4675 2464 4684
rect 2412 4641 2421 4675
rect 2421 4641 2455 4675
rect 2455 4641 2464 4675
rect 2412 4632 2464 4641
rect 3792 4675 3844 4684
rect 2320 4564 2372 4616
rect 3792 4641 3801 4675
rect 3801 4641 3835 4675
rect 3835 4641 3844 4675
rect 3792 4632 3844 4641
rect 4436 4632 4488 4684
rect 5172 4675 5224 4684
rect 5172 4641 5181 4675
rect 5181 4641 5215 4675
rect 5215 4641 5224 4675
rect 5172 4632 5224 4641
rect 5356 4675 5408 4684
rect 5356 4641 5365 4675
rect 5365 4641 5399 4675
rect 5399 4641 5408 4675
rect 5356 4632 5408 4641
rect 2964 4564 3016 4616
rect 7012 4675 7064 4684
rect 7012 4641 7021 4675
rect 7021 4641 7055 4675
rect 7055 4641 7064 4675
rect 7012 4632 7064 4641
rect 7288 4632 7340 4684
rect 11796 4675 11848 4684
rect 11796 4641 11805 4675
rect 11805 4641 11839 4675
rect 11839 4641 11848 4675
rect 12440 4700 12492 4752
rect 11796 4632 11848 4641
rect 12624 4700 12676 4752
rect 17684 4768 17736 4820
rect 18236 4768 18288 4820
rect 18328 4768 18380 4820
rect 19616 4811 19668 4820
rect 19616 4777 19625 4811
rect 19625 4777 19659 4811
rect 19659 4777 19668 4811
rect 19616 4768 19668 4777
rect 16764 4700 16816 4752
rect 18788 4743 18840 4752
rect 18788 4709 18797 4743
rect 18797 4709 18831 4743
rect 18831 4709 18840 4743
rect 18788 4700 18840 4709
rect 14832 4632 14884 4684
rect 7932 4564 7984 4616
rect 8116 4607 8168 4616
rect 8116 4573 8125 4607
rect 8125 4573 8159 4607
rect 8159 4573 8168 4607
rect 8116 4564 8168 4573
rect 9956 4564 10008 4616
rect 2228 4496 2280 4548
rect 9680 4496 9732 4548
rect 11520 4564 11572 4616
rect 12440 4607 12492 4616
rect 11888 4496 11940 4548
rect 12440 4573 12449 4607
rect 12449 4573 12483 4607
rect 12483 4573 12492 4607
rect 12440 4564 12492 4573
rect 14372 4607 14424 4616
rect 14372 4573 14381 4607
rect 14381 4573 14415 4607
rect 14415 4573 14424 4607
rect 14372 4564 14424 4573
rect 15384 4607 15436 4616
rect 15384 4573 15393 4607
rect 15393 4573 15427 4607
rect 15427 4573 15436 4607
rect 15384 4564 15436 4573
rect 16028 4607 16080 4616
rect 16028 4573 16037 4607
rect 16037 4573 16071 4607
rect 16071 4573 16080 4607
rect 16028 4564 16080 4573
rect 17132 4564 17184 4616
rect 18420 4564 18472 4616
rect 18972 4607 19024 4616
rect 18972 4573 18981 4607
rect 18981 4573 19015 4607
rect 19015 4573 19024 4607
rect 18972 4564 19024 4573
rect 15292 4496 15344 4548
rect 15476 4496 15528 4548
rect 1952 4428 2004 4480
rect 6644 4428 6696 4480
rect 7472 4471 7524 4480
rect 7472 4437 7481 4471
rect 7481 4437 7515 4471
rect 7515 4437 7524 4471
rect 7472 4428 7524 4437
rect 7564 4428 7616 4480
rect 11060 4428 11112 4480
rect 11428 4471 11480 4480
rect 11428 4437 11437 4471
rect 11437 4437 11471 4471
rect 11471 4437 11480 4471
rect 11428 4428 11480 4437
rect 4648 4326 4700 4378
rect 4712 4326 4764 4378
rect 4776 4326 4828 4378
rect 4840 4326 4892 4378
rect 11982 4326 12034 4378
rect 12046 4326 12098 4378
rect 12110 4326 12162 4378
rect 12174 4326 12226 4378
rect 19315 4326 19367 4378
rect 19379 4326 19431 4378
rect 19443 4326 19495 4378
rect 19507 4326 19559 4378
rect 2228 4156 2280 4208
rect 2504 4156 2556 4208
rect 2872 4156 2924 4208
rect 8668 4224 8720 4276
rect 9864 4224 9916 4276
rect 12716 4224 12768 4276
rect 14372 4224 14424 4276
rect 15844 4224 15896 4276
rect 18788 4224 18840 4276
rect 4988 4156 5040 4208
rect 9680 4156 9732 4208
rect 11888 4156 11940 4208
rect 12624 4156 12676 4208
rect 14832 4199 14884 4208
rect 14832 4165 14841 4199
rect 14841 4165 14875 4199
rect 14875 4165 14884 4199
rect 14832 4156 14884 4165
rect 2964 4088 3016 4140
rect 3148 4088 3200 4140
rect 2320 4063 2372 4072
rect 2320 4029 2329 4063
rect 2329 4029 2363 4063
rect 2363 4029 2372 4063
rect 2320 4020 2372 4029
rect 2504 4020 2556 4072
rect 3608 4020 3660 4072
rect 3884 4063 3936 4072
rect 3884 4029 3893 4063
rect 3893 4029 3927 4063
rect 3927 4029 3936 4063
rect 3884 4020 3936 4029
rect 4160 4063 4212 4072
rect 4160 4029 4169 4063
rect 4169 4029 4203 4063
rect 4203 4029 4212 4063
rect 4160 4020 4212 4029
rect 4436 4020 4488 4072
rect 4988 4020 5040 4072
rect 6184 4063 6236 4072
rect 6184 4029 6193 4063
rect 6193 4029 6227 4063
rect 6227 4029 6236 4063
rect 6184 4020 6236 4029
rect 7104 4063 7156 4072
rect 7104 4029 7113 4063
rect 7113 4029 7147 4063
rect 7147 4029 7156 4063
rect 7104 4020 7156 4029
rect 8208 4020 8260 4072
rect 3516 3952 3568 4004
rect 2412 3884 2464 3936
rect 4068 3884 4120 3936
rect 6644 3927 6696 3936
rect 6644 3893 6653 3927
rect 6653 3893 6687 3927
rect 6687 3893 6696 3927
rect 6644 3884 6696 3893
rect 7472 3927 7524 3936
rect 7472 3893 7481 3927
rect 7481 3893 7515 3927
rect 7515 3893 7524 3927
rect 7472 3884 7524 3893
rect 7656 3884 7708 3936
rect 8852 4020 8904 4072
rect 11428 4020 11480 4072
rect 13544 4088 13596 4140
rect 13452 4063 13504 4072
rect 13452 4029 13461 4063
rect 13461 4029 13495 4063
rect 13495 4029 13504 4063
rect 13452 4020 13504 4029
rect 12532 3995 12584 4004
rect 8760 3927 8812 3936
rect 8760 3893 8769 3927
rect 8769 3893 8803 3927
rect 8803 3893 8812 3927
rect 8760 3884 8812 3893
rect 8944 3884 8996 3936
rect 12532 3961 12541 3995
rect 12541 3961 12575 3995
rect 12575 3961 12584 3995
rect 12532 3952 12584 3961
rect 13912 4063 13964 4072
rect 13912 4029 13921 4063
rect 13921 4029 13955 4063
rect 13955 4029 13964 4063
rect 13912 4020 13964 4029
rect 18236 4020 18288 4072
rect 14924 3952 14976 4004
rect 15844 3995 15896 4004
rect 15844 3961 15853 3995
rect 15853 3961 15887 3995
rect 15887 3961 15896 3995
rect 15844 3952 15896 3961
rect 16028 3952 16080 4004
rect 16396 3995 16448 4004
rect 16396 3961 16405 3995
rect 16405 3961 16439 3995
rect 16439 3961 16448 3995
rect 16396 3952 16448 3961
rect 10416 3884 10468 3936
rect 12624 3884 12676 3936
rect 16764 3884 16816 3936
rect 16948 3927 17000 3936
rect 16948 3893 16957 3927
rect 16957 3893 16991 3927
rect 16991 3893 17000 3927
rect 16948 3884 17000 3893
rect 17132 3884 17184 3936
rect 8315 3782 8367 3834
rect 8379 3782 8431 3834
rect 8443 3782 8495 3834
rect 8507 3782 8559 3834
rect 15648 3782 15700 3834
rect 15712 3782 15764 3834
rect 15776 3782 15828 3834
rect 15840 3782 15892 3834
rect 2780 3680 2832 3732
rect 3516 3723 3568 3732
rect 3516 3689 3525 3723
rect 3525 3689 3559 3723
rect 3559 3689 3568 3723
rect 3516 3680 3568 3689
rect 3792 3723 3844 3732
rect 3792 3689 3801 3723
rect 3801 3689 3835 3723
rect 3835 3689 3844 3723
rect 3792 3680 3844 3689
rect 3884 3680 3936 3732
rect 4988 3680 5040 3732
rect 6184 3680 6236 3732
rect 4528 3612 4580 3664
rect 5264 3612 5316 3664
rect 2412 3587 2464 3596
rect 2412 3553 2421 3587
rect 2421 3553 2455 3587
rect 2455 3553 2464 3587
rect 2412 3544 2464 3553
rect 3424 3544 3476 3596
rect 5540 3587 5592 3596
rect 5540 3553 5549 3587
rect 5549 3553 5583 3587
rect 5583 3553 5592 3587
rect 5540 3544 5592 3553
rect 6460 3587 6512 3596
rect 6460 3553 6469 3587
rect 6469 3553 6503 3587
rect 6503 3553 6512 3587
rect 6460 3544 6512 3553
rect 7012 3680 7064 3732
rect 7288 3680 7340 3732
rect 7104 3612 7156 3664
rect 10140 3680 10192 3732
rect 11244 3680 11296 3732
rect 12532 3723 12584 3732
rect 12532 3689 12541 3723
rect 12541 3689 12575 3723
rect 12575 3689 12584 3723
rect 12532 3680 12584 3689
rect 13912 3680 13964 3732
rect 15384 3680 15436 3732
rect 8760 3612 8812 3664
rect 9864 3655 9916 3664
rect 9864 3621 9873 3655
rect 9873 3621 9907 3655
rect 9907 3621 9916 3655
rect 9864 3612 9916 3621
rect 9956 3612 10008 3664
rect 16396 3680 16448 3732
rect 18420 3680 18472 3732
rect 19064 3723 19116 3732
rect 19064 3689 19073 3723
rect 19073 3689 19107 3723
rect 19107 3689 19116 3723
rect 19064 3680 19116 3689
rect 7656 3544 7708 3596
rect 10784 3544 10836 3596
rect 11244 3544 11296 3596
rect 11888 3544 11940 3596
rect 12440 3544 12492 3596
rect 13176 3544 13228 3596
rect 13360 3544 13412 3596
rect 14280 3587 14332 3596
rect 14280 3553 14289 3587
rect 14289 3553 14323 3587
rect 14323 3553 14332 3587
rect 14280 3544 14332 3553
rect 7564 3476 7616 3528
rect 9588 3476 9640 3528
rect 12624 3476 12676 3528
rect 13636 3476 13688 3528
rect 1768 3408 1820 3460
rect 2504 3451 2556 3460
rect 2504 3417 2513 3451
rect 2513 3417 2547 3451
rect 2547 3417 2556 3451
rect 2504 3408 2556 3417
rect 9680 3408 9732 3460
rect 10324 3451 10376 3460
rect 10324 3417 10333 3451
rect 10333 3417 10367 3451
rect 10367 3417 10376 3451
rect 10324 3408 10376 3417
rect 10876 3451 10928 3460
rect 10876 3417 10885 3451
rect 10885 3417 10919 3451
rect 10919 3417 10928 3451
rect 10876 3408 10928 3417
rect 12348 3408 12400 3460
rect 15844 3655 15896 3664
rect 15844 3621 15853 3655
rect 15853 3621 15887 3655
rect 15887 3621 15896 3655
rect 15844 3612 15896 3621
rect 17224 3612 17276 3664
rect 17408 3612 17460 3664
rect 19156 3612 19208 3664
rect 16396 3587 16448 3596
rect 16396 3553 16405 3587
rect 16405 3553 16439 3587
rect 16439 3553 16448 3587
rect 17316 3587 17368 3596
rect 16396 3544 16448 3553
rect 17316 3553 17325 3587
rect 17325 3553 17359 3587
rect 17359 3553 17368 3587
rect 17316 3544 17368 3553
rect 14556 3476 14608 3528
rect 15844 3476 15896 3528
rect 16212 3476 16264 3528
rect 16764 3408 16816 3460
rect 16856 3408 16908 3460
rect 19064 3544 19116 3596
rect 2320 3340 2372 3392
rect 5540 3340 5592 3392
rect 9036 3383 9088 3392
rect 9036 3349 9045 3383
rect 9045 3349 9079 3383
rect 9079 3349 9088 3383
rect 9036 3340 9088 3349
rect 9312 3340 9364 3392
rect 14924 3340 14976 3392
rect 18236 3383 18288 3392
rect 18236 3349 18245 3383
rect 18245 3349 18279 3383
rect 18279 3349 18288 3383
rect 18236 3340 18288 3349
rect 4648 3238 4700 3290
rect 4712 3238 4764 3290
rect 4776 3238 4828 3290
rect 4840 3238 4892 3290
rect 11982 3238 12034 3290
rect 12046 3238 12098 3290
rect 12110 3238 12162 3290
rect 12174 3238 12226 3290
rect 19315 3238 19367 3290
rect 19379 3238 19431 3290
rect 19443 3238 19495 3290
rect 19507 3238 19559 3290
rect 2412 3136 2464 3188
rect 3424 3179 3476 3188
rect 3424 3145 3433 3179
rect 3433 3145 3467 3179
rect 3467 3145 3476 3179
rect 3424 3136 3476 3145
rect 5540 3136 5592 3188
rect 6184 3136 6236 3188
rect 7196 3136 7248 3188
rect 8852 3136 8904 3188
rect 9864 3179 9916 3188
rect 9864 3145 9873 3179
rect 9873 3145 9907 3179
rect 9907 3145 9916 3179
rect 9864 3136 9916 3145
rect 10140 3179 10192 3188
rect 10140 3145 10149 3179
rect 10149 3145 10183 3179
rect 10183 3145 10192 3179
rect 10140 3136 10192 3145
rect 11244 3136 11296 3188
rect 12348 3136 12400 3188
rect 12624 3179 12676 3188
rect 12624 3145 12633 3179
rect 12633 3145 12667 3179
rect 12667 3145 12676 3179
rect 12624 3136 12676 3145
rect 14280 3136 14332 3188
rect 15844 3136 15896 3188
rect 17316 3136 17368 3188
rect 19156 3179 19208 3188
rect 19156 3145 19165 3179
rect 19165 3145 19199 3179
rect 19199 3145 19208 3179
rect 19156 3136 19208 3145
rect 8760 3068 8812 3120
rect 10876 3111 10928 3120
rect 10876 3077 10885 3111
rect 10885 3077 10919 3111
rect 10919 3077 10928 3111
rect 10876 3068 10928 3077
rect 9036 3000 9088 3052
rect 13360 3068 13412 3120
rect 11520 3043 11572 3052
rect 11520 3009 11529 3043
rect 11529 3009 11563 3043
rect 11563 3009 11572 3043
rect 11520 3000 11572 3009
rect 3148 2932 3200 2984
rect 3792 2975 3844 2984
rect 3792 2941 3801 2975
rect 3801 2941 3835 2975
rect 3835 2941 3844 2975
rect 3792 2932 3844 2941
rect 4160 2975 4212 2984
rect 4160 2941 4169 2975
rect 4169 2941 4203 2975
rect 4203 2941 4212 2975
rect 4160 2932 4212 2941
rect 4988 2932 5040 2984
rect 5724 2975 5776 2984
rect 5724 2941 5733 2975
rect 5733 2941 5767 2975
rect 5767 2941 5776 2975
rect 5724 2932 5776 2941
rect 5908 2975 5960 2984
rect 5908 2941 5917 2975
rect 5917 2941 5951 2975
rect 5951 2941 5960 2975
rect 5908 2932 5960 2941
rect 6828 2932 6880 2984
rect 10784 2975 10836 2984
rect 3884 2864 3936 2916
rect 4344 2907 4396 2916
rect 4344 2873 4353 2907
rect 4353 2873 4387 2907
rect 4387 2873 4396 2907
rect 4344 2864 4396 2873
rect 4528 2864 4580 2916
rect 8576 2907 8628 2916
rect 1768 2796 1820 2848
rect 7288 2839 7340 2848
rect 7288 2805 7297 2839
rect 7297 2805 7331 2839
rect 7331 2805 7340 2839
rect 7288 2796 7340 2805
rect 7748 2796 7800 2848
rect 8576 2873 8579 2907
rect 8579 2873 8613 2907
rect 8613 2873 8628 2907
rect 8576 2864 8628 2873
rect 10784 2941 10793 2975
rect 10793 2941 10827 2975
rect 10827 2941 10836 2975
rect 10784 2932 10836 2941
rect 10876 2932 10928 2984
rect 11888 2932 11940 2984
rect 13176 2975 13228 2984
rect 13176 2941 13185 2975
rect 13185 2941 13219 2975
rect 13219 2941 13228 2975
rect 13176 2932 13228 2941
rect 13636 2975 13688 2984
rect 13636 2941 13645 2975
rect 13645 2941 13679 2975
rect 13679 2941 13688 2975
rect 13636 2932 13688 2941
rect 16396 3043 16448 3052
rect 16396 3009 16405 3043
rect 16405 3009 16439 3043
rect 16439 3009 16448 3043
rect 16396 3000 16448 3009
rect 17592 3068 17644 3120
rect 19064 3000 19116 3052
rect 16764 2932 16816 2984
rect 18696 2975 18748 2984
rect 18696 2941 18705 2975
rect 18705 2941 18739 2975
rect 18739 2941 18748 2975
rect 18696 2932 18748 2941
rect 19708 2975 19760 2984
rect 19708 2941 19726 2975
rect 19726 2941 19760 2975
rect 19708 2932 19760 2941
rect 16212 2907 16264 2916
rect 16212 2873 16221 2907
rect 16221 2873 16255 2907
rect 16255 2873 16264 2907
rect 16212 2864 16264 2873
rect 10784 2796 10836 2848
rect 11888 2839 11940 2848
rect 11888 2805 11897 2839
rect 11897 2805 11931 2839
rect 11931 2805 11940 2839
rect 11888 2796 11940 2805
rect 14280 2839 14332 2848
rect 14280 2805 14289 2839
rect 14289 2805 14323 2839
rect 14323 2805 14332 2839
rect 14280 2796 14332 2805
rect 8315 2694 8367 2746
rect 8379 2694 8431 2746
rect 8443 2694 8495 2746
rect 8507 2694 8559 2746
rect 15648 2694 15700 2746
rect 15712 2694 15764 2746
rect 15776 2694 15828 2746
rect 15840 2694 15892 2746
rect 1860 2635 1912 2644
rect 1860 2601 1869 2635
rect 1869 2601 1903 2635
rect 1903 2601 1912 2635
rect 1860 2592 1912 2601
rect 3148 2592 3200 2644
rect 3792 2635 3844 2644
rect 3792 2601 3801 2635
rect 3801 2601 3835 2635
rect 3835 2601 3844 2635
rect 3792 2592 3844 2601
rect 4160 2592 4212 2644
rect 5724 2592 5776 2644
rect 6460 2635 6512 2644
rect 6460 2601 6469 2635
rect 6469 2601 6503 2635
rect 6503 2601 6512 2635
rect 6460 2592 6512 2601
rect 10876 2635 10928 2644
rect 10876 2601 10885 2635
rect 10885 2601 10919 2635
rect 10919 2601 10928 2635
rect 10876 2592 10928 2601
rect 11244 2635 11296 2644
rect 11244 2601 11253 2635
rect 11253 2601 11287 2635
rect 11287 2601 11296 2635
rect 11244 2592 11296 2601
rect 13176 2635 13228 2644
rect 13176 2601 13185 2635
rect 13185 2601 13219 2635
rect 13219 2601 13228 2635
rect 13176 2592 13228 2601
rect 13544 2635 13596 2644
rect 13544 2601 13553 2635
rect 13553 2601 13587 2635
rect 13587 2601 13596 2635
rect 13544 2592 13596 2601
rect 5908 2524 5960 2576
rect 6368 2524 6420 2576
rect 3056 2456 3108 2508
rect 4068 2456 4120 2508
rect 1400 2431 1452 2440
rect 1400 2397 1409 2431
rect 1409 2397 1443 2431
rect 1443 2397 1452 2431
rect 1400 2388 1452 2397
rect 3976 2320 4028 2372
rect 5724 2456 5776 2508
rect 7656 2524 7708 2576
rect 7748 2524 7800 2576
rect 8668 2524 8720 2576
rect 11428 2499 11480 2508
rect 11428 2465 11437 2499
rect 11437 2465 11471 2499
rect 11471 2465 11480 2499
rect 11428 2456 11480 2465
rect 12440 2499 12492 2508
rect 12440 2465 12449 2499
rect 12449 2465 12483 2499
rect 12483 2465 12492 2499
rect 14280 2592 14332 2644
rect 18144 2592 18196 2644
rect 13820 2524 13872 2576
rect 12440 2456 12492 2465
rect 16580 2524 16632 2576
rect 9312 2388 9364 2440
rect 10324 2431 10376 2440
rect 10324 2397 10333 2431
rect 10333 2397 10367 2431
rect 10367 2397 10376 2431
rect 10324 2388 10376 2397
rect 15936 2499 15988 2508
rect 15936 2465 15945 2499
rect 15945 2465 15979 2499
rect 15979 2465 15988 2499
rect 15936 2456 15988 2465
rect 15016 2320 15068 2372
rect 16948 2524 17000 2576
rect 7748 2295 7800 2304
rect 7748 2261 7757 2295
rect 7757 2261 7791 2295
rect 7791 2261 7800 2295
rect 7748 2252 7800 2261
rect 14556 2295 14608 2304
rect 14556 2261 14565 2295
rect 14565 2261 14599 2295
rect 14599 2261 14608 2295
rect 14556 2252 14608 2261
rect 15200 2295 15252 2304
rect 15200 2261 15209 2295
rect 15209 2261 15243 2295
rect 15243 2261 15252 2295
rect 15200 2252 15252 2261
rect 18052 2295 18104 2304
rect 18052 2261 18061 2295
rect 18061 2261 18095 2295
rect 18095 2261 18104 2295
rect 18512 2388 18564 2440
rect 18788 2388 18840 2440
rect 18052 2252 18104 2261
rect 4648 2150 4700 2202
rect 4712 2150 4764 2202
rect 4776 2150 4828 2202
rect 4840 2150 4892 2202
rect 11982 2150 12034 2202
rect 12046 2150 12098 2202
rect 12110 2150 12162 2202
rect 12174 2150 12226 2202
rect 19315 2150 19367 2202
rect 19379 2150 19431 2202
rect 19443 2150 19495 2202
rect 19507 2150 19559 2202
rect 3148 2048 3200 2100
rect 6644 2048 6696 2100
rect 7748 2048 7800 2100
rect 12440 2048 12492 2100
rect 18512 2048 18564 2100
rect 940 76 992 128
rect 3976 76 4028 128
rect 7288 8 7340 60
rect 12900 8 12952 60
<< metal2 >>
rect 1214 21570 1270 22000
rect 3606 21570 3662 22000
rect 1214 21542 1532 21570
rect 1214 21520 1270 21542
rect 1504 16658 1532 21542
rect 3344 21542 3662 21570
rect 2502 20496 2558 20505
rect 2502 20431 2558 20440
rect 1582 18728 1638 18737
rect 1582 18663 1638 18672
rect 1596 18426 1624 18663
rect 1584 18420 1636 18426
rect 1584 18362 1636 18368
rect 1582 16824 1638 16833
rect 1582 16759 1638 16768
rect 1492 16652 1544 16658
rect 1492 16594 1544 16600
rect 1596 16250 1624 16759
rect 1584 16244 1636 16250
rect 1584 16186 1636 16192
rect 1308 16108 1360 16114
rect 1308 16050 1360 16056
rect 1320 13433 1348 16050
rect 2228 14952 2280 14958
rect 2228 14894 2280 14900
rect 1306 13424 1362 13433
rect 1306 13359 1362 13368
rect 1320 9518 1348 13359
rect 2044 12300 2096 12306
rect 2044 12242 2096 12248
rect 1860 12164 1912 12170
rect 1860 12106 1912 12112
rect 1872 11626 1900 12106
rect 1860 11620 1912 11626
rect 1860 11562 1912 11568
rect 2056 11558 2084 12242
rect 2044 11552 2096 11558
rect 1582 11520 1638 11529
rect 2044 11494 2096 11500
rect 1582 11455 1638 11464
rect 1596 11354 1624 11455
rect 1584 11348 1636 11354
rect 1584 11290 1636 11296
rect 1676 10600 1728 10606
rect 1676 10542 1728 10548
rect 1688 10266 1716 10542
rect 1952 10464 2004 10470
rect 1952 10406 2004 10412
rect 1676 10260 1728 10266
rect 1676 10202 1728 10208
rect 1964 10169 1992 10406
rect 1950 10160 2006 10169
rect 1950 10095 2006 10104
rect 1582 9752 1638 9761
rect 1582 9687 1638 9696
rect 1596 9654 1624 9687
rect 1584 9648 1636 9654
rect 1584 9590 1636 9596
rect 1308 9512 1360 9518
rect 1308 9454 1360 9460
rect 112 7540 164 7546
rect 112 7482 164 7488
rect 124 6361 152 7482
rect 110 6352 166 6361
rect 110 6287 166 6296
rect 1320 4690 1348 9454
rect 1952 9036 2004 9042
rect 1952 8978 2004 8984
rect 1964 8634 1992 8978
rect 1952 8628 2004 8634
rect 1952 8570 2004 8576
rect 1964 8537 1992 8570
rect 1950 8528 2006 8537
rect 1950 8463 2006 8472
rect 2056 8430 2084 11494
rect 2240 11218 2268 14894
rect 2410 13288 2466 13297
rect 2410 13223 2466 13232
rect 2228 11212 2280 11218
rect 2228 11154 2280 11160
rect 2240 10810 2268 11154
rect 2228 10804 2280 10810
rect 2228 10746 2280 10752
rect 2320 10124 2372 10130
rect 2320 10066 2372 10072
rect 2332 9722 2360 10066
rect 2320 9716 2372 9722
rect 2320 9658 2372 9664
rect 2228 9512 2280 9518
rect 2228 9454 2280 9460
rect 2044 8424 2096 8430
rect 2044 8366 2096 8372
rect 1952 7948 2004 7954
rect 1952 7890 2004 7896
rect 1964 7546 1992 7890
rect 1952 7540 2004 7546
rect 1952 7482 2004 7488
rect 1952 6724 2004 6730
rect 1952 6666 2004 6672
rect 1964 5370 1992 6666
rect 2044 6656 2096 6662
rect 2044 6598 2096 6604
rect 1952 5364 2004 5370
rect 1952 5306 2004 5312
rect 1308 4684 1360 4690
rect 1308 4626 1360 4632
rect 1860 4684 1912 4690
rect 1860 4626 1912 4632
rect 1768 3460 1820 3466
rect 1768 3402 1820 3408
rect 1780 2854 1808 3402
rect 1768 2848 1820 2854
rect 1768 2790 1820 2796
rect 1400 2440 1452 2446
rect 1400 2382 1452 2388
rect 1412 1737 1440 2382
rect 1398 1728 1454 1737
rect 1398 1663 1454 1672
rect 1780 1465 1808 2790
rect 1872 2650 1900 4626
rect 1952 4480 2004 4486
rect 2056 4457 2084 6598
rect 2240 5778 2268 9454
rect 2424 7954 2452 13223
rect 2516 9178 2544 20431
rect 3344 18426 3372 21542
rect 3606 21520 3662 21542
rect 6090 21570 6146 22000
rect 8482 21570 8538 22000
rect 10966 21570 11022 22000
rect 6090 21542 6408 21570
rect 6090 21520 6146 21542
rect 4622 19612 4918 19632
rect 4678 19610 4702 19612
rect 4758 19610 4782 19612
rect 4838 19610 4862 19612
rect 4700 19558 4702 19610
rect 4764 19558 4776 19610
rect 4838 19558 4840 19610
rect 4678 19556 4702 19558
rect 4758 19556 4782 19558
rect 4838 19556 4862 19558
rect 4622 19536 4918 19556
rect 4622 18524 4918 18544
rect 4678 18522 4702 18524
rect 4758 18522 4782 18524
rect 4838 18522 4862 18524
rect 4700 18470 4702 18522
rect 4764 18470 4776 18522
rect 4838 18470 4840 18522
rect 4678 18468 4702 18470
rect 4758 18468 4782 18470
rect 4838 18468 4862 18470
rect 4622 18448 4918 18468
rect 2780 18420 2832 18426
rect 2780 18362 2832 18368
rect 3332 18420 3384 18426
rect 3332 18362 3384 18368
rect 2688 13320 2740 13326
rect 2688 13262 2740 13268
rect 2596 11552 2648 11558
rect 2596 11494 2648 11500
rect 2608 11218 2636 11494
rect 2596 11212 2648 11218
rect 2596 11154 2648 11160
rect 2504 9172 2556 9178
rect 2504 9114 2556 9120
rect 2504 8900 2556 8906
rect 2504 8842 2556 8848
rect 2516 8090 2544 8842
rect 2596 8288 2648 8294
rect 2596 8230 2648 8236
rect 2504 8084 2556 8090
rect 2504 8026 2556 8032
rect 2412 7948 2464 7954
rect 2412 7890 2464 7896
rect 2320 7336 2372 7342
rect 2320 7278 2372 7284
rect 2332 6934 2360 7278
rect 2320 6928 2372 6934
rect 2320 6870 2372 6876
rect 2516 6866 2544 8026
rect 2608 7993 2636 8230
rect 2594 7984 2650 7993
rect 2594 7919 2650 7928
rect 2504 6860 2556 6866
rect 2504 6802 2556 6808
rect 2516 6361 2544 6802
rect 2502 6352 2558 6361
rect 2502 6287 2558 6296
rect 2320 6112 2372 6118
rect 2320 6054 2372 6060
rect 2332 5778 2360 6054
rect 2228 5772 2280 5778
rect 2228 5714 2280 5720
rect 2320 5772 2372 5778
rect 2320 5714 2372 5720
rect 2332 5574 2360 5714
rect 2504 5636 2556 5642
rect 2504 5578 2556 5584
rect 2320 5568 2372 5574
rect 2320 5510 2372 5516
rect 2332 5137 2360 5510
rect 2516 5234 2544 5578
rect 2700 5370 2728 13262
rect 2792 12986 2820 18362
rect 4622 17436 4918 17456
rect 4678 17434 4702 17436
rect 4758 17434 4782 17436
rect 4838 17434 4862 17436
rect 4700 17382 4702 17434
rect 4764 17382 4776 17434
rect 4838 17382 4840 17434
rect 4678 17380 4702 17382
rect 4758 17380 4782 17382
rect 4838 17380 4862 17382
rect 4622 17360 4918 17380
rect 4986 17232 5042 17241
rect 4986 17167 5042 17176
rect 2872 16652 2924 16658
rect 2872 16594 2924 16600
rect 2884 14482 2912 16594
rect 4622 16348 4918 16368
rect 4678 16346 4702 16348
rect 4758 16346 4782 16348
rect 4838 16346 4862 16348
rect 4700 16294 4702 16346
rect 4764 16294 4776 16346
rect 4838 16294 4840 16346
rect 4678 16292 4702 16294
rect 4758 16292 4782 16294
rect 4838 16292 4862 16294
rect 4622 16272 4918 16292
rect 2964 15904 3016 15910
rect 2964 15846 3016 15852
rect 2872 14476 2924 14482
rect 2872 14418 2924 14424
rect 2884 13326 2912 14418
rect 2872 13320 2924 13326
rect 2872 13262 2924 13268
rect 2872 13184 2924 13190
rect 2872 13126 2924 13132
rect 2884 12986 2912 13126
rect 2780 12980 2832 12986
rect 2780 12922 2832 12928
rect 2872 12980 2924 12986
rect 2872 12922 2924 12928
rect 2792 12306 2820 12922
rect 2976 12782 3004 15846
rect 4622 15260 4918 15280
rect 4678 15258 4702 15260
rect 4758 15258 4782 15260
rect 4838 15258 4862 15260
rect 4700 15206 4702 15258
rect 4764 15206 4776 15258
rect 4838 15206 4840 15258
rect 4678 15204 4702 15206
rect 4758 15204 4782 15206
rect 4838 15204 4862 15206
rect 4622 15184 4918 15204
rect 3330 15056 3386 15065
rect 3330 14991 3386 15000
rect 2964 12776 3016 12782
rect 2964 12718 3016 12724
rect 3056 12640 3108 12646
rect 3056 12582 3108 12588
rect 2780 12300 2832 12306
rect 2780 12242 2832 12248
rect 2792 11898 2820 12242
rect 2780 11892 2832 11898
rect 2780 11834 2832 11840
rect 3068 11121 3096 12582
rect 3148 12096 3200 12102
rect 3148 12038 3200 12044
rect 3160 11393 3188 12038
rect 3146 11384 3202 11393
rect 3146 11319 3202 11328
rect 3054 11112 3110 11121
rect 3054 11047 3110 11056
rect 3056 10804 3108 10810
rect 3056 10746 3108 10752
rect 3068 10470 3096 10746
rect 3344 10713 3372 14991
rect 4342 14920 4398 14929
rect 4342 14855 4398 14864
rect 4252 14272 4304 14278
rect 4252 14214 4304 14220
rect 4160 13864 4212 13870
rect 4160 13806 4212 13812
rect 3976 13456 4028 13462
rect 3976 13398 4028 13404
rect 3988 12986 4016 13398
rect 3976 12980 4028 12986
rect 3976 12922 4028 12928
rect 3516 12640 3568 12646
rect 3516 12582 3568 12588
rect 3528 11257 3556 12582
rect 3884 12232 3936 12238
rect 3884 12174 3936 12180
rect 3896 11694 3924 12174
rect 3884 11688 3936 11694
rect 3884 11630 3936 11636
rect 3514 11248 3570 11257
rect 3424 11212 3476 11218
rect 3514 11183 3570 11192
rect 3424 11154 3476 11160
rect 3330 10704 3386 10713
rect 3252 10662 3330 10690
rect 2964 10464 3016 10470
rect 2964 10406 3016 10412
rect 3056 10464 3108 10470
rect 3056 10406 3108 10412
rect 2976 9450 3004 10406
rect 3068 10130 3096 10406
rect 3056 10124 3108 10130
rect 3056 10066 3108 10072
rect 2964 9444 3016 9450
rect 2964 9386 3016 9392
rect 3068 9382 3096 10066
rect 3056 9376 3108 9382
rect 3056 9318 3108 9324
rect 3068 8809 3096 9318
rect 3054 8800 3110 8809
rect 3054 8735 3110 8744
rect 2964 8560 3016 8566
rect 2964 8502 3016 8508
rect 2976 8294 3004 8502
rect 2964 8288 3016 8294
rect 2964 8230 3016 8236
rect 3056 8288 3108 8294
rect 3056 8230 3108 8236
rect 2872 7812 2924 7818
rect 2872 7754 2924 7760
rect 2884 6866 2912 7754
rect 2976 7342 3004 8230
rect 3068 8090 3096 8230
rect 3056 8084 3108 8090
rect 3056 8026 3108 8032
rect 3068 7410 3096 8026
rect 3252 7954 3280 10662
rect 3330 10639 3386 10648
rect 3436 10470 3464 11154
rect 3896 10742 3924 11630
rect 4172 10810 4200 13806
rect 4160 10804 4212 10810
rect 4160 10746 4212 10752
rect 3884 10736 3936 10742
rect 3884 10678 3936 10684
rect 3896 10606 3924 10678
rect 3884 10600 3936 10606
rect 3884 10542 3936 10548
rect 4068 10600 4120 10606
rect 4068 10542 4120 10548
rect 3424 10464 3476 10470
rect 3424 10406 3476 10412
rect 3976 10464 4028 10470
rect 3976 10406 4028 10412
rect 3436 9518 3464 10406
rect 3516 10056 3568 10062
rect 3516 9998 3568 10004
rect 3528 9926 3556 9998
rect 3516 9920 3568 9926
rect 3516 9862 3568 9868
rect 3528 9674 3556 9862
rect 3528 9646 3740 9674
rect 3712 9518 3740 9646
rect 3424 9512 3476 9518
rect 3424 9454 3476 9460
rect 3608 9512 3660 9518
rect 3608 9454 3660 9460
rect 3700 9512 3752 9518
rect 3700 9454 3752 9460
rect 3436 9353 3464 9454
rect 3422 9344 3478 9353
rect 3422 9279 3478 9288
rect 3332 8424 3384 8430
rect 3332 8366 3384 8372
rect 3344 8090 3372 8366
rect 3332 8084 3384 8090
rect 3332 8026 3384 8032
rect 3240 7948 3292 7954
rect 3240 7890 3292 7896
rect 3252 7546 3280 7890
rect 3240 7540 3292 7546
rect 3240 7482 3292 7488
rect 3056 7404 3108 7410
rect 3056 7346 3108 7352
rect 2964 7336 3016 7342
rect 2964 7278 3016 7284
rect 2872 6860 2924 6866
rect 2924 6820 3004 6848
rect 2872 6802 2924 6808
rect 2778 6352 2834 6361
rect 2976 6322 3004 6820
rect 3148 6792 3200 6798
rect 3148 6734 3200 6740
rect 2778 6287 2834 6296
rect 2964 6316 3016 6322
rect 2688 5364 2740 5370
rect 2688 5306 2740 5312
rect 2504 5228 2556 5234
rect 2504 5170 2556 5176
rect 2700 5166 2728 5306
rect 2688 5160 2740 5166
rect 2318 5128 2374 5137
rect 2688 5102 2740 5108
rect 2318 5063 2374 5072
rect 2136 5024 2188 5030
rect 2136 4966 2188 4972
rect 1952 4422 2004 4428
rect 2042 4448 2098 4457
rect 1964 3097 1992 4422
rect 2042 4383 2098 4392
rect 2148 3777 2176 4966
rect 2412 4684 2464 4690
rect 2412 4626 2464 4632
rect 2320 4616 2372 4622
rect 2320 4558 2372 4564
rect 2228 4548 2280 4554
rect 2228 4490 2280 4496
rect 2240 4214 2268 4490
rect 2228 4208 2280 4214
rect 2228 4150 2280 4156
rect 2332 4078 2360 4558
rect 2320 4072 2372 4078
rect 2320 4014 2372 4020
rect 2134 3768 2190 3777
rect 2134 3703 2190 3712
rect 2332 3398 2360 4014
rect 2424 3942 2452 4626
rect 2504 4208 2556 4214
rect 2504 4150 2556 4156
rect 2516 4078 2544 4150
rect 2504 4072 2556 4078
rect 2504 4014 2556 4020
rect 2412 3936 2464 3942
rect 2412 3878 2464 3884
rect 2424 3602 2452 3878
rect 2412 3596 2464 3602
rect 2412 3538 2464 3544
rect 2320 3392 2372 3398
rect 2320 3334 2372 3340
rect 2424 3194 2452 3538
rect 2516 3466 2544 4014
rect 2792 3738 2820 6287
rect 2964 6258 3016 6264
rect 3160 5817 3188 6734
rect 3240 6248 3292 6254
rect 3240 6190 3292 6196
rect 3146 5808 3202 5817
rect 3146 5743 3202 5752
rect 3148 5704 3200 5710
rect 3148 5646 3200 5652
rect 2872 5024 2924 5030
rect 2872 4966 2924 4972
rect 2884 4214 2912 4966
rect 2964 4616 3016 4622
rect 2964 4558 3016 4564
rect 2872 4208 2924 4214
rect 2872 4150 2924 4156
rect 2976 4146 3004 4558
rect 3160 4146 3188 5646
rect 3252 4758 3280 6190
rect 3332 6112 3384 6118
rect 3332 6054 3384 6060
rect 3240 4752 3292 4758
rect 3240 4694 3292 4700
rect 2964 4140 3016 4146
rect 2964 4082 3016 4088
rect 3148 4140 3200 4146
rect 3148 4082 3200 4088
rect 2780 3732 2832 3738
rect 2780 3674 2832 3680
rect 2504 3460 2556 3466
rect 2504 3402 2556 3408
rect 2412 3188 2464 3194
rect 2412 3130 2464 3136
rect 1950 3088 2006 3097
rect 1950 3023 2006 3032
rect 3160 2990 3188 4082
rect 3148 2984 3200 2990
rect 3344 2961 3372 6054
rect 3620 4154 3648 9454
rect 3712 8838 3740 9454
rect 3884 9376 3936 9382
rect 3884 9318 3936 9324
rect 3700 8832 3752 8838
rect 3700 8774 3752 8780
rect 3712 8566 3740 8774
rect 3896 8566 3924 9318
rect 3988 8906 4016 10406
rect 4080 10062 4108 10542
rect 4068 10056 4120 10062
rect 4068 9998 4120 10004
rect 4264 9722 4292 14214
rect 4252 9716 4304 9722
rect 4252 9658 4304 9664
rect 4066 9072 4122 9081
rect 4066 9007 4122 9016
rect 3976 8900 4028 8906
rect 3976 8842 4028 8848
rect 3700 8560 3752 8566
rect 3700 8502 3752 8508
rect 3884 8560 3936 8566
rect 3884 8502 3936 8508
rect 4080 8294 4108 9007
rect 4160 8968 4212 8974
rect 4160 8910 4212 8916
rect 4068 8288 4120 8294
rect 4068 8230 4120 8236
rect 3790 7440 3846 7449
rect 3790 7375 3846 7384
rect 3804 7342 3832 7375
rect 3792 7336 3844 7342
rect 3792 7278 3844 7284
rect 3804 6934 3832 7278
rect 3884 7268 3936 7274
rect 3884 7210 3936 7216
rect 3792 6928 3844 6934
rect 3792 6870 3844 6876
rect 3698 5264 3754 5273
rect 3698 5199 3754 5208
rect 3712 5166 3740 5199
rect 3700 5160 3752 5166
rect 3700 5102 3752 5108
rect 3804 4690 3832 6870
rect 3896 6798 3924 7210
rect 4080 7018 4108 8230
rect 4172 8090 4200 8910
rect 4160 8084 4212 8090
rect 4160 8026 4212 8032
rect 3988 6990 4108 7018
rect 3884 6792 3936 6798
rect 3884 6734 3936 6740
rect 3988 6662 4016 6990
rect 4068 6928 4120 6934
rect 4068 6870 4120 6876
rect 3976 6656 4028 6662
rect 3896 6616 3976 6644
rect 3896 6254 3924 6616
rect 3976 6598 4028 6604
rect 3976 6316 4028 6322
rect 3976 6258 4028 6264
rect 3884 6248 3936 6254
rect 3884 6190 3936 6196
rect 3884 5772 3936 5778
rect 3884 5714 3936 5720
rect 3896 5166 3924 5714
rect 3988 5234 4016 6258
rect 3976 5228 4028 5234
rect 3976 5170 4028 5176
rect 3884 5160 3936 5166
rect 3884 5102 3936 5108
rect 3792 4684 3844 4690
rect 3844 4644 3924 4672
rect 3792 4626 3844 4632
rect 3620 4126 3832 4154
rect 3608 4072 3660 4078
rect 3514 4040 3570 4049
rect 3608 4014 3660 4020
rect 3514 3975 3516 3984
rect 3568 3975 3570 3984
rect 3516 3946 3568 3952
rect 3528 3738 3556 3946
rect 3516 3732 3568 3738
rect 3516 3674 3568 3680
rect 3620 3641 3648 4014
rect 3804 3738 3832 4126
rect 3896 4078 3924 4644
rect 3884 4072 3936 4078
rect 3884 4014 3936 4020
rect 3896 3738 3924 4014
rect 4080 3942 4108 6870
rect 4252 6384 4304 6390
rect 4252 6326 4304 6332
rect 4264 5370 4292 6326
rect 4356 5914 4384 14855
rect 5000 14482 5028 17167
rect 5262 15600 5318 15609
rect 5262 15535 5318 15544
rect 5170 15056 5226 15065
rect 5170 14991 5226 15000
rect 4988 14476 5040 14482
rect 4988 14418 5040 14424
rect 4622 14172 4918 14192
rect 4678 14170 4702 14172
rect 4758 14170 4782 14172
rect 4838 14170 4862 14172
rect 4700 14118 4702 14170
rect 4764 14118 4776 14170
rect 4838 14118 4840 14170
rect 4678 14116 4702 14118
rect 4758 14116 4782 14118
rect 4838 14116 4862 14118
rect 4622 14096 4918 14116
rect 5000 14074 5028 14418
rect 5184 14074 5212 14991
rect 4988 14068 5040 14074
rect 4988 14010 5040 14016
rect 5172 14068 5224 14074
rect 5172 14010 5224 14016
rect 5080 13864 5132 13870
rect 5080 13806 5132 13812
rect 5092 13394 5120 13806
rect 5170 13424 5226 13433
rect 5080 13388 5132 13394
rect 5170 13359 5226 13368
rect 5080 13330 5132 13336
rect 4988 13184 5040 13190
rect 4988 13126 5040 13132
rect 4622 13084 4918 13104
rect 4678 13082 4702 13084
rect 4758 13082 4782 13084
rect 4838 13082 4862 13084
rect 4700 13030 4702 13082
rect 4764 13030 4776 13082
rect 4838 13030 4840 13082
rect 4678 13028 4702 13030
rect 4758 13028 4782 13030
rect 4838 13028 4862 13030
rect 4622 13008 4918 13028
rect 4620 12912 4672 12918
rect 5000 12889 5028 13126
rect 4620 12854 4672 12860
rect 4986 12880 5042 12889
rect 4632 12442 4660 12854
rect 4986 12815 5042 12824
rect 4988 12640 5040 12646
rect 4988 12582 5040 12588
rect 4620 12436 4672 12442
rect 4620 12378 4672 12384
rect 4622 11996 4918 12016
rect 4678 11994 4702 11996
rect 4758 11994 4782 11996
rect 4838 11994 4862 11996
rect 4700 11942 4702 11994
rect 4764 11942 4776 11994
rect 4838 11942 4840 11994
rect 4678 11940 4702 11942
rect 4758 11940 4782 11942
rect 4838 11940 4862 11942
rect 4622 11920 4918 11940
rect 5000 11880 5028 12582
rect 4908 11852 5028 11880
rect 4908 11540 4936 11852
rect 5184 11778 5212 13359
rect 5276 12306 5304 15535
rect 6274 15464 6330 15473
rect 5356 15428 5408 15434
rect 6274 15399 6330 15408
rect 5356 15370 5408 15376
rect 5368 13394 5396 15370
rect 6288 15162 6316 15399
rect 6276 15156 6328 15162
rect 6276 15098 6328 15104
rect 6288 14958 6316 15098
rect 6276 14952 6328 14958
rect 6276 14894 6328 14900
rect 6092 14816 6144 14822
rect 6092 14758 6144 14764
rect 5448 14476 5500 14482
rect 5448 14418 5500 14424
rect 5908 14476 5960 14482
rect 5908 14418 5960 14424
rect 5460 13870 5488 14418
rect 5632 14272 5684 14278
rect 5632 14214 5684 14220
rect 5644 13870 5672 14214
rect 5448 13864 5500 13870
rect 5632 13864 5684 13870
rect 5448 13806 5500 13812
rect 5630 13832 5632 13841
rect 5684 13832 5686 13841
rect 5540 13796 5592 13802
rect 5630 13767 5686 13776
rect 5540 13738 5592 13744
rect 5552 13530 5580 13738
rect 5540 13524 5592 13530
rect 5540 13466 5592 13472
rect 5724 13524 5776 13530
rect 5724 13466 5776 13472
rect 5356 13388 5408 13394
rect 5408 13348 5488 13376
rect 5356 13330 5408 13336
rect 5264 12300 5316 12306
rect 5264 12242 5316 12248
rect 5092 11750 5212 11778
rect 4988 11688 5040 11694
rect 5092 11676 5120 11750
rect 5040 11648 5120 11676
rect 4988 11630 5040 11636
rect 4908 11512 5028 11540
rect 4436 11280 4488 11286
rect 4436 11222 4488 11228
rect 4448 10606 4476 11222
rect 4528 11144 4580 11150
rect 4528 11086 4580 11092
rect 4436 10600 4488 10606
rect 4436 10542 4488 10548
rect 4540 10130 4568 11086
rect 4622 10908 4918 10928
rect 4678 10906 4702 10908
rect 4758 10906 4782 10908
rect 4838 10906 4862 10908
rect 4700 10854 4702 10906
rect 4764 10854 4776 10906
rect 4838 10854 4840 10906
rect 4678 10852 4702 10854
rect 4758 10852 4782 10854
rect 4838 10852 4862 10854
rect 4622 10832 4918 10852
rect 4528 10124 4580 10130
rect 4528 10066 4580 10072
rect 4436 9716 4488 9722
rect 4436 9658 4488 9664
rect 4448 7954 4476 9658
rect 4540 9178 4568 10066
rect 4622 9820 4918 9840
rect 4678 9818 4702 9820
rect 4758 9818 4782 9820
rect 4838 9818 4862 9820
rect 4700 9766 4702 9818
rect 4764 9766 4776 9818
rect 4838 9766 4840 9818
rect 4678 9764 4702 9766
rect 4758 9764 4782 9766
rect 4838 9764 4862 9766
rect 4622 9744 4918 9764
rect 4528 9172 4580 9178
rect 4528 9114 4580 9120
rect 4622 8732 4918 8752
rect 4678 8730 4702 8732
rect 4758 8730 4782 8732
rect 4838 8730 4862 8732
rect 4700 8678 4702 8730
rect 4764 8678 4776 8730
rect 4838 8678 4840 8730
rect 4678 8676 4702 8678
rect 4758 8676 4782 8678
rect 4838 8676 4862 8678
rect 4622 8656 4918 8676
rect 4436 7948 4488 7954
rect 4488 7908 4568 7936
rect 4436 7890 4488 7896
rect 4436 7744 4488 7750
rect 4436 7686 4488 7692
rect 4448 6662 4476 7686
rect 4540 7546 4568 7908
rect 4622 7644 4918 7664
rect 4678 7642 4702 7644
rect 4758 7642 4782 7644
rect 4838 7642 4862 7644
rect 4700 7590 4702 7642
rect 4764 7590 4776 7642
rect 4838 7590 4840 7642
rect 4678 7588 4702 7590
rect 4758 7588 4782 7590
rect 4838 7588 4862 7590
rect 4622 7568 4918 7588
rect 4528 7540 4580 7546
rect 4528 7482 4580 7488
rect 4540 7342 4568 7482
rect 5000 7426 5028 11512
rect 5092 11218 5120 11648
rect 5172 11688 5224 11694
rect 5276 11676 5304 12242
rect 5356 12232 5408 12238
rect 5356 12174 5408 12180
rect 5368 11762 5396 12174
rect 5356 11756 5408 11762
rect 5356 11698 5408 11704
rect 5224 11648 5304 11676
rect 5172 11630 5224 11636
rect 5184 11354 5212 11630
rect 5172 11348 5224 11354
rect 5172 11290 5224 11296
rect 5356 11348 5408 11354
rect 5356 11290 5408 11296
rect 5080 11212 5132 11218
rect 5080 11154 5132 11160
rect 5092 10810 5120 11154
rect 5080 10804 5132 10810
rect 5080 10746 5132 10752
rect 5264 9444 5316 9450
rect 5264 9386 5316 9392
rect 5080 9376 5132 9382
rect 5080 9318 5132 9324
rect 5092 9178 5120 9318
rect 5276 9178 5304 9386
rect 5080 9172 5132 9178
rect 5080 9114 5132 9120
rect 5264 9172 5316 9178
rect 5264 9114 5316 9120
rect 5080 9036 5132 9042
rect 5080 8978 5132 8984
rect 5092 7818 5120 8978
rect 5368 8922 5396 11290
rect 5460 11218 5488 13348
rect 5540 13184 5592 13190
rect 5540 13126 5592 13132
rect 5552 12782 5580 13126
rect 5540 12776 5592 12782
rect 5540 12718 5592 12724
rect 5552 12374 5580 12718
rect 5632 12708 5684 12714
rect 5632 12650 5684 12656
rect 5540 12368 5592 12374
rect 5540 12310 5592 12316
rect 5552 12102 5580 12310
rect 5540 12096 5592 12102
rect 5540 12038 5592 12044
rect 5552 11898 5580 12038
rect 5540 11892 5592 11898
rect 5540 11834 5592 11840
rect 5448 11212 5500 11218
rect 5448 11154 5500 11160
rect 5460 10810 5488 11154
rect 5448 10804 5500 10810
rect 5448 10746 5500 10752
rect 5644 10606 5672 12650
rect 5736 11694 5764 13466
rect 5920 13190 5948 14418
rect 6000 13728 6052 13734
rect 6000 13670 6052 13676
rect 6012 13326 6040 13670
rect 6000 13320 6052 13326
rect 6000 13262 6052 13268
rect 5908 13184 5960 13190
rect 5814 13152 5870 13161
rect 5908 13126 5960 13132
rect 5814 13087 5870 13096
rect 5724 11688 5776 11694
rect 5724 11630 5776 11636
rect 5828 11200 5856 13087
rect 6012 12442 6040 13262
rect 6104 12850 6132 14758
rect 6380 14618 6408 21542
rect 8220 21542 8538 21570
rect 8220 18426 8248 21542
rect 8482 21520 8538 21542
rect 10888 21542 11022 21570
rect 8289 19068 8585 19088
rect 8345 19066 8369 19068
rect 8425 19066 8449 19068
rect 8505 19066 8529 19068
rect 8367 19014 8369 19066
rect 8431 19014 8443 19066
rect 8505 19014 8507 19066
rect 8345 19012 8369 19014
rect 8425 19012 8449 19014
rect 8505 19012 8529 19014
rect 8289 18992 8585 19012
rect 8208 18420 8260 18426
rect 8208 18362 8260 18368
rect 10888 18358 10916 21542
rect 10966 21520 11022 21542
rect 13358 21570 13414 22000
rect 15842 21570 15898 22000
rect 18234 21570 18290 22000
rect 20718 21570 20774 22000
rect 13358 21542 13584 21570
rect 13358 21520 13414 21542
rect 11956 19612 12252 19632
rect 12012 19610 12036 19612
rect 12092 19610 12116 19612
rect 12172 19610 12196 19612
rect 12034 19558 12036 19610
rect 12098 19558 12110 19610
rect 12172 19558 12174 19610
rect 12012 19556 12036 19558
rect 12092 19556 12116 19558
rect 12172 19556 12196 19558
rect 11956 19536 12252 19556
rect 11888 18828 11940 18834
rect 11888 18770 11940 18776
rect 13452 18828 13504 18834
rect 13452 18770 13504 18776
rect 7380 18352 7432 18358
rect 7380 18294 7432 18300
rect 10876 18352 10928 18358
rect 10876 18294 10928 18300
rect 7010 17776 7066 17785
rect 7010 17711 7066 17720
rect 6920 15360 6972 15366
rect 6920 15302 6972 15308
rect 6932 14958 6960 15302
rect 6828 14952 6880 14958
rect 6828 14894 6880 14900
rect 6920 14952 6972 14958
rect 6920 14894 6972 14900
rect 6368 14612 6420 14618
rect 6368 14554 6420 14560
rect 6840 14346 6868 14894
rect 6932 14550 6960 14894
rect 6920 14544 6972 14550
rect 6920 14486 6972 14492
rect 6736 14340 6788 14346
rect 6736 14282 6788 14288
rect 6828 14340 6880 14346
rect 6828 14282 6880 14288
rect 6274 13696 6330 13705
rect 6274 13631 6330 13640
rect 6288 13394 6316 13631
rect 6552 13456 6604 13462
rect 6552 13398 6604 13404
rect 6276 13388 6328 13394
rect 6276 13330 6328 13336
rect 6276 13184 6328 13190
rect 6276 13126 6328 13132
rect 6092 12844 6144 12850
rect 6092 12786 6144 12792
rect 6184 12776 6236 12782
rect 6184 12718 6236 12724
rect 6000 12436 6052 12442
rect 6000 12378 6052 12384
rect 6196 12238 6224 12718
rect 6184 12232 6236 12238
rect 6184 12174 6236 12180
rect 6092 11552 6144 11558
rect 6092 11494 6144 11500
rect 5828 11172 5948 11200
rect 5816 11076 5868 11082
rect 5816 11018 5868 11024
rect 5448 10600 5500 10606
rect 5448 10542 5500 10548
rect 5632 10600 5684 10606
rect 5632 10542 5684 10548
rect 5460 10266 5488 10542
rect 5632 10464 5684 10470
rect 5632 10406 5684 10412
rect 5448 10260 5500 10266
rect 5448 10202 5500 10208
rect 5460 9081 5488 10202
rect 5446 9072 5502 9081
rect 5644 9042 5672 10406
rect 5724 10192 5776 10198
rect 5724 10134 5776 10140
rect 5736 10033 5764 10134
rect 5722 10024 5778 10033
rect 5828 9994 5856 11018
rect 5722 9959 5778 9968
rect 5816 9988 5868 9994
rect 5816 9930 5868 9936
rect 5920 9722 5948 11172
rect 6104 10849 6132 11494
rect 6196 11354 6224 12174
rect 6184 11348 6236 11354
rect 6184 11290 6236 11296
rect 6184 11212 6236 11218
rect 6184 11154 6236 11160
rect 6090 10840 6146 10849
rect 6090 10775 6146 10784
rect 6196 10470 6224 11154
rect 6184 10464 6236 10470
rect 6184 10406 6236 10412
rect 6092 10192 6144 10198
rect 6092 10134 6144 10140
rect 6000 10056 6052 10062
rect 6000 9998 6052 10004
rect 5908 9716 5960 9722
rect 5908 9658 5960 9664
rect 5446 9007 5502 9016
rect 5632 9036 5684 9042
rect 5632 8978 5684 8984
rect 5276 8894 5396 8922
rect 5448 8968 5500 8974
rect 5448 8910 5500 8916
rect 5172 8560 5224 8566
rect 5172 8502 5224 8508
rect 5184 8362 5212 8502
rect 5172 8356 5224 8362
rect 5172 8298 5224 8304
rect 5080 7812 5132 7818
rect 5080 7754 5132 7760
rect 5000 7398 5120 7426
rect 4528 7336 4580 7342
rect 4528 7278 4580 7284
rect 4988 7336 5040 7342
rect 4988 7278 5040 7284
rect 4620 7200 4672 7206
rect 4620 7142 4672 7148
rect 4436 6656 4488 6662
rect 4632 6644 4660 7142
rect 4436 6598 4488 6604
rect 4540 6616 4660 6644
rect 4344 5908 4396 5914
rect 4344 5850 4396 5856
rect 4344 5772 4396 5778
rect 4448 5760 4476 6598
rect 4540 6100 4568 6616
rect 4622 6556 4918 6576
rect 4678 6554 4702 6556
rect 4758 6554 4782 6556
rect 4838 6554 4862 6556
rect 4700 6502 4702 6554
rect 4764 6502 4776 6554
rect 4838 6502 4840 6554
rect 4678 6500 4702 6502
rect 4758 6500 4782 6502
rect 4838 6500 4862 6502
rect 4622 6480 4918 6500
rect 4620 6112 4672 6118
rect 4540 6072 4620 6100
rect 4620 6054 4672 6060
rect 4396 5732 4476 5760
rect 4344 5714 4396 5720
rect 4252 5364 4304 5370
rect 4252 5306 4304 5312
rect 4160 5228 4212 5234
rect 4160 5170 4212 5176
rect 4172 4078 4200 5170
rect 4356 5098 4384 5714
rect 4526 5672 4582 5681
rect 4436 5636 4488 5642
rect 4526 5607 4582 5616
rect 4436 5578 4488 5584
rect 4448 5137 4476 5578
rect 4540 5166 4568 5607
rect 4622 5468 4918 5488
rect 4678 5466 4702 5468
rect 4758 5466 4782 5468
rect 4838 5466 4862 5468
rect 4700 5414 4702 5466
rect 4764 5414 4776 5466
rect 4838 5414 4840 5466
rect 4678 5412 4702 5414
rect 4758 5412 4782 5414
rect 4838 5412 4862 5414
rect 4622 5392 4918 5412
rect 4528 5160 4580 5166
rect 4434 5128 4490 5137
rect 4344 5092 4396 5098
rect 4528 5102 4580 5108
rect 4434 5063 4490 5072
rect 4344 5034 4396 5040
rect 4160 4072 4212 4078
rect 4160 4014 4212 4020
rect 4068 3936 4120 3942
rect 4068 3878 4120 3884
rect 3792 3732 3844 3738
rect 3792 3674 3844 3680
rect 3884 3732 3936 3738
rect 3884 3674 3936 3680
rect 3606 3632 3662 3641
rect 3424 3596 3476 3602
rect 3606 3567 3662 3576
rect 3424 3538 3476 3544
rect 3436 3194 3464 3538
rect 3424 3188 3476 3194
rect 3424 3130 3476 3136
rect 3804 2990 3832 3674
rect 3792 2984 3844 2990
rect 3148 2926 3200 2932
rect 3330 2952 3386 2961
rect 3160 2650 3188 2926
rect 3792 2926 3844 2932
rect 3330 2887 3386 2896
rect 3804 2650 3832 2926
rect 3896 2922 3924 3674
rect 3884 2916 3936 2922
rect 3884 2858 3936 2864
rect 1860 2644 1912 2650
rect 1860 2586 1912 2592
rect 3148 2644 3200 2650
rect 3148 2586 3200 2592
rect 3792 2644 3844 2650
rect 3792 2586 3844 2592
rect 3056 2508 3108 2514
rect 3160 2496 3188 2586
rect 4080 2514 4108 3878
rect 4172 2990 4200 4014
rect 4356 3505 4384 5034
rect 4448 4690 4476 5063
rect 4540 4826 4568 5102
rect 4528 4820 4580 4826
rect 4528 4762 4580 4768
rect 4436 4684 4488 4690
rect 4436 4626 4488 4632
rect 4622 4380 4918 4400
rect 4678 4378 4702 4380
rect 4758 4378 4782 4380
rect 4838 4378 4862 4380
rect 4700 4326 4702 4378
rect 4764 4326 4776 4378
rect 4838 4326 4840 4378
rect 4678 4324 4702 4326
rect 4758 4324 4782 4326
rect 4838 4324 4862 4326
rect 4622 4304 4918 4324
rect 5000 4214 5028 7278
rect 5092 6225 5120 7398
rect 5276 6866 5304 8894
rect 5356 8832 5408 8838
rect 5356 8774 5408 8780
rect 5368 8294 5396 8774
rect 5460 8634 5488 8910
rect 5448 8628 5500 8634
rect 5448 8570 5500 8576
rect 5356 8288 5408 8294
rect 5356 8230 5408 8236
rect 5460 7449 5488 8570
rect 5644 8294 5672 8978
rect 6012 8838 6040 9998
rect 6104 9722 6132 10134
rect 6092 9716 6144 9722
rect 6092 9658 6144 9664
rect 6104 9042 6132 9658
rect 6092 9036 6144 9042
rect 6092 8978 6144 8984
rect 6000 8832 6052 8838
rect 6000 8774 6052 8780
rect 6288 8634 6316 13126
rect 6366 12744 6422 12753
rect 6366 12679 6422 12688
rect 6380 12646 6408 12679
rect 6564 12646 6592 13398
rect 6368 12640 6420 12646
rect 6368 12582 6420 12588
rect 6552 12640 6604 12646
rect 6552 12582 6604 12588
rect 6460 12368 6512 12374
rect 6460 12310 6512 12316
rect 6472 11558 6500 12310
rect 6460 11552 6512 11558
rect 6460 11494 6512 11500
rect 6460 11144 6512 11150
rect 6460 11086 6512 11092
rect 6472 10577 6500 11086
rect 6458 10568 6514 10577
rect 6458 10503 6514 10512
rect 6644 9716 6696 9722
rect 6644 9658 6696 9664
rect 6368 9444 6420 9450
rect 6368 9386 6420 9392
rect 6380 9178 6408 9386
rect 6552 9376 6604 9382
rect 6472 9336 6552 9364
rect 6368 9172 6420 9178
rect 6368 9114 6420 9120
rect 6276 8628 6328 8634
rect 6276 8570 6328 8576
rect 6472 8566 6500 9336
rect 6552 9318 6604 9324
rect 6656 8974 6684 9658
rect 6644 8968 6696 8974
rect 6644 8910 6696 8916
rect 6460 8560 6512 8566
rect 6460 8502 6512 8508
rect 5540 8288 5592 8294
rect 5540 8230 5592 8236
rect 5632 8288 5684 8294
rect 5632 8230 5684 8236
rect 5552 8090 5580 8230
rect 5540 8084 5592 8090
rect 5540 8026 5592 8032
rect 5540 7472 5592 7478
rect 5446 7440 5502 7449
rect 5540 7414 5592 7420
rect 5446 7375 5502 7384
rect 5264 6860 5316 6866
rect 5264 6802 5316 6808
rect 5172 6656 5224 6662
rect 5172 6598 5224 6604
rect 5078 6216 5134 6225
rect 5078 6151 5134 6160
rect 4988 4208 5040 4214
rect 4988 4150 5040 4156
rect 5000 4078 5028 4150
rect 4436 4072 4488 4078
rect 4436 4014 4488 4020
rect 4988 4072 5040 4078
rect 4988 4014 5040 4020
rect 4342 3496 4398 3505
rect 4342 3431 4398 3440
rect 4160 2984 4212 2990
rect 4160 2926 4212 2932
rect 4172 2650 4200 2926
rect 4344 2916 4396 2922
rect 4344 2858 4396 2864
rect 4160 2644 4212 2650
rect 4160 2586 4212 2592
rect 3108 2468 3188 2496
rect 4068 2508 4120 2514
rect 3056 2450 3108 2456
rect 4068 2450 4120 2456
rect 3976 2372 4028 2378
rect 3976 2314 4028 2320
rect 3148 2100 3200 2106
rect 3148 2042 3200 2048
rect 1766 1456 1822 1465
rect 1766 1391 1822 1400
rect 938 128 994 480
rect 938 76 940 128
rect 992 76 994 128
rect 938 0 994 76
rect 2870 82 2926 480
rect 3160 82 3188 2042
rect 3988 134 4016 2314
rect 4356 1873 4384 2858
rect 4448 2553 4476 4014
rect 5000 3738 5028 4014
rect 4988 3732 5040 3738
rect 4988 3674 5040 3680
rect 4528 3664 4580 3670
rect 4528 3606 4580 3612
rect 4540 2922 4568 3606
rect 4622 3292 4918 3312
rect 4678 3290 4702 3292
rect 4758 3290 4782 3292
rect 4838 3290 4862 3292
rect 4700 3238 4702 3290
rect 4764 3238 4776 3290
rect 4838 3238 4840 3290
rect 4678 3236 4702 3238
rect 4758 3236 4782 3238
rect 4838 3236 4862 3238
rect 4622 3216 4918 3236
rect 5000 2990 5028 3674
rect 4988 2984 5040 2990
rect 4988 2926 5040 2932
rect 4528 2916 4580 2922
rect 4528 2858 4580 2864
rect 4434 2544 4490 2553
rect 4434 2479 4490 2488
rect 4622 2204 4918 2224
rect 4678 2202 4702 2204
rect 4758 2202 4782 2204
rect 4838 2202 4862 2204
rect 4700 2150 4702 2202
rect 4764 2150 4776 2202
rect 4838 2150 4840 2202
rect 4678 2148 4702 2150
rect 4758 2148 4782 2150
rect 4838 2148 4862 2150
rect 4622 2128 4918 2148
rect 4342 1864 4398 1873
rect 4342 1799 4398 1808
rect 2870 54 3188 82
rect 3976 128 4028 134
rect 3976 70 4028 76
rect 4894 82 4950 480
rect 5092 82 5120 6151
rect 5184 5574 5212 6598
rect 5276 5914 5304 6802
rect 5448 6112 5500 6118
rect 5448 6054 5500 6060
rect 5264 5908 5316 5914
rect 5264 5850 5316 5856
rect 5172 5568 5224 5574
rect 5172 5510 5224 5516
rect 5184 5166 5212 5510
rect 5172 5160 5224 5166
rect 5172 5102 5224 5108
rect 5172 4684 5224 4690
rect 5276 4672 5304 5850
rect 5356 5228 5408 5234
rect 5356 5170 5408 5176
rect 5368 4690 5396 5170
rect 5460 5166 5488 6054
rect 5552 5234 5580 7414
rect 5644 7342 5672 8230
rect 5814 7848 5870 7857
rect 5814 7783 5870 7792
rect 5828 7750 5856 7783
rect 5816 7744 5868 7750
rect 5816 7686 5868 7692
rect 5632 7336 5684 7342
rect 5632 7278 5684 7284
rect 5644 7206 5672 7278
rect 6472 7206 6500 8502
rect 5632 7200 5684 7206
rect 5632 7142 5684 7148
rect 6460 7200 6512 7206
rect 6460 7142 6512 7148
rect 5644 6866 5672 7142
rect 6472 6934 6500 7142
rect 6460 6928 6512 6934
rect 6460 6870 6512 6876
rect 5632 6860 5684 6866
rect 5632 6802 5684 6808
rect 5644 6769 5672 6802
rect 5630 6760 5686 6769
rect 5630 6695 5686 6704
rect 6276 6452 6328 6458
rect 6276 6394 6328 6400
rect 6182 6352 6238 6361
rect 6182 6287 6238 6296
rect 6196 6254 6224 6287
rect 6184 6248 6236 6254
rect 6184 6190 6236 6196
rect 5908 5772 5960 5778
rect 5908 5714 5960 5720
rect 5920 5302 5948 5714
rect 6184 5636 6236 5642
rect 6184 5578 6236 5584
rect 5908 5296 5960 5302
rect 5908 5238 5960 5244
rect 5540 5228 5592 5234
rect 5540 5170 5592 5176
rect 5448 5160 5500 5166
rect 5448 5102 5500 5108
rect 6196 4826 6224 5578
rect 6288 5574 6316 6394
rect 6368 6180 6420 6186
rect 6368 6122 6420 6128
rect 6380 5710 6408 6122
rect 6472 6118 6500 6870
rect 6550 6760 6606 6769
rect 6550 6695 6606 6704
rect 6460 6112 6512 6118
rect 6460 6054 6512 6060
rect 6564 5914 6592 6695
rect 6748 6458 6776 14282
rect 6920 13864 6972 13870
rect 6840 13824 6920 13852
rect 6840 13705 6868 13824
rect 6920 13806 6972 13812
rect 6826 13696 6882 13705
rect 6826 13631 6882 13640
rect 6840 13462 6868 13631
rect 6828 13456 6880 13462
rect 6828 13398 6880 13404
rect 6828 9920 6880 9926
rect 6828 9862 6880 9868
rect 6840 9586 6868 9862
rect 6828 9580 6880 9586
rect 6828 9522 6880 9528
rect 6920 9580 6972 9586
rect 6920 9522 6972 9528
rect 6932 9110 6960 9522
rect 6920 9104 6972 9110
rect 6920 9046 6972 9052
rect 7024 7392 7052 17711
rect 7392 16046 7420 18294
rect 10600 18216 10652 18222
rect 10600 18158 10652 18164
rect 9588 18148 9640 18154
rect 9588 18090 9640 18096
rect 9312 18080 9364 18086
rect 9312 18022 9364 18028
rect 8289 17980 8585 18000
rect 8345 17978 8369 17980
rect 8425 17978 8449 17980
rect 8505 17978 8529 17980
rect 8367 17926 8369 17978
rect 8431 17926 8443 17978
rect 8505 17926 8507 17978
rect 8345 17924 8369 17926
rect 8425 17924 8449 17926
rect 8505 17924 8529 17926
rect 8289 17904 8585 17924
rect 8668 16992 8720 16998
rect 8668 16934 8720 16940
rect 8289 16892 8585 16912
rect 8345 16890 8369 16892
rect 8425 16890 8449 16892
rect 8505 16890 8529 16892
rect 8367 16838 8369 16890
rect 8431 16838 8443 16890
rect 8505 16838 8507 16890
rect 8345 16836 8369 16838
rect 8425 16836 8449 16838
rect 8505 16836 8529 16838
rect 8289 16816 8585 16836
rect 8484 16652 8536 16658
rect 8484 16594 8536 16600
rect 8116 16448 8168 16454
rect 8116 16390 8168 16396
rect 7380 16040 7432 16046
rect 7380 15982 7432 15988
rect 8128 15978 8156 16390
rect 8496 15978 8524 16594
rect 8680 15978 8708 16934
rect 9036 16720 9088 16726
rect 9036 16662 9088 16668
rect 8760 16584 8812 16590
rect 8760 16526 8812 16532
rect 7472 15972 7524 15978
rect 7472 15914 7524 15920
rect 8024 15972 8076 15978
rect 8024 15914 8076 15920
rect 8116 15972 8168 15978
rect 8116 15914 8168 15920
rect 8484 15972 8536 15978
rect 8484 15914 8536 15920
rect 8668 15972 8720 15978
rect 8668 15914 8720 15920
rect 7196 14000 7248 14006
rect 7196 13942 7248 13948
rect 7208 13734 7236 13942
rect 7196 13728 7248 13734
rect 7196 13670 7248 13676
rect 7380 12844 7432 12850
rect 7380 12786 7432 12792
rect 7392 12442 7420 12786
rect 7380 12436 7432 12442
rect 7380 12378 7432 12384
rect 7484 12102 7512 15914
rect 7748 15904 7800 15910
rect 7748 15846 7800 15852
rect 7564 15496 7616 15502
rect 7564 15438 7616 15444
rect 7576 15026 7604 15438
rect 7564 15020 7616 15026
rect 7564 14962 7616 14968
rect 7760 14006 7788 15846
rect 8036 15706 8064 15914
rect 8128 15706 8156 15914
rect 8289 15804 8585 15824
rect 8345 15802 8369 15804
rect 8425 15802 8449 15804
rect 8505 15802 8529 15804
rect 8367 15750 8369 15802
rect 8431 15750 8443 15802
rect 8505 15750 8507 15802
rect 8345 15748 8369 15750
rect 8425 15748 8449 15750
rect 8505 15748 8529 15750
rect 8289 15728 8585 15748
rect 8024 15700 8076 15706
rect 8024 15642 8076 15648
rect 8116 15700 8168 15706
rect 8116 15642 8168 15648
rect 7932 15632 7984 15638
rect 7932 15574 7984 15580
rect 7944 15162 7972 15574
rect 7932 15156 7984 15162
rect 7932 15098 7984 15104
rect 7944 14550 7972 15098
rect 8289 14716 8585 14736
rect 8345 14714 8369 14716
rect 8425 14714 8449 14716
rect 8505 14714 8529 14716
rect 8367 14662 8369 14714
rect 8431 14662 8443 14714
rect 8505 14662 8507 14714
rect 8345 14660 8369 14662
rect 8425 14660 8449 14662
rect 8505 14660 8529 14662
rect 8289 14640 8585 14660
rect 7932 14544 7984 14550
rect 7932 14486 7984 14492
rect 8024 14408 8076 14414
rect 8024 14350 8076 14356
rect 7840 14272 7892 14278
rect 7840 14214 7892 14220
rect 7748 14000 7800 14006
rect 7748 13942 7800 13948
rect 7656 13728 7708 13734
rect 7656 13670 7708 13676
rect 7564 13320 7616 13326
rect 7564 13262 7616 13268
rect 7576 12850 7604 13262
rect 7564 12844 7616 12850
rect 7564 12786 7616 12792
rect 7668 12646 7696 13670
rect 7852 13462 7880 14214
rect 8036 14074 8064 14350
rect 8024 14068 8076 14074
rect 8024 14010 8076 14016
rect 8289 13628 8585 13648
rect 8345 13626 8369 13628
rect 8425 13626 8449 13628
rect 8505 13626 8529 13628
rect 8367 13574 8369 13626
rect 8431 13574 8443 13626
rect 8505 13574 8507 13626
rect 8345 13572 8369 13574
rect 8425 13572 8449 13574
rect 8505 13572 8529 13574
rect 8289 13552 8585 13572
rect 7840 13456 7892 13462
rect 7840 13398 7892 13404
rect 7748 13184 7800 13190
rect 7748 13126 7800 13132
rect 7760 12714 7788 13126
rect 7748 12708 7800 12714
rect 7748 12650 7800 12656
rect 7656 12640 7708 12646
rect 7656 12582 7708 12588
rect 7852 12442 7880 13398
rect 8680 13326 8708 15914
rect 8772 15570 8800 16526
rect 9048 16017 9076 16662
rect 9034 16008 9090 16017
rect 9034 15943 9090 15952
rect 9048 15910 9076 15943
rect 9036 15904 9088 15910
rect 9036 15846 9088 15852
rect 8760 15564 8812 15570
rect 8760 15506 8812 15512
rect 8944 15360 8996 15366
rect 8944 15302 8996 15308
rect 8956 14822 8984 15302
rect 8944 14816 8996 14822
rect 8944 14758 8996 14764
rect 9048 14482 9076 15846
rect 9324 15026 9352 18022
rect 9496 17128 9548 17134
rect 9496 17070 9548 17076
rect 9508 16454 9536 17070
rect 9496 16448 9548 16454
rect 9496 16390 9548 16396
rect 9312 15020 9364 15026
rect 9312 14962 9364 14968
rect 9220 14884 9272 14890
rect 9220 14826 9272 14832
rect 9036 14476 9088 14482
rect 9036 14418 9088 14424
rect 9232 14414 9260 14826
rect 9324 14618 9352 14962
rect 9312 14612 9364 14618
rect 9312 14554 9364 14560
rect 9220 14408 9272 14414
rect 9220 14350 9272 14356
rect 8760 14272 8812 14278
rect 8760 14214 8812 14220
rect 8772 13938 8800 14214
rect 8760 13932 8812 13938
rect 8760 13874 8812 13880
rect 9508 13841 9536 16390
rect 9600 16046 9628 18090
rect 10612 17678 10640 18158
rect 10692 17740 10744 17746
rect 10692 17682 10744 17688
rect 10600 17672 10652 17678
rect 10600 17614 10652 17620
rect 10612 17066 10640 17614
rect 10140 17060 10192 17066
rect 10140 17002 10192 17008
rect 10600 17060 10652 17066
rect 10600 17002 10652 17008
rect 9864 16992 9916 16998
rect 9864 16934 9916 16940
rect 9876 16658 9904 16934
rect 9680 16652 9732 16658
rect 9680 16594 9732 16600
rect 9864 16652 9916 16658
rect 9864 16594 9916 16600
rect 9692 16182 9720 16594
rect 9680 16176 9732 16182
rect 9680 16118 9732 16124
rect 9588 16040 9640 16046
rect 9588 15982 9640 15988
rect 9600 13938 9628 15982
rect 9692 15434 9720 16118
rect 9876 15978 9904 16594
rect 9864 15972 9916 15978
rect 9864 15914 9916 15920
rect 9956 15904 10008 15910
rect 9956 15846 10008 15852
rect 9864 15564 9916 15570
rect 9864 15506 9916 15512
rect 9680 15428 9732 15434
rect 9680 15370 9732 15376
rect 9876 14618 9904 15506
rect 9864 14612 9916 14618
rect 9864 14554 9916 14560
rect 9864 14340 9916 14346
rect 9864 14282 9916 14288
rect 9588 13932 9640 13938
rect 9588 13874 9640 13880
rect 9680 13864 9732 13870
rect 9494 13832 9550 13841
rect 9680 13806 9732 13812
rect 9494 13767 9550 13776
rect 8668 13320 8720 13326
rect 8668 13262 8720 13268
rect 8680 12850 8708 13262
rect 8668 12844 8720 12850
rect 8668 12786 8720 12792
rect 9692 12714 9720 13806
rect 9876 13161 9904 14282
rect 9968 13326 9996 15846
rect 10152 15026 10180 17002
rect 10508 16584 10560 16590
rect 10508 16526 10560 16532
rect 10232 15972 10284 15978
rect 10232 15914 10284 15920
rect 10244 15638 10272 15914
rect 10232 15632 10284 15638
rect 10232 15574 10284 15580
rect 10244 15162 10272 15574
rect 10232 15156 10284 15162
rect 10232 15098 10284 15104
rect 10140 15020 10192 15026
rect 10140 14962 10192 14968
rect 10244 14890 10272 15098
rect 10232 14884 10284 14890
rect 10232 14826 10284 14832
rect 10244 14618 10272 14826
rect 10232 14612 10284 14618
rect 10232 14554 10284 14560
rect 10324 14476 10376 14482
rect 10324 14418 10376 14424
rect 10232 14000 10284 14006
rect 10232 13942 10284 13948
rect 10140 13932 10192 13938
rect 10140 13874 10192 13880
rect 10046 13832 10102 13841
rect 10046 13767 10102 13776
rect 9956 13320 10008 13326
rect 9956 13262 10008 13268
rect 9862 13152 9918 13161
rect 9862 13087 9918 13096
rect 9772 12980 9824 12986
rect 9772 12922 9824 12928
rect 8208 12708 8260 12714
rect 8208 12650 8260 12656
rect 8852 12708 8904 12714
rect 8852 12650 8904 12656
rect 9680 12708 9732 12714
rect 9680 12650 9732 12656
rect 7840 12436 7892 12442
rect 7840 12378 7892 12384
rect 8220 12238 8248 12650
rect 8289 12540 8585 12560
rect 8345 12538 8369 12540
rect 8425 12538 8449 12540
rect 8505 12538 8529 12540
rect 8367 12486 8369 12538
rect 8431 12486 8443 12538
rect 8505 12486 8507 12538
rect 8345 12484 8369 12486
rect 8425 12484 8449 12486
rect 8505 12484 8529 12486
rect 8289 12464 8585 12484
rect 8864 12442 8892 12650
rect 8852 12436 8904 12442
rect 8852 12378 8904 12384
rect 8208 12232 8260 12238
rect 8208 12174 8260 12180
rect 7196 12096 7248 12102
rect 7196 12038 7248 12044
rect 7472 12096 7524 12102
rect 7472 12038 7524 12044
rect 7104 11756 7156 11762
rect 7104 11698 7156 11704
rect 7116 11354 7144 11698
rect 7104 11348 7156 11354
rect 7104 11290 7156 11296
rect 7102 10840 7158 10849
rect 7102 10775 7158 10784
rect 7116 7954 7144 10775
rect 7208 8838 7236 12038
rect 8024 11892 8076 11898
rect 8024 11834 8076 11840
rect 7472 11552 7524 11558
rect 7472 11494 7524 11500
rect 7378 11384 7434 11393
rect 7378 11319 7434 11328
rect 7392 11150 7420 11319
rect 7484 11286 7512 11494
rect 7472 11280 7524 11286
rect 7472 11222 7524 11228
rect 7380 11144 7432 11150
rect 7380 11086 7432 11092
rect 7392 10266 7420 11086
rect 7484 10538 7512 11222
rect 7564 10600 7616 10606
rect 7564 10542 7616 10548
rect 7472 10532 7524 10538
rect 7472 10474 7524 10480
rect 7576 10266 7604 10542
rect 8036 10538 8064 11834
rect 8116 11756 8168 11762
rect 8116 11698 8168 11704
rect 8128 10713 8156 11698
rect 8220 11286 8248 12174
rect 8668 12164 8720 12170
rect 8668 12106 8720 12112
rect 8289 11452 8585 11472
rect 8345 11450 8369 11452
rect 8425 11450 8449 11452
rect 8505 11450 8529 11452
rect 8367 11398 8369 11450
rect 8431 11398 8443 11450
rect 8505 11398 8507 11450
rect 8345 11396 8369 11398
rect 8425 11396 8449 11398
rect 8505 11396 8529 11398
rect 8289 11376 8585 11396
rect 8680 11286 8708 12106
rect 8208 11280 8260 11286
rect 8208 11222 8260 11228
rect 8668 11280 8720 11286
rect 8668 11222 8720 11228
rect 8392 11008 8444 11014
rect 8392 10950 8444 10956
rect 8404 10810 8432 10950
rect 8392 10804 8444 10810
rect 8392 10746 8444 10752
rect 8114 10704 8170 10713
rect 8114 10639 8170 10648
rect 8758 10704 8814 10713
rect 8864 10674 8892 12378
rect 9036 12368 9088 12374
rect 9036 12310 9088 12316
rect 9048 11898 9076 12310
rect 9784 12238 9812 12922
rect 9772 12232 9824 12238
rect 9772 12174 9824 12180
rect 9128 12096 9180 12102
rect 9128 12038 9180 12044
rect 9036 11892 9088 11898
rect 9036 11834 9088 11840
rect 8758 10639 8814 10648
rect 8852 10668 8904 10674
rect 8024 10532 8076 10538
rect 8024 10474 8076 10480
rect 8289 10364 8585 10384
rect 8345 10362 8369 10364
rect 8425 10362 8449 10364
rect 8505 10362 8529 10364
rect 8367 10310 8369 10362
rect 8431 10310 8443 10362
rect 8505 10310 8507 10362
rect 8345 10308 8369 10310
rect 8425 10308 8449 10310
rect 8505 10308 8529 10310
rect 8289 10288 8585 10308
rect 7380 10260 7432 10266
rect 7380 10202 7432 10208
rect 7564 10260 7616 10266
rect 7564 10202 7616 10208
rect 7656 10192 7708 10198
rect 7562 10160 7618 10169
rect 7656 10134 7708 10140
rect 7562 10095 7618 10104
rect 7576 10062 7604 10095
rect 7564 10056 7616 10062
rect 7564 9998 7616 10004
rect 7576 9110 7604 9998
rect 7668 9518 7696 10134
rect 8668 9920 8720 9926
rect 8668 9862 8720 9868
rect 8680 9586 8708 9862
rect 8668 9580 8720 9586
rect 8668 9522 8720 9528
rect 7656 9512 7708 9518
rect 7656 9454 7708 9460
rect 8208 9376 8260 9382
rect 8114 9344 8170 9353
rect 8208 9318 8260 9324
rect 8114 9279 8170 9288
rect 7748 9172 7800 9178
rect 7748 9114 7800 9120
rect 7472 9104 7524 9110
rect 7472 9046 7524 9052
rect 7564 9104 7616 9110
rect 7564 9046 7616 9052
rect 7380 8900 7432 8906
rect 7380 8842 7432 8848
rect 7196 8832 7248 8838
rect 7196 8774 7248 8780
rect 7392 8634 7420 8842
rect 7484 8634 7512 9046
rect 7380 8628 7432 8634
rect 7380 8570 7432 8576
rect 7472 8628 7524 8634
rect 7472 8570 7524 8576
rect 7760 8498 7788 9114
rect 8128 8974 8156 9279
rect 8220 9042 8248 9318
rect 8289 9276 8585 9296
rect 8345 9274 8369 9276
rect 8425 9274 8449 9276
rect 8505 9274 8529 9276
rect 8367 9222 8369 9274
rect 8431 9222 8443 9274
rect 8505 9222 8507 9274
rect 8345 9220 8369 9222
rect 8425 9220 8449 9222
rect 8505 9220 8529 9222
rect 8289 9200 8585 9220
rect 8772 9110 8800 10639
rect 8852 10610 8904 10616
rect 8852 9988 8904 9994
rect 8852 9930 8904 9936
rect 8760 9104 8812 9110
rect 8760 9046 8812 9052
rect 8208 9036 8260 9042
rect 8208 8978 8260 8984
rect 8668 9036 8720 9042
rect 8668 8978 8720 8984
rect 8116 8968 8168 8974
rect 8116 8910 8168 8916
rect 7748 8492 7800 8498
rect 7748 8434 7800 8440
rect 7932 8492 7984 8498
rect 7932 8434 7984 8440
rect 7654 8120 7710 8129
rect 7654 8055 7710 8064
rect 7668 7954 7696 8055
rect 7104 7948 7156 7954
rect 7104 7890 7156 7896
rect 7656 7948 7708 7954
rect 7656 7890 7708 7896
rect 7116 7546 7144 7890
rect 7760 7818 7788 8434
rect 7944 8022 7972 8434
rect 8024 8356 8076 8362
rect 8024 8298 8076 8304
rect 7932 8016 7984 8022
rect 7932 7958 7984 7964
rect 7932 7880 7984 7886
rect 7932 7822 7984 7828
rect 7748 7812 7800 7818
rect 7748 7754 7800 7760
rect 7288 7744 7340 7750
rect 7288 7686 7340 7692
rect 7104 7540 7156 7546
rect 7104 7482 7156 7488
rect 7300 7410 7328 7686
rect 6840 7364 7052 7392
rect 7288 7404 7340 7410
rect 6736 6452 6788 6458
rect 6736 6394 6788 6400
rect 6552 5908 6604 5914
rect 6552 5850 6604 5856
rect 6368 5704 6420 5710
rect 6368 5646 6420 5652
rect 6276 5568 6328 5574
rect 6276 5510 6328 5516
rect 6288 4826 6316 5510
rect 6380 5234 6408 5646
rect 6368 5228 6420 5234
rect 6368 5170 6420 5176
rect 6184 4820 6236 4826
rect 6184 4762 6236 4768
rect 6276 4820 6328 4826
rect 6276 4762 6328 4768
rect 5224 4644 5304 4672
rect 5172 4626 5224 4632
rect 5276 3670 5304 4644
rect 5356 4684 5408 4690
rect 5356 4626 5408 4632
rect 6288 4593 6316 4762
rect 6368 4752 6420 4758
rect 6420 4712 6500 4740
rect 6368 4694 6420 4700
rect 6274 4584 6330 4593
rect 6274 4519 6330 4528
rect 6288 4154 6316 4519
rect 6288 4126 6408 4154
rect 6184 4072 6236 4078
rect 6184 4014 6236 4020
rect 6196 3738 6224 4014
rect 6184 3732 6236 3738
rect 6184 3674 6236 3680
rect 5264 3664 5316 3670
rect 5264 3606 5316 3612
rect 5540 3596 5592 3602
rect 5540 3538 5592 3544
rect 5552 3398 5580 3538
rect 5540 3392 5592 3398
rect 5540 3334 5592 3340
rect 5552 3194 5580 3334
rect 6196 3194 6224 3674
rect 5540 3188 5592 3194
rect 5540 3130 5592 3136
rect 6184 3188 6236 3194
rect 6184 3130 6236 3136
rect 5552 2961 5580 3130
rect 5906 3088 5962 3097
rect 5906 3023 5962 3032
rect 5920 2990 5948 3023
rect 5724 2984 5776 2990
rect 5538 2952 5594 2961
rect 5724 2926 5776 2932
rect 5908 2984 5960 2990
rect 5908 2926 5960 2932
rect 5538 2887 5594 2896
rect 5736 2650 5764 2926
rect 5724 2644 5776 2650
rect 5724 2586 5776 2592
rect 5736 2514 5764 2586
rect 6380 2582 6408 4126
rect 6472 3602 6500 4712
rect 6644 4480 6696 4486
rect 6644 4422 6696 4428
rect 6656 3942 6684 4422
rect 6840 4185 6868 7364
rect 7288 7346 7340 7352
rect 7944 6798 7972 7822
rect 7380 6792 7432 6798
rect 7380 6734 7432 6740
rect 7932 6792 7984 6798
rect 7932 6734 7984 6740
rect 7288 6248 7340 6254
rect 7288 6190 7340 6196
rect 7300 5914 7328 6190
rect 7392 5914 7420 6734
rect 7472 6180 7524 6186
rect 7472 6122 7524 6128
rect 7288 5908 7340 5914
rect 7288 5850 7340 5856
rect 7380 5908 7432 5914
rect 7380 5850 7432 5856
rect 7300 4690 7328 5850
rect 7484 5710 7512 6122
rect 7840 6112 7892 6118
rect 7840 6054 7892 6060
rect 7852 5914 7880 6054
rect 7840 5908 7892 5914
rect 7840 5850 7892 5856
rect 7472 5704 7524 5710
rect 7472 5646 7524 5652
rect 7484 5370 7512 5646
rect 7472 5364 7524 5370
rect 7472 5306 7524 5312
rect 7380 5160 7432 5166
rect 7380 5102 7432 5108
rect 7392 4758 7420 5102
rect 7852 5098 7880 5850
rect 7840 5092 7892 5098
rect 7840 5034 7892 5040
rect 7472 5024 7524 5030
rect 8036 5001 8064 8298
rect 8680 8294 8708 8978
rect 8116 8288 8168 8294
rect 8116 8230 8168 8236
rect 8668 8288 8720 8294
rect 8668 8230 8720 8236
rect 8128 8129 8156 8230
rect 8289 8188 8585 8208
rect 8345 8186 8369 8188
rect 8425 8186 8449 8188
rect 8505 8186 8529 8188
rect 8367 8134 8369 8186
rect 8431 8134 8443 8186
rect 8505 8134 8507 8186
rect 8345 8132 8369 8134
rect 8425 8132 8449 8134
rect 8505 8132 8529 8134
rect 8114 8120 8170 8129
rect 8289 8112 8585 8132
rect 8114 8055 8170 8064
rect 8116 8016 8168 8022
rect 8680 7993 8708 8230
rect 8864 8090 8892 9930
rect 8944 9580 8996 9586
rect 8944 9522 8996 9528
rect 8956 9178 8984 9522
rect 8944 9172 8996 9178
rect 8944 9114 8996 9120
rect 8852 8084 8904 8090
rect 8852 8026 8904 8032
rect 8116 7958 8168 7964
rect 8666 7984 8722 7993
rect 8128 7410 8156 7958
rect 8666 7919 8722 7928
rect 8300 7880 8352 7886
rect 8220 7840 8300 7868
rect 8116 7404 8168 7410
rect 8116 7346 8168 7352
rect 8128 7206 8156 7346
rect 8116 7200 8168 7206
rect 8116 7142 8168 7148
rect 8128 7002 8156 7142
rect 8116 6996 8168 7002
rect 8116 6938 8168 6944
rect 8220 6866 8248 7840
rect 8300 7822 8352 7828
rect 8680 7154 8708 7919
rect 8864 7546 8892 8026
rect 8852 7540 8904 7546
rect 8852 7482 8904 7488
rect 8760 7268 8812 7274
rect 8864 7256 8892 7482
rect 8812 7228 8892 7256
rect 8760 7210 8812 7216
rect 8680 7126 8892 7154
rect 8289 7100 8585 7120
rect 8345 7098 8369 7100
rect 8425 7098 8449 7100
rect 8505 7098 8529 7100
rect 8367 7046 8369 7098
rect 8431 7046 8443 7098
rect 8505 7046 8507 7098
rect 8345 7044 8369 7046
rect 8425 7044 8449 7046
rect 8505 7044 8529 7046
rect 8289 7024 8585 7044
rect 8208 6860 8260 6866
rect 8208 6802 8260 6808
rect 8760 6860 8812 6866
rect 8760 6802 8812 6808
rect 8116 6452 8168 6458
rect 8116 6394 8168 6400
rect 7472 4966 7524 4972
rect 8022 4992 8078 5001
rect 7380 4752 7432 4758
rect 7380 4694 7432 4700
rect 7012 4684 7064 4690
rect 7012 4626 7064 4632
rect 7288 4684 7340 4690
rect 7288 4626 7340 4632
rect 6826 4176 6882 4185
rect 6826 4111 6882 4120
rect 6644 3936 6696 3942
rect 6644 3878 6696 3884
rect 6460 3596 6512 3602
rect 6460 3538 6512 3544
rect 6472 2650 6500 3538
rect 6460 2644 6512 2650
rect 6460 2586 6512 2592
rect 5908 2576 5960 2582
rect 5908 2518 5960 2524
rect 6368 2576 6420 2582
rect 6368 2518 6420 2524
rect 5724 2508 5776 2514
rect 5724 2450 5776 2456
rect 5920 2417 5948 2518
rect 5906 2408 5962 2417
rect 5906 2343 5962 2352
rect 6656 2106 6684 3878
rect 6840 2990 6868 4111
rect 7024 3738 7052 4626
rect 7484 4486 7512 4966
rect 8022 4927 8078 4936
rect 7930 4720 7986 4729
rect 7930 4655 7986 4664
rect 7944 4622 7972 4655
rect 8128 4622 8156 6394
rect 8772 6225 8800 6802
rect 8758 6216 8814 6225
rect 8758 6151 8814 6160
rect 8772 6118 8800 6151
rect 8760 6112 8812 6118
rect 8666 6080 8722 6089
rect 8289 6012 8585 6032
rect 8760 6054 8812 6060
rect 8666 6015 8722 6024
rect 8345 6010 8369 6012
rect 8425 6010 8449 6012
rect 8505 6010 8529 6012
rect 8367 5958 8369 6010
rect 8431 5958 8443 6010
rect 8505 5958 8507 6010
rect 8345 5956 8369 5958
rect 8425 5956 8449 5958
rect 8505 5956 8529 5958
rect 8289 5936 8585 5956
rect 8680 5234 8708 6015
rect 8668 5228 8720 5234
rect 8668 5170 8720 5176
rect 8289 4924 8585 4944
rect 8345 4922 8369 4924
rect 8425 4922 8449 4924
rect 8505 4922 8529 4924
rect 8367 4870 8369 4922
rect 8431 4870 8443 4922
rect 8505 4870 8507 4922
rect 8345 4868 8369 4870
rect 8425 4868 8449 4870
rect 8505 4868 8529 4870
rect 8289 4848 8585 4868
rect 8208 4752 8260 4758
rect 8208 4694 8260 4700
rect 7932 4616 7984 4622
rect 7932 4558 7984 4564
rect 8116 4616 8168 4622
rect 8116 4558 8168 4564
rect 7472 4480 7524 4486
rect 7472 4422 7524 4428
rect 7564 4480 7616 4486
rect 7564 4422 7616 4428
rect 7104 4072 7156 4078
rect 7104 4014 7156 4020
rect 7194 4040 7250 4049
rect 7012 3732 7064 3738
rect 7012 3674 7064 3680
rect 7116 3670 7144 4014
rect 7194 3975 7250 3984
rect 7104 3664 7156 3670
rect 7104 3606 7156 3612
rect 7208 3369 7236 3975
rect 7484 3942 7512 4422
rect 7472 3936 7524 3942
rect 7286 3904 7342 3913
rect 7472 3878 7524 3884
rect 7286 3839 7342 3848
rect 7300 3738 7328 3839
rect 7288 3732 7340 3738
rect 7288 3674 7340 3680
rect 7576 3534 7604 4422
rect 8220 4078 8248 4694
rect 8668 4276 8720 4282
rect 8668 4218 8720 4224
rect 8208 4072 8260 4078
rect 8208 4014 8260 4020
rect 7656 3936 7708 3942
rect 8680 3913 8708 4218
rect 8864 4078 8892 7126
rect 8944 6928 8996 6934
rect 8944 6870 8996 6876
rect 8956 6186 8984 6870
rect 9036 6316 9088 6322
rect 9036 6258 9088 6264
rect 9048 6225 9076 6258
rect 9034 6216 9090 6225
rect 8944 6180 8996 6186
rect 9034 6151 9090 6160
rect 8944 6122 8996 6128
rect 9140 5914 9168 12038
rect 9784 11898 9812 12174
rect 9876 12102 9904 13087
rect 9864 12096 9916 12102
rect 9864 12038 9916 12044
rect 9772 11892 9824 11898
rect 9772 11834 9824 11840
rect 9864 11212 9916 11218
rect 9864 11154 9916 11160
rect 9770 10840 9826 10849
rect 9770 10775 9826 10784
rect 9784 10606 9812 10775
rect 9772 10600 9824 10606
rect 9772 10542 9824 10548
rect 9876 10266 9904 11154
rect 9954 10432 10010 10441
rect 9954 10367 10010 10376
rect 9588 10260 9640 10266
rect 9588 10202 9640 10208
rect 9864 10260 9916 10266
rect 9864 10202 9916 10208
rect 9600 9586 9628 10202
rect 9968 10130 9996 10367
rect 9956 10124 10008 10130
rect 9956 10066 10008 10072
rect 9864 9988 9916 9994
rect 9864 9930 9916 9936
rect 9588 9580 9640 9586
rect 9588 9522 9640 9528
rect 9312 8968 9364 8974
rect 9312 8910 9364 8916
rect 9220 8492 9272 8498
rect 9220 8434 9272 8440
rect 9232 8090 9260 8434
rect 9220 8084 9272 8090
rect 9220 8026 9272 8032
rect 9324 5930 9352 8910
rect 9496 8628 9548 8634
rect 9496 8570 9548 8576
rect 9508 8362 9536 8570
rect 9496 8356 9548 8362
rect 9496 8298 9548 8304
rect 9404 8016 9456 8022
rect 9404 7958 9456 7964
rect 9416 7342 9444 7958
rect 9772 7948 9824 7954
rect 9772 7890 9824 7896
rect 9680 7540 9732 7546
rect 9680 7482 9732 7488
rect 9692 7449 9720 7482
rect 9784 7478 9812 7890
rect 9876 7750 9904 9930
rect 9968 9382 9996 10066
rect 9956 9376 10008 9382
rect 9956 9318 10008 9324
rect 9968 8537 9996 9318
rect 9954 8528 10010 8537
rect 9954 8463 10010 8472
rect 9864 7744 9916 7750
rect 9864 7686 9916 7692
rect 9772 7472 9824 7478
rect 9678 7440 9734 7449
rect 9772 7414 9824 7420
rect 9678 7375 9734 7384
rect 9404 7336 9456 7342
rect 9404 7278 9456 7284
rect 9496 7200 9548 7206
rect 9496 7142 9548 7148
rect 9404 6112 9456 6118
rect 9404 6054 9456 6060
rect 9128 5908 9180 5914
rect 9128 5850 9180 5856
rect 9232 5902 9352 5930
rect 9140 5302 9168 5850
rect 9128 5296 9180 5302
rect 9128 5238 9180 5244
rect 9232 4154 9260 5902
rect 9312 5840 9364 5846
rect 9312 5782 9364 5788
rect 9324 5098 9352 5782
rect 9416 5710 9444 6054
rect 9508 5778 9536 7142
rect 10060 6984 10088 13767
rect 10152 9994 10180 13874
rect 10244 13433 10272 13942
rect 10336 13870 10364 14418
rect 10416 14272 10468 14278
rect 10416 14214 10468 14220
rect 10324 13864 10376 13870
rect 10324 13806 10376 13812
rect 10230 13424 10286 13433
rect 10230 13359 10286 13368
rect 10140 9988 10192 9994
rect 10140 9930 10192 9936
rect 10244 8566 10272 13359
rect 10428 13258 10456 14214
rect 10520 13938 10548 16526
rect 10612 14346 10640 17002
rect 10704 16998 10732 17682
rect 10784 17672 10836 17678
rect 10784 17614 10836 17620
rect 10692 16992 10744 16998
rect 10692 16934 10744 16940
rect 10796 16794 10824 17614
rect 10784 16788 10836 16794
rect 10784 16730 10836 16736
rect 10796 16114 10824 16730
rect 10784 16108 10836 16114
rect 10784 16050 10836 16056
rect 10692 14816 10744 14822
rect 10692 14758 10744 14764
rect 10600 14340 10652 14346
rect 10600 14282 10652 14288
rect 10508 13932 10560 13938
rect 10508 13874 10560 13880
rect 10704 13462 10732 14758
rect 10888 13814 10916 18294
rect 11900 18086 11928 18770
rect 12624 18624 12676 18630
rect 12624 18566 12676 18572
rect 11956 18524 12252 18544
rect 12012 18522 12036 18524
rect 12092 18522 12116 18524
rect 12172 18522 12196 18524
rect 12034 18470 12036 18522
rect 12098 18470 12110 18522
rect 12172 18470 12174 18522
rect 12012 18468 12036 18470
rect 12092 18468 12116 18470
rect 12172 18468 12196 18470
rect 11956 18448 12252 18468
rect 12636 18222 12664 18566
rect 13464 18426 13492 18770
rect 13452 18420 13504 18426
rect 13452 18362 13504 18368
rect 12624 18216 12676 18222
rect 12624 18158 12676 18164
rect 13176 18216 13228 18222
rect 13176 18158 13228 18164
rect 10968 18080 11020 18086
rect 10968 18022 11020 18028
rect 11888 18080 11940 18086
rect 11888 18022 11940 18028
rect 12348 18080 12400 18086
rect 12348 18022 12400 18028
rect 10980 15065 11008 18022
rect 11060 17196 11112 17202
rect 11060 17138 11112 17144
rect 11072 17105 11100 17138
rect 11058 17096 11114 17105
rect 11058 17031 11114 17040
rect 11704 16992 11756 16998
rect 11704 16934 11756 16940
rect 11716 16590 11744 16934
rect 11796 16720 11848 16726
rect 11796 16662 11848 16668
rect 11704 16584 11756 16590
rect 11704 16526 11756 16532
rect 11716 16250 11744 16526
rect 11704 16244 11756 16250
rect 11704 16186 11756 16192
rect 11808 16182 11836 16662
rect 11900 16590 11928 18022
rect 11956 17436 12252 17456
rect 12012 17434 12036 17436
rect 12092 17434 12116 17436
rect 12172 17434 12196 17436
rect 12034 17382 12036 17434
rect 12098 17382 12110 17434
rect 12172 17382 12174 17434
rect 12012 17380 12036 17382
rect 12092 17380 12116 17382
rect 12172 17380 12196 17382
rect 11956 17360 12252 17380
rect 12360 17202 12388 18022
rect 12636 17270 12664 18158
rect 13188 17746 13216 18158
rect 13268 18148 13320 18154
rect 13268 18090 13320 18096
rect 12808 17740 12860 17746
rect 12808 17682 12860 17688
rect 13176 17740 13228 17746
rect 13176 17682 13228 17688
rect 12820 17610 12848 17682
rect 12808 17604 12860 17610
rect 12808 17546 12860 17552
rect 12716 17536 12768 17542
rect 12716 17478 12768 17484
rect 12728 17377 12756 17478
rect 12714 17368 12770 17377
rect 12714 17303 12770 17312
rect 12624 17264 12676 17270
rect 12624 17206 12676 17212
rect 12348 17196 12400 17202
rect 12348 17138 12400 17144
rect 12360 16998 12388 17138
rect 12728 17134 12756 17303
rect 12716 17128 12768 17134
rect 12716 17070 12768 17076
rect 12348 16992 12400 16998
rect 12348 16934 12400 16940
rect 12716 16992 12768 16998
rect 12716 16934 12768 16940
rect 11888 16584 11940 16590
rect 11888 16526 11940 16532
rect 11796 16176 11848 16182
rect 11796 16118 11848 16124
rect 11704 15632 11756 15638
rect 11704 15574 11756 15580
rect 11612 15496 11664 15502
rect 11612 15438 11664 15444
rect 11336 15360 11388 15366
rect 11336 15302 11388 15308
rect 10966 15056 11022 15065
rect 10966 14991 11022 15000
rect 11152 14884 11204 14890
rect 11152 14826 11204 14832
rect 10968 14816 11020 14822
rect 10968 14758 11020 14764
rect 10980 14550 11008 14758
rect 10968 14544 11020 14550
rect 10968 14486 11020 14492
rect 10796 13786 10916 13814
rect 10692 13456 10744 13462
rect 10692 13398 10744 13404
rect 10692 13320 10744 13326
rect 10692 13262 10744 13268
rect 10416 13252 10468 13258
rect 10416 13194 10468 13200
rect 10324 13184 10376 13190
rect 10324 13126 10376 13132
rect 10336 12918 10364 13126
rect 10324 12912 10376 12918
rect 10324 12854 10376 12860
rect 10508 12708 10560 12714
rect 10508 12650 10560 12656
rect 10520 11694 10548 12650
rect 10704 12442 10732 13262
rect 10692 12436 10744 12442
rect 10692 12378 10744 12384
rect 10508 11688 10560 11694
rect 10508 11630 10560 11636
rect 10416 11552 10468 11558
rect 10416 11494 10468 11500
rect 10428 11286 10456 11494
rect 10416 11280 10468 11286
rect 10416 11222 10468 11228
rect 10322 11112 10378 11121
rect 10322 11047 10378 11056
rect 10232 8560 10284 8566
rect 10232 8502 10284 8508
rect 10336 8480 10364 11047
rect 10428 10470 10456 11222
rect 10416 10464 10468 10470
rect 10796 10441 10824 13786
rect 11164 13258 11192 14826
rect 11348 13530 11376 15302
rect 11624 14890 11652 15438
rect 11716 15162 11744 15574
rect 11900 15502 11928 16526
rect 11956 16348 12252 16368
rect 12012 16346 12036 16348
rect 12092 16346 12116 16348
rect 12172 16346 12196 16348
rect 12034 16294 12036 16346
rect 12098 16294 12110 16346
rect 12172 16294 12174 16346
rect 12012 16292 12036 16294
rect 12092 16292 12116 16294
rect 12172 16292 12196 16294
rect 11956 16272 12252 16292
rect 11888 15496 11940 15502
rect 11888 15438 11940 15444
rect 11704 15156 11756 15162
rect 11704 15098 11756 15104
rect 11612 14884 11664 14890
rect 11612 14826 11664 14832
rect 11900 14550 11928 15438
rect 12360 15366 12388 16934
rect 12532 16788 12584 16794
rect 12532 16730 12584 16736
rect 12348 15360 12400 15366
rect 12348 15302 12400 15308
rect 11956 15260 12252 15280
rect 12012 15258 12036 15260
rect 12092 15258 12116 15260
rect 12172 15258 12196 15260
rect 12034 15206 12036 15258
rect 12098 15206 12110 15258
rect 12172 15206 12174 15258
rect 12012 15204 12036 15206
rect 12092 15204 12116 15206
rect 12172 15204 12196 15206
rect 11956 15184 12252 15204
rect 12544 14618 12572 16730
rect 12624 16652 12676 16658
rect 12624 16594 12676 16600
rect 12636 16114 12664 16594
rect 12624 16108 12676 16114
rect 12624 16050 12676 16056
rect 12532 14612 12584 14618
rect 12532 14554 12584 14560
rect 11520 14544 11572 14550
rect 11520 14486 11572 14492
rect 11888 14544 11940 14550
rect 11888 14486 11940 14492
rect 11428 13728 11480 13734
rect 11428 13670 11480 13676
rect 11336 13524 11388 13530
rect 11336 13466 11388 13472
rect 11440 13462 11468 13670
rect 11532 13530 11560 14486
rect 11796 14408 11848 14414
rect 11796 14350 11848 14356
rect 11520 13524 11572 13530
rect 11520 13466 11572 13472
rect 11428 13456 11480 13462
rect 11428 13398 11480 13404
rect 11152 13252 11204 13258
rect 11152 13194 11204 13200
rect 11164 12714 11192 13194
rect 11440 12986 11468 13398
rect 11808 13190 11836 14350
rect 11956 14172 12252 14192
rect 12012 14170 12036 14172
rect 12092 14170 12116 14172
rect 12172 14170 12196 14172
rect 12034 14118 12036 14170
rect 12098 14118 12110 14170
rect 12172 14118 12174 14170
rect 12012 14116 12036 14118
rect 12092 14116 12116 14118
rect 12172 14116 12196 14118
rect 11956 14096 12252 14116
rect 12544 13938 12572 14554
rect 12532 13932 12584 13938
rect 12532 13874 12584 13880
rect 12624 13728 12676 13734
rect 12624 13670 12676 13676
rect 11888 13456 11940 13462
rect 11888 13398 11940 13404
rect 11520 13184 11572 13190
rect 11520 13126 11572 13132
rect 11796 13184 11848 13190
rect 11796 13126 11848 13132
rect 11428 12980 11480 12986
rect 11428 12922 11480 12928
rect 11152 12708 11204 12714
rect 11152 12650 11204 12656
rect 11532 12238 11560 13126
rect 11900 12918 11928 13398
rect 12348 13320 12400 13326
rect 12348 13262 12400 13268
rect 11956 13084 12252 13104
rect 12012 13082 12036 13084
rect 12092 13082 12116 13084
rect 12172 13082 12196 13084
rect 12034 13030 12036 13082
rect 12098 13030 12110 13082
rect 12172 13030 12174 13082
rect 12012 13028 12036 13030
rect 12092 13028 12116 13030
rect 12172 13028 12196 13030
rect 11956 13008 12252 13028
rect 11888 12912 11940 12918
rect 11888 12854 11940 12860
rect 11888 12708 11940 12714
rect 11888 12650 11940 12656
rect 11612 12368 11664 12374
rect 11612 12310 11664 12316
rect 11520 12232 11572 12238
rect 11520 12174 11572 12180
rect 11244 12164 11296 12170
rect 11244 12106 11296 12112
rect 11060 12096 11112 12102
rect 11060 12038 11112 12044
rect 10876 11688 10928 11694
rect 10876 11630 10928 11636
rect 10888 10538 10916 11630
rect 10876 10532 10928 10538
rect 10876 10474 10928 10480
rect 10416 10406 10468 10412
rect 10782 10432 10838 10441
rect 10428 9926 10456 10406
rect 10782 10367 10838 10376
rect 10888 10266 10916 10474
rect 10876 10260 10928 10266
rect 10876 10202 10928 10208
rect 10416 9920 10468 9926
rect 10416 9862 10468 9868
rect 10692 9920 10744 9926
rect 10692 9862 10744 9868
rect 10600 9580 10652 9586
rect 10600 9522 10652 9528
rect 10612 9178 10640 9522
rect 10704 9450 10732 9862
rect 10692 9444 10744 9450
rect 10692 9386 10744 9392
rect 10600 9172 10652 9178
rect 10600 9114 10652 9120
rect 10416 8968 10468 8974
rect 10416 8910 10468 8916
rect 10968 8968 11020 8974
rect 10968 8910 11020 8916
rect 10428 8634 10456 8910
rect 10980 8838 11008 8910
rect 10508 8832 10560 8838
rect 10508 8774 10560 8780
rect 10968 8832 11020 8838
rect 10968 8774 11020 8780
rect 10416 8628 10468 8634
rect 10416 8570 10468 8576
rect 10336 8452 10456 8480
rect 10324 8356 10376 8362
rect 10324 8298 10376 8304
rect 10060 6956 10272 6984
rect 10140 6860 10192 6866
rect 10140 6802 10192 6808
rect 9772 6724 9824 6730
rect 9772 6666 9824 6672
rect 10048 6724 10100 6730
rect 10048 6666 10100 6672
rect 9588 6180 9640 6186
rect 9588 6122 9640 6128
rect 9496 5772 9548 5778
rect 9496 5714 9548 5720
rect 9404 5704 9456 5710
rect 9404 5646 9456 5652
rect 9312 5092 9364 5098
rect 9312 5034 9364 5040
rect 9324 4826 9352 5034
rect 9600 4826 9628 6122
rect 9784 5710 9812 6666
rect 9956 6656 10008 6662
rect 9956 6598 10008 6604
rect 9968 6458 9996 6598
rect 9956 6452 10008 6458
rect 9956 6394 10008 6400
rect 10060 6390 10088 6666
rect 10048 6384 10100 6390
rect 10048 6326 10100 6332
rect 9956 6316 10008 6322
rect 9956 6258 10008 6264
rect 9772 5704 9824 5710
rect 9772 5646 9824 5652
rect 9968 5234 9996 6258
rect 10060 5914 10088 6326
rect 10152 6254 10180 6802
rect 10140 6248 10192 6254
rect 10140 6190 10192 6196
rect 10152 6089 10180 6190
rect 10138 6080 10194 6089
rect 10138 6015 10194 6024
rect 10048 5908 10100 5914
rect 10048 5850 10100 5856
rect 9956 5228 10008 5234
rect 9956 5170 10008 5176
rect 9312 4820 9364 4826
rect 9312 4762 9364 4768
rect 9588 4820 9640 4826
rect 9588 4762 9640 4768
rect 9140 4126 9260 4154
rect 8852 4072 8904 4078
rect 8852 4014 8904 4020
rect 8760 3936 8812 3942
rect 7656 3878 7708 3884
rect 8666 3904 8722 3913
rect 7668 3602 7696 3878
rect 8289 3836 8585 3856
rect 8760 3878 8812 3884
rect 8666 3839 8722 3848
rect 8345 3834 8369 3836
rect 8425 3834 8449 3836
rect 8505 3834 8529 3836
rect 8367 3782 8369 3834
rect 8431 3782 8443 3834
rect 8505 3782 8507 3834
rect 8345 3780 8369 3782
rect 8425 3780 8449 3782
rect 8505 3780 8529 3782
rect 8289 3760 8585 3780
rect 8772 3670 8800 3878
rect 8760 3664 8812 3670
rect 8760 3606 8812 3612
rect 7656 3596 7708 3602
rect 7656 3538 7708 3544
rect 7564 3528 7616 3534
rect 7564 3470 7616 3476
rect 7194 3360 7250 3369
rect 7194 3295 7250 3304
rect 7196 3188 7248 3194
rect 7196 3130 7248 3136
rect 6828 2984 6880 2990
rect 6828 2926 6880 2932
rect 6644 2100 6696 2106
rect 6644 2042 6696 2048
rect 4894 54 5120 82
rect 6918 82 6974 480
rect 7208 82 7236 3130
rect 7288 2848 7340 2854
rect 7288 2790 7340 2796
rect 6918 54 7236 82
rect 7300 66 7328 2790
rect 7668 2582 7696 3538
rect 8772 3126 8800 3606
rect 8864 3194 8892 4014
rect 8944 3936 8996 3942
rect 8944 3878 8996 3884
rect 8852 3188 8904 3194
rect 8852 3130 8904 3136
rect 8760 3120 8812 3126
rect 8760 3062 8812 3068
rect 8576 2916 8628 2922
rect 8956 2904 8984 3878
rect 9036 3392 9088 3398
rect 9036 3334 9088 3340
rect 9048 3058 9076 3334
rect 9036 3052 9088 3058
rect 9036 2994 9088 3000
rect 8628 2876 8984 2904
rect 8576 2858 8628 2864
rect 7748 2848 7800 2854
rect 7748 2790 7800 2796
rect 7760 2582 7788 2790
rect 8289 2748 8585 2768
rect 8345 2746 8369 2748
rect 8425 2746 8449 2748
rect 8505 2746 8529 2748
rect 8367 2694 8369 2746
rect 8431 2694 8443 2746
rect 8505 2694 8507 2746
rect 8345 2692 8369 2694
rect 8425 2692 8449 2694
rect 8505 2692 8529 2694
rect 8289 2672 8585 2692
rect 8680 2582 8708 2876
rect 7656 2576 7708 2582
rect 7656 2518 7708 2524
rect 7748 2576 7800 2582
rect 7748 2518 7800 2524
rect 8668 2576 8720 2582
rect 8668 2518 8720 2524
rect 7760 2310 7788 2518
rect 7748 2304 7800 2310
rect 7748 2246 7800 2252
rect 7760 2106 7788 2246
rect 7748 2100 7800 2106
rect 7748 2042 7800 2048
rect 8850 82 8906 480
rect 9140 82 9168 4126
rect 9600 3534 9628 4762
rect 9864 4752 9916 4758
rect 9864 4694 9916 4700
rect 9680 4548 9732 4554
rect 9680 4490 9732 4496
rect 9692 4214 9720 4490
rect 9876 4282 9904 4694
rect 9968 4622 9996 5170
rect 10244 5030 10272 6956
rect 10336 5370 10364 8298
rect 10428 6168 10456 8452
rect 10520 6798 10548 8774
rect 10692 7744 10744 7750
rect 10692 7686 10744 7692
rect 10600 7540 10652 7546
rect 10600 7482 10652 7488
rect 10612 7449 10640 7482
rect 10598 7440 10654 7449
rect 10598 7375 10654 7384
rect 10508 6792 10560 6798
rect 10508 6734 10560 6740
rect 10508 6180 10560 6186
rect 10428 6140 10508 6168
rect 10508 6122 10560 6128
rect 10520 5710 10548 6122
rect 10416 5704 10468 5710
rect 10416 5646 10468 5652
rect 10508 5704 10560 5710
rect 10508 5646 10560 5652
rect 10324 5364 10376 5370
rect 10324 5306 10376 5312
rect 10232 5024 10284 5030
rect 10232 4966 10284 4972
rect 9956 4616 10008 4622
rect 9956 4558 10008 4564
rect 9864 4276 9916 4282
rect 9864 4218 9916 4224
rect 9680 4208 9732 4214
rect 9680 4150 9732 4156
rect 9588 3528 9640 3534
rect 9588 3470 9640 3476
rect 9692 3466 9720 4150
rect 9968 3670 9996 4558
rect 10336 4154 10364 5306
rect 10428 4826 10456 5646
rect 10600 5092 10652 5098
rect 10600 5034 10652 5040
rect 10416 4820 10468 4826
rect 10416 4762 10468 4768
rect 10336 4126 10456 4154
rect 10428 3942 10456 4126
rect 10416 3936 10468 3942
rect 10416 3878 10468 3884
rect 10140 3732 10192 3738
rect 10140 3674 10192 3680
rect 9864 3664 9916 3670
rect 9864 3606 9916 3612
rect 9956 3664 10008 3670
rect 9956 3606 10008 3612
rect 9680 3460 9732 3466
rect 9680 3402 9732 3408
rect 9312 3392 9364 3398
rect 9312 3334 9364 3340
rect 9324 2446 9352 3334
rect 9876 3194 9904 3606
rect 10152 3194 10180 3674
rect 10612 3641 10640 5034
rect 10598 3632 10654 3641
rect 10598 3567 10654 3576
rect 10324 3460 10376 3466
rect 10324 3402 10376 3408
rect 9864 3188 9916 3194
rect 9864 3130 9916 3136
rect 10140 3188 10192 3194
rect 10140 3130 10192 3136
rect 10336 2446 10364 3402
rect 9312 2440 9364 2446
rect 9312 2382 9364 2388
rect 10324 2440 10376 2446
rect 10324 2382 10376 2388
rect 7288 60 7340 66
rect 2870 0 2926 54
rect 4894 0 4950 54
rect 6918 0 6974 54
rect 7288 2 7340 8
rect 8850 54 9168 82
rect 10704 82 10732 7686
rect 10980 7002 11008 8774
rect 11072 7002 11100 12038
rect 11256 11354 11284 12106
rect 11244 11348 11296 11354
rect 11244 11290 11296 11296
rect 11256 11257 11284 11290
rect 11242 11248 11298 11257
rect 11242 11183 11298 11192
rect 11428 11144 11480 11150
rect 11428 11086 11480 11092
rect 11440 10198 11468 11086
rect 11532 10674 11560 12174
rect 11624 11558 11652 12310
rect 11796 11824 11848 11830
rect 11796 11766 11848 11772
rect 11808 11626 11836 11766
rect 11796 11620 11848 11626
rect 11796 11562 11848 11568
rect 11612 11552 11664 11558
rect 11612 11494 11664 11500
rect 11624 11286 11652 11494
rect 11612 11280 11664 11286
rect 11612 11222 11664 11228
rect 11624 10810 11652 11222
rect 11900 11150 11928 12650
rect 12360 12442 12388 13262
rect 12636 12696 12664 13670
rect 12728 12850 12756 16934
rect 12820 16454 12848 17546
rect 13188 17134 13216 17682
rect 13176 17128 13228 17134
rect 13176 17070 13228 17076
rect 12808 16448 12860 16454
rect 12808 16390 12860 16396
rect 13280 16114 13308 18090
rect 13556 17814 13584 21542
rect 15842 21542 15976 21570
rect 15842 21520 15898 21542
rect 14462 20904 14518 20913
rect 14462 20839 14518 20848
rect 13820 19304 13872 19310
rect 13820 19246 13872 19252
rect 13636 18624 13688 18630
rect 13636 18566 13688 18572
rect 13544 17808 13596 17814
rect 13544 17750 13596 17756
rect 13360 17672 13412 17678
rect 13360 17614 13412 17620
rect 13268 16108 13320 16114
rect 13268 16050 13320 16056
rect 13372 15570 13400 17614
rect 13544 17128 13596 17134
rect 13544 17070 13596 17076
rect 13452 16788 13504 16794
rect 13452 16730 13504 16736
rect 13360 15564 13412 15570
rect 13360 15506 13412 15512
rect 12900 14952 12952 14958
rect 12900 14894 12952 14900
rect 12808 14816 12860 14822
rect 12808 14758 12860 14764
rect 12820 13326 12848 14758
rect 12912 14328 12940 14894
rect 13372 14618 13400 15506
rect 13464 15026 13492 16730
rect 13556 16658 13584 17070
rect 13544 16652 13596 16658
rect 13544 16594 13596 16600
rect 13452 15020 13504 15026
rect 13452 14962 13504 14968
rect 13360 14612 13412 14618
rect 13360 14554 13412 14560
rect 12992 14340 13044 14346
rect 12912 14300 12992 14328
rect 12808 13320 12860 13326
rect 12912 13297 12940 14300
rect 12992 14282 13044 14288
rect 13464 14278 13492 14962
rect 13544 14544 13596 14550
rect 13544 14486 13596 14492
rect 13452 14272 13504 14278
rect 13452 14214 13504 14220
rect 13452 14068 13504 14074
rect 13452 14010 13504 14016
rect 13360 13728 13412 13734
rect 13360 13670 13412 13676
rect 13372 13462 13400 13670
rect 13464 13530 13492 14010
rect 13556 13734 13584 14486
rect 13544 13728 13596 13734
rect 13544 13670 13596 13676
rect 13452 13524 13504 13530
rect 13452 13466 13504 13472
rect 13360 13456 13412 13462
rect 13360 13398 13412 13404
rect 13452 13320 13504 13326
rect 12808 13262 12860 13268
rect 12898 13288 12954 13297
rect 13452 13262 13504 13268
rect 12898 13223 12954 13232
rect 12716 12844 12768 12850
rect 12716 12786 12768 12792
rect 12716 12708 12768 12714
rect 12636 12668 12716 12696
rect 12716 12650 12768 12656
rect 12348 12436 12400 12442
rect 12348 12378 12400 12384
rect 12728 12102 12756 12650
rect 13464 12442 13492 13262
rect 13452 12436 13504 12442
rect 13452 12378 13504 12384
rect 12716 12096 12768 12102
rect 12716 12038 12768 12044
rect 12808 12096 12860 12102
rect 12808 12038 12860 12044
rect 11956 11996 12252 12016
rect 12012 11994 12036 11996
rect 12092 11994 12116 11996
rect 12172 11994 12196 11996
rect 12034 11942 12036 11994
rect 12098 11942 12110 11994
rect 12172 11942 12174 11994
rect 12012 11940 12036 11942
rect 12092 11940 12116 11942
rect 12172 11940 12196 11942
rect 11956 11920 12252 11940
rect 12728 11558 12756 12038
rect 12716 11552 12768 11558
rect 12716 11494 12768 11500
rect 11888 11144 11940 11150
rect 11888 11086 11940 11092
rect 12440 11144 12492 11150
rect 12440 11086 12492 11092
rect 11956 10908 12252 10928
rect 12012 10906 12036 10908
rect 12092 10906 12116 10908
rect 12172 10906 12196 10908
rect 12034 10854 12036 10906
rect 12098 10854 12110 10906
rect 12172 10854 12174 10906
rect 12012 10852 12036 10854
rect 12092 10852 12116 10854
rect 12172 10852 12196 10854
rect 11956 10832 12252 10852
rect 11612 10804 11664 10810
rect 11612 10746 11664 10752
rect 11520 10668 11572 10674
rect 11520 10610 11572 10616
rect 11520 10464 11572 10470
rect 11520 10406 11572 10412
rect 11244 10192 11296 10198
rect 11244 10134 11296 10140
rect 11428 10192 11480 10198
rect 11532 10169 11560 10406
rect 11428 10134 11480 10140
rect 11518 10160 11574 10169
rect 11152 10056 11204 10062
rect 11152 9998 11204 10004
rect 11164 9654 11192 9998
rect 11152 9648 11204 9654
rect 11152 9590 11204 9596
rect 11256 9382 11284 10134
rect 12452 10130 12480 11086
rect 12532 11076 12584 11082
rect 12532 11018 12584 11024
rect 12544 10674 12572 11018
rect 12532 10668 12584 10674
rect 12532 10610 12584 10616
rect 12622 10568 12678 10577
rect 12622 10503 12678 10512
rect 12636 10130 12664 10503
rect 12820 10266 12848 12038
rect 12900 11688 12952 11694
rect 12900 11630 12952 11636
rect 12912 11354 12940 11630
rect 13360 11552 13412 11558
rect 13360 11494 13412 11500
rect 12900 11348 12952 11354
rect 12900 11290 12952 11296
rect 12808 10260 12860 10266
rect 12808 10202 12860 10208
rect 13372 10198 13400 11494
rect 13544 11280 13596 11286
rect 13544 11222 13596 11228
rect 13452 10532 13504 10538
rect 13452 10474 13504 10480
rect 13360 10192 13412 10198
rect 13360 10134 13412 10140
rect 11518 10095 11574 10104
rect 12440 10124 12492 10130
rect 11336 9444 11388 9450
rect 11336 9386 11388 9392
rect 11244 9376 11296 9382
rect 11244 9318 11296 9324
rect 11348 8022 11376 9386
rect 11336 8016 11388 8022
rect 11336 7958 11388 7964
rect 11348 7274 11376 7958
rect 11428 7812 11480 7818
rect 11428 7754 11480 7760
rect 11336 7268 11388 7274
rect 11336 7210 11388 7216
rect 10968 6996 11020 7002
rect 10968 6938 11020 6944
rect 11060 6996 11112 7002
rect 11060 6938 11112 6944
rect 11336 6996 11388 7002
rect 11336 6938 11388 6944
rect 10968 6656 11020 6662
rect 10968 6598 11020 6604
rect 10980 6186 11008 6598
rect 10968 6180 11020 6186
rect 10968 6122 11020 6128
rect 11244 5568 11296 5574
rect 11244 5510 11296 5516
rect 10784 5160 10836 5166
rect 10784 5102 10836 5108
rect 11060 5160 11112 5166
rect 11060 5102 11112 5108
rect 10796 3602 10824 5102
rect 11072 4486 11100 5102
rect 11256 5030 11284 5510
rect 11244 5024 11296 5030
rect 11244 4966 11296 4972
rect 11060 4480 11112 4486
rect 11060 4422 11112 4428
rect 11348 4154 11376 6938
rect 11440 6934 11468 7754
rect 11532 7342 11560 10095
rect 12440 10066 12492 10072
rect 12624 10124 12676 10130
rect 12624 10066 12676 10072
rect 12452 10033 12480 10066
rect 12438 10024 12494 10033
rect 12438 9959 12494 9968
rect 11956 9820 12252 9840
rect 12012 9818 12036 9820
rect 12092 9818 12116 9820
rect 12172 9818 12196 9820
rect 12034 9766 12036 9818
rect 12098 9766 12110 9818
rect 12172 9766 12174 9818
rect 12012 9764 12036 9766
rect 12092 9764 12116 9766
rect 12172 9764 12196 9766
rect 11956 9744 12252 9764
rect 11888 9376 11940 9382
rect 11888 9318 11940 9324
rect 11900 9110 11928 9318
rect 12636 9178 12664 10066
rect 13084 9988 13136 9994
rect 13084 9930 13136 9936
rect 12806 9888 12862 9897
rect 12806 9823 12862 9832
rect 12820 9722 12848 9823
rect 12808 9716 12860 9722
rect 12808 9658 12860 9664
rect 12624 9172 12676 9178
rect 12624 9114 12676 9120
rect 11888 9104 11940 9110
rect 11888 9046 11940 9052
rect 11794 8936 11850 8945
rect 11704 8900 11756 8906
rect 11756 8880 11794 8888
rect 11756 8871 11850 8880
rect 11756 8860 11836 8871
rect 11704 8842 11756 8848
rect 11900 8566 11928 9046
rect 12348 8968 12400 8974
rect 12348 8910 12400 8916
rect 11956 8732 12252 8752
rect 12012 8730 12036 8732
rect 12092 8730 12116 8732
rect 12172 8730 12196 8732
rect 12034 8678 12036 8730
rect 12098 8678 12110 8730
rect 12172 8678 12174 8730
rect 12012 8676 12036 8678
rect 12092 8676 12116 8678
rect 12172 8676 12196 8678
rect 11956 8656 12252 8676
rect 11888 8560 11940 8566
rect 11888 8502 11940 8508
rect 11612 7880 11664 7886
rect 11612 7822 11664 7828
rect 11624 7546 11652 7822
rect 11796 7744 11848 7750
rect 11796 7686 11848 7692
rect 11612 7540 11664 7546
rect 11612 7482 11664 7488
rect 11520 7336 11572 7342
rect 11520 7278 11572 7284
rect 11808 6934 11836 7686
rect 11956 7644 12252 7664
rect 12012 7642 12036 7644
rect 12092 7642 12116 7644
rect 12172 7642 12196 7644
rect 12034 7590 12036 7642
rect 12098 7590 12110 7642
rect 12172 7590 12174 7642
rect 12012 7588 12036 7590
rect 12092 7588 12116 7590
rect 12172 7588 12196 7590
rect 11956 7568 12252 7588
rect 12360 6934 12388 8910
rect 13096 8566 13124 9930
rect 13372 9450 13400 10134
rect 13360 9444 13412 9450
rect 13360 9386 13412 9392
rect 13464 8974 13492 10474
rect 13556 10470 13584 11222
rect 13544 10464 13596 10470
rect 13544 10406 13596 10412
rect 13556 10266 13584 10406
rect 13544 10260 13596 10266
rect 13544 10202 13596 10208
rect 13452 8968 13504 8974
rect 13452 8910 13504 8916
rect 13084 8560 13136 8566
rect 13084 8502 13136 8508
rect 12716 8492 12768 8498
rect 12716 8434 12768 8440
rect 12532 8356 12584 8362
rect 12532 8298 12584 8304
rect 12624 8356 12676 8362
rect 12624 8298 12676 8304
rect 11428 6928 11480 6934
rect 11428 6870 11480 6876
rect 11796 6928 11848 6934
rect 11796 6870 11848 6876
rect 12348 6928 12400 6934
rect 12348 6870 12400 6876
rect 11440 6390 11468 6870
rect 11808 6458 11836 6870
rect 12544 6866 12572 8298
rect 12636 7750 12664 8298
rect 12728 7750 12756 8434
rect 13268 8356 13320 8362
rect 13268 8298 13320 8304
rect 13280 8090 13308 8298
rect 13268 8084 13320 8090
rect 13268 8026 13320 8032
rect 13544 8084 13596 8090
rect 13544 8026 13596 8032
rect 13452 7948 13504 7954
rect 13452 7890 13504 7896
rect 12624 7744 12676 7750
rect 12624 7686 12676 7692
rect 12716 7744 12768 7750
rect 12716 7686 12768 7692
rect 12532 6860 12584 6866
rect 12532 6802 12584 6808
rect 11956 6556 12252 6576
rect 12012 6554 12036 6556
rect 12092 6554 12116 6556
rect 12172 6554 12196 6556
rect 12034 6502 12036 6554
rect 12098 6502 12110 6554
rect 12172 6502 12174 6554
rect 12012 6500 12036 6502
rect 12092 6500 12116 6502
rect 12172 6500 12196 6502
rect 11956 6480 12252 6500
rect 11612 6452 11664 6458
rect 11612 6394 11664 6400
rect 11796 6452 11848 6458
rect 11796 6394 11848 6400
rect 11428 6384 11480 6390
rect 11428 6326 11480 6332
rect 11624 5098 11652 6394
rect 12348 6248 12400 6254
rect 12348 6190 12400 6196
rect 11796 5772 11848 5778
rect 11796 5714 11848 5720
rect 11808 5370 11836 5714
rect 11956 5468 12252 5488
rect 12012 5466 12036 5468
rect 12092 5466 12116 5468
rect 12172 5466 12196 5468
rect 12034 5414 12036 5466
rect 12098 5414 12110 5466
rect 12172 5414 12174 5466
rect 12012 5412 12036 5414
rect 12092 5412 12116 5414
rect 12172 5412 12196 5414
rect 11956 5392 12252 5412
rect 11796 5364 11848 5370
rect 11848 5324 11928 5352
rect 11796 5306 11848 5312
rect 11612 5092 11664 5098
rect 11612 5034 11664 5040
rect 11796 4684 11848 4690
rect 11796 4626 11848 4632
rect 11520 4616 11572 4622
rect 11808 4593 11836 4626
rect 11520 4558 11572 4564
rect 11794 4584 11850 4593
rect 11428 4480 11480 4486
rect 11428 4422 11480 4428
rect 11256 4126 11376 4154
rect 11256 3738 11284 4126
rect 11440 4078 11468 4422
rect 11428 4072 11480 4078
rect 11428 4014 11480 4020
rect 11244 3732 11296 3738
rect 11244 3674 11296 3680
rect 10784 3596 10836 3602
rect 10784 3538 10836 3544
rect 11244 3596 11296 3602
rect 11244 3538 11296 3544
rect 10796 3369 10824 3538
rect 10876 3460 10928 3466
rect 10876 3402 10928 3408
rect 10782 3360 10838 3369
rect 10782 3295 10838 3304
rect 10888 3126 10916 3402
rect 11256 3194 11284 3538
rect 11244 3188 11296 3194
rect 11244 3130 11296 3136
rect 10876 3120 10928 3126
rect 10876 3062 10928 3068
rect 10784 2984 10836 2990
rect 10876 2984 10928 2990
rect 10784 2926 10836 2932
rect 10874 2952 10876 2961
rect 10928 2952 10930 2961
rect 10796 2854 10824 2926
rect 10874 2887 10930 2896
rect 10784 2848 10836 2854
rect 10784 2790 10836 2796
rect 10888 2650 10916 2887
rect 11256 2650 11284 3130
rect 10876 2644 10928 2650
rect 10876 2586 10928 2592
rect 11244 2644 11296 2650
rect 11244 2586 11296 2592
rect 11440 2514 11468 4014
rect 11532 3058 11560 4558
rect 11900 4570 11928 5324
rect 12360 5273 12388 6190
rect 12532 6180 12584 6186
rect 12532 6122 12584 6128
rect 12440 5568 12492 5574
rect 12440 5510 12492 5516
rect 12346 5264 12402 5273
rect 12346 5199 12348 5208
rect 12400 5199 12402 5208
rect 12348 5170 12400 5176
rect 12360 5139 12388 5170
rect 12452 5166 12480 5510
rect 12440 5160 12492 5166
rect 12544 5137 12572 6122
rect 12622 6080 12678 6089
rect 12622 6015 12678 6024
rect 12440 5102 12492 5108
rect 12530 5128 12586 5137
rect 12348 5092 12400 5098
rect 12348 5034 12400 5040
rect 11978 4584 12034 4593
rect 11900 4554 11978 4570
rect 11794 4519 11850 4528
rect 11888 4548 11978 4554
rect 11940 4542 11978 4548
rect 11978 4519 12034 4528
rect 11888 4490 11940 4496
rect 11900 4214 11928 4490
rect 11956 4380 12252 4400
rect 12012 4378 12036 4380
rect 12092 4378 12116 4380
rect 12172 4378 12196 4380
rect 12034 4326 12036 4378
rect 12098 4326 12110 4378
rect 12172 4326 12174 4378
rect 12012 4324 12036 4326
rect 12092 4324 12116 4326
rect 12172 4324 12196 4326
rect 11956 4304 12252 4324
rect 11888 4208 11940 4214
rect 11888 4150 11940 4156
rect 11888 3596 11940 3602
rect 11888 3538 11940 3544
rect 11520 3052 11572 3058
rect 11520 2994 11572 3000
rect 11900 2990 11928 3538
rect 12360 3466 12388 5034
rect 12452 4758 12480 5102
rect 12530 5063 12586 5072
rect 12440 4752 12492 4758
rect 12440 4694 12492 4700
rect 12440 4616 12492 4622
rect 12440 4558 12492 4564
rect 12452 3602 12480 4558
rect 12544 4010 12572 5063
rect 12636 4758 12664 6015
rect 12624 4752 12676 4758
rect 12624 4694 12676 4700
rect 12636 4214 12664 4694
rect 12728 4282 12756 7686
rect 13464 7478 13492 7890
rect 13452 7472 13504 7478
rect 13452 7414 13504 7420
rect 13556 7206 13584 8026
rect 12808 7200 12860 7206
rect 12808 7142 12860 7148
rect 13544 7200 13596 7206
rect 13544 7142 13596 7148
rect 12820 5817 12848 7142
rect 13452 6860 13504 6866
rect 13452 6802 13504 6808
rect 13176 6792 13228 6798
rect 13176 6734 13228 6740
rect 13188 6118 13216 6734
rect 13464 6458 13492 6802
rect 13556 6662 13584 7142
rect 13544 6656 13596 6662
rect 13544 6598 13596 6604
rect 13452 6452 13504 6458
rect 13452 6394 13504 6400
rect 13176 6112 13228 6118
rect 13176 6054 13228 6060
rect 13188 5846 13216 6054
rect 13176 5840 13228 5846
rect 12806 5808 12862 5817
rect 13176 5782 13228 5788
rect 12806 5743 12862 5752
rect 13188 5681 13216 5782
rect 13452 5772 13504 5778
rect 13452 5714 13504 5720
rect 13174 5672 13230 5681
rect 13174 5607 13230 5616
rect 13464 5166 13492 5714
rect 13452 5160 13504 5166
rect 13452 5102 13504 5108
rect 13464 5030 13492 5102
rect 13452 5024 13504 5030
rect 13452 4966 13504 4972
rect 12716 4276 12768 4282
rect 12716 4218 12768 4224
rect 12624 4208 12676 4214
rect 12624 4150 12676 4156
rect 13464 4078 13492 4966
rect 13556 4146 13584 6598
rect 13648 5710 13676 18566
rect 13832 17785 13860 19246
rect 14004 19236 14056 19242
rect 14004 19178 14056 19184
rect 13818 17776 13874 17785
rect 13818 17711 13874 17720
rect 13728 17536 13780 17542
rect 13728 17478 13780 17484
rect 13740 14414 13768 17478
rect 13912 16040 13964 16046
rect 13912 15982 13964 15988
rect 13820 15904 13872 15910
rect 13820 15846 13872 15852
rect 13832 15706 13860 15846
rect 13820 15700 13872 15706
rect 13820 15642 13872 15648
rect 13832 15162 13860 15642
rect 13820 15156 13872 15162
rect 13820 15098 13872 15104
rect 13728 14408 13780 14414
rect 13728 14350 13780 14356
rect 13740 14074 13768 14350
rect 13728 14068 13780 14074
rect 13728 14010 13780 14016
rect 13820 13456 13872 13462
rect 13820 13398 13872 13404
rect 13832 12986 13860 13398
rect 13820 12980 13872 12986
rect 13820 12922 13872 12928
rect 13820 12368 13872 12374
rect 13820 12310 13872 12316
rect 13832 11898 13860 12310
rect 13820 11892 13872 11898
rect 13820 11834 13872 11840
rect 13728 9920 13780 9926
rect 13728 9862 13780 9868
rect 13740 9586 13768 9862
rect 13728 9580 13780 9586
rect 13728 9522 13780 9528
rect 13820 9376 13872 9382
rect 13820 9318 13872 9324
rect 13728 9104 13780 9110
rect 13728 9046 13780 9052
rect 13740 8634 13768 9046
rect 13728 8628 13780 8634
rect 13728 8570 13780 8576
rect 13740 8090 13768 8570
rect 13728 8084 13780 8090
rect 13728 8026 13780 8032
rect 13728 6724 13780 6730
rect 13728 6666 13780 6672
rect 13740 6186 13768 6666
rect 13728 6180 13780 6186
rect 13728 6122 13780 6128
rect 13636 5704 13688 5710
rect 13636 5646 13688 5652
rect 13832 4457 13860 9318
rect 13924 7954 13952 15982
rect 14016 11830 14044 19178
rect 14280 19168 14332 19174
rect 14280 19110 14332 19116
rect 14096 17808 14148 17814
rect 14096 17750 14148 17756
rect 14108 16998 14136 17750
rect 14096 16992 14148 16998
rect 14096 16934 14148 16940
rect 14108 15473 14136 16934
rect 14094 15464 14150 15473
rect 14094 15399 14150 15408
rect 14188 14272 14240 14278
rect 14188 14214 14240 14220
rect 14200 13802 14228 14214
rect 14188 13796 14240 13802
rect 14188 13738 14240 13744
rect 14094 12336 14150 12345
rect 14094 12271 14150 12280
rect 14292 12288 14320 19110
rect 14476 18970 14504 20839
rect 15750 19952 15806 19961
rect 15750 19887 15806 19896
rect 15764 19514 15792 19887
rect 15752 19508 15804 19514
rect 15752 19450 15804 19456
rect 15108 19304 15160 19310
rect 15108 19246 15160 19252
rect 14832 19168 14884 19174
rect 14832 19110 14884 19116
rect 14464 18964 14516 18970
rect 14464 18906 14516 18912
rect 14556 18828 14608 18834
rect 14556 18770 14608 18776
rect 14372 18216 14424 18222
rect 14372 18158 14424 18164
rect 14384 17241 14412 18158
rect 14568 18086 14596 18770
rect 14844 18222 14872 19110
rect 14832 18216 14884 18222
rect 14832 18158 14884 18164
rect 14556 18080 14608 18086
rect 14556 18022 14608 18028
rect 14370 17232 14426 17241
rect 14370 17167 14426 17176
rect 14464 17196 14516 17202
rect 14464 17138 14516 17144
rect 14476 16454 14504 17138
rect 14464 16448 14516 16454
rect 14464 16390 14516 16396
rect 14476 16114 14504 16390
rect 14568 16130 14596 18022
rect 14924 17740 14976 17746
rect 14924 17682 14976 17688
rect 14648 17060 14700 17066
rect 14648 17002 14700 17008
rect 14660 16454 14688 17002
rect 14936 16454 14964 17682
rect 15120 17066 15148 19246
rect 15622 19068 15918 19088
rect 15678 19066 15702 19068
rect 15758 19066 15782 19068
rect 15838 19066 15862 19068
rect 15700 19014 15702 19066
rect 15764 19014 15776 19066
rect 15838 19014 15840 19066
rect 15678 19012 15702 19014
rect 15758 19012 15782 19014
rect 15838 19012 15862 19014
rect 15622 18992 15918 19012
rect 15568 18624 15620 18630
rect 15568 18566 15620 18572
rect 15580 18222 15608 18566
rect 15948 18426 15976 21542
rect 18234 21542 18368 21570
rect 18234 21520 18290 21542
rect 17868 19304 17920 19310
rect 17868 19246 17920 19252
rect 17132 19236 17184 19242
rect 17132 19178 17184 19184
rect 16028 18828 16080 18834
rect 16028 18770 16080 18776
rect 16304 18828 16356 18834
rect 16304 18770 16356 18776
rect 15936 18420 15988 18426
rect 15936 18362 15988 18368
rect 15568 18216 15620 18222
rect 15568 18158 15620 18164
rect 15936 18216 15988 18222
rect 15936 18158 15988 18164
rect 15476 18080 15528 18086
rect 15476 18022 15528 18028
rect 15384 17876 15436 17882
rect 15384 17818 15436 17824
rect 15200 17672 15252 17678
rect 15252 17632 15332 17660
rect 15200 17614 15252 17620
rect 15200 17332 15252 17338
rect 15200 17274 15252 17280
rect 15108 17060 15160 17066
rect 15108 17002 15160 17008
rect 14648 16448 14700 16454
rect 14648 16390 14700 16396
rect 14924 16448 14976 16454
rect 14924 16390 14976 16396
rect 14660 16250 14688 16390
rect 14648 16244 14700 16250
rect 14648 16186 14700 16192
rect 14832 16244 14884 16250
rect 14832 16186 14884 16192
rect 14464 16108 14516 16114
rect 14568 16102 14688 16130
rect 14464 16050 14516 16056
rect 14372 15360 14424 15366
rect 14372 15302 14424 15308
rect 14556 15360 14608 15366
rect 14556 15302 14608 15308
rect 14384 14074 14412 15302
rect 14372 14068 14424 14074
rect 14424 14028 14504 14056
rect 14372 14010 14424 14016
rect 14476 13802 14504 14028
rect 14372 13796 14424 13802
rect 14372 13738 14424 13744
rect 14464 13796 14516 13802
rect 14464 13738 14516 13744
rect 14384 13326 14412 13738
rect 14372 13320 14424 13326
rect 14372 13262 14424 13268
rect 14464 12912 14516 12918
rect 14464 12854 14516 12860
rect 14004 11824 14056 11830
rect 14004 11766 14056 11772
rect 14004 11144 14056 11150
rect 14004 11086 14056 11092
rect 14016 10674 14044 11086
rect 14004 10668 14056 10674
rect 14004 10610 14056 10616
rect 14016 10266 14044 10610
rect 14004 10260 14056 10266
rect 14004 10202 14056 10208
rect 14016 9994 14044 10202
rect 14004 9988 14056 9994
rect 14004 9930 14056 9936
rect 14108 9674 14136 12271
rect 14292 12260 14412 12288
rect 14188 12232 14240 12238
rect 14240 12192 14320 12220
rect 14188 12174 14240 12180
rect 14292 11014 14320 12192
rect 14280 11008 14332 11014
rect 14280 10950 14332 10956
rect 14292 10713 14320 10950
rect 14278 10704 14334 10713
rect 14278 10639 14334 10648
rect 14108 9646 14228 9674
rect 14200 9382 14228 9646
rect 14188 9376 14240 9382
rect 14188 9318 14240 9324
rect 13912 7948 13964 7954
rect 13912 7890 13964 7896
rect 14384 7274 14412 12260
rect 14476 11694 14504 12854
rect 14568 12850 14596 15302
rect 14556 12844 14608 12850
rect 14556 12786 14608 12792
rect 14568 12442 14596 12786
rect 14556 12436 14608 12442
rect 14556 12378 14608 12384
rect 14464 11688 14516 11694
rect 14464 11630 14516 11636
rect 14556 11620 14608 11626
rect 14556 11562 14608 11568
rect 14568 11286 14596 11562
rect 14556 11280 14608 11286
rect 14556 11222 14608 11228
rect 14660 10674 14688 16102
rect 14844 16017 14872 16186
rect 14830 16008 14886 16017
rect 14830 15943 14886 15952
rect 14740 15564 14792 15570
rect 14740 15506 14792 15512
rect 14752 14822 14780 15506
rect 14844 15450 14872 15943
rect 14936 15609 14964 16390
rect 15016 15904 15068 15910
rect 15016 15846 15068 15852
rect 14922 15600 14978 15609
rect 14922 15535 14978 15544
rect 14844 15422 14964 15450
rect 14740 14816 14792 14822
rect 14740 14758 14792 14764
rect 14752 13841 14780 14758
rect 14832 14612 14884 14618
rect 14832 14554 14884 14560
rect 14738 13832 14794 13841
rect 14738 13767 14794 13776
rect 14844 12850 14872 14554
rect 14832 12844 14884 12850
rect 14832 12786 14884 12792
rect 14844 12374 14872 12786
rect 14832 12368 14884 12374
rect 14832 12310 14884 12316
rect 14740 11756 14792 11762
rect 14740 11698 14792 11704
rect 14752 11150 14780 11698
rect 14740 11144 14792 11150
rect 14740 11086 14792 11092
rect 14648 10668 14700 10674
rect 14648 10610 14700 10616
rect 14464 10532 14516 10538
rect 14464 10474 14516 10480
rect 14476 9722 14504 10474
rect 14464 9716 14516 9722
rect 14464 9658 14516 9664
rect 14660 9110 14688 10610
rect 14648 9104 14700 9110
rect 14648 9046 14700 9052
rect 14660 8498 14688 9046
rect 14936 8498 14964 15422
rect 15028 14074 15056 15846
rect 15120 15026 15148 17002
rect 15108 15020 15160 15026
rect 15108 14962 15160 14968
rect 15016 14068 15068 14074
rect 15016 14010 15068 14016
rect 15120 13938 15148 14962
rect 15108 13932 15160 13938
rect 15108 13874 15160 13880
rect 15106 13832 15162 13841
rect 15016 13796 15068 13802
rect 15106 13767 15162 13776
rect 15016 13738 15068 13744
rect 15028 9178 15056 13738
rect 15120 10130 15148 13767
rect 15212 11762 15240 17274
rect 15304 16998 15332 17632
rect 15292 16992 15344 16998
rect 15292 16934 15344 16940
rect 15304 15910 15332 16934
rect 15292 15904 15344 15910
rect 15292 15846 15344 15852
rect 15292 14884 15344 14890
rect 15292 14826 15344 14832
rect 15304 14618 15332 14826
rect 15292 14612 15344 14618
rect 15292 14554 15344 14560
rect 15200 11756 15252 11762
rect 15200 11698 15252 11704
rect 15212 11354 15240 11698
rect 15200 11348 15252 11354
rect 15200 11290 15252 11296
rect 15396 11218 15424 17818
rect 15488 16998 15516 18022
rect 15622 17980 15918 18000
rect 15678 17978 15702 17980
rect 15758 17978 15782 17980
rect 15838 17978 15862 17980
rect 15700 17926 15702 17978
rect 15764 17926 15776 17978
rect 15838 17926 15840 17978
rect 15678 17924 15702 17926
rect 15758 17924 15782 17926
rect 15838 17924 15862 17926
rect 15622 17904 15918 17924
rect 15948 17377 15976 18158
rect 16040 17610 16068 18770
rect 16120 18148 16172 18154
rect 16120 18090 16172 18096
rect 16028 17604 16080 17610
rect 16028 17546 16080 17552
rect 15934 17368 15990 17377
rect 15934 17303 15990 17312
rect 15476 16992 15528 16998
rect 15476 16934 15528 16940
rect 15488 14929 15516 16934
rect 15622 16892 15918 16912
rect 15678 16890 15702 16892
rect 15758 16890 15782 16892
rect 15838 16890 15862 16892
rect 15700 16838 15702 16890
rect 15764 16838 15776 16890
rect 15838 16838 15840 16890
rect 15678 16836 15702 16838
rect 15758 16836 15782 16838
rect 15838 16836 15862 16838
rect 15622 16816 15918 16836
rect 15568 16652 15620 16658
rect 15568 16594 15620 16600
rect 15752 16652 15804 16658
rect 15752 16594 15804 16600
rect 15580 16522 15608 16594
rect 15568 16516 15620 16522
rect 15568 16458 15620 16464
rect 15580 16250 15608 16458
rect 15568 16244 15620 16250
rect 15568 16186 15620 16192
rect 15764 16114 15792 16594
rect 15752 16108 15804 16114
rect 15752 16050 15804 16056
rect 15622 15804 15918 15824
rect 15678 15802 15702 15804
rect 15758 15802 15782 15804
rect 15838 15802 15862 15804
rect 15700 15750 15702 15802
rect 15764 15750 15776 15802
rect 15838 15750 15840 15802
rect 15678 15748 15702 15750
rect 15758 15748 15782 15750
rect 15838 15748 15862 15750
rect 15622 15728 15918 15748
rect 15948 15026 15976 17303
rect 15936 15020 15988 15026
rect 15936 14962 15988 14968
rect 15474 14920 15530 14929
rect 15474 14855 15530 14864
rect 15476 14816 15528 14822
rect 15476 14758 15528 14764
rect 15488 14618 15516 14758
rect 15622 14716 15918 14736
rect 15678 14714 15702 14716
rect 15758 14714 15782 14716
rect 15838 14714 15862 14716
rect 15700 14662 15702 14714
rect 15764 14662 15776 14714
rect 15838 14662 15840 14714
rect 15678 14660 15702 14662
rect 15758 14660 15782 14662
rect 15838 14660 15862 14662
rect 15622 14640 15918 14660
rect 16026 14648 16082 14657
rect 15948 14618 16026 14634
rect 15476 14612 15528 14618
rect 15476 14554 15528 14560
rect 15936 14612 16026 14618
rect 15988 14606 16026 14612
rect 16026 14583 16082 14592
rect 15936 14554 15988 14560
rect 15660 14476 15712 14482
rect 15660 14418 15712 14424
rect 15672 14074 15700 14418
rect 15660 14068 15712 14074
rect 15660 14010 15712 14016
rect 15476 13728 15528 13734
rect 15476 13670 15528 13676
rect 15488 13394 15516 13670
rect 15622 13628 15918 13648
rect 15678 13626 15702 13628
rect 15758 13626 15782 13628
rect 15838 13626 15862 13628
rect 15700 13574 15702 13626
rect 15764 13574 15776 13626
rect 15838 13574 15840 13626
rect 15678 13572 15702 13574
rect 15758 13572 15782 13574
rect 15838 13572 15862 13574
rect 15622 13552 15918 13572
rect 15476 13388 15528 13394
rect 15476 13330 15528 13336
rect 15488 12986 15516 13330
rect 16132 13326 16160 18090
rect 16316 18086 16344 18770
rect 16488 18760 16540 18766
rect 16488 18702 16540 18708
rect 16396 18148 16448 18154
rect 16396 18090 16448 18096
rect 16304 18080 16356 18086
rect 16304 18022 16356 18028
rect 16304 17876 16356 17882
rect 16304 17818 16356 17824
rect 16212 17128 16264 17134
rect 16212 17070 16264 17076
rect 16224 16794 16252 17070
rect 16212 16788 16264 16794
rect 16212 16730 16264 16736
rect 16224 16046 16252 16730
rect 16212 16040 16264 16046
rect 16212 15982 16264 15988
rect 16224 15706 16252 15982
rect 16212 15700 16264 15706
rect 16212 15642 16264 15648
rect 16212 14408 16264 14414
rect 16212 14350 16264 14356
rect 16224 13938 16252 14350
rect 16212 13932 16264 13938
rect 16212 13874 16264 13880
rect 16316 13530 16344 17818
rect 16408 14482 16436 18090
rect 16500 14482 16528 18702
rect 16948 18692 17000 18698
rect 16948 18634 17000 18640
rect 16580 17060 16632 17066
rect 16580 17002 16632 17008
rect 16592 15570 16620 17002
rect 16672 15972 16724 15978
rect 16672 15914 16724 15920
rect 16580 15564 16632 15570
rect 16580 15506 16632 15512
rect 16592 15162 16620 15506
rect 16580 15156 16632 15162
rect 16580 15098 16632 15104
rect 16396 14476 16448 14482
rect 16396 14418 16448 14424
rect 16488 14476 16540 14482
rect 16488 14418 16540 14424
rect 16580 13796 16632 13802
rect 16580 13738 16632 13744
rect 16304 13524 16356 13530
rect 16304 13466 16356 13472
rect 16028 13320 16080 13326
rect 16028 13262 16080 13268
rect 16120 13320 16172 13326
rect 16120 13262 16172 13268
rect 15476 12980 15528 12986
rect 15476 12922 15528 12928
rect 15936 12640 15988 12646
rect 15936 12582 15988 12588
rect 15622 12540 15918 12560
rect 15678 12538 15702 12540
rect 15758 12538 15782 12540
rect 15838 12538 15862 12540
rect 15700 12486 15702 12538
rect 15764 12486 15776 12538
rect 15838 12486 15840 12538
rect 15678 12484 15702 12486
rect 15758 12484 15782 12486
rect 15838 12484 15862 12486
rect 15622 12464 15918 12484
rect 15476 12368 15528 12374
rect 15476 12310 15528 12316
rect 15488 11898 15516 12310
rect 15948 12084 15976 12582
rect 16040 12374 16068 13262
rect 16212 13252 16264 13258
rect 16212 13194 16264 13200
rect 16028 12368 16080 12374
rect 16028 12310 16080 12316
rect 16028 12096 16080 12102
rect 15948 12056 16028 12084
rect 16028 12038 16080 12044
rect 15476 11892 15528 11898
rect 15476 11834 15528 11840
rect 15622 11452 15918 11472
rect 15678 11450 15702 11452
rect 15758 11450 15782 11452
rect 15838 11450 15862 11452
rect 15700 11398 15702 11450
rect 15764 11398 15776 11450
rect 15838 11398 15840 11450
rect 15678 11396 15702 11398
rect 15758 11396 15782 11398
rect 15838 11396 15862 11398
rect 15622 11376 15918 11396
rect 16040 11286 16068 12038
rect 16224 11762 16252 13194
rect 16316 12850 16344 13466
rect 16592 13462 16620 13738
rect 16396 13456 16448 13462
rect 16396 13398 16448 13404
rect 16580 13456 16632 13462
rect 16580 13398 16632 13404
rect 16684 13410 16712 15914
rect 16854 15056 16910 15065
rect 16854 14991 16910 15000
rect 16868 14958 16896 14991
rect 16856 14952 16908 14958
rect 16856 14894 16908 14900
rect 16764 14476 16816 14482
rect 16764 14418 16816 14424
rect 16776 13530 16804 14418
rect 16960 13814 16988 18634
rect 17038 15464 17094 15473
rect 17038 15399 17094 15408
rect 17052 15162 17080 15399
rect 17040 15156 17092 15162
rect 17040 15098 17092 15104
rect 17040 15020 17092 15026
rect 17040 14962 17092 14968
rect 16868 13786 16988 13814
rect 16764 13524 16816 13530
rect 16764 13466 16816 13472
rect 16304 12844 16356 12850
rect 16304 12786 16356 12792
rect 16408 12714 16436 13398
rect 16684 13382 16804 13410
rect 16672 13320 16724 13326
rect 16672 13262 16724 13268
rect 16488 13184 16540 13190
rect 16488 13126 16540 13132
rect 16580 13184 16632 13190
rect 16580 13126 16632 13132
rect 16396 12708 16448 12714
rect 16396 12650 16448 12656
rect 16500 12238 16528 13126
rect 16488 12232 16540 12238
rect 16488 12174 16540 12180
rect 16212 11756 16264 11762
rect 16212 11698 16264 11704
rect 16592 11626 16620 13126
rect 16684 12442 16712 13262
rect 16672 12436 16724 12442
rect 16672 12378 16724 12384
rect 16776 12306 16804 13382
rect 16764 12300 16816 12306
rect 16764 12242 16816 12248
rect 16868 11762 16896 13786
rect 17052 12753 17080 14962
rect 17144 13814 17172 19178
rect 17880 19174 17908 19246
rect 17592 19168 17644 19174
rect 17592 19110 17644 19116
rect 17868 19168 17920 19174
rect 17868 19110 17920 19116
rect 18144 19168 18196 19174
rect 18144 19110 18196 19116
rect 17500 18828 17552 18834
rect 17500 18770 17552 18776
rect 17512 18154 17540 18770
rect 17500 18148 17552 18154
rect 17500 18090 17552 18096
rect 17224 17740 17276 17746
rect 17224 17682 17276 17688
rect 17316 17740 17368 17746
rect 17316 17682 17368 17688
rect 17236 17338 17264 17682
rect 17224 17332 17276 17338
rect 17224 17274 17276 17280
rect 17328 16998 17356 17682
rect 17316 16992 17368 16998
rect 17316 16934 17368 16940
rect 17500 16788 17552 16794
rect 17500 16730 17552 16736
rect 17512 16250 17540 16730
rect 17500 16244 17552 16250
rect 17500 16186 17552 16192
rect 17316 16108 17368 16114
rect 17316 16050 17368 16056
rect 17224 15088 17276 15094
rect 17224 15030 17276 15036
rect 17236 14550 17264 15030
rect 17224 14544 17276 14550
rect 17224 14486 17276 14492
rect 17236 14006 17264 14486
rect 17224 14000 17276 14006
rect 17224 13942 17276 13948
rect 17144 13786 17264 13814
rect 17038 12744 17094 12753
rect 17038 12679 17094 12688
rect 16856 11756 16908 11762
rect 16856 11698 16908 11704
rect 16580 11620 16632 11626
rect 16580 11562 16632 11568
rect 16394 11384 16450 11393
rect 16868 11354 16896 11698
rect 16394 11319 16450 11328
rect 16856 11348 16908 11354
rect 16028 11280 16080 11286
rect 16028 11222 16080 11228
rect 15384 11212 15436 11218
rect 15384 11154 15436 11160
rect 15396 10266 15424 11154
rect 15934 10568 15990 10577
rect 15934 10503 15990 10512
rect 15474 10432 15530 10441
rect 15474 10367 15530 10376
rect 15384 10260 15436 10266
rect 15384 10202 15436 10208
rect 15108 10124 15160 10130
rect 15108 10066 15160 10072
rect 15120 9722 15148 10066
rect 15108 9716 15160 9722
rect 15108 9658 15160 9664
rect 15016 9172 15068 9178
rect 15016 9114 15068 9120
rect 15488 9042 15516 10367
rect 15622 10364 15918 10384
rect 15678 10362 15702 10364
rect 15758 10362 15782 10364
rect 15838 10362 15862 10364
rect 15700 10310 15702 10362
rect 15764 10310 15776 10362
rect 15838 10310 15840 10362
rect 15678 10308 15702 10310
rect 15758 10308 15782 10310
rect 15838 10308 15862 10310
rect 15622 10288 15918 10308
rect 15948 9994 15976 10503
rect 16040 10470 16068 11222
rect 16304 11008 16356 11014
rect 16304 10950 16356 10956
rect 16316 10810 16344 10950
rect 16304 10804 16356 10810
rect 16304 10746 16356 10752
rect 16316 10538 16344 10746
rect 16304 10532 16356 10538
rect 16304 10474 16356 10480
rect 16028 10464 16080 10470
rect 16028 10406 16080 10412
rect 16408 10169 16436 11319
rect 16856 11290 16908 11296
rect 17052 11234 17080 12679
rect 16868 11206 17080 11234
rect 16488 11144 16540 11150
rect 16488 11086 16540 11092
rect 16500 10674 16528 11086
rect 16488 10668 16540 10674
rect 16488 10610 16540 10616
rect 16394 10160 16450 10169
rect 16394 10095 16450 10104
rect 16304 10056 16356 10062
rect 16304 9998 16356 10004
rect 15936 9988 15988 9994
rect 15936 9930 15988 9936
rect 16316 9722 16344 9998
rect 16488 9920 16540 9926
rect 16488 9862 16540 9868
rect 16028 9716 16080 9722
rect 16028 9658 16080 9664
rect 16304 9716 16356 9722
rect 16304 9658 16356 9664
rect 15622 9276 15918 9296
rect 15678 9274 15702 9276
rect 15758 9274 15782 9276
rect 15838 9274 15862 9276
rect 15700 9222 15702 9274
rect 15764 9222 15776 9274
rect 15838 9222 15840 9274
rect 15678 9220 15702 9222
rect 15758 9220 15782 9222
rect 15838 9220 15862 9222
rect 15622 9200 15918 9220
rect 15476 9036 15528 9042
rect 15476 8978 15528 8984
rect 15488 8634 15516 8978
rect 15476 8628 15528 8634
rect 15476 8570 15528 8576
rect 14648 8492 14700 8498
rect 14648 8434 14700 8440
rect 14924 8492 14976 8498
rect 14924 8434 14976 8440
rect 15292 8424 15344 8430
rect 15292 8366 15344 8372
rect 14648 8356 14700 8362
rect 14648 8298 14700 8304
rect 14660 7750 14688 8298
rect 14648 7744 14700 7750
rect 14648 7686 14700 7692
rect 14660 7546 14688 7686
rect 14648 7540 14700 7546
rect 14648 7482 14700 7488
rect 14372 7268 14424 7274
rect 14372 7210 14424 7216
rect 15016 6792 15068 6798
rect 15016 6734 15068 6740
rect 15028 6322 15056 6734
rect 15016 6316 15068 6322
rect 15016 6258 15068 6264
rect 15028 6225 15056 6258
rect 15108 6248 15160 6254
rect 15014 6216 15070 6225
rect 14188 6180 14240 6186
rect 15108 6190 15160 6196
rect 15014 6151 15070 6160
rect 14188 6122 14240 6128
rect 14200 5914 14228 6122
rect 14188 5908 14240 5914
rect 14188 5850 14240 5856
rect 14832 4684 14884 4690
rect 14832 4626 14884 4632
rect 14372 4616 14424 4622
rect 14372 4558 14424 4564
rect 13818 4448 13874 4457
rect 13818 4383 13874 4392
rect 14384 4282 14412 4558
rect 14372 4276 14424 4282
rect 14372 4218 14424 4224
rect 14844 4214 14872 4626
rect 14832 4208 14884 4214
rect 14832 4150 14884 4156
rect 13544 4140 13596 4146
rect 13544 4082 13596 4088
rect 13452 4072 13504 4078
rect 13450 4040 13452 4049
rect 13504 4040 13506 4049
rect 12532 4004 12584 4010
rect 13450 3975 13506 3984
rect 12532 3946 12584 3952
rect 13464 3949 13492 3975
rect 12544 3738 12572 3946
rect 12624 3936 12676 3942
rect 12624 3878 12676 3884
rect 12532 3732 12584 3738
rect 12532 3674 12584 3680
rect 12440 3596 12492 3602
rect 12440 3538 12492 3544
rect 12452 3505 12480 3538
rect 12636 3534 12664 3878
rect 13176 3596 13228 3602
rect 13176 3538 13228 3544
rect 13360 3596 13412 3602
rect 13360 3538 13412 3544
rect 12624 3528 12676 3534
rect 12438 3496 12494 3505
rect 12348 3460 12400 3466
rect 12624 3470 12676 3476
rect 12438 3431 12494 3440
rect 12348 3402 12400 3408
rect 11956 3292 12252 3312
rect 12012 3290 12036 3292
rect 12092 3290 12116 3292
rect 12172 3290 12196 3292
rect 12034 3238 12036 3290
rect 12098 3238 12110 3290
rect 12172 3238 12174 3290
rect 12012 3236 12036 3238
rect 12092 3236 12116 3238
rect 12172 3236 12196 3238
rect 11956 3216 12252 3236
rect 12360 3194 12388 3402
rect 12636 3194 12664 3470
rect 12348 3188 12400 3194
rect 12348 3130 12400 3136
rect 12624 3188 12676 3194
rect 12624 3130 12676 3136
rect 13188 2990 13216 3538
rect 13372 3126 13400 3538
rect 13360 3120 13412 3126
rect 13360 3062 13412 3068
rect 11888 2984 11940 2990
rect 11888 2926 11940 2932
rect 13176 2984 13228 2990
rect 13176 2926 13228 2932
rect 11900 2854 11928 2926
rect 11888 2848 11940 2854
rect 11888 2790 11940 2796
rect 11428 2508 11480 2514
rect 11428 2450 11480 2456
rect 11900 2009 11928 2790
rect 13188 2650 13216 2926
rect 13556 2666 13584 4082
rect 13912 4072 13964 4078
rect 13912 4014 13964 4020
rect 13924 3738 13952 4014
rect 14924 4004 14976 4010
rect 14924 3946 14976 3952
rect 13912 3732 13964 3738
rect 13912 3674 13964 3680
rect 14280 3596 14332 3602
rect 14280 3538 14332 3544
rect 13636 3528 13688 3534
rect 13636 3470 13688 3476
rect 13648 2990 13676 3470
rect 14292 3194 14320 3538
rect 14556 3528 14608 3534
rect 14556 3470 14608 3476
rect 14280 3188 14332 3194
rect 14280 3130 14332 3136
rect 13636 2984 13688 2990
rect 13636 2926 13688 2932
rect 14280 2848 14332 2854
rect 14280 2790 14332 2796
rect 13556 2650 13860 2666
rect 14292 2650 14320 2790
rect 13176 2644 13228 2650
rect 13176 2586 13228 2592
rect 13544 2644 13860 2650
rect 13596 2638 13860 2644
rect 13544 2586 13596 2592
rect 13832 2582 13860 2638
rect 14280 2644 14332 2650
rect 14280 2586 14332 2592
rect 13820 2576 13872 2582
rect 13820 2518 13872 2524
rect 12440 2508 12492 2514
rect 12440 2450 12492 2456
rect 11956 2204 12252 2224
rect 12012 2202 12036 2204
rect 12092 2202 12116 2204
rect 12172 2202 12196 2204
rect 12034 2150 12036 2202
rect 12098 2150 12110 2202
rect 12172 2150 12174 2202
rect 12012 2148 12036 2150
rect 12092 2148 12116 2150
rect 12172 2148 12196 2150
rect 11956 2128 12252 2148
rect 12452 2106 12480 2450
rect 14568 2310 14596 3470
rect 14936 3398 14964 3946
rect 14924 3392 14976 3398
rect 14924 3334 14976 3340
rect 14936 3097 14964 3334
rect 15120 3097 15148 6190
rect 15304 4554 15332 8366
rect 15622 8188 15918 8208
rect 15678 8186 15702 8188
rect 15758 8186 15782 8188
rect 15838 8186 15862 8188
rect 15700 8134 15702 8186
rect 15764 8134 15776 8186
rect 15838 8134 15840 8186
rect 15678 8132 15702 8134
rect 15758 8132 15782 8134
rect 15838 8132 15862 8134
rect 15622 8112 15918 8132
rect 15384 8084 15436 8090
rect 15384 8026 15436 8032
rect 15396 7546 15424 8026
rect 15384 7540 15436 7546
rect 15384 7482 15436 7488
rect 15476 7472 15528 7478
rect 15476 7414 15528 7420
rect 15488 6934 15516 7414
rect 15622 7100 15918 7120
rect 15678 7098 15702 7100
rect 15758 7098 15782 7100
rect 15838 7098 15862 7100
rect 15700 7046 15702 7098
rect 15764 7046 15776 7098
rect 15838 7046 15840 7098
rect 15678 7044 15702 7046
rect 15758 7044 15782 7046
rect 15838 7044 15862 7046
rect 15622 7024 15918 7044
rect 15476 6928 15528 6934
rect 15476 6870 15528 6876
rect 15488 6458 15516 6870
rect 15476 6452 15528 6458
rect 15476 6394 15528 6400
rect 16040 6390 16068 9658
rect 16212 8832 16264 8838
rect 16212 8774 16264 8780
rect 16224 8430 16252 8774
rect 16212 8424 16264 8430
rect 16212 8366 16264 8372
rect 16120 7948 16172 7954
rect 16120 7890 16172 7896
rect 16132 7546 16160 7890
rect 16120 7540 16172 7546
rect 16120 7482 16172 7488
rect 16028 6384 16080 6390
rect 16028 6326 16080 6332
rect 16316 6322 16344 9658
rect 16500 9450 16528 9862
rect 16580 9648 16632 9654
rect 16580 9590 16632 9596
rect 16592 9450 16620 9590
rect 16488 9444 16540 9450
rect 16488 9386 16540 9392
rect 16580 9444 16632 9450
rect 16580 9386 16632 9392
rect 16396 9172 16448 9178
rect 16396 9114 16448 9120
rect 16408 8430 16436 9114
rect 16500 9042 16528 9386
rect 16488 9036 16540 9042
rect 16488 8978 16540 8984
rect 16396 8424 16448 8430
rect 16396 8366 16448 8372
rect 16408 7954 16436 8366
rect 16580 8016 16632 8022
rect 16580 7958 16632 7964
rect 16396 7948 16448 7954
rect 16396 7890 16448 7896
rect 16408 7478 16436 7890
rect 16396 7472 16448 7478
rect 16396 7414 16448 7420
rect 16488 7404 16540 7410
rect 16488 7346 16540 7352
rect 16500 7002 16528 7346
rect 16592 7274 16620 7958
rect 16672 7472 16724 7478
rect 16672 7414 16724 7420
rect 16580 7268 16632 7274
rect 16580 7210 16632 7216
rect 16592 7002 16620 7210
rect 16488 6996 16540 7002
rect 16488 6938 16540 6944
rect 16580 6996 16632 7002
rect 16580 6938 16632 6944
rect 16580 6860 16632 6866
rect 16580 6802 16632 6808
rect 16304 6316 16356 6322
rect 16304 6258 16356 6264
rect 15476 6248 15528 6254
rect 15476 6190 15528 6196
rect 15488 5642 15516 6190
rect 16592 6118 16620 6802
rect 16580 6112 16632 6118
rect 16580 6054 16632 6060
rect 15622 6012 15918 6032
rect 15678 6010 15702 6012
rect 15758 6010 15782 6012
rect 15838 6010 15862 6012
rect 15700 5958 15702 6010
rect 15764 5958 15776 6010
rect 15838 5958 15840 6010
rect 15678 5956 15702 5958
rect 15758 5956 15782 5958
rect 15838 5956 15862 5958
rect 15622 5936 15918 5956
rect 16120 5840 16172 5846
rect 16120 5782 16172 5788
rect 15476 5636 15528 5642
rect 15476 5578 15528 5584
rect 16132 5370 16160 5782
rect 16120 5364 16172 5370
rect 16120 5306 16172 5312
rect 15476 5160 15528 5166
rect 15476 5102 15528 5108
rect 15488 4729 15516 5102
rect 16592 5098 16620 6054
rect 16684 5846 16712 7414
rect 16672 5840 16724 5846
rect 16672 5782 16724 5788
rect 16684 5234 16712 5782
rect 16764 5636 16816 5642
rect 16764 5578 16816 5584
rect 16776 5302 16804 5578
rect 16764 5296 16816 5302
rect 16764 5238 16816 5244
rect 16672 5228 16724 5234
rect 16672 5170 16724 5176
rect 16580 5092 16632 5098
rect 16580 5034 16632 5040
rect 16764 5092 16816 5098
rect 16764 5034 16816 5040
rect 15622 4924 15918 4944
rect 15678 4922 15702 4924
rect 15758 4922 15782 4924
rect 15838 4922 15862 4924
rect 15700 4870 15702 4922
rect 15764 4870 15776 4922
rect 15838 4870 15840 4922
rect 15678 4868 15702 4870
rect 15758 4868 15782 4870
rect 15838 4868 15862 4870
rect 15622 4848 15918 4868
rect 16776 4758 16804 5034
rect 16764 4752 16816 4758
rect 15474 4720 15530 4729
rect 16764 4694 16816 4700
rect 15474 4655 15530 4664
rect 15384 4616 15436 4622
rect 15384 4558 15436 4564
rect 15292 4548 15344 4554
rect 15292 4490 15344 4496
rect 15396 3913 15424 4558
rect 15488 4554 15516 4655
rect 16028 4616 16080 4622
rect 16028 4558 16080 4564
rect 15476 4548 15528 4554
rect 15476 4490 15528 4496
rect 15934 4448 15990 4457
rect 15934 4383 15990 4392
rect 15844 4276 15896 4282
rect 15844 4218 15896 4224
rect 15856 4010 15884 4218
rect 15844 4004 15896 4010
rect 15844 3946 15896 3952
rect 15382 3904 15438 3913
rect 15382 3839 15438 3848
rect 15396 3738 15424 3839
rect 15622 3836 15918 3856
rect 15678 3834 15702 3836
rect 15758 3834 15782 3836
rect 15838 3834 15862 3836
rect 15700 3782 15702 3834
rect 15764 3782 15776 3834
rect 15838 3782 15840 3834
rect 15678 3780 15702 3782
rect 15758 3780 15782 3782
rect 15838 3780 15862 3782
rect 15622 3760 15918 3780
rect 15384 3732 15436 3738
rect 15384 3674 15436 3680
rect 15844 3664 15896 3670
rect 15844 3606 15896 3612
rect 15856 3534 15884 3606
rect 15844 3528 15896 3534
rect 15844 3470 15896 3476
rect 15856 3194 15884 3470
rect 15844 3188 15896 3194
rect 15844 3130 15896 3136
rect 14922 3088 14978 3097
rect 14922 3023 14978 3032
rect 15106 3088 15162 3097
rect 15106 3023 15162 3032
rect 15622 2748 15918 2768
rect 15678 2746 15702 2748
rect 15758 2746 15782 2748
rect 15838 2746 15862 2748
rect 15700 2694 15702 2746
rect 15764 2694 15776 2746
rect 15838 2694 15840 2746
rect 15678 2692 15702 2694
rect 15758 2692 15782 2694
rect 15838 2692 15862 2694
rect 15622 2672 15918 2692
rect 15948 2514 15976 4383
rect 16040 4010 16068 4558
rect 16028 4004 16080 4010
rect 16028 3946 16080 3952
rect 16396 4004 16448 4010
rect 16396 3946 16448 3952
rect 16408 3738 16436 3946
rect 16776 3942 16804 4694
rect 16764 3936 16816 3942
rect 16764 3878 16816 3884
rect 16396 3732 16448 3738
rect 16396 3674 16448 3680
rect 16396 3596 16448 3602
rect 16396 3538 16448 3544
rect 16212 3528 16264 3534
rect 16212 3470 16264 3476
rect 16224 2922 16252 3470
rect 16408 3058 16436 3538
rect 16868 3466 16896 11206
rect 17132 10532 17184 10538
rect 17132 10474 17184 10480
rect 16948 10464 17000 10470
rect 16948 10406 17000 10412
rect 16960 10198 16988 10406
rect 16948 10192 17000 10198
rect 16948 10134 17000 10140
rect 16960 9586 16988 10134
rect 17144 9586 17172 10474
rect 16948 9580 17000 9586
rect 16948 9522 17000 9528
rect 17132 9580 17184 9586
rect 17132 9522 17184 9528
rect 16960 9178 16988 9522
rect 16948 9172 17000 9178
rect 16948 9114 17000 9120
rect 16960 8294 16988 9114
rect 16948 8288 17000 8294
rect 16948 8230 17000 8236
rect 16960 6866 16988 8230
rect 17132 7880 17184 7886
rect 17130 7848 17132 7857
rect 17184 7848 17186 7857
rect 17130 7783 17186 7792
rect 17144 7750 17172 7783
rect 17132 7744 17184 7750
rect 17132 7686 17184 7692
rect 17040 7200 17092 7206
rect 17040 7142 17092 7148
rect 17052 7002 17080 7142
rect 17040 6996 17092 7002
rect 17040 6938 17092 6944
rect 16948 6860 17000 6866
rect 16948 6802 17000 6808
rect 16948 5704 17000 5710
rect 16948 5646 17000 5652
rect 16960 5302 16988 5646
rect 16948 5296 17000 5302
rect 16948 5238 17000 5244
rect 17132 4616 17184 4622
rect 17132 4558 17184 4564
rect 17144 3942 17172 4558
rect 16948 3936 17000 3942
rect 16948 3878 17000 3884
rect 17132 3936 17184 3942
rect 17132 3878 17184 3884
rect 16764 3460 16816 3466
rect 16764 3402 16816 3408
rect 16856 3460 16908 3466
rect 16856 3402 16908 3408
rect 16396 3052 16448 3058
rect 16396 2994 16448 3000
rect 16776 2990 16804 3402
rect 16764 2984 16816 2990
rect 16764 2926 16816 2932
rect 16212 2916 16264 2922
rect 16212 2858 16264 2864
rect 16960 2582 16988 3878
rect 17144 3233 17172 3878
rect 17236 3670 17264 13786
rect 17328 8106 17356 16050
rect 17408 15904 17460 15910
rect 17408 15846 17460 15852
rect 17420 13394 17448 15846
rect 17512 14074 17540 16186
rect 17500 14068 17552 14074
rect 17500 14010 17552 14016
rect 17408 13388 17460 13394
rect 17408 13330 17460 13336
rect 17408 12436 17460 12442
rect 17408 12378 17460 12384
rect 17420 11558 17448 12378
rect 17408 11552 17460 11558
rect 17408 11494 17460 11500
rect 17420 11286 17448 11494
rect 17408 11280 17460 11286
rect 17408 11222 17460 11228
rect 17604 9586 17632 19110
rect 17776 17536 17828 17542
rect 17776 17478 17828 17484
rect 17788 17134 17816 17478
rect 17880 17202 17908 19110
rect 17960 18624 18012 18630
rect 17960 18566 18012 18572
rect 17868 17196 17920 17202
rect 17868 17138 17920 17144
rect 17776 17128 17828 17134
rect 17776 17070 17828 17076
rect 17788 16726 17816 17070
rect 17868 16992 17920 16998
rect 17868 16934 17920 16940
rect 17776 16720 17828 16726
rect 17776 16662 17828 16668
rect 17776 16584 17828 16590
rect 17776 16526 17828 16532
rect 17788 16250 17816 16526
rect 17776 16244 17828 16250
rect 17776 16186 17828 16192
rect 17880 14414 17908 16934
rect 17972 16726 18000 18566
rect 17960 16720 18012 16726
rect 17960 16662 18012 16668
rect 17972 16046 18000 16662
rect 17960 16040 18012 16046
rect 17960 15982 18012 15988
rect 17868 14408 17920 14414
rect 17868 14350 17920 14356
rect 18156 13938 18184 19110
rect 18340 18426 18368 21542
rect 20456 21542 20774 21570
rect 19289 19612 19585 19632
rect 19345 19610 19369 19612
rect 19425 19610 19449 19612
rect 19505 19610 19529 19612
rect 19367 19558 19369 19610
rect 19431 19558 19443 19610
rect 19505 19558 19507 19610
rect 19345 19556 19369 19558
rect 19425 19556 19449 19558
rect 19505 19556 19529 19558
rect 19289 19536 19585 19556
rect 19800 19168 19852 19174
rect 19800 19110 19852 19116
rect 18604 18828 18656 18834
rect 18604 18770 18656 18776
rect 18328 18420 18380 18426
rect 18328 18362 18380 18368
rect 18616 18358 18644 18770
rect 19289 18524 19585 18544
rect 19345 18522 19369 18524
rect 19425 18522 19449 18524
rect 19505 18522 19529 18524
rect 19367 18470 19369 18522
rect 19431 18470 19443 18522
rect 19505 18470 19507 18522
rect 19345 18468 19369 18470
rect 19425 18468 19449 18470
rect 19505 18468 19529 18470
rect 19289 18448 19585 18468
rect 18604 18352 18656 18358
rect 18604 18294 18656 18300
rect 18420 18080 18472 18086
rect 18420 18022 18472 18028
rect 19156 18080 19208 18086
rect 19156 18022 19208 18028
rect 19616 18080 19668 18086
rect 19616 18022 19668 18028
rect 18328 16108 18380 16114
rect 18328 16050 18380 16056
rect 18236 15972 18288 15978
rect 18236 15914 18288 15920
rect 18248 15706 18276 15914
rect 18236 15700 18288 15706
rect 18236 15642 18288 15648
rect 18144 13932 18196 13938
rect 18144 13874 18196 13880
rect 18156 13530 18184 13874
rect 18144 13524 18196 13530
rect 18144 13466 18196 13472
rect 18340 13326 18368 16050
rect 18432 13814 18460 18022
rect 18512 17876 18564 17882
rect 18512 17818 18564 17824
rect 18524 15570 18552 17818
rect 18696 17740 18748 17746
rect 18696 17682 18748 17688
rect 18880 17740 18932 17746
rect 18880 17682 18932 17688
rect 18708 16794 18736 17682
rect 18892 17134 18920 17682
rect 18880 17128 18932 17134
rect 18880 17070 18932 17076
rect 18696 16788 18748 16794
rect 18696 16730 18748 16736
rect 18604 16584 18656 16590
rect 18604 16526 18656 16532
rect 18512 15564 18564 15570
rect 18512 15506 18564 15512
rect 18524 15162 18552 15506
rect 18512 15156 18564 15162
rect 18512 15098 18564 15104
rect 18616 14550 18644 16526
rect 18708 16522 18736 16730
rect 18696 16516 18748 16522
rect 18696 16458 18748 16464
rect 19064 16176 19116 16182
rect 19064 16118 19116 16124
rect 18880 16040 18932 16046
rect 18880 15982 18932 15988
rect 18788 15700 18840 15706
rect 18788 15642 18840 15648
rect 18696 15360 18748 15366
rect 18696 15302 18748 15308
rect 18708 14890 18736 15302
rect 18800 15094 18828 15642
rect 18788 15088 18840 15094
rect 18788 15030 18840 15036
rect 18696 14884 18748 14890
rect 18696 14826 18748 14832
rect 18604 14544 18656 14550
rect 18604 14486 18656 14492
rect 18432 13786 18552 13814
rect 18420 13456 18472 13462
rect 18420 13398 18472 13404
rect 18328 13320 18380 13326
rect 18328 13262 18380 13268
rect 18052 12980 18104 12986
rect 18052 12922 18104 12928
rect 17776 12300 17828 12306
rect 17776 12242 17828 12248
rect 17788 11898 17816 12242
rect 17776 11892 17828 11898
rect 17776 11834 17828 11840
rect 17684 11144 17736 11150
rect 17684 11086 17736 11092
rect 17696 10470 17724 11086
rect 17684 10464 17736 10470
rect 17684 10406 17736 10412
rect 17592 9580 17644 9586
rect 17592 9522 17644 9528
rect 17500 9376 17552 9382
rect 17500 9318 17552 9324
rect 17512 9178 17540 9318
rect 17500 9172 17552 9178
rect 17500 9114 17552 9120
rect 17408 8968 17460 8974
rect 17408 8910 17460 8916
rect 17420 8294 17448 8910
rect 17512 8634 17540 9114
rect 17592 9036 17644 9042
rect 17592 8978 17644 8984
rect 17500 8628 17552 8634
rect 17500 8570 17552 8576
rect 17408 8288 17460 8294
rect 17408 8230 17460 8236
rect 17328 8078 17448 8106
rect 17316 6656 17368 6662
rect 17316 6598 17368 6604
rect 17328 5137 17356 6598
rect 17420 5914 17448 8078
rect 17500 8016 17552 8022
rect 17500 7958 17552 7964
rect 17512 7546 17540 7958
rect 17604 7546 17632 8978
rect 17696 8498 17724 10406
rect 17776 10192 17828 10198
rect 17776 10134 17828 10140
rect 17788 9722 17816 10134
rect 17776 9716 17828 9722
rect 17776 9658 17828 9664
rect 17788 9450 17816 9658
rect 17776 9444 17828 9450
rect 17776 9386 17828 9392
rect 17684 8492 17736 8498
rect 17684 8434 17736 8440
rect 17500 7540 17552 7546
rect 17500 7482 17552 7488
rect 17592 7540 17644 7546
rect 17592 7482 17644 7488
rect 18064 6866 18092 12922
rect 18340 12442 18368 13262
rect 18432 12782 18460 13398
rect 18420 12776 18472 12782
rect 18420 12718 18472 12724
rect 18328 12436 18380 12442
rect 18328 12378 18380 12384
rect 18524 11914 18552 13786
rect 18616 13326 18644 14486
rect 18892 13814 18920 15982
rect 19076 15094 19104 16118
rect 19064 15088 19116 15094
rect 19064 15030 19116 15036
rect 18972 15020 19024 15026
rect 18972 14962 19024 14968
rect 18708 13786 18920 13814
rect 18604 13320 18656 13326
rect 18604 13262 18656 13268
rect 18708 12986 18736 13786
rect 18880 13728 18932 13734
rect 18984 13716 19012 14962
rect 19064 14544 19116 14550
rect 19064 14486 19116 14492
rect 19076 14074 19104 14486
rect 19064 14068 19116 14074
rect 19064 14010 19116 14016
rect 18932 13688 19012 13716
rect 18880 13670 18932 13676
rect 18696 12980 18748 12986
rect 18696 12922 18748 12928
rect 18788 12912 18840 12918
rect 18788 12854 18840 12860
rect 18800 12442 18828 12854
rect 18892 12850 18920 13670
rect 19168 12918 19196 18022
rect 19289 17436 19585 17456
rect 19345 17434 19369 17436
rect 19425 17434 19449 17436
rect 19505 17434 19529 17436
rect 19367 17382 19369 17434
rect 19431 17382 19443 17434
rect 19505 17382 19507 17434
rect 19345 17380 19369 17382
rect 19425 17380 19449 17382
rect 19505 17380 19529 17382
rect 19289 17360 19585 17380
rect 19628 16658 19656 18022
rect 19616 16652 19668 16658
rect 19616 16594 19668 16600
rect 19289 16348 19585 16368
rect 19345 16346 19369 16348
rect 19425 16346 19449 16348
rect 19505 16346 19529 16348
rect 19367 16294 19369 16346
rect 19431 16294 19443 16346
rect 19505 16294 19507 16346
rect 19345 16292 19369 16294
rect 19425 16292 19449 16294
rect 19505 16292 19529 16294
rect 19289 16272 19585 16292
rect 19628 15910 19656 16594
rect 19616 15904 19668 15910
rect 19616 15846 19668 15852
rect 19289 15260 19585 15280
rect 19345 15258 19369 15260
rect 19425 15258 19449 15260
rect 19505 15258 19529 15260
rect 19367 15206 19369 15258
rect 19431 15206 19443 15258
rect 19505 15206 19507 15258
rect 19345 15204 19369 15206
rect 19425 15204 19449 15206
rect 19505 15204 19529 15206
rect 19289 15184 19585 15204
rect 19248 15088 19300 15094
rect 19248 15030 19300 15036
rect 19260 14550 19288 15030
rect 19248 14544 19300 14550
rect 19248 14486 19300 14492
rect 19289 14172 19585 14192
rect 19345 14170 19369 14172
rect 19425 14170 19449 14172
rect 19505 14170 19529 14172
rect 19367 14118 19369 14170
rect 19431 14118 19443 14170
rect 19505 14118 19507 14170
rect 19345 14116 19369 14118
rect 19425 14116 19449 14118
rect 19505 14116 19529 14118
rect 19289 14096 19585 14116
rect 19616 14000 19668 14006
rect 19616 13942 19668 13948
rect 19628 13870 19656 13942
rect 19628 13864 19703 13870
rect 19628 13812 19651 13864
rect 19812 13841 19840 19110
rect 19890 19000 19946 19009
rect 19890 18935 19946 18944
rect 19904 14074 19932 18935
rect 19984 18828 20036 18834
rect 19984 18770 20036 18776
rect 19996 18426 20024 18770
rect 19984 18420 20036 18426
rect 19984 18362 20036 18368
rect 19996 16182 20024 18362
rect 20456 17105 20484 21542
rect 20718 21520 20774 21542
rect 20628 19236 20680 19242
rect 20628 19178 20680 19184
rect 20442 17096 20498 17105
rect 20442 17031 20498 17040
rect 19984 16176 20036 16182
rect 19984 16118 20036 16124
rect 19892 14068 19944 14074
rect 19892 14010 19944 14016
rect 19628 13806 19703 13812
rect 19798 13832 19854 13841
rect 19432 13728 19484 13734
rect 19432 13670 19484 13676
rect 19444 13326 19472 13670
rect 19432 13320 19484 13326
rect 19432 13262 19484 13268
rect 19289 13084 19585 13104
rect 19345 13082 19369 13084
rect 19425 13082 19449 13084
rect 19505 13082 19529 13084
rect 19367 13030 19369 13082
rect 19431 13030 19443 13082
rect 19505 13030 19507 13082
rect 19345 13028 19369 13030
rect 19425 13028 19449 13030
rect 19505 13028 19529 13030
rect 19289 13008 19585 13028
rect 19156 12912 19208 12918
rect 19156 12854 19208 12860
rect 18880 12844 18932 12850
rect 18880 12786 18932 12792
rect 18788 12436 18840 12442
rect 18788 12378 18840 12384
rect 18788 12164 18840 12170
rect 18788 12106 18840 12112
rect 18432 11886 18552 11914
rect 18328 10464 18380 10470
rect 18328 10406 18380 10412
rect 18340 10266 18368 10406
rect 18328 10260 18380 10266
rect 18328 10202 18380 10208
rect 18144 9580 18196 9586
rect 18144 9522 18196 9528
rect 18156 9178 18184 9522
rect 18144 9172 18196 9178
rect 18144 9114 18196 9120
rect 18236 8968 18288 8974
rect 18236 8910 18288 8916
rect 18144 8016 18196 8022
rect 18144 7958 18196 7964
rect 18156 7274 18184 7958
rect 18248 7886 18276 8910
rect 18328 8628 18380 8634
rect 18328 8570 18380 8576
rect 18340 8362 18368 8570
rect 18328 8356 18380 8362
rect 18328 8298 18380 8304
rect 18432 8242 18460 11886
rect 18512 11824 18564 11830
rect 18512 11766 18564 11772
rect 18340 8214 18460 8242
rect 18236 7880 18288 7886
rect 18236 7822 18288 7828
rect 18340 7274 18368 8214
rect 18524 8022 18552 11766
rect 18800 11626 18828 12106
rect 18892 11762 18920 12786
rect 19064 12368 19116 12374
rect 19064 12310 19116 12316
rect 18972 12232 19024 12238
rect 18972 12174 19024 12180
rect 18984 11830 19012 12174
rect 19076 11898 19104 12310
rect 19156 12232 19208 12238
rect 19156 12174 19208 12180
rect 19064 11892 19116 11898
rect 19064 11834 19116 11840
rect 18972 11824 19024 11830
rect 18972 11766 19024 11772
rect 18880 11756 18932 11762
rect 18880 11698 18932 11704
rect 18696 11620 18748 11626
rect 18696 11562 18748 11568
rect 18788 11620 18840 11626
rect 18788 11562 18840 11568
rect 18604 10532 18656 10538
rect 18604 10474 18656 10480
rect 18616 10266 18644 10474
rect 18604 10260 18656 10266
rect 18604 10202 18656 10208
rect 18708 9654 18736 11562
rect 18800 11354 18828 11562
rect 18788 11348 18840 11354
rect 18788 11290 18840 11296
rect 18788 11144 18840 11150
rect 18788 11086 18840 11092
rect 18800 10470 18828 11086
rect 19076 11014 19104 11834
rect 19168 11150 19196 12174
rect 19289 11996 19585 12016
rect 19345 11994 19369 11996
rect 19425 11994 19449 11996
rect 19505 11994 19529 11996
rect 19367 11942 19369 11994
rect 19431 11942 19443 11994
rect 19505 11942 19507 11994
rect 19345 11940 19369 11942
rect 19425 11940 19449 11942
rect 19505 11940 19529 11942
rect 19289 11920 19585 11940
rect 19628 11762 19656 13806
rect 19798 13767 19854 13776
rect 19616 11756 19668 11762
rect 19536 11716 19616 11744
rect 19536 11150 19564 11716
rect 19616 11698 19668 11704
rect 19616 11280 19668 11286
rect 19616 11222 19668 11228
rect 19156 11144 19208 11150
rect 19156 11086 19208 11092
rect 19524 11144 19576 11150
rect 19524 11086 19576 11092
rect 19064 11008 19116 11014
rect 19064 10950 19116 10956
rect 19289 10908 19585 10928
rect 19345 10906 19369 10908
rect 19425 10906 19449 10908
rect 19505 10906 19529 10908
rect 19367 10854 19369 10906
rect 19431 10854 19443 10906
rect 19505 10854 19507 10906
rect 19345 10852 19369 10854
rect 19425 10852 19449 10854
rect 19505 10852 19529 10854
rect 19289 10832 19585 10852
rect 19628 10810 19656 11222
rect 19708 11076 19760 11082
rect 19708 11018 19760 11024
rect 19616 10804 19668 10810
rect 19616 10746 19668 10752
rect 19720 10674 19748 11018
rect 19708 10668 19760 10674
rect 19708 10610 19760 10616
rect 18788 10464 18840 10470
rect 18788 10406 18840 10412
rect 18800 10062 18828 10406
rect 18788 10056 18840 10062
rect 18788 9998 18840 10004
rect 18696 9648 18748 9654
rect 18696 9590 18748 9596
rect 18800 8566 18828 9998
rect 19616 9988 19668 9994
rect 19616 9930 19668 9936
rect 19289 9820 19585 9840
rect 19345 9818 19369 9820
rect 19425 9818 19449 9820
rect 19505 9818 19529 9820
rect 19367 9766 19369 9818
rect 19431 9766 19443 9818
rect 19505 9766 19507 9818
rect 19345 9764 19369 9766
rect 19425 9764 19449 9766
rect 19505 9764 19529 9766
rect 19289 9744 19585 9764
rect 19064 9716 19116 9722
rect 19064 9658 19116 9664
rect 19076 9178 19104 9658
rect 19628 9382 19656 9930
rect 19616 9376 19668 9382
rect 19616 9318 19668 9324
rect 19064 9172 19116 9178
rect 19064 9114 19116 9120
rect 19156 9104 19208 9110
rect 19156 9046 19208 9052
rect 19168 8634 19196 9046
rect 19289 8732 19585 8752
rect 19345 8730 19369 8732
rect 19425 8730 19449 8732
rect 19505 8730 19529 8732
rect 19367 8678 19369 8730
rect 19431 8678 19443 8730
rect 19505 8678 19507 8730
rect 19345 8676 19369 8678
rect 19425 8676 19449 8678
rect 19505 8676 19529 8678
rect 19289 8656 19585 8676
rect 19156 8628 19208 8634
rect 19156 8570 19208 8576
rect 18788 8560 18840 8566
rect 18788 8502 18840 8508
rect 18972 8288 19024 8294
rect 18972 8230 19024 8236
rect 18512 8016 18564 8022
rect 18512 7958 18564 7964
rect 18880 7948 18932 7954
rect 18880 7890 18932 7896
rect 18420 7812 18472 7818
rect 18420 7754 18472 7760
rect 18144 7268 18196 7274
rect 18144 7210 18196 7216
rect 18328 7268 18380 7274
rect 18328 7210 18380 7216
rect 18052 6860 18104 6866
rect 18052 6802 18104 6808
rect 18432 6322 18460 7754
rect 18892 7410 18920 7890
rect 18880 7404 18932 7410
rect 18880 7346 18932 7352
rect 18512 7200 18564 7206
rect 18512 7142 18564 7148
rect 18524 6662 18552 7142
rect 18512 6656 18564 6662
rect 18512 6598 18564 6604
rect 18420 6316 18472 6322
rect 18420 6258 18472 6264
rect 17500 6248 17552 6254
rect 17500 6190 17552 6196
rect 17408 5908 17460 5914
rect 17408 5850 17460 5856
rect 17314 5128 17370 5137
rect 17314 5063 17370 5072
rect 17512 4154 17540 6190
rect 18144 6180 18196 6186
rect 18144 6122 18196 6128
rect 17684 5840 17736 5846
rect 17684 5782 17736 5788
rect 17592 5704 17644 5710
rect 17592 5646 17644 5652
rect 17420 4126 17540 4154
rect 17420 3670 17448 4126
rect 17224 3664 17276 3670
rect 17224 3606 17276 3612
rect 17408 3664 17460 3670
rect 17408 3606 17460 3612
rect 17316 3596 17368 3602
rect 17316 3538 17368 3544
rect 17130 3224 17186 3233
rect 17328 3194 17356 3538
rect 17130 3159 17186 3168
rect 17316 3188 17368 3194
rect 17316 3130 17368 3136
rect 17604 3126 17632 5646
rect 17696 5370 17724 5782
rect 18156 5556 18184 6122
rect 18432 5846 18460 6258
rect 18524 6186 18552 6598
rect 18512 6180 18564 6186
rect 18512 6122 18564 6128
rect 18420 5840 18472 5846
rect 18420 5782 18472 5788
rect 18236 5568 18288 5574
rect 18156 5528 18236 5556
rect 17684 5364 17736 5370
rect 17684 5306 17736 5312
rect 17684 5024 17736 5030
rect 17684 4966 17736 4972
rect 17696 4826 17724 4966
rect 17684 4820 17736 4826
rect 17684 4762 17736 4768
rect 17592 3120 17644 3126
rect 17592 3062 17644 3068
rect 18156 2650 18184 5528
rect 18236 5510 18288 5516
rect 18328 5228 18380 5234
rect 18328 5170 18380 5176
rect 18236 5092 18288 5098
rect 18236 5034 18288 5040
rect 18248 4826 18276 5034
rect 18340 4826 18368 5170
rect 18236 4820 18288 4826
rect 18236 4762 18288 4768
rect 18328 4820 18380 4826
rect 18328 4762 18380 4768
rect 18432 4622 18460 5782
rect 18984 5250 19012 8230
rect 19064 7948 19116 7954
rect 19064 7890 19116 7896
rect 19076 7206 19104 7890
rect 19289 7644 19585 7664
rect 19345 7642 19369 7644
rect 19425 7642 19449 7644
rect 19505 7642 19529 7644
rect 19367 7590 19369 7642
rect 19431 7590 19443 7642
rect 19505 7590 19507 7642
rect 19345 7588 19369 7590
rect 19425 7588 19449 7590
rect 19505 7588 19529 7590
rect 19289 7568 19585 7588
rect 19064 7200 19116 7206
rect 19064 7142 19116 7148
rect 19522 7168 19578 7177
rect 19076 6769 19104 7142
rect 19522 7103 19578 7112
rect 19536 7002 19564 7103
rect 19524 6996 19576 7002
rect 19524 6938 19576 6944
rect 19156 6860 19208 6866
rect 19156 6802 19208 6808
rect 19062 6760 19118 6769
rect 19062 6695 19118 6704
rect 19168 6458 19196 6802
rect 19289 6556 19585 6576
rect 19345 6554 19369 6556
rect 19425 6554 19449 6556
rect 19505 6554 19529 6556
rect 19367 6502 19369 6554
rect 19431 6502 19443 6554
rect 19505 6502 19507 6554
rect 19345 6500 19369 6502
rect 19425 6500 19449 6502
rect 19505 6500 19529 6502
rect 19289 6480 19585 6500
rect 19628 6458 19656 9318
rect 19892 8288 19944 8294
rect 19892 8230 19944 8236
rect 19708 7200 19760 7206
rect 19708 7142 19760 7148
rect 19156 6452 19208 6458
rect 19156 6394 19208 6400
rect 19616 6452 19668 6458
rect 19616 6394 19668 6400
rect 19156 5772 19208 5778
rect 19156 5714 19208 5720
rect 19064 5636 19116 5642
rect 19064 5578 19116 5584
rect 19076 5370 19104 5578
rect 19064 5364 19116 5370
rect 19064 5306 19116 5312
rect 18512 5228 18564 5234
rect 18984 5222 19104 5250
rect 18512 5170 18564 5176
rect 18420 4616 18472 4622
rect 18420 4558 18472 4564
rect 18236 4072 18288 4078
rect 18236 4014 18288 4020
rect 18248 3398 18276 4014
rect 18432 3738 18460 4558
rect 18524 4457 18552 5170
rect 18972 5092 19024 5098
rect 18972 5034 19024 5040
rect 18788 4752 18840 4758
rect 18788 4694 18840 4700
rect 18510 4448 18566 4457
rect 18510 4383 18566 4392
rect 18800 4282 18828 4694
rect 18984 4622 19012 5034
rect 18972 4616 19024 4622
rect 18972 4558 19024 4564
rect 18788 4276 18840 4282
rect 18788 4218 18840 4224
rect 18984 4154 19012 4558
rect 18800 4126 19012 4154
rect 18420 3732 18472 3738
rect 18420 3674 18472 3680
rect 18236 3392 18288 3398
rect 18236 3334 18288 3340
rect 18144 2644 18196 2650
rect 18144 2586 18196 2592
rect 16580 2576 16632 2582
rect 16580 2518 16632 2524
rect 16948 2576 17000 2582
rect 18248 2553 18276 3334
rect 18696 2984 18748 2990
rect 18696 2926 18748 2932
rect 16948 2518 17000 2524
rect 18234 2544 18290 2553
rect 15936 2508 15988 2514
rect 15936 2450 15988 2456
rect 15016 2372 15068 2378
rect 15016 2314 15068 2320
rect 14556 2304 14608 2310
rect 14556 2246 14608 2252
rect 12440 2100 12492 2106
rect 12440 2042 12492 2048
rect 11886 2000 11942 2009
rect 11886 1935 11942 1944
rect 10874 82 10930 480
rect 10704 54 10930 82
rect 8850 0 8906 54
rect 10874 0 10930 54
rect 12898 60 12954 480
rect 12898 8 12900 60
rect 12952 8 12954 60
rect 12898 0 12954 8
rect 14922 82 14978 480
rect 15028 82 15056 2314
rect 15200 2304 15252 2310
rect 15200 2246 15252 2252
rect 15212 1873 15240 2246
rect 15198 1864 15254 1873
rect 15198 1799 15254 1808
rect 14922 54 15056 82
rect 16592 82 16620 2518
rect 18234 2479 18290 2488
rect 18512 2440 18564 2446
rect 18512 2382 18564 2388
rect 18602 2408 18658 2417
rect 18052 2304 18104 2310
rect 18052 2246 18104 2252
rect 18064 1737 18092 2246
rect 18524 2106 18552 2382
rect 18602 2343 18658 2352
rect 18512 2100 18564 2106
rect 18512 2042 18564 2048
rect 18050 1728 18106 1737
rect 18050 1663 18106 1672
rect 16854 82 16910 480
rect 16592 54 16910 82
rect 18616 82 18644 2343
rect 18708 1057 18736 2926
rect 18800 2446 18828 4126
rect 19076 3738 19104 5222
rect 19168 5030 19196 5714
rect 19616 5636 19668 5642
rect 19616 5578 19668 5584
rect 19289 5468 19585 5488
rect 19345 5466 19369 5468
rect 19425 5466 19449 5468
rect 19505 5466 19529 5468
rect 19367 5414 19369 5466
rect 19431 5414 19443 5466
rect 19505 5414 19507 5466
rect 19345 5412 19369 5414
rect 19425 5412 19449 5414
rect 19505 5412 19529 5414
rect 19289 5392 19585 5412
rect 19156 5024 19208 5030
rect 19156 4966 19208 4972
rect 19628 4826 19656 5578
rect 19616 4820 19668 4826
rect 19616 4762 19668 4768
rect 19289 4380 19585 4400
rect 19345 4378 19369 4380
rect 19425 4378 19449 4380
rect 19505 4378 19529 4380
rect 19367 4326 19369 4378
rect 19431 4326 19443 4378
rect 19505 4326 19507 4378
rect 19345 4324 19369 4326
rect 19425 4324 19449 4326
rect 19505 4324 19529 4326
rect 19289 4304 19585 4324
rect 19720 4185 19748 7142
rect 19904 5370 19932 8230
rect 19892 5364 19944 5370
rect 19892 5306 19944 5312
rect 19706 4176 19762 4185
rect 19706 4111 19762 4120
rect 19064 3732 19116 3738
rect 19064 3674 19116 3680
rect 19156 3664 19208 3670
rect 19156 3606 19208 3612
rect 19064 3596 19116 3602
rect 19064 3538 19116 3544
rect 19076 3058 19104 3538
rect 19168 3194 19196 3606
rect 19289 3292 19585 3312
rect 19345 3290 19369 3292
rect 19425 3290 19449 3292
rect 19505 3290 19529 3292
rect 19367 3238 19369 3290
rect 19431 3238 19443 3290
rect 19505 3238 19507 3290
rect 19345 3236 19369 3238
rect 19425 3236 19449 3238
rect 19505 3236 19529 3238
rect 19289 3216 19585 3236
rect 19156 3188 19208 3194
rect 19156 3130 19208 3136
rect 19064 3052 19116 3058
rect 19064 2994 19116 3000
rect 19720 2990 19748 4111
rect 19708 2984 19760 2990
rect 19708 2926 19760 2932
rect 18788 2440 18840 2446
rect 18788 2382 18840 2388
rect 19289 2204 19585 2224
rect 19345 2202 19369 2204
rect 19425 2202 19449 2204
rect 19505 2202 19529 2204
rect 19367 2150 19369 2202
rect 19431 2150 19443 2202
rect 19505 2150 19507 2202
rect 19345 2148 19369 2150
rect 19425 2148 19449 2150
rect 19505 2148 19529 2150
rect 19289 2128 19585 2148
rect 18694 1048 18750 1057
rect 18694 983 18750 992
rect 18878 82 18934 480
rect 18616 54 18934 82
rect 20640 82 20668 19178
rect 21640 18896 21692 18902
rect 21640 18838 21692 18844
rect 21548 18624 21600 18630
rect 21652 18601 21680 18838
rect 21548 18566 21600 18572
rect 21638 18592 21694 18601
rect 21560 17649 21588 18566
rect 21638 18527 21694 18536
rect 21546 17640 21602 17649
rect 21546 17575 21602 17584
rect 21548 16788 21600 16794
rect 21548 16730 21600 16736
rect 21560 16697 21588 16730
rect 21546 16688 21602 16697
rect 21546 16623 21602 16632
rect 21548 8900 21600 8906
rect 21548 8842 21600 8848
rect 21560 8129 21588 8842
rect 21546 8120 21602 8129
rect 21546 8055 21602 8064
rect 20902 82 20958 480
rect 20640 54 20958 82
rect 14922 0 14978 54
rect 16854 0 16910 54
rect 18878 0 18934 54
rect 20902 0 20958 54
<< via2 >>
rect 2502 20440 2558 20496
rect 1582 18672 1638 18728
rect 1582 16768 1638 16824
rect 1306 13368 1362 13424
rect 1582 11464 1638 11520
rect 1950 10104 2006 10160
rect 1582 9696 1638 9752
rect 110 6296 166 6352
rect 1950 8472 2006 8528
rect 2410 13232 2466 13288
rect 1398 1672 1454 1728
rect 4622 19610 4678 19612
rect 4702 19610 4758 19612
rect 4782 19610 4838 19612
rect 4862 19610 4918 19612
rect 4622 19558 4648 19610
rect 4648 19558 4678 19610
rect 4702 19558 4712 19610
rect 4712 19558 4758 19610
rect 4782 19558 4828 19610
rect 4828 19558 4838 19610
rect 4862 19558 4892 19610
rect 4892 19558 4918 19610
rect 4622 19556 4678 19558
rect 4702 19556 4758 19558
rect 4782 19556 4838 19558
rect 4862 19556 4918 19558
rect 4622 18522 4678 18524
rect 4702 18522 4758 18524
rect 4782 18522 4838 18524
rect 4862 18522 4918 18524
rect 4622 18470 4648 18522
rect 4648 18470 4678 18522
rect 4702 18470 4712 18522
rect 4712 18470 4758 18522
rect 4782 18470 4828 18522
rect 4828 18470 4838 18522
rect 4862 18470 4892 18522
rect 4892 18470 4918 18522
rect 4622 18468 4678 18470
rect 4702 18468 4758 18470
rect 4782 18468 4838 18470
rect 4862 18468 4918 18470
rect 2594 7928 2650 7984
rect 2502 6296 2558 6352
rect 4622 17434 4678 17436
rect 4702 17434 4758 17436
rect 4782 17434 4838 17436
rect 4862 17434 4918 17436
rect 4622 17382 4648 17434
rect 4648 17382 4678 17434
rect 4702 17382 4712 17434
rect 4712 17382 4758 17434
rect 4782 17382 4828 17434
rect 4828 17382 4838 17434
rect 4862 17382 4892 17434
rect 4892 17382 4918 17434
rect 4622 17380 4678 17382
rect 4702 17380 4758 17382
rect 4782 17380 4838 17382
rect 4862 17380 4918 17382
rect 4986 17176 5042 17232
rect 4622 16346 4678 16348
rect 4702 16346 4758 16348
rect 4782 16346 4838 16348
rect 4862 16346 4918 16348
rect 4622 16294 4648 16346
rect 4648 16294 4678 16346
rect 4702 16294 4712 16346
rect 4712 16294 4758 16346
rect 4782 16294 4828 16346
rect 4828 16294 4838 16346
rect 4862 16294 4892 16346
rect 4892 16294 4918 16346
rect 4622 16292 4678 16294
rect 4702 16292 4758 16294
rect 4782 16292 4838 16294
rect 4862 16292 4918 16294
rect 4622 15258 4678 15260
rect 4702 15258 4758 15260
rect 4782 15258 4838 15260
rect 4862 15258 4918 15260
rect 4622 15206 4648 15258
rect 4648 15206 4678 15258
rect 4702 15206 4712 15258
rect 4712 15206 4758 15258
rect 4782 15206 4828 15258
rect 4828 15206 4838 15258
rect 4862 15206 4892 15258
rect 4892 15206 4918 15258
rect 4622 15204 4678 15206
rect 4702 15204 4758 15206
rect 4782 15204 4838 15206
rect 4862 15204 4918 15206
rect 3330 15000 3386 15056
rect 3146 11328 3202 11384
rect 3054 11056 3110 11112
rect 4342 14864 4398 14920
rect 3514 11192 3570 11248
rect 3054 8744 3110 8800
rect 3330 10648 3386 10704
rect 3422 9288 3478 9344
rect 2778 6296 2834 6352
rect 2318 5072 2374 5128
rect 2042 4392 2098 4448
rect 2134 3712 2190 3768
rect 3146 5752 3202 5808
rect 1950 3032 2006 3088
rect 4066 9016 4122 9072
rect 3790 7384 3846 7440
rect 3698 5208 3754 5264
rect 3514 4004 3570 4040
rect 3514 3984 3516 4004
rect 3516 3984 3568 4004
rect 3568 3984 3570 4004
rect 5262 15544 5318 15600
rect 5170 15000 5226 15056
rect 4622 14170 4678 14172
rect 4702 14170 4758 14172
rect 4782 14170 4838 14172
rect 4862 14170 4918 14172
rect 4622 14118 4648 14170
rect 4648 14118 4678 14170
rect 4702 14118 4712 14170
rect 4712 14118 4758 14170
rect 4782 14118 4828 14170
rect 4828 14118 4838 14170
rect 4862 14118 4892 14170
rect 4892 14118 4918 14170
rect 4622 14116 4678 14118
rect 4702 14116 4758 14118
rect 4782 14116 4838 14118
rect 4862 14116 4918 14118
rect 5170 13368 5226 13424
rect 4622 13082 4678 13084
rect 4702 13082 4758 13084
rect 4782 13082 4838 13084
rect 4862 13082 4918 13084
rect 4622 13030 4648 13082
rect 4648 13030 4678 13082
rect 4702 13030 4712 13082
rect 4712 13030 4758 13082
rect 4782 13030 4828 13082
rect 4828 13030 4838 13082
rect 4862 13030 4892 13082
rect 4892 13030 4918 13082
rect 4622 13028 4678 13030
rect 4702 13028 4758 13030
rect 4782 13028 4838 13030
rect 4862 13028 4918 13030
rect 4986 12824 5042 12880
rect 4622 11994 4678 11996
rect 4702 11994 4758 11996
rect 4782 11994 4838 11996
rect 4862 11994 4918 11996
rect 4622 11942 4648 11994
rect 4648 11942 4678 11994
rect 4702 11942 4712 11994
rect 4712 11942 4758 11994
rect 4782 11942 4828 11994
rect 4828 11942 4838 11994
rect 4862 11942 4892 11994
rect 4892 11942 4918 11994
rect 4622 11940 4678 11942
rect 4702 11940 4758 11942
rect 4782 11940 4838 11942
rect 4862 11940 4918 11942
rect 6274 15408 6330 15464
rect 5630 13812 5632 13832
rect 5632 13812 5684 13832
rect 5684 13812 5686 13832
rect 5630 13776 5686 13812
rect 4622 10906 4678 10908
rect 4702 10906 4758 10908
rect 4782 10906 4838 10908
rect 4862 10906 4918 10908
rect 4622 10854 4648 10906
rect 4648 10854 4678 10906
rect 4702 10854 4712 10906
rect 4712 10854 4758 10906
rect 4782 10854 4828 10906
rect 4828 10854 4838 10906
rect 4862 10854 4892 10906
rect 4892 10854 4918 10906
rect 4622 10852 4678 10854
rect 4702 10852 4758 10854
rect 4782 10852 4838 10854
rect 4862 10852 4918 10854
rect 4622 9818 4678 9820
rect 4702 9818 4758 9820
rect 4782 9818 4838 9820
rect 4862 9818 4918 9820
rect 4622 9766 4648 9818
rect 4648 9766 4678 9818
rect 4702 9766 4712 9818
rect 4712 9766 4758 9818
rect 4782 9766 4828 9818
rect 4828 9766 4838 9818
rect 4862 9766 4892 9818
rect 4892 9766 4918 9818
rect 4622 9764 4678 9766
rect 4702 9764 4758 9766
rect 4782 9764 4838 9766
rect 4862 9764 4918 9766
rect 4622 8730 4678 8732
rect 4702 8730 4758 8732
rect 4782 8730 4838 8732
rect 4862 8730 4918 8732
rect 4622 8678 4648 8730
rect 4648 8678 4678 8730
rect 4702 8678 4712 8730
rect 4712 8678 4758 8730
rect 4782 8678 4828 8730
rect 4828 8678 4838 8730
rect 4862 8678 4892 8730
rect 4892 8678 4918 8730
rect 4622 8676 4678 8678
rect 4702 8676 4758 8678
rect 4782 8676 4838 8678
rect 4862 8676 4918 8678
rect 4622 7642 4678 7644
rect 4702 7642 4758 7644
rect 4782 7642 4838 7644
rect 4862 7642 4918 7644
rect 4622 7590 4648 7642
rect 4648 7590 4678 7642
rect 4702 7590 4712 7642
rect 4712 7590 4758 7642
rect 4782 7590 4828 7642
rect 4828 7590 4838 7642
rect 4862 7590 4892 7642
rect 4892 7590 4918 7642
rect 4622 7588 4678 7590
rect 4702 7588 4758 7590
rect 4782 7588 4838 7590
rect 4862 7588 4918 7590
rect 5814 13096 5870 13152
rect 8289 19066 8345 19068
rect 8369 19066 8425 19068
rect 8449 19066 8505 19068
rect 8529 19066 8585 19068
rect 8289 19014 8315 19066
rect 8315 19014 8345 19066
rect 8369 19014 8379 19066
rect 8379 19014 8425 19066
rect 8449 19014 8495 19066
rect 8495 19014 8505 19066
rect 8529 19014 8559 19066
rect 8559 19014 8585 19066
rect 8289 19012 8345 19014
rect 8369 19012 8425 19014
rect 8449 19012 8505 19014
rect 8529 19012 8585 19014
rect 11956 19610 12012 19612
rect 12036 19610 12092 19612
rect 12116 19610 12172 19612
rect 12196 19610 12252 19612
rect 11956 19558 11982 19610
rect 11982 19558 12012 19610
rect 12036 19558 12046 19610
rect 12046 19558 12092 19610
rect 12116 19558 12162 19610
rect 12162 19558 12172 19610
rect 12196 19558 12226 19610
rect 12226 19558 12252 19610
rect 11956 19556 12012 19558
rect 12036 19556 12092 19558
rect 12116 19556 12172 19558
rect 12196 19556 12252 19558
rect 7010 17720 7066 17776
rect 6274 13640 6330 13696
rect 5446 9016 5502 9072
rect 5722 9968 5778 10024
rect 6090 10784 6146 10840
rect 4622 6554 4678 6556
rect 4702 6554 4758 6556
rect 4782 6554 4838 6556
rect 4862 6554 4918 6556
rect 4622 6502 4648 6554
rect 4648 6502 4678 6554
rect 4702 6502 4712 6554
rect 4712 6502 4758 6554
rect 4782 6502 4828 6554
rect 4828 6502 4838 6554
rect 4862 6502 4892 6554
rect 4892 6502 4918 6554
rect 4622 6500 4678 6502
rect 4702 6500 4758 6502
rect 4782 6500 4838 6502
rect 4862 6500 4918 6502
rect 4526 5616 4582 5672
rect 4622 5466 4678 5468
rect 4702 5466 4758 5468
rect 4782 5466 4838 5468
rect 4862 5466 4918 5468
rect 4622 5414 4648 5466
rect 4648 5414 4678 5466
rect 4702 5414 4712 5466
rect 4712 5414 4758 5466
rect 4782 5414 4828 5466
rect 4828 5414 4838 5466
rect 4862 5414 4892 5466
rect 4892 5414 4918 5466
rect 4622 5412 4678 5414
rect 4702 5412 4758 5414
rect 4782 5412 4838 5414
rect 4862 5412 4918 5414
rect 4434 5072 4490 5128
rect 3606 3576 3662 3632
rect 3330 2896 3386 2952
rect 4622 4378 4678 4380
rect 4702 4378 4758 4380
rect 4782 4378 4838 4380
rect 4862 4378 4918 4380
rect 4622 4326 4648 4378
rect 4648 4326 4678 4378
rect 4702 4326 4712 4378
rect 4712 4326 4758 4378
rect 4782 4326 4828 4378
rect 4828 4326 4838 4378
rect 4862 4326 4892 4378
rect 4892 4326 4918 4378
rect 4622 4324 4678 4326
rect 4702 4324 4758 4326
rect 4782 4324 4838 4326
rect 4862 4324 4918 4326
rect 6366 12688 6422 12744
rect 6458 10512 6514 10568
rect 5446 7384 5502 7440
rect 5078 6160 5134 6216
rect 4342 3440 4398 3496
rect 1766 1400 1822 1456
rect 4622 3290 4678 3292
rect 4702 3290 4758 3292
rect 4782 3290 4838 3292
rect 4862 3290 4918 3292
rect 4622 3238 4648 3290
rect 4648 3238 4678 3290
rect 4702 3238 4712 3290
rect 4712 3238 4758 3290
rect 4782 3238 4828 3290
rect 4828 3238 4838 3290
rect 4862 3238 4892 3290
rect 4892 3238 4918 3290
rect 4622 3236 4678 3238
rect 4702 3236 4758 3238
rect 4782 3236 4838 3238
rect 4862 3236 4918 3238
rect 4434 2488 4490 2544
rect 4622 2202 4678 2204
rect 4702 2202 4758 2204
rect 4782 2202 4838 2204
rect 4862 2202 4918 2204
rect 4622 2150 4648 2202
rect 4648 2150 4678 2202
rect 4702 2150 4712 2202
rect 4712 2150 4758 2202
rect 4782 2150 4828 2202
rect 4828 2150 4838 2202
rect 4862 2150 4892 2202
rect 4892 2150 4918 2202
rect 4622 2148 4678 2150
rect 4702 2148 4758 2150
rect 4782 2148 4838 2150
rect 4862 2148 4918 2150
rect 4342 1808 4398 1864
rect 5814 7792 5870 7848
rect 5630 6704 5686 6760
rect 6182 6296 6238 6352
rect 6550 6704 6606 6760
rect 6826 13640 6882 13696
rect 8289 17978 8345 17980
rect 8369 17978 8425 17980
rect 8449 17978 8505 17980
rect 8529 17978 8585 17980
rect 8289 17926 8315 17978
rect 8315 17926 8345 17978
rect 8369 17926 8379 17978
rect 8379 17926 8425 17978
rect 8449 17926 8495 17978
rect 8495 17926 8505 17978
rect 8529 17926 8559 17978
rect 8559 17926 8585 17978
rect 8289 17924 8345 17926
rect 8369 17924 8425 17926
rect 8449 17924 8505 17926
rect 8529 17924 8585 17926
rect 8289 16890 8345 16892
rect 8369 16890 8425 16892
rect 8449 16890 8505 16892
rect 8529 16890 8585 16892
rect 8289 16838 8315 16890
rect 8315 16838 8345 16890
rect 8369 16838 8379 16890
rect 8379 16838 8425 16890
rect 8449 16838 8495 16890
rect 8495 16838 8505 16890
rect 8529 16838 8559 16890
rect 8559 16838 8585 16890
rect 8289 16836 8345 16838
rect 8369 16836 8425 16838
rect 8449 16836 8505 16838
rect 8529 16836 8585 16838
rect 8289 15802 8345 15804
rect 8369 15802 8425 15804
rect 8449 15802 8505 15804
rect 8529 15802 8585 15804
rect 8289 15750 8315 15802
rect 8315 15750 8345 15802
rect 8369 15750 8379 15802
rect 8379 15750 8425 15802
rect 8449 15750 8495 15802
rect 8495 15750 8505 15802
rect 8529 15750 8559 15802
rect 8559 15750 8585 15802
rect 8289 15748 8345 15750
rect 8369 15748 8425 15750
rect 8449 15748 8505 15750
rect 8529 15748 8585 15750
rect 8289 14714 8345 14716
rect 8369 14714 8425 14716
rect 8449 14714 8505 14716
rect 8529 14714 8585 14716
rect 8289 14662 8315 14714
rect 8315 14662 8345 14714
rect 8369 14662 8379 14714
rect 8379 14662 8425 14714
rect 8449 14662 8495 14714
rect 8495 14662 8505 14714
rect 8529 14662 8559 14714
rect 8559 14662 8585 14714
rect 8289 14660 8345 14662
rect 8369 14660 8425 14662
rect 8449 14660 8505 14662
rect 8529 14660 8585 14662
rect 8289 13626 8345 13628
rect 8369 13626 8425 13628
rect 8449 13626 8505 13628
rect 8529 13626 8585 13628
rect 8289 13574 8315 13626
rect 8315 13574 8345 13626
rect 8369 13574 8379 13626
rect 8379 13574 8425 13626
rect 8449 13574 8495 13626
rect 8495 13574 8505 13626
rect 8529 13574 8559 13626
rect 8559 13574 8585 13626
rect 8289 13572 8345 13574
rect 8369 13572 8425 13574
rect 8449 13572 8505 13574
rect 8529 13572 8585 13574
rect 9034 15952 9090 16008
rect 9494 13776 9550 13832
rect 10046 13776 10102 13832
rect 9862 13096 9918 13152
rect 8289 12538 8345 12540
rect 8369 12538 8425 12540
rect 8449 12538 8505 12540
rect 8529 12538 8585 12540
rect 8289 12486 8315 12538
rect 8315 12486 8345 12538
rect 8369 12486 8379 12538
rect 8379 12486 8425 12538
rect 8449 12486 8495 12538
rect 8495 12486 8505 12538
rect 8529 12486 8559 12538
rect 8559 12486 8585 12538
rect 8289 12484 8345 12486
rect 8369 12484 8425 12486
rect 8449 12484 8505 12486
rect 8529 12484 8585 12486
rect 7102 10784 7158 10840
rect 7378 11328 7434 11384
rect 8289 11450 8345 11452
rect 8369 11450 8425 11452
rect 8449 11450 8505 11452
rect 8529 11450 8585 11452
rect 8289 11398 8315 11450
rect 8315 11398 8345 11450
rect 8369 11398 8379 11450
rect 8379 11398 8425 11450
rect 8449 11398 8495 11450
rect 8495 11398 8505 11450
rect 8529 11398 8559 11450
rect 8559 11398 8585 11450
rect 8289 11396 8345 11398
rect 8369 11396 8425 11398
rect 8449 11396 8505 11398
rect 8529 11396 8585 11398
rect 8114 10648 8170 10704
rect 8758 10648 8814 10704
rect 8289 10362 8345 10364
rect 8369 10362 8425 10364
rect 8449 10362 8505 10364
rect 8529 10362 8585 10364
rect 8289 10310 8315 10362
rect 8315 10310 8345 10362
rect 8369 10310 8379 10362
rect 8379 10310 8425 10362
rect 8449 10310 8495 10362
rect 8495 10310 8505 10362
rect 8529 10310 8559 10362
rect 8559 10310 8585 10362
rect 8289 10308 8345 10310
rect 8369 10308 8425 10310
rect 8449 10308 8505 10310
rect 8529 10308 8585 10310
rect 7562 10104 7618 10160
rect 8114 9288 8170 9344
rect 8289 9274 8345 9276
rect 8369 9274 8425 9276
rect 8449 9274 8505 9276
rect 8529 9274 8585 9276
rect 8289 9222 8315 9274
rect 8315 9222 8345 9274
rect 8369 9222 8379 9274
rect 8379 9222 8425 9274
rect 8449 9222 8495 9274
rect 8495 9222 8505 9274
rect 8529 9222 8559 9274
rect 8559 9222 8585 9274
rect 8289 9220 8345 9222
rect 8369 9220 8425 9222
rect 8449 9220 8505 9222
rect 8529 9220 8585 9222
rect 7654 8064 7710 8120
rect 6274 4528 6330 4584
rect 5906 3032 5962 3088
rect 5538 2896 5594 2952
rect 8289 8186 8345 8188
rect 8369 8186 8425 8188
rect 8449 8186 8505 8188
rect 8529 8186 8585 8188
rect 8289 8134 8315 8186
rect 8315 8134 8345 8186
rect 8369 8134 8379 8186
rect 8379 8134 8425 8186
rect 8449 8134 8495 8186
rect 8495 8134 8505 8186
rect 8529 8134 8559 8186
rect 8559 8134 8585 8186
rect 8289 8132 8345 8134
rect 8369 8132 8425 8134
rect 8449 8132 8505 8134
rect 8529 8132 8585 8134
rect 8114 8064 8170 8120
rect 8666 7928 8722 7984
rect 8289 7098 8345 7100
rect 8369 7098 8425 7100
rect 8449 7098 8505 7100
rect 8529 7098 8585 7100
rect 8289 7046 8315 7098
rect 8315 7046 8345 7098
rect 8369 7046 8379 7098
rect 8379 7046 8425 7098
rect 8449 7046 8495 7098
rect 8495 7046 8505 7098
rect 8529 7046 8559 7098
rect 8559 7046 8585 7098
rect 8289 7044 8345 7046
rect 8369 7044 8425 7046
rect 8449 7044 8505 7046
rect 8529 7044 8585 7046
rect 6826 4120 6882 4176
rect 5906 2352 5962 2408
rect 8022 4936 8078 4992
rect 7930 4664 7986 4720
rect 8758 6160 8814 6216
rect 8666 6024 8722 6080
rect 8289 6010 8345 6012
rect 8369 6010 8425 6012
rect 8449 6010 8505 6012
rect 8529 6010 8585 6012
rect 8289 5958 8315 6010
rect 8315 5958 8345 6010
rect 8369 5958 8379 6010
rect 8379 5958 8425 6010
rect 8449 5958 8495 6010
rect 8495 5958 8505 6010
rect 8529 5958 8559 6010
rect 8559 5958 8585 6010
rect 8289 5956 8345 5958
rect 8369 5956 8425 5958
rect 8449 5956 8505 5958
rect 8529 5956 8585 5958
rect 8289 4922 8345 4924
rect 8369 4922 8425 4924
rect 8449 4922 8505 4924
rect 8529 4922 8585 4924
rect 8289 4870 8315 4922
rect 8315 4870 8345 4922
rect 8369 4870 8379 4922
rect 8379 4870 8425 4922
rect 8449 4870 8495 4922
rect 8495 4870 8505 4922
rect 8529 4870 8559 4922
rect 8559 4870 8585 4922
rect 8289 4868 8345 4870
rect 8369 4868 8425 4870
rect 8449 4868 8505 4870
rect 8529 4868 8585 4870
rect 7194 3984 7250 4040
rect 7286 3848 7342 3904
rect 9034 6160 9090 6216
rect 9770 10784 9826 10840
rect 9954 10376 10010 10432
rect 9954 8472 10010 8528
rect 9678 7384 9734 7440
rect 10230 13368 10286 13424
rect 11956 18522 12012 18524
rect 12036 18522 12092 18524
rect 12116 18522 12172 18524
rect 12196 18522 12252 18524
rect 11956 18470 11982 18522
rect 11982 18470 12012 18522
rect 12036 18470 12046 18522
rect 12046 18470 12092 18522
rect 12116 18470 12162 18522
rect 12162 18470 12172 18522
rect 12196 18470 12226 18522
rect 12226 18470 12252 18522
rect 11956 18468 12012 18470
rect 12036 18468 12092 18470
rect 12116 18468 12172 18470
rect 12196 18468 12252 18470
rect 11058 17040 11114 17096
rect 11956 17434 12012 17436
rect 12036 17434 12092 17436
rect 12116 17434 12172 17436
rect 12196 17434 12252 17436
rect 11956 17382 11982 17434
rect 11982 17382 12012 17434
rect 12036 17382 12046 17434
rect 12046 17382 12092 17434
rect 12116 17382 12162 17434
rect 12162 17382 12172 17434
rect 12196 17382 12226 17434
rect 12226 17382 12252 17434
rect 11956 17380 12012 17382
rect 12036 17380 12092 17382
rect 12116 17380 12172 17382
rect 12196 17380 12252 17382
rect 12714 17312 12770 17368
rect 10966 15000 11022 15056
rect 10322 11056 10378 11112
rect 11956 16346 12012 16348
rect 12036 16346 12092 16348
rect 12116 16346 12172 16348
rect 12196 16346 12252 16348
rect 11956 16294 11982 16346
rect 11982 16294 12012 16346
rect 12036 16294 12046 16346
rect 12046 16294 12092 16346
rect 12116 16294 12162 16346
rect 12162 16294 12172 16346
rect 12196 16294 12226 16346
rect 12226 16294 12252 16346
rect 11956 16292 12012 16294
rect 12036 16292 12092 16294
rect 12116 16292 12172 16294
rect 12196 16292 12252 16294
rect 11956 15258 12012 15260
rect 12036 15258 12092 15260
rect 12116 15258 12172 15260
rect 12196 15258 12252 15260
rect 11956 15206 11982 15258
rect 11982 15206 12012 15258
rect 12036 15206 12046 15258
rect 12046 15206 12092 15258
rect 12116 15206 12162 15258
rect 12162 15206 12172 15258
rect 12196 15206 12226 15258
rect 12226 15206 12252 15258
rect 11956 15204 12012 15206
rect 12036 15204 12092 15206
rect 12116 15204 12172 15206
rect 12196 15204 12252 15206
rect 11956 14170 12012 14172
rect 12036 14170 12092 14172
rect 12116 14170 12172 14172
rect 12196 14170 12252 14172
rect 11956 14118 11982 14170
rect 11982 14118 12012 14170
rect 12036 14118 12046 14170
rect 12046 14118 12092 14170
rect 12116 14118 12162 14170
rect 12162 14118 12172 14170
rect 12196 14118 12226 14170
rect 12226 14118 12252 14170
rect 11956 14116 12012 14118
rect 12036 14116 12092 14118
rect 12116 14116 12172 14118
rect 12196 14116 12252 14118
rect 11956 13082 12012 13084
rect 12036 13082 12092 13084
rect 12116 13082 12172 13084
rect 12196 13082 12252 13084
rect 11956 13030 11982 13082
rect 11982 13030 12012 13082
rect 12036 13030 12046 13082
rect 12046 13030 12092 13082
rect 12116 13030 12162 13082
rect 12162 13030 12172 13082
rect 12196 13030 12226 13082
rect 12226 13030 12252 13082
rect 11956 13028 12012 13030
rect 12036 13028 12092 13030
rect 12116 13028 12172 13030
rect 12196 13028 12252 13030
rect 10782 10376 10838 10432
rect 10138 6024 10194 6080
rect 8666 3848 8722 3904
rect 8289 3834 8345 3836
rect 8369 3834 8425 3836
rect 8449 3834 8505 3836
rect 8529 3834 8585 3836
rect 8289 3782 8315 3834
rect 8315 3782 8345 3834
rect 8369 3782 8379 3834
rect 8379 3782 8425 3834
rect 8449 3782 8495 3834
rect 8495 3782 8505 3834
rect 8529 3782 8559 3834
rect 8559 3782 8585 3834
rect 8289 3780 8345 3782
rect 8369 3780 8425 3782
rect 8449 3780 8505 3782
rect 8529 3780 8585 3782
rect 7194 3304 7250 3360
rect 8289 2746 8345 2748
rect 8369 2746 8425 2748
rect 8449 2746 8505 2748
rect 8529 2746 8585 2748
rect 8289 2694 8315 2746
rect 8315 2694 8345 2746
rect 8369 2694 8379 2746
rect 8379 2694 8425 2746
rect 8449 2694 8495 2746
rect 8495 2694 8505 2746
rect 8529 2694 8559 2746
rect 8559 2694 8585 2746
rect 8289 2692 8345 2694
rect 8369 2692 8425 2694
rect 8449 2692 8505 2694
rect 8529 2692 8585 2694
rect 10598 7384 10654 7440
rect 10598 3576 10654 3632
rect 11242 11192 11298 11248
rect 14462 20848 14518 20904
rect 12898 13232 12954 13288
rect 11956 11994 12012 11996
rect 12036 11994 12092 11996
rect 12116 11994 12172 11996
rect 12196 11994 12252 11996
rect 11956 11942 11982 11994
rect 11982 11942 12012 11994
rect 12036 11942 12046 11994
rect 12046 11942 12092 11994
rect 12116 11942 12162 11994
rect 12162 11942 12172 11994
rect 12196 11942 12226 11994
rect 12226 11942 12252 11994
rect 11956 11940 12012 11942
rect 12036 11940 12092 11942
rect 12116 11940 12172 11942
rect 12196 11940 12252 11942
rect 11956 10906 12012 10908
rect 12036 10906 12092 10908
rect 12116 10906 12172 10908
rect 12196 10906 12252 10908
rect 11956 10854 11982 10906
rect 11982 10854 12012 10906
rect 12036 10854 12046 10906
rect 12046 10854 12092 10906
rect 12116 10854 12162 10906
rect 12162 10854 12172 10906
rect 12196 10854 12226 10906
rect 12226 10854 12252 10906
rect 11956 10852 12012 10854
rect 12036 10852 12092 10854
rect 12116 10852 12172 10854
rect 12196 10852 12252 10854
rect 11518 10104 11574 10160
rect 12622 10512 12678 10568
rect 12438 9968 12494 10024
rect 11956 9818 12012 9820
rect 12036 9818 12092 9820
rect 12116 9818 12172 9820
rect 12196 9818 12252 9820
rect 11956 9766 11982 9818
rect 11982 9766 12012 9818
rect 12036 9766 12046 9818
rect 12046 9766 12092 9818
rect 12116 9766 12162 9818
rect 12162 9766 12172 9818
rect 12196 9766 12226 9818
rect 12226 9766 12252 9818
rect 11956 9764 12012 9766
rect 12036 9764 12092 9766
rect 12116 9764 12172 9766
rect 12196 9764 12252 9766
rect 12806 9832 12862 9888
rect 11794 8880 11850 8936
rect 11956 8730 12012 8732
rect 12036 8730 12092 8732
rect 12116 8730 12172 8732
rect 12196 8730 12252 8732
rect 11956 8678 11982 8730
rect 11982 8678 12012 8730
rect 12036 8678 12046 8730
rect 12046 8678 12092 8730
rect 12116 8678 12162 8730
rect 12162 8678 12172 8730
rect 12196 8678 12226 8730
rect 12226 8678 12252 8730
rect 11956 8676 12012 8678
rect 12036 8676 12092 8678
rect 12116 8676 12172 8678
rect 12196 8676 12252 8678
rect 11956 7642 12012 7644
rect 12036 7642 12092 7644
rect 12116 7642 12172 7644
rect 12196 7642 12252 7644
rect 11956 7590 11982 7642
rect 11982 7590 12012 7642
rect 12036 7590 12046 7642
rect 12046 7590 12092 7642
rect 12116 7590 12162 7642
rect 12162 7590 12172 7642
rect 12196 7590 12226 7642
rect 12226 7590 12252 7642
rect 11956 7588 12012 7590
rect 12036 7588 12092 7590
rect 12116 7588 12172 7590
rect 12196 7588 12252 7590
rect 11956 6554 12012 6556
rect 12036 6554 12092 6556
rect 12116 6554 12172 6556
rect 12196 6554 12252 6556
rect 11956 6502 11982 6554
rect 11982 6502 12012 6554
rect 12036 6502 12046 6554
rect 12046 6502 12092 6554
rect 12116 6502 12162 6554
rect 12162 6502 12172 6554
rect 12196 6502 12226 6554
rect 12226 6502 12252 6554
rect 11956 6500 12012 6502
rect 12036 6500 12092 6502
rect 12116 6500 12172 6502
rect 12196 6500 12252 6502
rect 11956 5466 12012 5468
rect 12036 5466 12092 5468
rect 12116 5466 12172 5468
rect 12196 5466 12252 5468
rect 11956 5414 11982 5466
rect 11982 5414 12012 5466
rect 12036 5414 12046 5466
rect 12046 5414 12092 5466
rect 12116 5414 12162 5466
rect 12162 5414 12172 5466
rect 12196 5414 12226 5466
rect 12226 5414 12252 5466
rect 11956 5412 12012 5414
rect 12036 5412 12092 5414
rect 12116 5412 12172 5414
rect 12196 5412 12252 5414
rect 10782 3304 10838 3360
rect 10874 2932 10876 2952
rect 10876 2932 10928 2952
rect 10928 2932 10930 2952
rect 10874 2896 10930 2932
rect 11794 4528 11850 4584
rect 12346 5228 12402 5264
rect 12346 5208 12348 5228
rect 12348 5208 12400 5228
rect 12400 5208 12402 5228
rect 12622 6024 12678 6080
rect 11978 4528 12034 4584
rect 11956 4378 12012 4380
rect 12036 4378 12092 4380
rect 12116 4378 12172 4380
rect 12196 4378 12252 4380
rect 11956 4326 11982 4378
rect 11982 4326 12012 4378
rect 12036 4326 12046 4378
rect 12046 4326 12092 4378
rect 12116 4326 12162 4378
rect 12162 4326 12172 4378
rect 12196 4326 12226 4378
rect 12226 4326 12252 4378
rect 11956 4324 12012 4326
rect 12036 4324 12092 4326
rect 12116 4324 12172 4326
rect 12196 4324 12252 4326
rect 12530 5072 12586 5128
rect 12806 5752 12862 5808
rect 13174 5616 13230 5672
rect 13818 17720 13874 17776
rect 14094 15408 14150 15464
rect 14094 12280 14150 12336
rect 15750 19896 15806 19952
rect 14370 17176 14426 17232
rect 15622 19066 15678 19068
rect 15702 19066 15758 19068
rect 15782 19066 15838 19068
rect 15862 19066 15918 19068
rect 15622 19014 15648 19066
rect 15648 19014 15678 19066
rect 15702 19014 15712 19066
rect 15712 19014 15758 19066
rect 15782 19014 15828 19066
rect 15828 19014 15838 19066
rect 15862 19014 15892 19066
rect 15892 19014 15918 19066
rect 15622 19012 15678 19014
rect 15702 19012 15758 19014
rect 15782 19012 15838 19014
rect 15862 19012 15918 19014
rect 14278 10648 14334 10704
rect 14830 15952 14886 16008
rect 14922 15544 14978 15600
rect 14738 13776 14794 13832
rect 15106 13776 15162 13832
rect 15622 17978 15678 17980
rect 15702 17978 15758 17980
rect 15782 17978 15838 17980
rect 15862 17978 15918 17980
rect 15622 17926 15648 17978
rect 15648 17926 15678 17978
rect 15702 17926 15712 17978
rect 15712 17926 15758 17978
rect 15782 17926 15828 17978
rect 15828 17926 15838 17978
rect 15862 17926 15892 17978
rect 15892 17926 15918 17978
rect 15622 17924 15678 17926
rect 15702 17924 15758 17926
rect 15782 17924 15838 17926
rect 15862 17924 15918 17926
rect 15934 17312 15990 17368
rect 15622 16890 15678 16892
rect 15702 16890 15758 16892
rect 15782 16890 15838 16892
rect 15862 16890 15918 16892
rect 15622 16838 15648 16890
rect 15648 16838 15678 16890
rect 15702 16838 15712 16890
rect 15712 16838 15758 16890
rect 15782 16838 15828 16890
rect 15828 16838 15838 16890
rect 15862 16838 15892 16890
rect 15892 16838 15918 16890
rect 15622 16836 15678 16838
rect 15702 16836 15758 16838
rect 15782 16836 15838 16838
rect 15862 16836 15918 16838
rect 15622 15802 15678 15804
rect 15702 15802 15758 15804
rect 15782 15802 15838 15804
rect 15862 15802 15918 15804
rect 15622 15750 15648 15802
rect 15648 15750 15678 15802
rect 15702 15750 15712 15802
rect 15712 15750 15758 15802
rect 15782 15750 15828 15802
rect 15828 15750 15838 15802
rect 15862 15750 15892 15802
rect 15892 15750 15918 15802
rect 15622 15748 15678 15750
rect 15702 15748 15758 15750
rect 15782 15748 15838 15750
rect 15862 15748 15918 15750
rect 15474 14864 15530 14920
rect 15622 14714 15678 14716
rect 15702 14714 15758 14716
rect 15782 14714 15838 14716
rect 15862 14714 15918 14716
rect 15622 14662 15648 14714
rect 15648 14662 15678 14714
rect 15702 14662 15712 14714
rect 15712 14662 15758 14714
rect 15782 14662 15828 14714
rect 15828 14662 15838 14714
rect 15862 14662 15892 14714
rect 15892 14662 15918 14714
rect 15622 14660 15678 14662
rect 15702 14660 15758 14662
rect 15782 14660 15838 14662
rect 15862 14660 15918 14662
rect 16026 14592 16082 14648
rect 15622 13626 15678 13628
rect 15702 13626 15758 13628
rect 15782 13626 15838 13628
rect 15862 13626 15918 13628
rect 15622 13574 15648 13626
rect 15648 13574 15678 13626
rect 15702 13574 15712 13626
rect 15712 13574 15758 13626
rect 15782 13574 15828 13626
rect 15828 13574 15838 13626
rect 15862 13574 15892 13626
rect 15892 13574 15918 13626
rect 15622 13572 15678 13574
rect 15702 13572 15758 13574
rect 15782 13572 15838 13574
rect 15862 13572 15918 13574
rect 15622 12538 15678 12540
rect 15702 12538 15758 12540
rect 15782 12538 15838 12540
rect 15862 12538 15918 12540
rect 15622 12486 15648 12538
rect 15648 12486 15678 12538
rect 15702 12486 15712 12538
rect 15712 12486 15758 12538
rect 15782 12486 15828 12538
rect 15828 12486 15838 12538
rect 15862 12486 15892 12538
rect 15892 12486 15918 12538
rect 15622 12484 15678 12486
rect 15702 12484 15758 12486
rect 15782 12484 15838 12486
rect 15862 12484 15918 12486
rect 15622 11450 15678 11452
rect 15702 11450 15758 11452
rect 15782 11450 15838 11452
rect 15862 11450 15918 11452
rect 15622 11398 15648 11450
rect 15648 11398 15678 11450
rect 15702 11398 15712 11450
rect 15712 11398 15758 11450
rect 15782 11398 15828 11450
rect 15828 11398 15838 11450
rect 15862 11398 15892 11450
rect 15892 11398 15918 11450
rect 15622 11396 15678 11398
rect 15702 11396 15758 11398
rect 15782 11396 15838 11398
rect 15862 11396 15918 11398
rect 16854 15000 16910 15056
rect 17038 15408 17094 15464
rect 17038 12688 17094 12744
rect 16394 11328 16450 11384
rect 15934 10512 15990 10568
rect 15474 10376 15530 10432
rect 15622 10362 15678 10364
rect 15702 10362 15758 10364
rect 15782 10362 15838 10364
rect 15862 10362 15918 10364
rect 15622 10310 15648 10362
rect 15648 10310 15678 10362
rect 15702 10310 15712 10362
rect 15712 10310 15758 10362
rect 15782 10310 15828 10362
rect 15828 10310 15838 10362
rect 15862 10310 15892 10362
rect 15892 10310 15918 10362
rect 15622 10308 15678 10310
rect 15702 10308 15758 10310
rect 15782 10308 15838 10310
rect 15862 10308 15918 10310
rect 16394 10104 16450 10160
rect 15622 9274 15678 9276
rect 15702 9274 15758 9276
rect 15782 9274 15838 9276
rect 15862 9274 15918 9276
rect 15622 9222 15648 9274
rect 15648 9222 15678 9274
rect 15702 9222 15712 9274
rect 15712 9222 15758 9274
rect 15782 9222 15828 9274
rect 15828 9222 15838 9274
rect 15862 9222 15892 9274
rect 15892 9222 15918 9274
rect 15622 9220 15678 9222
rect 15702 9220 15758 9222
rect 15782 9220 15838 9222
rect 15862 9220 15918 9222
rect 15014 6160 15070 6216
rect 13818 4392 13874 4448
rect 13450 4020 13452 4040
rect 13452 4020 13504 4040
rect 13504 4020 13506 4040
rect 13450 3984 13506 4020
rect 12438 3440 12494 3496
rect 11956 3290 12012 3292
rect 12036 3290 12092 3292
rect 12116 3290 12172 3292
rect 12196 3290 12252 3292
rect 11956 3238 11982 3290
rect 11982 3238 12012 3290
rect 12036 3238 12046 3290
rect 12046 3238 12092 3290
rect 12116 3238 12162 3290
rect 12162 3238 12172 3290
rect 12196 3238 12226 3290
rect 12226 3238 12252 3290
rect 11956 3236 12012 3238
rect 12036 3236 12092 3238
rect 12116 3236 12172 3238
rect 12196 3236 12252 3238
rect 11956 2202 12012 2204
rect 12036 2202 12092 2204
rect 12116 2202 12172 2204
rect 12196 2202 12252 2204
rect 11956 2150 11982 2202
rect 11982 2150 12012 2202
rect 12036 2150 12046 2202
rect 12046 2150 12092 2202
rect 12116 2150 12162 2202
rect 12162 2150 12172 2202
rect 12196 2150 12226 2202
rect 12226 2150 12252 2202
rect 11956 2148 12012 2150
rect 12036 2148 12092 2150
rect 12116 2148 12172 2150
rect 12196 2148 12252 2150
rect 15622 8186 15678 8188
rect 15702 8186 15758 8188
rect 15782 8186 15838 8188
rect 15862 8186 15918 8188
rect 15622 8134 15648 8186
rect 15648 8134 15678 8186
rect 15702 8134 15712 8186
rect 15712 8134 15758 8186
rect 15782 8134 15828 8186
rect 15828 8134 15838 8186
rect 15862 8134 15892 8186
rect 15892 8134 15918 8186
rect 15622 8132 15678 8134
rect 15702 8132 15758 8134
rect 15782 8132 15838 8134
rect 15862 8132 15918 8134
rect 15622 7098 15678 7100
rect 15702 7098 15758 7100
rect 15782 7098 15838 7100
rect 15862 7098 15918 7100
rect 15622 7046 15648 7098
rect 15648 7046 15678 7098
rect 15702 7046 15712 7098
rect 15712 7046 15758 7098
rect 15782 7046 15828 7098
rect 15828 7046 15838 7098
rect 15862 7046 15892 7098
rect 15892 7046 15918 7098
rect 15622 7044 15678 7046
rect 15702 7044 15758 7046
rect 15782 7044 15838 7046
rect 15862 7044 15918 7046
rect 15622 6010 15678 6012
rect 15702 6010 15758 6012
rect 15782 6010 15838 6012
rect 15862 6010 15918 6012
rect 15622 5958 15648 6010
rect 15648 5958 15678 6010
rect 15702 5958 15712 6010
rect 15712 5958 15758 6010
rect 15782 5958 15828 6010
rect 15828 5958 15838 6010
rect 15862 5958 15892 6010
rect 15892 5958 15918 6010
rect 15622 5956 15678 5958
rect 15702 5956 15758 5958
rect 15782 5956 15838 5958
rect 15862 5956 15918 5958
rect 15622 4922 15678 4924
rect 15702 4922 15758 4924
rect 15782 4922 15838 4924
rect 15862 4922 15918 4924
rect 15622 4870 15648 4922
rect 15648 4870 15678 4922
rect 15702 4870 15712 4922
rect 15712 4870 15758 4922
rect 15782 4870 15828 4922
rect 15828 4870 15838 4922
rect 15862 4870 15892 4922
rect 15892 4870 15918 4922
rect 15622 4868 15678 4870
rect 15702 4868 15758 4870
rect 15782 4868 15838 4870
rect 15862 4868 15918 4870
rect 15474 4664 15530 4720
rect 15934 4392 15990 4448
rect 15382 3848 15438 3904
rect 15622 3834 15678 3836
rect 15702 3834 15758 3836
rect 15782 3834 15838 3836
rect 15862 3834 15918 3836
rect 15622 3782 15648 3834
rect 15648 3782 15678 3834
rect 15702 3782 15712 3834
rect 15712 3782 15758 3834
rect 15782 3782 15828 3834
rect 15828 3782 15838 3834
rect 15862 3782 15892 3834
rect 15892 3782 15918 3834
rect 15622 3780 15678 3782
rect 15702 3780 15758 3782
rect 15782 3780 15838 3782
rect 15862 3780 15918 3782
rect 14922 3032 14978 3088
rect 15106 3032 15162 3088
rect 15622 2746 15678 2748
rect 15702 2746 15758 2748
rect 15782 2746 15838 2748
rect 15862 2746 15918 2748
rect 15622 2694 15648 2746
rect 15648 2694 15678 2746
rect 15702 2694 15712 2746
rect 15712 2694 15758 2746
rect 15782 2694 15828 2746
rect 15828 2694 15838 2746
rect 15862 2694 15892 2746
rect 15892 2694 15918 2746
rect 15622 2692 15678 2694
rect 15702 2692 15758 2694
rect 15782 2692 15838 2694
rect 15862 2692 15918 2694
rect 17130 7828 17132 7848
rect 17132 7828 17184 7848
rect 17184 7828 17186 7848
rect 17130 7792 17186 7828
rect 19289 19610 19345 19612
rect 19369 19610 19425 19612
rect 19449 19610 19505 19612
rect 19529 19610 19585 19612
rect 19289 19558 19315 19610
rect 19315 19558 19345 19610
rect 19369 19558 19379 19610
rect 19379 19558 19425 19610
rect 19449 19558 19495 19610
rect 19495 19558 19505 19610
rect 19529 19558 19559 19610
rect 19559 19558 19585 19610
rect 19289 19556 19345 19558
rect 19369 19556 19425 19558
rect 19449 19556 19505 19558
rect 19529 19556 19585 19558
rect 19289 18522 19345 18524
rect 19369 18522 19425 18524
rect 19449 18522 19505 18524
rect 19529 18522 19585 18524
rect 19289 18470 19315 18522
rect 19315 18470 19345 18522
rect 19369 18470 19379 18522
rect 19379 18470 19425 18522
rect 19449 18470 19495 18522
rect 19495 18470 19505 18522
rect 19529 18470 19559 18522
rect 19559 18470 19585 18522
rect 19289 18468 19345 18470
rect 19369 18468 19425 18470
rect 19449 18468 19505 18470
rect 19529 18468 19585 18470
rect 19289 17434 19345 17436
rect 19369 17434 19425 17436
rect 19449 17434 19505 17436
rect 19529 17434 19585 17436
rect 19289 17382 19315 17434
rect 19315 17382 19345 17434
rect 19369 17382 19379 17434
rect 19379 17382 19425 17434
rect 19449 17382 19495 17434
rect 19495 17382 19505 17434
rect 19529 17382 19559 17434
rect 19559 17382 19585 17434
rect 19289 17380 19345 17382
rect 19369 17380 19425 17382
rect 19449 17380 19505 17382
rect 19529 17380 19585 17382
rect 19289 16346 19345 16348
rect 19369 16346 19425 16348
rect 19449 16346 19505 16348
rect 19529 16346 19585 16348
rect 19289 16294 19315 16346
rect 19315 16294 19345 16346
rect 19369 16294 19379 16346
rect 19379 16294 19425 16346
rect 19449 16294 19495 16346
rect 19495 16294 19505 16346
rect 19529 16294 19559 16346
rect 19559 16294 19585 16346
rect 19289 16292 19345 16294
rect 19369 16292 19425 16294
rect 19449 16292 19505 16294
rect 19529 16292 19585 16294
rect 19289 15258 19345 15260
rect 19369 15258 19425 15260
rect 19449 15258 19505 15260
rect 19529 15258 19585 15260
rect 19289 15206 19315 15258
rect 19315 15206 19345 15258
rect 19369 15206 19379 15258
rect 19379 15206 19425 15258
rect 19449 15206 19495 15258
rect 19495 15206 19505 15258
rect 19529 15206 19559 15258
rect 19559 15206 19585 15258
rect 19289 15204 19345 15206
rect 19369 15204 19425 15206
rect 19449 15204 19505 15206
rect 19529 15204 19585 15206
rect 19289 14170 19345 14172
rect 19369 14170 19425 14172
rect 19449 14170 19505 14172
rect 19529 14170 19585 14172
rect 19289 14118 19315 14170
rect 19315 14118 19345 14170
rect 19369 14118 19379 14170
rect 19379 14118 19425 14170
rect 19449 14118 19495 14170
rect 19495 14118 19505 14170
rect 19529 14118 19559 14170
rect 19559 14118 19585 14170
rect 19289 14116 19345 14118
rect 19369 14116 19425 14118
rect 19449 14116 19505 14118
rect 19529 14116 19585 14118
rect 19890 18944 19946 19000
rect 20442 17040 20498 17096
rect 19289 13082 19345 13084
rect 19369 13082 19425 13084
rect 19449 13082 19505 13084
rect 19529 13082 19585 13084
rect 19289 13030 19315 13082
rect 19315 13030 19345 13082
rect 19369 13030 19379 13082
rect 19379 13030 19425 13082
rect 19449 13030 19495 13082
rect 19495 13030 19505 13082
rect 19529 13030 19559 13082
rect 19559 13030 19585 13082
rect 19289 13028 19345 13030
rect 19369 13028 19425 13030
rect 19449 13028 19505 13030
rect 19529 13028 19585 13030
rect 19289 11994 19345 11996
rect 19369 11994 19425 11996
rect 19449 11994 19505 11996
rect 19529 11994 19585 11996
rect 19289 11942 19315 11994
rect 19315 11942 19345 11994
rect 19369 11942 19379 11994
rect 19379 11942 19425 11994
rect 19449 11942 19495 11994
rect 19495 11942 19505 11994
rect 19529 11942 19559 11994
rect 19559 11942 19585 11994
rect 19289 11940 19345 11942
rect 19369 11940 19425 11942
rect 19449 11940 19505 11942
rect 19529 11940 19585 11942
rect 19798 13776 19854 13832
rect 19289 10906 19345 10908
rect 19369 10906 19425 10908
rect 19449 10906 19505 10908
rect 19529 10906 19585 10908
rect 19289 10854 19315 10906
rect 19315 10854 19345 10906
rect 19369 10854 19379 10906
rect 19379 10854 19425 10906
rect 19449 10854 19495 10906
rect 19495 10854 19505 10906
rect 19529 10854 19559 10906
rect 19559 10854 19585 10906
rect 19289 10852 19345 10854
rect 19369 10852 19425 10854
rect 19449 10852 19505 10854
rect 19529 10852 19585 10854
rect 19289 9818 19345 9820
rect 19369 9818 19425 9820
rect 19449 9818 19505 9820
rect 19529 9818 19585 9820
rect 19289 9766 19315 9818
rect 19315 9766 19345 9818
rect 19369 9766 19379 9818
rect 19379 9766 19425 9818
rect 19449 9766 19495 9818
rect 19495 9766 19505 9818
rect 19529 9766 19559 9818
rect 19559 9766 19585 9818
rect 19289 9764 19345 9766
rect 19369 9764 19425 9766
rect 19449 9764 19505 9766
rect 19529 9764 19585 9766
rect 19289 8730 19345 8732
rect 19369 8730 19425 8732
rect 19449 8730 19505 8732
rect 19529 8730 19585 8732
rect 19289 8678 19315 8730
rect 19315 8678 19345 8730
rect 19369 8678 19379 8730
rect 19379 8678 19425 8730
rect 19449 8678 19495 8730
rect 19495 8678 19505 8730
rect 19529 8678 19559 8730
rect 19559 8678 19585 8730
rect 19289 8676 19345 8678
rect 19369 8676 19425 8678
rect 19449 8676 19505 8678
rect 19529 8676 19585 8678
rect 17314 5072 17370 5128
rect 17130 3168 17186 3224
rect 19289 7642 19345 7644
rect 19369 7642 19425 7644
rect 19449 7642 19505 7644
rect 19529 7642 19585 7644
rect 19289 7590 19315 7642
rect 19315 7590 19345 7642
rect 19369 7590 19379 7642
rect 19379 7590 19425 7642
rect 19449 7590 19495 7642
rect 19495 7590 19505 7642
rect 19529 7590 19559 7642
rect 19559 7590 19585 7642
rect 19289 7588 19345 7590
rect 19369 7588 19425 7590
rect 19449 7588 19505 7590
rect 19529 7588 19585 7590
rect 19522 7112 19578 7168
rect 19062 6704 19118 6760
rect 19289 6554 19345 6556
rect 19369 6554 19425 6556
rect 19449 6554 19505 6556
rect 19529 6554 19585 6556
rect 19289 6502 19315 6554
rect 19315 6502 19345 6554
rect 19369 6502 19379 6554
rect 19379 6502 19425 6554
rect 19449 6502 19495 6554
rect 19495 6502 19505 6554
rect 19529 6502 19559 6554
rect 19559 6502 19585 6554
rect 19289 6500 19345 6502
rect 19369 6500 19425 6502
rect 19449 6500 19505 6502
rect 19529 6500 19585 6502
rect 18510 4392 18566 4448
rect 11886 1944 11942 2000
rect 15198 1808 15254 1864
rect 18234 2488 18290 2544
rect 18602 2352 18658 2408
rect 18050 1672 18106 1728
rect 19289 5466 19345 5468
rect 19369 5466 19425 5468
rect 19449 5466 19505 5468
rect 19529 5466 19585 5468
rect 19289 5414 19315 5466
rect 19315 5414 19345 5466
rect 19369 5414 19379 5466
rect 19379 5414 19425 5466
rect 19449 5414 19495 5466
rect 19495 5414 19505 5466
rect 19529 5414 19559 5466
rect 19559 5414 19585 5466
rect 19289 5412 19345 5414
rect 19369 5412 19425 5414
rect 19449 5412 19505 5414
rect 19529 5412 19585 5414
rect 19289 4378 19345 4380
rect 19369 4378 19425 4380
rect 19449 4378 19505 4380
rect 19529 4378 19585 4380
rect 19289 4326 19315 4378
rect 19315 4326 19345 4378
rect 19369 4326 19379 4378
rect 19379 4326 19425 4378
rect 19449 4326 19495 4378
rect 19495 4326 19505 4378
rect 19529 4326 19559 4378
rect 19559 4326 19585 4378
rect 19289 4324 19345 4326
rect 19369 4324 19425 4326
rect 19449 4324 19505 4326
rect 19529 4324 19585 4326
rect 19706 4120 19762 4176
rect 19289 3290 19345 3292
rect 19369 3290 19425 3292
rect 19449 3290 19505 3292
rect 19529 3290 19585 3292
rect 19289 3238 19315 3290
rect 19315 3238 19345 3290
rect 19369 3238 19379 3290
rect 19379 3238 19425 3290
rect 19449 3238 19495 3290
rect 19495 3238 19505 3290
rect 19529 3238 19559 3290
rect 19559 3238 19585 3290
rect 19289 3236 19345 3238
rect 19369 3236 19425 3238
rect 19449 3236 19505 3238
rect 19529 3236 19585 3238
rect 19289 2202 19345 2204
rect 19369 2202 19425 2204
rect 19449 2202 19505 2204
rect 19529 2202 19585 2204
rect 19289 2150 19315 2202
rect 19315 2150 19345 2202
rect 19369 2150 19379 2202
rect 19379 2150 19425 2202
rect 19449 2150 19495 2202
rect 19495 2150 19505 2202
rect 19529 2150 19559 2202
rect 19559 2150 19585 2202
rect 19289 2148 19345 2150
rect 19369 2148 19425 2150
rect 19449 2148 19505 2150
rect 19529 2148 19585 2150
rect 18694 992 18750 1048
rect 21638 18536 21694 18592
rect 21546 17584 21602 17640
rect 21546 16632 21602 16688
rect 21546 8064 21602 8120
<< metal3 >>
rect 21520 21360 22000 21480
rect 0 20952 480 21072
rect 62 20498 122 20952
rect 14457 20906 14523 20909
rect 21590 20906 21650 21360
rect 14457 20904 21650 20906
rect 14457 20848 14462 20904
rect 14518 20848 21650 20904
rect 14457 20846 21650 20848
rect 14457 20843 14523 20846
rect 2497 20498 2563 20501
rect 62 20496 2563 20498
rect 62 20440 2502 20496
rect 2558 20440 2563 20496
rect 62 20438 2563 20440
rect 2497 20435 2563 20438
rect 21520 20408 22000 20528
rect 15745 19954 15811 19957
rect 21590 19954 21650 20408
rect 15745 19952 21650 19954
rect 15745 19896 15750 19952
rect 15806 19896 21650 19952
rect 15745 19894 21650 19896
rect 15745 19891 15811 19894
rect 4610 19616 4930 19617
rect 4610 19552 4618 19616
rect 4682 19552 4698 19616
rect 4762 19552 4778 19616
rect 4842 19552 4858 19616
rect 4922 19552 4930 19616
rect 4610 19551 4930 19552
rect 11944 19616 12264 19617
rect 11944 19552 11952 19616
rect 12016 19552 12032 19616
rect 12096 19552 12112 19616
rect 12176 19552 12192 19616
rect 12256 19552 12264 19616
rect 11944 19551 12264 19552
rect 19277 19616 19597 19617
rect 19277 19552 19285 19616
rect 19349 19552 19365 19616
rect 19429 19552 19445 19616
rect 19509 19552 19525 19616
rect 19589 19552 19597 19616
rect 19277 19551 19597 19552
rect 21520 19456 22000 19576
rect 0 19184 480 19304
rect 62 18730 122 19184
rect 8277 19072 8597 19073
rect 8277 19008 8285 19072
rect 8349 19008 8365 19072
rect 8429 19008 8445 19072
rect 8509 19008 8525 19072
rect 8589 19008 8597 19072
rect 8277 19007 8597 19008
rect 15610 19072 15930 19073
rect 15610 19008 15618 19072
rect 15682 19008 15698 19072
rect 15762 19008 15778 19072
rect 15842 19008 15858 19072
rect 15922 19008 15930 19072
rect 15610 19007 15930 19008
rect 19885 19002 19951 19005
rect 21590 19002 21650 19456
rect 19885 19000 21650 19002
rect 19885 18944 19890 19000
rect 19946 18944 21650 19000
rect 19885 18942 21650 18944
rect 19885 18939 19951 18942
rect 1577 18730 1643 18733
rect 62 18728 1643 18730
rect 62 18672 1582 18728
rect 1638 18672 1643 18728
rect 62 18670 1643 18672
rect 1577 18667 1643 18670
rect 21520 18592 22000 18624
rect 21520 18536 21638 18592
rect 21694 18536 22000 18592
rect 4610 18528 4930 18529
rect 4610 18464 4618 18528
rect 4682 18464 4698 18528
rect 4762 18464 4778 18528
rect 4842 18464 4858 18528
rect 4922 18464 4930 18528
rect 4610 18463 4930 18464
rect 11944 18528 12264 18529
rect 11944 18464 11952 18528
rect 12016 18464 12032 18528
rect 12096 18464 12112 18528
rect 12176 18464 12192 18528
rect 12256 18464 12264 18528
rect 11944 18463 12264 18464
rect 19277 18528 19597 18529
rect 19277 18464 19285 18528
rect 19349 18464 19365 18528
rect 19429 18464 19445 18528
rect 19509 18464 19525 18528
rect 19589 18464 19597 18528
rect 21520 18504 22000 18536
rect 19277 18463 19597 18464
rect 8277 17984 8597 17985
rect 8277 17920 8285 17984
rect 8349 17920 8365 17984
rect 8429 17920 8445 17984
rect 8509 17920 8525 17984
rect 8589 17920 8597 17984
rect 8277 17919 8597 17920
rect 15610 17984 15930 17985
rect 15610 17920 15618 17984
rect 15682 17920 15698 17984
rect 15762 17920 15778 17984
rect 15842 17920 15858 17984
rect 15922 17920 15930 17984
rect 15610 17919 15930 17920
rect 7005 17778 7071 17781
rect 13813 17778 13879 17781
rect 7005 17776 13879 17778
rect 7005 17720 7010 17776
rect 7066 17720 13818 17776
rect 13874 17720 13879 17776
rect 7005 17718 13879 17720
rect 7005 17715 7071 17718
rect 13813 17715 13879 17718
rect 21520 17642 22000 17672
rect 21460 17640 22000 17642
rect 21460 17584 21546 17640
rect 21602 17584 22000 17640
rect 21460 17582 22000 17584
rect 21520 17552 22000 17582
rect 4610 17440 4930 17441
rect 0 17280 480 17400
rect 4610 17376 4618 17440
rect 4682 17376 4698 17440
rect 4762 17376 4778 17440
rect 4842 17376 4858 17440
rect 4922 17376 4930 17440
rect 4610 17375 4930 17376
rect 11944 17440 12264 17441
rect 11944 17376 11952 17440
rect 12016 17376 12032 17440
rect 12096 17376 12112 17440
rect 12176 17376 12192 17440
rect 12256 17376 12264 17440
rect 11944 17375 12264 17376
rect 19277 17440 19597 17441
rect 19277 17376 19285 17440
rect 19349 17376 19365 17440
rect 19429 17376 19445 17440
rect 19509 17376 19525 17440
rect 19589 17376 19597 17440
rect 19277 17375 19597 17376
rect 12709 17370 12775 17373
rect 15929 17370 15995 17373
rect 12709 17368 15995 17370
rect 12709 17312 12714 17368
rect 12770 17312 15934 17368
rect 15990 17312 15995 17368
rect 12709 17310 15995 17312
rect 12709 17307 12775 17310
rect 15929 17307 15995 17310
rect 62 16826 122 17280
rect 4981 17234 5047 17237
rect 14365 17234 14431 17237
rect 4981 17232 14431 17234
rect 4981 17176 4986 17232
rect 5042 17176 14370 17232
rect 14426 17176 14431 17232
rect 4981 17174 14431 17176
rect 4981 17171 5047 17174
rect 14365 17171 14431 17174
rect 11053 17098 11119 17101
rect 20437 17098 20503 17101
rect 11053 17096 20503 17098
rect 11053 17040 11058 17096
rect 11114 17040 20442 17096
rect 20498 17040 20503 17096
rect 11053 17038 20503 17040
rect 11053 17035 11119 17038
rect 20437 17035 20503 17038
rect 8277 16896 8597 16897
rect 8277 16832 8285 16896
rect 8349 16832 8365 16896
rect 8429 16832 8445 16896
rect 8509 16832 8525 16896
rect 8589 16832 8597 16896
rect 8277 16831 8597 16832
rect 15610 16896 15930 16897
rect 15610 16832 15618 16896
rect 15682 16832 15698 16896
rect 15762 16832 15778 16896
rect 15842 16832 15858 16896
rect 15922 16832 15930 16896
rect 15610 16831 15930 16832
rect 1577 16826 1643 16829
rect 62 16824 1643 16826
rect 62 16768 1582 16824
rect 1638 16768 1643 16824
rect 62 16766 1643 16768
rect 1577 16763 1643 16766
rect 21520 16690 22000 16720
rect 21460 16688 22000 16690
rect 21460 16632 21546 16688
rect 21602 16632 22000 16688
rect 21460 16630 22000 16632
rect 21520 16600 22000 16630
rect 4610 16352 4930 16353
rect 4610 16288 4618 16352
rect 4682 16288 4698 16352
rect 4762 16288 4778 16352
rect 4842 16288 4858 16352
rect 4922 16288 4930 16352
rect 4610 16287 4930 16288
rect 11944 16352 12264 16353
rect 11944 16288 11952 16352
rect 12016 16288 12032 16352
rect 12096 16288 12112 16352
rect 12176 16288 12192 16352
rect 12256 16288 12264 16352
rect 11944 16287 12264 16288
rect 19277 16352 19597 16353
rect 19277 16288 19285 16352
rect 19349 16288 19365 16352
rect 19429 16288 19445 16352
rect 19509 16288 19525 16352
rect 19589 16288 19597 16352
rect 19277 16287 19597 16288
rect 9029 16010 9095 16013
rect 14825 16010 14891 16013
rect 9029 16008 14891 16010
rect 9029 15952 9034 16008
rect 9090 15952 14830 16008
rect 14886 15952 14891 16008
rect 9029 15950 14891 15952
rect 9029 15947 9095 15950
rect 14825 15947 14891 15950
rect 8277 15808 8597 15809
rect 8277 15744 8285 15808
rect 8349 15744 8365 15808
rect 8429 15744 8445 15808
rect 8509 15744 8525 15808
rect 8589 15744 8597 15808
rect 8277 15743 8597 15744
rect 15610 15808 15930 15809
rect 15610 15744 15618 15808
rect 15682 15744 15698 15808
rect 15762 15744 15778 15808
rect 15842 15744 15858 15808
rect 15922 15744 15930 15808
rect 15610 15743 15930 15744
rect 21520 15648 22000 15768
rect 0 15512 480 15632
rect 5257 15602 5323 15605
rect 14917 15602 14983 15605
rect 5257 15600 14983 15602
rect 5257 15544 5262 15600
rect 5318 15544 14922 15600
rect 14978 15544 14983 15600
rect 5257 15542 14983 15544
rect 5257 15539 5323 15542
rect 14917 15539 14983 15542
rect 62 15058 122 15512
rect 6269 15466 6335 15469
rect 14089 15466 14155 15469
rect 6269 15464 14155 15466
rect 6269 15408 6274 15464
rect 6330 15408 14094 15464
rect 14150 15408 14155 15464
rect 6269 15406 14155 15408
rect 6269 15403 6335 15406
rect 14089 15403 14155 15406
rect 17033 15466 17099 15469
rect 21590 15466 21650 15648
rect 17033 15464 21650 15466
rect 17033 15408 17038 15464
rect 17094 15408 21650 15464
rect 17033 15406 21650 15408
rect 17033 15403 17099 15406
rect 4610 15264 4930 15265
rect 4610 15200 4618 15264
rect 4682 15200 4698 15264
rect 4762 15200 4778 15264
rect 4842 15200 4858 15264
rect 4922 15200 4930 15264
rect 4610 15199 4930 15200
rect 11944 15264 12264 15265
rect 11944 15200 11952 15264
rect 12016 15200 12032 15264
rect 12096 15200 12112 15264
rect 12176 15200 12192 15264
rect 12256 15200 12264 15264
rect 11944 15199 12264 15200
rect 19277 15264 19597 15265
rect 19277 15200 19285 15264
rect 19349 15200 19365 15264
rect 19429 15200 19445 15264
rect 19509 15200 19525 15264
rect 19589 15200 19597 15264
rect 19277 15199 19597 15200
rect 3325 15058 3391 15061
rect 62 15056 3391 15058
rect 62 15000 3330 15056
rect 3386 15000 3391 15056
rect 62 14998 3391 15000
rect 3325 14995 3391 14998
rect 5165 15058 5231 15061
rect 10961 15058 11027 15061
rect 16849 15058 16915 15061
rect 5165 15056 16915 15058
rect 5165 15000 5170 15056
rect 5226 15000 10966 15056
rect 11022 15000 16854 15056
rect 16910 15000 16915 15056
rect 5165 14998 16915 15000
rect 5165 14995 5231 14998
rect 10961 14995 11027 14998
rect 16849 14995 16915 14998
rect 4337 14922 4403 14925
rect 15469 14922 15535 14925
rect 4337 14920 15535 14922
rect 4337 14864 4342 14920
rect 4398 14864 15474 14920
rect 15530 14864 15535 14920
rect 4337 14862 15535 14864
rect 4337 14859 4403 14862
rect 15469 14859 15535 14862
rect 21520 14788 22000 14816
rect 21520 14786 21588 14788
rect 21460 14726 21588 14786
rect 21520 14724 21588 14726
rect 21652 14724 22000 14788
rect 8277 14720 8597 14721
rect 8277 14656 8285 14720
rect 8349 14656 8365 14720
rect 8429 14656 8445 14720
rect 8509 14656 8525 14720
rect 8589 14656 8597 14720
rect 8277 14655 8597 14656
rect 15610 14720 15930 14721
rect 15610 14656 15618 14720
rect 15682 14656 15698 14720
rect 15762 14656 15778 14720
rect 15842 14656 15858 14720
rect 15922 14656 15930 14720
rect 21520 14696 22000 14724
rect 15610 14655 15930 14656
rect 16021 14650 16087 14653
rect 21398 14650 21404 14652
rect 16021 14648 21404 14650
rect 16021 14592 16026 14648
rect 16082 14592 21404 14648
rect 16021 14590 21404 14592
rect 16021 14587 16087 14590
rect 21398 14588 21404 14590
rect 21468 14588 21474 14652
rect 4610 14176 4930 14177
rect 4610 14112 4618 14176
rect 4682 14112 4698 14176
rect 4762 14112 4778 14176
rect 4842 14112 4858 14176
rect 4922 14112 4930 14176
rect 4610 14111 4930 14112
rect 11944 14176 12264 14177
rect 11944 14112 11952 14176
rect 12016 14112 12032 14176
rect 12096 14112 12112 14176
rect 12176 14112 12192 14176
rect 12256 14112 12264 14176
rect 11944 14111 12264 14112
rect 19277 14176 19597 14177
rect 19277 14112 19285 14176
rect 19349 14112 19365 14176
rect 19429 14112 19445 14176
rect 19509 14112 19525 14176
rect 19589 14112 19597 14176
rect 19277 14111 19597 14112
rect 5625 13834 5691 13837
rect 9489 13834 9555 13837
rect 10041 13834 10107 13837
rect 5625 13832 10107 13834
rect 5625 13776 5630 13832
rect 5686 13776 9494 13832
rect 9550 13776 10046 13832
rect 10102 13776 10107 13832
rect 5625 13774 10107 13776
rect 5625 13771 5691 13774
rect 9489 13771 9555 13774
rect 10041 13771 10107 13774
rect 14733 13834 14799 13837
rect 15101 13834 15167 13837
rect 19793 13834 19859 13837
rect 21520 13834 22000 13864
rect 14733 13832 22000 13834
rect 14733 13776 14738 13832
rect 14794 13776 15106 13832
rect 15162 13776 19798 13832
rect 19854 13776 22000 13832
rect 14733 13774 22000 13776
rect 14733 13771 14799 13774
rect 15101 13771 15167 13774
rect 19793 13771 19859 13774
rect 21520 13744 22000 13774
rect 0 13700 480 13728
rect 0 13636 60 13700
rect 124 13636 480 13700
rect 0 13608 480 13636
rect 6269 13698 6335 13701
rect 6821 13698 6887 13701
rect 6269 13696 6887 13698
rect 6269 13640 6274 13696
rect 6330 13640 6826 13696
rect 6882 13640 6887 13696
rect 6269 13638 6887 13640
rect 6269 13635 6335 13638
rect 6821 13635 6887 13638
rect 8277 13632 8597 13633
rect 8277 13568 8285 13632
rect 8349 13568 8365 13632
rect 8429 13568 8445 13632
rect 8509 13568 8525 13632
rect 8589 13568 8597 13632
rect 8277 13567 8597 13568
rect 15610 13632 15930 13633
rect 15610 13568 15618 13632
rect 15682 13568 15698 13632
rect 15762 13568 15778 13632
rect 15842 13568 15858 13632
rect 15922 13568 15930 13632
rect 15610 13567 15930 13568
rect 54 13364 60 13428
rect 124 13426 130 13428
rect 1301 13426 1367 13429
rect 124 13424 1367 13426
rect 124 13368 1306 13424
rect 1362 13368 1367 13424
rect 124 13366 1367 13368
rect 124 13364 130 13366
rect 1301 13363 1367 13366
rect 5165 13426 5231 13429
rect 10225 13426 10291 13429
rect 5165 13424 10291 13426
rect 5165 13368 5170 13424
rect 5226 13368 10230 13424
rect 10286 13368 10291 13424
rect 5165 13366 10291 13368
rect 5165 13363 5231 13366
rect 10225 13363 10291 13366
rect 2405 13290 2471 13293
rect 12893 13290 12959 13293
rect 2405 13288 12959 13290
rect 2405 13232 2410 13288
rect 2466 13232 12898 13288
rect 12954 13232 12959 13288
rect 2405 13230 12959 13232
rect 2405 13227 2471 13230
rect 12893 13227 12959 13230
rect 5809 13154 5875 13157
rect 9857 13154 9923 13157
rect 5682 13152 9923 13154
rect 5682 13096 5814 13152
rect 5870 13096 9862 13152
rect 9918 13096 9923 13152
rect 5682 13094 9923 13096
rect 5809 13091 5875 13094
rect 9857 13091 9923 13094
rect 4610 13088 4930 13089
rect 4610 13024 4618 13088
rect 4682 13024 4698 13088
rect 4762 13024 4778 13088
rect 4842 13024 4858 13088
rect 4922 13024 4930 13088
rect 4610 13023 4930 13024
rect 11944 13088 12264 13089
rect 11944 13024 11952 13088
rect 12016 13024 12032 13088
rect 12096 13024 12112 13088
rect 12176 13024 12192 13088
rect 12256 13024 12264 13088
rect 11944 13023 12264 13024
rect 19277 13088 19597 13089
rect 19277 13024 19285 13088
rect 19349 13024 19365 13088
rect 19429 13024 19445 13088
rect 19509 13024 19525 13088
rect 19589 13024 19597 13088
rect 19277 13023 19597 13024
rect 4981 12882 5047 12885
rect 6126 12882 6132 12884
rect 4981 12880 6132 12882
rect 4981 12824 4986 12880
rect 5042 12824 6132 12880
rect 4981 12822 6132 12824
rect 4981 12819 5047 12822
rect 6126 12820 6132 12822
rect 6196 12820 6202 12884
rect 21520 12792 22000 12912
rect 6361 12746 6427 12749
rect 17033 12746 17099 12749
rect 6361 12744 17099 12746
rect 6361 12688 6366 12744
rect 6422 12688 17038 12744
rect 17094 12688 17099 12744
rect 6361 12686 17099 12688
rect 6361 12683 6427 12686
rect 17033 12683 17099 12686
rect 8277 12544 8597 12545
rect 8277 12480 8285 12544
rect 8349 12480 8365 12544
rect 8429 12480 8445 12544
rect 8509 12480 8525 12544
rect 8589 12480 8597 12544
rect 8277 12479 8597 12480
rect 15610 12544 15930 12545
rect 15610 12480 15618 12544
rect 15682 12480 15698 12544
rect 15762 12480 15778 12544
rect 15842 12480 15858 12544
rect 15922 12480 15930 12544
rect 15610 12479 15930 12480
rect 14089 12338 14155 12341
rect 21590 12338 21650 12792
rect 14089 12336 21650 12338
rect 14089 12280 14094 12336
rect 14150 12280 21650 12336
rect 14089 12278 21650 12280
rect 14089 12275 14155 12278
rect 4610 12000 4930 12001
rect 0 11840 480 11960
rect 4610 11936 4618 12000
rect 4682 11936 4698 12000
rect 4762 11936 4778 12000
rect 4842 11936 4858 12000
rect 4922 11936 4930 12000
rect 4610 11935 4930 11936
rect 11944 12000 12264 12001
rect 11944 11936 11952 12000
rect 12016 11936 12032 12000
rect 12096 11936 12112 12000
rect 12176 11936 12192 12000
rect 12256 11936 12264 12000
rect 11944 11935 12264 11936
rect 19277 12000 19597 12001
rect 19277 11936 19285 12000
rect 19349 11936 19365 12000
rect 19429 11936 19445 12000
rect 19509 11936 19525 12000
rect 19589 11936 19597 12000
rect 19277 11935 19597 11936
rect 21520 11840 22000 11960
rect 62 11522 122 11840
rect 1577 11522 1643 11525
rect 62 11520 1643 11522
rect 62 11464 1582 11520
rect 1638 11464 1643 11520
rect 62 11462 1643 11464
rect 1577 11459 1643 11462
rect 8277 11456 8597 11457
rect 8277 11392 8285 11456
rect 8349 11392 8365 11456
rect 8429 11392 8445 11456
rect 8509 11392 8525 11456
rect 8589 11392 8597 11456
rect 8277 11391 8597 11392
rect 15610 11456 15930 11457
rect 15610 11392 15618 11456
rect 15682 11392 15698 11456
rect 15762 11392 15778 11456
rect 15842 11392 15858 11456
rect 15922 11392 15930 11456
rect 15610 11391 15930 11392
rect 3141 11386 3207 11389
rect 7373 11386 7439 11389
rect 3141 11384 7439 11386
rect 3141 11328 3146 11384
rect 3202 11328 7378 11384
rect 7434 11328 7439 11384
rect 3141 11326 7439 11328
rect 3141 11323 3207 11326
rect 7373 11323 7439 11326
rect 16389 11386 16455 11389
rect 21590 11386 21650 11840
rect 16389 11384 21650 11386
rect 16389 11328 16394 11384
rect 16450 11328 21650 11384
rect 16389 11326 21650 11328
rect 16389 11323 16455 11326
rect 3509 11250 3575 11253
rect 11237 11250 11303 11253
rect 3509 11248 11303 11250
rect 3509 11192 3514 11248
rect 3570 11192 11242 11248
rect 11298 11192 11303 11248
rect 3509 11190 11303 11192
rect 3509 11187 3575 11190
rect 11237 11187 11303 11190
rect 3049 11114 3115 11117
rect 10317 11114 10383 11117
rect 3049 11112 10383 11114
rect 3049 11056 3054 11112
rect 3110 11056 10322 11112
rect 10378 11056 10383 11112
rect 3049 11054 10383 11056
rect 3049 11051 3115 11054
rect 10317 11051 10383 11054
rect 4610 10912 4930 10913
rect 4610 10848 4618 10912
rect 4682 10848 4698 10912
rect 4762 10848 4778 10912
rect 4842 10848 4858 10912
rect 4922 10848 4930 10912
rect 4610 10847 4930 10848
rect 11944 10912 12264 10913
rect 11944 10848 11952 10912
rect 12016 10848 12032 10912
rect 12096 10848 12112 10912
rect 12176 10848 12192 10912
rect 12256 10848 12264 10912
rect 11944 10847 12264 10848
rect 19277 10912 19597 10913
rect 19277 10848 19285 10912
rect 19349 10848 19365 10912
rect 19429 10848 19445 10912
rect 19509 10848 19525 10912
rect 19589 10848 19597 10912
rect 21520 10888 22000 11008
rect 19277 10847 19597 10848
rect 6085 10842 6151 10845
rect 7097 10842 7163 10845
rect 9765 10842 9831 10845
rect 6085 10840 9831 10842
rect 6085 10784 6090 10840
rect 6146 10784 7102 10840
rect 7158 10784 9770 10840
rect 9826 10784 9831 10840
rect 6085 10782 9831 10784
rect 6085 10779 6151 10782
rect 7097 10779 7163 10782
rect 9765 10779 9831 10782
rect 3325 10706 3391 10709
rect 8109 10706 8175 10709
rect 3325 10704 8175 10706
rect 3325 10648 3330 10704
rect 3386 10648 8114 10704
rect 8170 10648 8175 10704
rect 3325 10646 8175 10648
rect 3325 10643 3391 10646
rect 8109 10643 8175 10646
rect 8753 10706 8819 10709
rect 14273 10706 14339 10709
rect 8753 10704 14339 10706
rect 8753 10648 8758 10704
rect 8814 10648 14278 10704
rect 14334 10648 14339 10704
rect 8753 10646 14339 10648
rect 8753 10643 8819 10646
rect 14273 10643 14339 10646
rect 6453 10570 6519 10573
rect 12617 10570 12683 10573
rect 6453 10568 12683 10570
rect 6453 10512 6458 10568
rect 6514 10512 12622 10568
rect 12678 10512 12683 10568
rect 6453 10510 12683 10512
rect 6453 10507 6519 10510
rect 12617 10507 12683 10510
rect 15929 10570 15995 10573
rect 21590 10570 21650 10888
rect 15929 10568 21650 10570
rect 15929 10512 15934 10568
rect 15990 10512 21650 10568
rect 15929 10510 21650 10512
rect 15929 10507 15995 10510
rect 9949 10434 10015 10437
rect 10777 10434 10843 10437
rect 15469 10434 15535 10437
rect 9949 10432 15535 10434
rect 9949 10376 9954 10432
rect 10010 10376 10782 10432
rect 10838 10376 15474 10432
rect 15530 10376 15535 10432
rect 9949 10374 15535 10376
rect 9949 10371 10015 10374
rect 10777 10371 10843 10374
rect 15469 10371 15535 10374
rect 8277 10368 8597 10369
rect 8277 10304 8285 10368
rect 8349 10304 8365 10368
rect 8429 10304 8445 10368
rect 8509 10304 8525 10368
rect 8589 10304 8597 10368
rect 8277 10303 8597 10304
rect 15610 10368 15930 10369
rect 15610 10304 15618 10368
rect 15682 10304 15698 10368
rect 15762 10304 15778 10368
rect 15842 10304 15858 10368
rect 15922 10304 15930 10368
rect 15610 10303 15930 10304
rect 1945 10162 2011 10165
rect 7557 10162 7623 10165
rect 1945 10160 7623 10162
rect 1945 10104 1950 10160
rect 2006 10104 7562 10160
rect 7618 10104 7623 10160
rect 1945 10102 7623 10104
rect 1945 10099 2011 10102
rect 7557 10099 7623 10102
rect 11513 10162 11579 10165
rect 16389 10162 16455 10165
rect 11513 10160 16455 10162
rect 11513 10104 11518 10160
rect 11574 10104 16394 10160
rect 16450 10104 16455 10160
rect 11513 10102 16455 10104
rect 11513 10099 11579 10102
rect 16389 10099 16455 10102
rect 0 9936 480 10056
rect 5717 10026 5783 10029
rect 12433 10026 12499 10029
rect 21520 10026 22000 10056
rect 5717 10024 12499 10026
rect 5717 9968 5722 10024
rect 5778 9968 12438 10024
rect 12494 9968 12499 10024
rect 5717 9966 12499 9968
rect 5717 9963 5783 9966
rect 12433 9963 12499 9966
rect 13770 9966 22000 10026
rect 62 9754 122 9936
rect 12801 9890 12867 9893
rect 13770 9890 13830 9966
rect 21520 9936 22000 9966
rect 12801 9888 13830 9890
rect 12801 9832 12806 9888
rect 12862 9832 13830 9888
rect 12801 9830 13830 9832
rect 12801 9827 12867 9830
rect 4610 9824 4930 9825
rect 4610 9760 4618 9824
rect 4682 9760 4698 9824
rect 4762 9760 4778 9824
rect 4842 9760 4858 9824
rect 4922 9760 4930 9824
rect 4610 9759 4930 9760
rect 11944 9824 12264 9825
rect 11944 9760 11952 9824
rect 12016 9760 12032 9824
rect 12096 9760 12112 9824
rect 12176 9760 12192 9824
rect 12256 9760 12264 9824
rect 11944 9759 12264 9760
rect 19277 9824 19597 9825
rect 19277 9760 19285 9824
rect 19349 9760 19365 9824
rect 19429 9760 19445 9824
rect 19509 9760 19525 9824
rect 19589 9760 19597 9824
rect 19277 9759 19597 9760
rect 1577 9754 1643 9757
rect 62 9752 1643 9754
rect 62 9696 1582 9752
rect 1638 9696 1643 9752
rect 62 9694 1643 9696
rect 1577 9691 1643 9694
rect 3417 9346 3483 9349
rect 8109 9346 8175 9349
rect 3417 9344 8175 9346
rect 3417 9288 3422 9344
rect 3478 9288 8114 9344
rect 8170 9288 8175 9344
rect 3417 9286 8175 9288
rect 3417 9283 3483 9286
rect 8109 9283 8175 9286
rect 8277 9280 8597 9281
rect 8277 9216 8285 9280
rect 8349 9216 8365 9280
rect 8429 9216 8445 9280
rect 8509 9216 8525 9280
rect 8589 9216 8597 9280
rect 8277 9215 8597 9216
rect 15610 9280 15930 9281
rect 15610 9216 15618 9280
rect 15682 9216 15698 9280
rect 15762 9216 15778 9280
rect 15842 9216 15858 9280
rect 15922 9216 15930 9280
rect 15610 9215 15930 9216
rect 4061 9074 4127 9077
rect 5441 9074 5507 9077
rect 21520 9076 22000 9104
rect 21520 9074 21588 9076
rect 4061 9072 5507 9074
rect 4061 9016 4066 9072
rect 4122 9016 5446 9072
rect 5502 9016 5507 9072
rect 4061 9014 5507 9016
rect 21460 9014 21588 9074
rect 4061 9011 4127 9014
rect 5441 9011 5507 9014
rect 21520 9012 21588 9014
rect 21652 9012 22000 9076
rect 21520 8984 22000 9012
rect 11789 8938 11855 8941
rect 11789 8936 21466 8938
rect 11789 8880 11794 8936
rect 11850 8904 21466 8936
rect 21582 8904 21588 8906
rect 11850 8880 21588 8904
rect 11789 8878 21588 8880
rect 11789 8875 11855 8878
rect 21406 8844 21588 8878
rect 21582 8842 21588 8844
rect 21652 8842 21658 8906
rect 3049 8802 3115 8805
rect 62 8800 3115 8802
rect 62 8744 3054 8800
rect 3110 8744 3115 8800
rect 62 8742 3115 8744
rect 62 8288 122 8742
rect 3049 8739 3115 8742
rect 4610 8736 4930 8737
rect 4610 8672 4618 8736
rect 4682 8672 4698 8736
rect 4762 8672 4778 8736
rect 4842 8672 4858 8736
rect 4922 8672 4930 8736
rect 4610 8671 4930 8672
rect 11944 8736 12264 8737
rect 11944 8672 11952 8736
rect 12016 8672 12032 8736
rect 12096 8672 12112 8736
rect 12176 8672 12192 8736
rect 12256 8672 12264 8736
rect 11944 8671 12264 8672
rect 19277 8736 19597 8737
rect 19277 8672 19285 8736
rect 19349 8672 19365 8736
rect 19429 8672 19445 8736
rect 19509 8672 19525 8736
rect 19589 8672 19597 8736
rect 19277 8671 19597 8672
rect 1945 8530 2011 8533
rect 9949 8530 10015 8533
rect 1945 8528 10015 8530
rect 1945 8472 1950 8528
rect 2006 8472 9954 8528
rect 10010 8472 10015 8528
rect 1945 8470 10015 8472
rect 1945 8467 2011 8470
rect 9949 8467 10015 8470
rect 0 8168 480 8288
rect 8277 8192 8597 8193
rect 8277 8128 8285 8192
rect 8349 8128 8365 8192
rect 8429 8128 8445 8192
rect 8509 8128 8525 8192
rect 8589 8128 8597 8192
rect 8277 8127 8597 8128
rect 15610 8192 15930 8193
rect 15610 8128 15618 8192
rect 15682 8128 15698 8192
rect 15762 8128 15778 8192
rect 15842 8128 15858 8192
rect 15922 8128 15930 8192
rect 15610 8127 15930 8128
rect 7649 8122 7715 8125
rect 8109 8122 8175 8125
rect 21520 8122 22000 8152
rect 7649 8120 8175 8122
rect 7649 8064 7654 8120
rect 7710 8064 8114 8120
rect 8170 8064 8175 8120
rect 7649 8062 8175 8064
rect 21460 8120 22000 8122
rect 21460 8064 21546 8120
rect 21602 8064 22000 8120
rect 21460 8062 22000 8064
rect 7649 8059 7715 8062
rect 8109 8059 8175 8062
rect 21520 8032 22000 8062
rect 2589 7986 2655 7989
rect 8661 7986 8727 7989
rect 2589 7984 8727 7986
rect 2589 7928 2594 7984
rect 2650 7928 8666 7984
rect 8722 7928 8727 7984
rect 2589 7926 8727 7928
rect 2589 7923 2655 7926
rect 8661 7923 8727 7926
rect 5809 7850 5875 7853
rect 17125 7850 17191 7853
rect 5809 7848 17191 7850
rect 5809 7792 5814 7848
rect 5870 7792 17130 7848
rect 17186 7792 17191 7848
rect 5809 7790 17191 7792
rect 5809 7787 5875 7790
rect 17125 7787 17191 7790
rect 4610 7648 4930 7649
rect 4610 7584 4618 7648
rect 4682 7584 4698 7648
rect 4762 7584 4778 7648
rect 4842 7584 4858 7648
rect 4922 7584 4930 7648
rect 4610 7583 4930 7584
rect 11944 7648 12264 7649
rect 11944 7584 11952 7648
rect 12016 7584 12032 7648
rect 12096 7584 12112 7648
rect 12176 7584 12192 7648
rect 12256 7584 12264 7648
rect 11944 7583 12264 7584
rect 19277 7648 19597 7649
rect 19277 7584 19285 7648
rect 19349 7584 19365 7648
rect 19429 7584 19445 7648
rect 19509 7584 19525 7648
rect 19589 7584 19597 7648
rect 19277 7583 19597 7584
rect 3785 7442 3851 7445
rect 5441 7442 5507 7445
rect 3785 7440 5507 7442
rect 3785 7384 3790 7440
rect 3846 7384 5446 7440
rect 5502 7384 5507 7440
rect 3785 7382 5507 7384
rect 3785 7379 3851 7382
rect 5441 7379 5507 7382
rect 9673 7442 9739 7445
rect 10593 7442 10659 7445
rect 9673 7440 10659 7442
rect 9673 7384 9678 7440
rect 9734 7384 10598 7440
rect 10654 7384 10659 7440
rect 9673 7382 10659 7384
rect 9673 7379 9739 7382
rect 10593 7379 10659 7382
rect 19517 7170 19583 7173
rect 21520 7170 22000 7200
rect 19517 7168 22000 7170
rect 19517 7112 19522 7168
rect 19578 7112 22000 7168
rect 19517 7110 22000 7112
rect 19517 7107 19583 7110
rect 8277 7104 8597 7105
rect 8277 7040 8285 7104
rect 8349 7040 8365 7104
rect 8429 7040 8445 7104
rect 8509 7040 8525 7104
rect 8589 7040 8597 7104
rect 8277 7039 8597 7040
rect 15610 7104 15930 7105
rect 15610 7040 15618 7104
rect 15682 7040 15698 7104
rect 15762 7040 15778 7104
rect 15842 7040 15858 7104
rect 15922 7040 15930 7104
rect 21520 7080 22000 7110
rect 15610 7039 15930 7040
rect 5625 6762 5691 6765
rect 6545 6762 6611 6765
rect 19057 6762 19123 6765
rect 5625 6760 19123 6762
rect 5625 6704 5630 6760
rect 5686 6704 6550 6760
rect 6606 6704 19062 6760
rect 19118 6704 19123 6760
rect 5625 6702 19123 6704
rect 5625 6699 5691 6702
rect 6545 6699 6611 6702
rect 19057 6699 19123 6702
rect 4610 6560 4930 6561
rect 4610 6496 4618 6560
rect 4682 6496 4698 6560
rect 4762 6496 4778 6560
rect 4842 6496 4858 6560
rect 4922 6496 4930 6560
rect 4610 6495 4930 6496
rect 11944 6560 12264 6561
rect 11944 6496 11952 6560
rect 12016 6496 12032 6560
rect 12096 6496 12112 6560
rect 12176 6496 12192 6560
rect 12256 6496 12264 6560
rect 11944 6495 12264 6496
rect 19277 6560 19597 6561
rect 19277 6496 19285 6560
rect 19349 6496 19365 6560
rect 19429 6496 19445 6560
rect 19509 6496 19525 6560
rect 19589 6496 19597 6560
rect 19277 6495 19597 6496
rect 0 6352 480 6384
rect 0 6296 110 6352
rect 166 6296 480 6352
rect 0 6264 480 6296
rect 2497 6354 2563 6357
rect 2773 6354 2839 6357
rect 6177 6354 6243 6357
rect 2497 6352 6243 6354
rect 2497 6296 2502 6352
rect 2558 6296 2778 6352
rect 2834 6296 6182 6352
rect 6238 6296 6243 6352
rect 2497 6294 6243 6296
rect 2497 6291 2563 6294
rect 2773 6291 2839 6294
rect 6177 6291 6243 6294
rect 5073 6218 5139 6221
rect 8753 6218 8819 6221
rect 5073 6216 8819 6218
rect 5073 6160 5078 6216
rect 5134 6160 8758 6216
rect 8814 6160 8819 6216
rect 5073 6158 8819 6160
rect 5073 6155 5139 6158
rect 8753 6155 8819 6158
rect 9029 6218 9095 6221
rect 15009 6218 15075 6221
rect 9029 6216 15075 6218
rect 9029 6160 9034 6216
rect 9090 6160 15014 6216
rect 15070 6160 15075 6216
rect 9029 6158 15075 6160
rect 9029 6155 9095 6158
rect 15009 6155 15075 6158
rect 21520 6128 22000 6248
rect 8661 6082 8727 6085
rect 10133 6082 10199 6085
rect 12617 6082 12683 6085
rect 8661 6080 12683 6082
rect 8661 6024 8666 6080
rect 8722 6024 10138 6080
rect 10194 6024 12622 6080
rect 12678 6024 12683 6080
rect 8661 6022 12683 6024
rect 8661 6019 8727 6022
rect 10133 6019 10199 6022
rect 12617 6019 12683 6022
rect 8277 6016 8597 6017
rect 8277 5952 8285 6016
rect 8349 5952 8365 6016
rect 8429 5952 8445 6016
rect 8509 5952 8525 6016
rect 8589 5952 8597 6016
rect 8277 5951 8597 5952
rect 15610 6016 15930 6017
rect 15610 5952 15618 6016
rect 15682 5952 15698 6016
rect 15762 5952 15778 6016
rect 15842 5952 15858 6016
rect 15922 5952 15930 6016
rect 15610 5951 15930 5952
rect 3141 5810 3207 5813
rect 4102 5810 4108 5812
rect 3141 5808 4108 5810
rect 3141 5752 3146 5808
rect 3202 5752 4108 5808
rect 3141 5750 4108 5752
rect 3141 5747 3207 5750
rect 4102 5748 4108 5750
rect 4172 5748 4178 5812
rect 12801 5810 12867 5813
rect 21590 5810 21650 6128
rect 12801 5808 21650 5810
rect 12801 5752 12806 5808
rect 12862 5752 21650 5808
rect 12801 5750 21650 5752
rect 12801 5747 12867 5750
rect 4521 5674 4587 5677
rect 13169 5674 13235 5677
rect 4521 5672 13235 5674
rect 4521 5616 4526 5672
rect 4582 5616 13174 5672
rect 13230 5616 13235 5672
rect 4521 5614 13235 5616
rect 4521 5611 4587 5614
rect 13169 5611 13235 5614
rect 4610 5472 4930 5473
rect 4610 5408 4618 5472
rect 4682 5408 4698 5472
rect 4762 5408 4778 5472
rect 4842 5408 4858 5472
rect 4922 5408 4930 5472
rect 4610 5407 4930 5408
rect 11944 5472 12264 5473
rect 11944 5408 11952 5472
rect 12016 5408 12032 5472
rect 12096 5408 12112 5472
rect 12176 5408 12192 5472
rect 12256 5408 12264 5472
rect 11944 5407 12264 5408
rect 19277 5472 19597 5473
rect 19277 5408 19285 5472
rect 19349 5408 19365 5472
rect 19429 5408 19445 5472
rect 19509 5408 19525 5472
rect 19589 5408 19597 5472
rect 19277 5407 19597 5408
rect 3693 5266 3759 5269
rect 12341 5266 12407 5269
rect 21520 5268 22000 5296
rect 21520 5266 21588 5268
rect 3693 5264 12407 5266
rect 3693 5208 3698 5264
rect 3754 5208 12346 5264
rect 12402 5208 12407 5264
rect 3693 5206 12407 5208
rect 21460 5206 21588 5266
rect 3693 5203 3759 5206
rect 12341 5203 12407 5206
rect 21520 5204 21588 5206
rect 21652 5204 22000 5268
rect 21520 5176 22000 5204
rect 2313 5130 2379 5133
rect 4429 5130 4495 5133
rect 12525 5130 12591 5133
rect 2313 5128 4170 5130
rect 2313 5072 2318 5128
rect 2374 5072 4170 5128
rect 2313 5070 4170 5072
rect 2313 5067 2379 5070
rect 4110 4994 4170 5070
rect 4429 5128 12591 5130
rect 4429 5072 4434 5128
rect 4490 5072 12530 5128
rect 12586 5072 12591 5128
rect 4429 5070 12591 5072
rect 4429 5067 4495 5070
rect 12525 5067 12591 5070
rect 17166 5068 17172 5132
rect 17236 5130 17242 5132
rect 17309 5130 17375 5133
rect 17236 5128 17375 5130
rect 17236 5072 17314 5128
rect 17370 5072 17375 5128
rect 17236 5070 17375 5072
rect 17236 5068 17242 5070
rect 17309 5067 17375 5070
rect 8017 4994 8083 4997
rect 4110 4992 8083 4994
rect 4110 4936 8022 4992
rect 8078 4936 8083 4992
rect 4110 4934 8083 4936
rect 8017 4931 8083 4934
rect 8277 4928 8597 4929
rect 8277 4864 8285 4928
rect 8349 4864 8365 4928
rect 8429 4864 8445 4928
rect 8509 4864 8525 4928
rect 8589 4864 8597 4928
rect 8277 4863 8597 4864
rect 15610 4928 15930 4929
rect 15610 4864 15618 4928
rect 15682 4864 15698 4928
rect 15762 4864 15778 4928
rect 15842 4864 15858 4928
rect 15922 4864 15930 4928
rect 15610 4863 15930 4864
rect 7925 4722 7991 4725
rect 15469 4722 15535 4725
rect 7925 4720 15535 4722
rect 7925 4664 7930 4720
rect 7986 4664 15474 4720
rect 15530 4664 15535 4720
rect 7925 4662 15535 4664
rect 7925 4659 7991 4662
rect 15469 4659 15535 4662
rect 0 4496 480 4616
rect 6269 4586 6335 4589
rect 11789 4586 11855 4589
rect 6269 4584 11855 4586
rect 6269 4528 6274 4584
rect 6330 4528 11794 4584
rect 11850 4528 11855 4584
rect 6269 4526 11855 4528
rect 6269 4523 6335 4526
rect 11789 4523 11855 4526
rect 11973 4586 12039 4589
rect 11973 4584 21650 4586
rect 11973 4528 11978 4584
rect 12034 4528 21650 4584
rect 11973 4526 21650 4528
rect 11973 4523 12039 4526
rect 62 4178 122 4496
rect 2037 4450 2103 4453
rect 4102 4450 4108 4452
rect 2037 4448 4108 4450
rect 2037 4392 2042 4448
rect 2098 4392 4108 4448
rect 2037 4390 4108 4392
rect 2037 4387 2103 4390
rect 4102 4388 4108 4390
rect 4172 4388 4178 4452
rect 13813 4450 13879 4453
rect 15326 4450 15332 4452
rect 13813 4448 15332 4450
rect 13813 4392 13818 4448
rect 13874 4392 15332 4448
rect 13813 4390 15332 4392
rect 13813 4387 13879 4390
rect 15326 4388 15332 4390
rect 15396 4450 15402 4452
rect 15929 4450 15995 4453
rect 18505 4450 18571 4453
rect 15396 4448 18571 4450
rect 15396 4392 15934 4448
rect 15990 4392 18510 4448
rect 18566 4392 18571 4448
rect 15396 4390 18571 4392
rect 15396 4388 15402 4390
rect 15929 4387 15995 4390
rect 18505 4387 18571 4390
rect 4610 4384 4930 4385
rect 4610 4320 4618 4384
rect 4682 4320 4698 4384
rect 4762 4320 4778 4384
rect 4842 4320 4858 4384
rect 4922 4320 4930 4384
rect 4610 4319 4930 4320
rect 11944 4384 12264 4385
rect 11944 4320 11952 4384
rect 12016 4320 12032 4384
rect 12096 4320 12112 4384
rect 12176 4320 12192 4384
rect 12256 4320 12264 4384
rect 11944 4319 12264 4320
rect 19277 4384 19597 4385
rect 19277 4320 19285 4384
rect 19349 4320 19365 4384
rect 19429 4320 19445 4384
rect 19509 4320 19525 4384
rect 19589 4320 19597 4384
rect 21590 4344 21650 4526
rect 19277 4319 19597 4320
rect 21520 4224 22000 4344
rect 6821 4178 6887 4181
rect 62 4176 6887 4178
rect 62 4120 6826 4176
rect 6882 4120 6887 4176
rect 62 4118 6887 4120
rect 6821 4115 6887 4118
rect 9622 4116 9628 4180
rect 9692 4178 9698 4180
rect 19701 4178 19767 4181
rect 21398 4178 21404 4180
rect 9692 4176 21404 4178
rect 9692 4120 19706 4176
rect 19762 4120 21404 4176
rect 9692 4118 21404 4120
rect 9692 4116 9698 4118
rect 19701 4115 19767 4118
rect 21398 4116 21404 4118
rect 21468 4116 21474 4180
rect 3509 4042 3575 4045
rect 7189 4042 7255 4045
rect 9622 4042 9628 4044
rect 3509 4040 7255 4042
rect 3509 3984 3514 4040
rect 3570 3984 7194 4040
rect 7250 3984 7255 4040
rect 3509 3982 7255 3984
rect 3509 3979 3575 3982
rect 7189 3979 7255 3982
rect 7422 3982 9628 4042
rect 6126 3844 6132 3908
rect 6196 3906 6202 3908
rect 7281 3906 7347 3909
rect 6196 3904 7347 3906
rect 6196 3848 7286 3904
rect 7342 3848 7347 3904
rect 6196 3846 7347 3848
rect 6196 3844 6202 3846
rect 7281 3843 7347 3846
rect 2129 3770 2195 3773
rect 7422 3770 7482 3982
rect 9622 3980 9628 3982
rect 9692 3980 9698 4044
rect 13445 4042 13511 4045
rect 13445 4040 21650 4042
rect 13445 3984 13450 4040
rect 13506 3984 21650 4040
rect 13445 3982 21650 3984
rect 13445 3979 13511 3982
rect 8661 3906 8727 3909
rect 15377 3906 15443 3909
rect 8661 3904 15443 3906
rect 8661 3848 8666 3904
rect 8722 3848 15382 3904
rect 15438 3848 15443 3904
rect 8661 3846 15443 3848
rect 8661 3843 8727 3846
rect 15377 3843 15443 3846
rect 8277 3840 8597 3841
rect 8277 3776 8285 3840
rect 8349 3776 8365 3840
rect 8429 3776 8445 3840
rect 8509 3776 8525 3840
rect 8589 3776 8597 3840
rect 8277 3775 8597 3776
rect 15610 3840 15930 3841
rect 15610 3776 15618 3840
rect 15682 3776 15698 3840
rect 15762 3776 15778 3840
rect 15842 3776 15858 3840
rect 15922 3776 15930 3840
rect 15610 3775 15930 3776
rect 2129 3768 7482 3770
rect 2129 3712 2134 3768
rect 2190 3712 7482 3768
rect 2129 3710 7482 3712
rect 2129 3707 2195 3710
rect 3601 3634 3667 3637
rect 10593 3634 10659 3637
rect 3601 3632 10659 3634
rect 3601 3576 3606 3632
rect 3662 3576 10598 3632
rect 10654 3576 10659 3632
rect 3601 3574 10659 3576
rect 3601 3571 3667 3574
rect 10593 3571 10659 3574
rect 4337 3498 4403 3501
rect 12433 3498 12499 3501
rect 4337 3496 12499 3498
rect 4337 3440 4342 3496
rect 4398 3440 12438 3496
rect 12494 3440 12499 3496
rect 4337 3438 12499 3440
rect 4337 3435 4403 3438
rect 12433 3435 12499 3438
rect 21590 3392 21650 3982
rect 7189 3362 7255 3365
rect 10777 3362 10843 3365
rect 7189 3360 10843 3362
rect 7189 3304 7194 3360
rect 7250 3304 10782 3360
rect 10838 3304 10843 3360
rect 7189 3302 10843 3304
rect 7189 3299 7255 3302
rect 10777 3299 10843 3302
rect 4610 3296 4930 3297
rect 4610 3232 4618 3296
rect 4682 3232 4698 3296
rect 4762 3232 4778 3296
rect 4842 3232 4858 3296
rect 4922 3232 4930 3296
rect 4610 3231 4930 3232
rect 11944 3296 12264 3297
rect 11944 3232 11952 3296
rect 12016 3232 12032 3296
rect 12096 3232 12112 3296
rect 12176 3232 12192 3296
rect 12256 3232 12264 3296
rect 11944 3231 12264 3232
rect 19277 3296 19597 3297
rect 19277 3232 19285 3296
rect 19349 3232 19365 3296
rect 19429 3232 19445 3296
rect 19509 3232 19525 3296
rect 19589 3232 19597 3296
rect 21520 3272 22000 3392
rect 19277 3231 19597 3232
rect 17125 3226 17191 3229
rect 13770 3224 17191 3226
rect 13770 3168 17130 3224
rect 17186 3168 17191 3224
rect 13770 3166 17191 3168
rect 1945 3090 2011 3093
rect 4102 3090 4108 3092
rect 1945 3088 4108 3090
rect 1945 3032 1950 3088
rect 2006 3032 4108 3088
rect 1945 3030 4108 3032
rect 1945 3027 2011 3030
rect 4102 3028 4108 3030
rect 4172 3028 4178 3092
rect 5901 3090 5967 3093
rect 13770 3090 13830 3166
rect 17125 3163 17191 3166
rect 5901 3088 13830 3090
rect 5901 3032 5906 3088
rect 5962 3032 13830 3088
rect 5901 3030 13830 3032
rect 5901 3027 5967 3030
rect 14774 3028 14780 3092
rect 14844 3090 14850 3092
rect 14917 3090 14983 3093
rect 14844 3088 14983 3090
rect 14844 3032 14922 3088
rect 14978 3032 14983 3088
rect 14844 3030 14983 3032
rect 14844 3028 14850 3030
rect 14917 3027 14983 3030
rect 15101 3090 15167 3093
rect 15101 3088 21650 3090
rect 15101 3032 15106 3088
rect 15162 3032 21650 3088
rect 15101 3030 21650 3032
rect 15101 3027 15167 3030
rect 3325 2954 3391 2957
rect 62 2952 3391 2954
rect 62 2896 3330 2952
rect 3386 2896 3391 2952
rect 62 2894 3391 2896
rect 62 2712 122 2894
rect 3325 2891 3391 2894
rect 5533 2954 5599 2957
rect 10869 2954 10935 2957
rect 5533 2952 10935 2954
rect 5533 2896 5538 2952
rect 5594 2896 10874 2952
rect 10930 2896 10935 2952
rect 5533 2894 10935 2896
rect 5533 2891 5599 2894
rect 10869 2891 10935 2894
rect 8277 2752 8597 2753
rect 0 2592 480 2712
rect 8277 2688 8285 2752
rect 8349 2688 8365 2752
rect 8429 2688 8445 2752
rect 8509 2688 8525 2752
rect 8589 2688 8597 2752
rect 8277 2687 8597 2688
rect 15610 2752 15930 2753
rect 15610 2688 15618 2752
rect 15682 2688 15698 2752
rect 15762 2688 15778 2752
rect 15842 2688 15858 2752
rect 15922 2688 15930 2752
rect 15610 2687 15930 2688
rect 4429 2546 4495 2549
rect 18229 2546 18295 2549
rect 4429 2544 18295 2546
rect 4429 2488 4434 2544
rect 4490 2488 18234 2544
rect 18290 2488 18295 2544
rect 4429 2486 18295 2488
rect 4429 2483 4495 2486
rect 18229 2483 18295 2486
rect 21590 2440 21650 3030
rect 5901 2410 5967 2413
rect 18597 2410 18663 2413
rect 5901 2408 18663 2410
rect 5901 2352 5906 2408
rect 5962 2352 18602 2408
rect 18658 2352 18663 2408
rect 5901 2350 18663 2352
rect 5901 2347 5967 2350
rect 18597 2347 18663 2350
rect 21520 2320 22000 2440
rect 4610 2208 4930 2209
rect 4610 2144 4618 2208
rect 4682 2144 4698 2208
rect 4762 2144 4778 2208
rect 4842 2144 4858 2208
rect 4922 2144 4930 2208
rect 4610 2143 4930 2144
rect 11944 2208 12264 2209
rect 11944 2144 11952 2208
rect 12016 2144 12032 2208
rect 12096 2144 12112 2208
rect 12176 2144 12192 2208
rect 12256 2144 12264 2208
rect 11944 2143 12264 2144
rect 19277 2208 19597 2209
rect 19277 2144 19285 2208
rect 19349 2144 19365 2208
rect 19429 2144 19445 2208
rect 19509 2144 19525 2208
rect 19589 2144 19597 2208
rect 19277 2143 19597 2144
rect 11881 2002 11947 2005
rect 11881 2000 21650 2002
rect 11881 1944 11886 2000
rect 11942 1944 21650 2000
rect 11881 1942 21650 1944
rect 11881 1939 11947 1942
rect 4337 1866 4403 1869
rect 15193 1866 15259 1869
rect 4337 1864 15259 1866
rect 4337 1808 4342 1864
rect 4398 1808 15198 1864
rect 15254 1808 15259 1864
rect 4337 1806 15259 1808
rect 4337 1803 4403 1806
rect 15193 1803 15259 1806
rect 1393 1730 1459 1733
rect 18045 1730 18111 1733
rect 1393 1728 18111 1730
rect 1393 1672 1398 1728
rect 1454 1672 18050 1728
rect 18106 1672 18111 1728
rect 1393 1670 18111 1672
rect 1393 1667 1459 1670
rect 18045 1667 18111 1670
rect 21590 1488 21650 1942
rect 1761 1458 1827 1461
rect 62 1456 1827 1458
rect 62 1400 1766 1456
rect 1822 1400 1827 1456
rect 62 1398 1827 1400
rect 62 944 122 1398
rect 1761 1395 1827 1398
rect 21520 1368 22000 1488
rect 18689 1050 18755 1053
rect 18689 1048 21650 1050
rect 18689 992 18694 1048
rect 18750 992 21650 1048
rect 18689 990 21650 992
rect 18689 987 18755 990
rect 0 824 480 944
rect 21590 536 21650 990
rect 21520 416 22000 536
<< via3 >>
rect 4618 19612 4682 19616
rect 4618 19556 4622 19612
rect 4622 19556 4678 19612
rect 4678 19556 4682 19612
rect 4618 19552 4682 19556
rect 4698 19612 4762 19616
rect 4698 19556 4702 19612
rect 4702 19556 4758 19612
rect 4758 19556 4762 19612
rect 4698 19552 4762 19556
rect 4778 19612 4842 19616
rect 4778 19556 4782 19612
rect 4782 19556 4838 19612
rect 4838 19556 4842 19612
rect 4778 19552 4842 19556
rect 4858 19612 4922 19616
rect 4858 19556 4862 19612
rect 4862 19556 4918 19612
rect 4918 19556 4922 19612
rect 4858 19552 4922 19556
rect 11952 19612 12016 19616
rect 11952 19556 11956 19612
rect 11956 19556 12012 19612
rect 12012 19556 12016 19612
rect 11952 19552 12016 19556
rect 12032 19612 12096 19616
rect 12032 19556 12036 19612
rect 12036 19556 12092 19612
rect 12092 19556 12096 19612
rect 12032 19552 12096 19556
rect 12112 19612 12176 19616
rect 12112 19556 12116 19612
rect 12116 19556 12172 19612
rect 12172 19556 12176 19612
rect 12112 19552 12176 19556
rect 12192 19612 12256 19616
rect 12192 19556 12196 19612
rect 12196 19556 12252 19612
rect 12252 19556 12256 19612
rect 12192 19552 12256 19556
rect 19285 19612 19349 19616
rect 19285 19556 19289 19612
rect 19289 19556 19345 19612
rect 19345 19556 19349 19612
rect 19285 19552 19349 19556
rect 19365 19612 19429 19616
rect 19365 19556 19369 19612
rect 19369 19556 19425 19612
rect 19425 19556 19429 19612
rect 19365 19552 19429 19556
rect 19445 19612 19509 19616
rect 19445 19556 19449 19612
rect 19449 19556 19505 19612
rect 19505 19556 19509 19612
rect 19445 19552 19509 19556
rect 19525 19612 19589 19616
rect 19525 19556 19529 19612
rect 19529 19556 19585 19612
rect 19585 19556 19589 19612
rect 19525 19552 19589 19556
rect 8285 19068 8349 19072
rect 8285 19012 8289 19068
rect 8289 19012 8345 19068
rect 8345 19012 8349 19068
rect 8285 19008 8349 19012
rect 8365 19068 8429 19072
rect 8365 19012 8369 19068
rect 8369 19012 8425 19068
rect 8425 19012 8429 19068
rect 8365 19008 8429 19012
rect 8445 19068 8509 19072
rect 8445 19012 8449 19068
rect 8449 19012 8505 19068
rect 8505 19012 8509 19068
rect 8445 19008 8509 19012
rect 8525 19068 8589 19072
rect 8525 19012 8529 19068
rect 8529 19012 8585 19068
rect 8585 19012 8589 19068
rect 8525 19008 8589 19012
rect 15618 19068 15682 19072
rect 15618 19012 15622 19068
rect 15622 19012 15678 19068
rect 15678 19012 15682 19068
rect 15618 19008 15682 19012
rect 15698 19068 15762 19072
rect 15698 19012 15702 19068
rect 15702 19012 15758 19068
rect 15758 19012 15762 19068
rect 15698 19008 15762 19012
rect 15778 19068 15842 19072
rect 15778 19012 15782 19068
rect 15782 19012 15838 19068
rect 15838 19012 15842 19068
rect 15778 19008 15842 19012
rect 15858 19068 15922 19072
rect 15858 19012 15862 19068
rect 15862 19012 15918 19068
rect 15918 19012 15922 19068
rect 15858 19008 15922 19012
rect 4618 18524 4682 18528
rect 4618 18468 4622 18524
rect 4622 18468 4678 18524
rect 4678 18468 4682 18524
rect 4618 18464 4682 18468
rect 4698 18524 4762 18528
rect 4698 18468 4702 18524
rect 4702 18468 4758 18524
rect 4758 18468 4762 18524
rect 4698 18464 4762 18468
rect 4778 18524 4842 18528
rect 4778 18468 4782 18524
rect 4782 18468 4838 18524
rect 4838 18468 4842 18524
rect 4778 18464 4842 18468
rect 4858 18524 4922 18528
rect 4858 18468 4862 18524
rect 4862 18468 4918 18524
rect 4918 18468 4922 18524
rect 4858 18464 4922 18468
rect 11952 18524 12016 18528
rect 11952 18468 11956 18524
rect 11956 18468 12012 18524
rect 12012 18468 12016 18524
rect 11952 18464 12016 18468
rect 12032 18524 12096 18528
rect 12032 18468 12036 18524
rect 12036 18468 12092 18524
rect 12092 18468 12096 18524
rect 12032 18464 12096 18468
rect 12112 18524 12176 18528
rect 12112 18468 12116 18524
rect 12116 18468 12172 18524
rect 12172 18468 12176 18524
rect 12112 18464 12176 18468
rect 12192 18524 12256 18528
rect 12192 18468 12196 18524
rect 12196 18468 12252 18524
rect 12252 18468 12256 18524
rect 12192 18464 12256 18468
rect 19285 18524 19349 18528
rect 19285 18468 19289 18524
rect 19289 18468 19345 18524
rect 19345 18468 19349 18524
rect 19285 18464 19349 18468
rect 19365 18524 19429 18528
rect 19365 18468 19369 18524
rect 19369 18468 19425 18524
rect 19425 18468 19429 18524
rect 19365 18464 19429 18468
rect 19445 18524 19509 18528
rect 19445 18468 19449 18524
rect 19449 18468 19505 18524
rect 19505 18468 19509 18524
rect 19445 18464 19509 18468
rect 19525 18524 19589 18528
rect 19525 18468 19529 18524
rect 19529 18468 19585 18524
rect 19585 18468 19589 18524
rect 19525 18464 19589 18468
rect 8285 17980 8349 17984
rect 8285 17924 8289 17980
rect 8289 17924 8345 17980
rect 8345 17924 8349 17980
rect 8285 17920 8349 17924
rect 8365 17980 8429 17984
rect 8365 17924 8369 17980
rect 8369 17924 8425 17980
rect 8425 17924 8429 17980
rect 8365 17920 8429 17924
rect 8445 17980 8509 17984
rect 8445 17924 8449 17980
rect 8449 17924 8505 17980
rect 8505 17924 8509 17980
rect 8445 17920 8509 17924
rect 8525 17980 8589 17984
rect 8525 17924 8529 17980
rect 8529 17924 8585 17980
rect 8585 17924 8589 17980
rect 8525 17920 8589 17924
rect 15618 17980 15682 17984
rect 15618 17924 15622 17980
rect 15622 17924 15678 17980
rect 15678 17924 15682 17980
rect 15618 17920 15682 17924
rect 15698 17980 15762 17984
rect 15698 17924 15702 17980
rect 15702 17924 15758 17980
rect 15758 17924 15762 17980
rect 15698 17920 15762 17924
rect 15778 17980 15842 17984
rect 15778 17924 15782 17980
rect 15782 17924 15838 17980
rect 15838 17924 15842 17980
rect 15778 17920 15842 17924
rect 15858 17980 15922 17984
rect 15858 17924 15862 17980
rect 15862 17924 15918 17980
rect 15918 17924 15922 17980
rect 15858 17920 15922 17924
rect 4618 17436 4682 17440
rect 4618 17380 4622 17436
rect 4622 17380 4678 17436
rect 4678 17380 4682 17436
rect 4618 17376 4682 17380
rect 4698 17436 4762 17440
rect 4698 17380 4702 17436
rect 4702 17380 4758 17436
rect 4758 17380 4762 17436
rect 4698 17376 4762 17380
rect 4778 17436 4842 17440
rect 4778 17380 4782 17436
rect 4782 17380 4838 17436
rect 4838 17380 4842 17436
rect 4778 17376 4842 17380
rect 4858 17436 4922 17440
rect 4858 17380 4862 17436
rect 4862 17380 4918 17436
rect 4918 17380 4922 17436
rect 4858 17376 4922 17380
rect 11952 17436 12016 17440
rect 11952 17380 11956 17436
rect 11956 17380 12012 17436
rect 12012 17380 12016 17436
rect 11952 17376 12016 17380
rect 12032 17436 12096 17440
rect 12032 17380 12036 17436
rect 12036 17380 12092 17436
rect 12092 17380 12096 17436
rect 12032 17376 12096 17380
rect 12112 17436 12176 17440
rect 12112 17380 12116 17436
rect 12116 17380 12172 17436
rect 12172 17380 12176 17436
rect 12112 17376 12176 17380
rect 12192 17436 12256 17440
rect 12192 17380 12196 17436
rect 12196 17380 12252 17436
rect 12252 17380 12256 17436
rect 12192 17376 12256 17380
rect 19285 17436 19349 17440
rect 19285 17380 19289 17436
rect 19289 17380 19345 17436
rect 19345 17380 19349 17436
rect 19285 17376 19349 17380
rect 19365 17436 19429 17440
rect 19365 17380 19369 17436
rect 19369 17380 19425 17436
rect 19425 17380 19429 17436
rect 19365 17376 19429 17380
rect 19445 17436 19509 17440
rect 19445 17380 19449 17436
rect 19449 17380 19505 17436
rect 19505 17380 19509 17436
rect 19445 17376 19509 17380
rect 19525 17436 19589 17440
rect 19525 17380 19529 17436
rect 19529 17380 19585 17436
rect 19585 17380 19589 17436
rect 19525 17376 19589 17380
rect 8285 16892 8349 16896
rect 8285 16836 8289 16892
rect 8289 16836 8345 16892
rect 8345 16836 8349 16892
rect 8285 16832 8349 16836
rect 8365 16892 8429 16896
rect 8365 16836 8369 16892
rect 8369 16836 8425 16892
rect 8425 16836 8429 16892
rect 8365 16832 8429 16836
rect 8445 16892 8509 16896
rect 8445 16836 8449 16892
rect 8449 16836 8505 16892
rect 8505 16836 8509 16892
rect 8445 16832 8509 16836
rect 8525 16892 8589 16896
rect 8525 16836 8529 16892
rect 8529 16836 8585 16892
rect 8585 16836 8589 16892
rect 8525 16832 8589 16836
rect 15618 16892 15682 16896
rect 15618 16836 15622 16892
rect 15622 16836 15678 16892
rect 15678 16836 15682 16892
rect 15618 16832 15682 16836
rect 15698 16892 15762 16896
rect 15698 16836 15702 16892
rect 15702 16836 15758 16892
rect 15758 16836 15762 16892
rect 15698 16832 15762 16836
rect 15778 16892 15842 16896
rect 15778 16836 15782 16892
rect 15782 16836 15838 16892
rect 15838 16836 15842 16892
rect 15778 16832 15842 16836
rect 15858 16892 15922 16896
rect 15858 16836 15862 16892
rect 15862 16836 15918 16892
rect 15918 16836 15922 16892
rect 15858 16832 15922 16836
rect 4618 16348 4682 16352
rect 4618 16292 4622 16348
rect 4622 16292 4678 16348
rect 4678 16292 4682 16348
rect 4618 16288 4682 16292
rect 4698 16348 4762 16352
rect 4698 16292 4702 16348
rect 4702 16292 4758 16348
rect 4758 16292 4762 16348
rect 4698 16288 4762 16292
rect 4778 16348 4842 16352
rect 4778 16292 4782 16348
rect 4782 16292 4838 16348
rect 4838 16292 4842 16348
rect 4778 16288 4842 16292
rect 4858 16348 4922 16352
rect 4858 16292 4862 16348
rect 4862 16292 4918 16348
rect 4918 16292 4922 16348
rect 4858 16288 4922 16292
rect 11952 16348 12016 16352
rect 11952 16292 11956 16348
rect 11956 16292 12012 16348
rect 12012 16292 12016 16348
rect 11952 16288 12016 16292
rect 12032 16348 12096 16352
rect 12032 16292 12036 16348
rect 12036 16292 12092 16348
rect 12092 16292 12096 16348
rect 12032 16288 12096 16292
rect 12112 16348 12176 16352
rect 12112 16292 12116 16348
rect 12116 16292 12172 16348
rect 12172 16292 12176 16348
rect 12112 16288 12176 16292
rect 12192 16348 12256 16352
rect 12192 16292 12196 16348
rect 12196 16292 12252 16348
rect 12252 16292 12256 16348
rect 12192 16288 12256 16292
rect 19285 16348 19349 16352
rect 19285 16292 19289 16348
rect 19289 16292 19345 16348
rect 19345 16292 19349 16348
rect 19285 16288 19349 16292
rect 19365 16348 19429 16352
rect 19365 16292 19369 16348
rect 19369 16292 19425 16348
rect 19425 16292 19429 16348
rect 19365 16288 19429 16292
rect 19445 16348 19509 16352
rect 19445 16292 19449 16348
rect 19449 16292 19505 16348
rect 19505 16292 19509 16348
rect 19445 16288 19509 16292
rect 19525 16348 19589 16352
rect 19525 16292 19529 16348
rect 19529 16292 19585 16348
rect 19585 16292 19589 16348
rect 19525 16288 19589 16292
rect 8285 15804 8349 15808
rect 8285 15748 8289 15804
rect 8289 15748 8345 15804
rect 8345 15748 8349 15804
rect 8285 15744 8349 15748
rect 8365 15804 8429 15808
rect 8365 15748 8369 15804
rect 8369 15748 8425 15804
rect 8425 15748 8429 15804
rect 8365 15744 8429 15748
rect 8445 15804 8509 15808
rect 8445 15748 8449 15804
rect 8449 15748 8505 15804
rect 8505 15748 8509 15804
rect 8445 15744 8509 15748
rect 8525 15804 8589 15808
rect 8525 15748 8529 15804
rect 8529 15748 8585 15804
rect 8585 15748 8589 15804
rect 8525 15744 8589 15748
rect 15618 15804 15682 15808
rect 15618 15748 15622 15804
rect 15622 15748 15678 15804
rect 15678 15748 15682 15804
rect 15618 15744 15682 15748
rect 15698 15804 15762 15808
rect 15698 15748 15702 15804
rect 15702 15748 15758 15804
rect 15758 15748 15762 15804
rect 15698 15744 15762 15748
rect 15778 15804 15842 15808
rect 15778 15748 15782 15804
rect 15782 15748 15838 15804
rect 15838 15748 15842 15804
rect 15778 15744 15842 15748
rect 15858 15804 15922 15808
rect 15858 15748 15862 15804
rect 15862 15748 15918 15804
rect 15918 15748 15922 15804
rect 15858 15744 15922 15748
rect 4618 15260 4682 15264
rect 4618 15204 4622 15260
rect 4622 15204 4678 15260
rect 4678 15204 4682 15260
rect 4618 15200 4682 15204
rect 4698 15260 4762 15264
rect 4698 15204 4702 15260
rect 4702 15204 4758 15260
rect 4758 15204 4762 15260
rect 4698 15200 4762 15204
rect 4778 15260 4842 15264
rect 4778 15204 4782 15260
rect 4782 15204 4838 15260
rect 4838 15204 4842 15260
rect 4778 15200 4842 15204
rect 4858 15260 4922 15264
rect 4858 15204 4862 15260
rect 4862 15204 4918 15260
rect 4918 15204 4922 15260
rect 4858 15200 4922 15204
rect 11952 15260 12016 15264
rect 11952 15204 11956 15260
rect 11956 15204 12012 15260
rect 12012 15204 12016 15260
rect 11952 15200 12016 15204
rect 12032 15260 12096 15264
rect 12032 15204 12036 15260
rect 12036 15204 12092 15260
rect 12092 15204 12096 15260
rect 12032 15200 12096 15204
rect 12112 15260 12176 15264
rect 12112 15204 12116 15260
rect 12116 15204 12172 15260
rect 12172 15204 12176 15260
rect 12112 15200 12176 15204
rect 12192 15260 12256 15264
rect 12192 15204 12196 15260
rect 12196 15204 12252 15260
rect 12252 15204 12256 15260
rect 12192 15200 12256 15204
rect 19285 15260 19349 15264
rect 19285 15204 19289 15260
rect 19289 15204 19345 15260
rect 19345 15204 19349 15260
rect 19285 15200 19349 15204
rect 19365 15260 19429 15264
rect 19365 15204 19369 15260
rect 19369 15204 19425 15260
rect 19425 15204 19429 15260
rect 19365 15200 19429 15204
rect 19445 15260 19509 15264
rect 19445 15204 19449 15260
rect 19449 15204 19505 15260
rect 19505 15204 19509 15260
rect 19445 15200 19509 15204
rect 19525 15260 19589 15264
rect 19525 15204 19529 15260
rect 19529 15204 19585 15260
rect 19585 15204 19589 15260
rect 19525 15200 19589 15204
rect 21588 14724 21652 14788
rect 8285 14716 8349 14720
rect 8285 14660 8289 14716
rect 8289 14660 8345 14716
rect 8345 14660 8349 14716
rect 8285 14656 8349 14660
rect 8365 14716 8429 14720
rect 8365 14660 8369 14716
rect 8369 14660 8425 14716
rect 8425 14660 8429 14716
rect 8365 14656 8429 14660
rect 8445 14716 8509 14720
rect 8445 14660 8449 14716
rect 8449 14660 8505 14716
rect 8505 14660 8509 14716
rect 8445 14656 8509 14660
rect 8525 14716 8589 14720
rect 8525 14660 8529 14716
rect 8529 14660 8585 14716
rect 8585 14660 8589 14716
rect 8525 14656 8589 14660
rect 15618 14716 15682 14720
rect 15618 14660 15622 14716
rect 15622 14660 15678 14716
rect 15678 14660 15682 14716
rect 15618 14656 15682 14660
rect 15698 14716 15762 14720
rect 15698 14660 15702 14716
rect 15702 14660 15758 14716
rect 15758 14660 15762 14716
rect 15698 14656 15762 14660
rect 15778 14716 15842 14720
rect 15778 14660 15782 14716
rect 15782 14660 15838 14716
rect 15838 14660 15842 14716
rect 15778 14656 15842 14660
rect 15858 14716 15922 14720
rect 15858 14660 15862 14716
rect 15862 14660 15918 14716
rect 15918 14660 15922 14716
rect 15858 14656 15922 14660
rect 21404 14588 21468 14652
rect 4618 14172 4682 14176
rect 4618 14116 4622 14172
rect 4622 14116 4678 14172
rect 4678 14116 4682 14172
rect 4618 14112 4682 14116
rect 4698 14172 4762 14176
rect 4698 14116 4702 14172
rect 4702 14116 4758 14172
rect 4758 14116 4762 14172
rect 4698 14112 4762 14116
rect 4778 14172 4842 14176
rect 4778 14116 4782 14172
rect 4782 14116 4838 14172
rect 4838 14116 4842 14172
rect 4778 14112 4842 14116
rect 4858 14172 4922 14176
rect 4858 14116 4862 14172
rect 4862 14116 4918 14172
rect 4918 14116 4922 14172
rect 4858 14112 4922 14116
rect 11952 14172 12016 14176
rect 11952 14116 11956 14172
rect 11956 14116 12012 14172
rect 12012 14116 12016 14172
rect 11952 14112 12016 14116
rect 12032 14172 12096 14176
rect 12032 14116 12036 14172
rect 12036 14116 12092 14172
rect 12092 14116 12096 14172
rect 12032 14112 12096 14116
rect 12112 14172 12176 14176
rect 12112 14116 12116 14172
rect 12116 14116 12172 14172
rect 12172 14116 12176 14172
rect 12112 14112 12176 14116
rect 12192 14172 12256 14176
rect 12192 14116 12196 14172
rect 12196 14116 12252 14172
rect 12252 14116 12256 14172
rect 12192 14112 12256 14116
rect 19285 14172 19349 14176
rect 19285 14116 19289 14172
rect 19289 14116 19345 14172
rect 19345 14116 19349 14172
rect 19285 14112 19349 14116
rect 19365 14172 19429 14176
rect 19365 14116 19369 14172
rect 19369 14116 19425 14172
rect 19425 14116 19429 14172
rect 19365 14112 19429 14116
rect 19445 14172 19509 14176
rect 19445 14116 19449 14172
rect 19449 14116 19505 14172
rect 19505 14116 19509 14172
rect 19445 14112 19509 14116
rect 19525 14172 19589 14176
rect 19525 14116 19529 14172
rect 19529 14116 19585 14172
rect 19585 14116 19589 14172
rect 19525 14112 19589 14116
rect 60 13636 124 13700
rect 8285 13628 8349 13632
rect 8285 13572 8289 13628
rect 8289 13572 8345 13628
rect 8345 13572 8349 13628
rect 8285 13568 8349 13572
rect 8365 13628 8429 13632
rect 8365 13572 8369 13628
rect 8369 13572 8425 13628
rect 8425 13572 8429 13628
rect 8365 13568 8429 13572
rect 8445 13628 8509 13632
rect 8445 13572 8449 13628
rect 8449 13572 8505 13628
rect 8505 13572 8509 13628
rect 8445 13568 8509 13572
rect 8525 13628 8589 13632
rect 8525 13572 8529 13628
rect 8529 13572 8585 13628
rect 8585 13572 8589 13628
rect 8525 13568 8589 13572
rect 15618 13628 15682 13632
rect 15618 13572 15622 13628
rect 15622 13572 15678 13628
rect 15678 13572 15682 13628
rect 15618 13568 15682 13572
rect 15698 13628 15762 13632
rect 15698 13572 15702 13628
rect 15702 13572 15758 13628
rect 15758 13572 15762 13628
rect 15698 13568 15762 13572
rect 15778 13628 15842 13632
rect 15778 13572 15782 13628
rect 15782 13572 15838 13628
rect 15838 13572 15842 13628
rect 15778 13568 15842 13572
rect 15858 13628 15922 13632
rect 15858 13572 15862 13628
rect 15862 13572 15918 13628
rect 15918 13572 15922 13628
rect 15858 13568 15922 13572
rect 60 13364 124 13428
rect 4618 13084 4682 13088
rect 4618 13028 4622 13084
rect 4622 13028 4678 13084
rect 4678 13028 4682 13084
rect 4618 13024 4682 13028
rect 4698 13084 4762 13088
rect 4698 13028 4702 13084
rect 4702 13028 4758 13084
rect 4758 13028 4762 13084
rect 4698 13024 4762 13028
rect 4778 13084 4842 13088
rect 4778 13028 4782 13084
rect 4782 13028 4838 13084
rect 4838 13028 4842 13084
rect 4778 13024 4842 13028
rect 4858 13084 4922 13088
rect 4858 13028 4862 13084
rect 4862 13028 4918 13084
rect 4918 13028 4922 13084
rect 4858 13024 4922 13028
rect 11952 13084 12016 13088
rect 11952 13028 11956 13084
rect 11956 13028 12012 13084
rect 12012 13028 12016 13084
rect 11952 13024 12016 13028
rect 12032 13084 12096 13088
rect 12032 13028 12036 13084
rect 12036 13028 12092 13084
rect 12092 13028 12096 13084
rect 12032 13024 12096 13028
rect 12112 13084 12176 13088
rect 12112 13028 12116 13084
rect 12116 13028 12172 13084
rect 12172 13028 12176 13084
rect 12112 13024 12176 13028
rect 12192 13084 12256 13088
rect 12192 13028 12196 13084
rect 12196 13028 12252 13084
rect 12252 13028 12256 13084
rect 12192 13024 12256 13028
rect 19285 13084 19349 13088
rect 19285 13028 19289 13084
rect 19289 13028 19345 13084
rect 19345 13028 19349 13084
rect 19285 13024 19349 13028
rect 19365 13084 19429 13088
rect 19365 13028 19369 13084
rect 19369 13028 19425 13084
rect 19425 13028 19429 13084
rect 19365 13024 19429 13028
rect 19445 13084 19509 13088
rect 19445 13028 19449 13084
rect 19449 13028 19505 13084
rect 19505 13028 19509 13084
rect 19445 13024 19509 13028
rect 19525 13084 19589 13088
rect 19525 13028 19529 13084
rect 19529 13028 19585 13084
rect 19585 13028 19589 13084
rect 19525 13024 19589 13028
rect 6132 12820 6196 12884
rect 8285 12540 8349 12544
rect 8285 12484 8289 12540
rect 8289 12484 8345 12540
rect 8345 12484 8349 12540
rect 8285 12480 8349 12484
rect 8365 12540 8429 12544
rect 8365 12484 8369 12540
rect 8369 12484 8425 12540
rect 8425 12484 8429 12540
rect 8365 12480 8429 12484
rect 8445 12540 8509 12544
rect 8445 12484 8449 12540
rect 8449 12484 8505 12540
rect 8505 12484 8509 12540
rect 8445 12480 8509 12484
rect 8525 12540 8589 12544
rect 8525 12484 8529 12540
rect 8529 12484 8585 12540
rect 8585 12484 8589 12540
rect 8525 12480 8589 12484
rect 15618 12540 15682 12544
rect 15618 12484 15622 12540
rect 15622 12484 15678 12540
rect 15678 12484 15682 12540
rect 15618 12480 15682 12484
rect 15698 12540 15762 12544
rect 15698 12484 15702 12540
rect 15702 12484 15758 12540
rect 15758 12484 15762 12540
rect 15698 12480 15762 12484
rect 15778 12540 15842 12544
rect 15778 12484 15782 12540
rect 15782 12484 15838 12540
rect 15838 12484 15842 12540
rect 15778 12480 15842 12484
rect 15858 12540 15922 12544
rect 15858 12484 15862 12540
rect 15862 12484 15918 12540
rect 15918 12484 15922 12540
rect 15858 12480 15922 12484
rect 4618 11996 4682 12000
rect 4618 11940 4622 11996
rect 4622 11940 4678 11996
rect 4678 11940 4682 11996
rect 4618 11936 4682 11940
rect 4698 11996 4762 12000
rect 4698 11940 4702 11996
rect 4702 11940 4758 11996
rect 4758 11940 4762 11996
rect 4698 11936 4762 11940
rect 4778 11996 4842 12000
rect 4778 11940 4782 11996
rect 4782 11940 4838 11996
rect 4838 11940 4842 11996
rect 4778 11936 4842 11940
rect 4858 11996 4922 12000
rect 4858 11940 4862 11996
rect 4862 11940 4918 11996
rect 4918 11940 4922 11996
rect 4858 11936 4922 11940
rect 11952 11996 12016 12000
rect 11952 11940 11956 11996
rect 11956 11940 12012 11996
rect 12012 11940 12016 11996
rect 11952 11936 12016 11940
rect 12032 11996 12096 12000
rect 12032 11940 12036 11996
rect 12036 11940 12092 11996
rect 12092 11940 12096 11996
rect 12032 11936 12096 11940
rect 12112 11996 12176 12000
rect 12112 11940 12116 11996
rect 12116 11940 12172 11996
rect 12172 11940 12176 11996
rect 12112 11936 12176 11940
rect 12192 11996 12256 12000
rect 12192 11940 12196 11996
rect 12196 11940 12252 11996
rect 12252 11940 12256 11996
rect 12192 11936 12256 11940
rect 19285 11996 19349 12000
rect 19285 11940 19289 11996
rect 19289 11940 19345 11996
rect 19345 11940 19349 11996
rect 19285 11936 19349 11940
rect 19365 11996 19429 12000
rect 19365 11940 19369 11996
rect 19369 11940 19425 11996
rect 19425 11940 19429 11996
rect 19365 11936 19429 11940
rect 19445 11996 19509 12000
rect 19445 11940 19449 11996
rect 19449 11940 19505 11996
rect 19505 11940 19509 11996
rect 19445 11936 19509 11940
rect 19525 11996 19589 12000
rect 19525 11940 19529 11996
rect 19529 11940 19585 11996
rect 19585 11940 19589 11996
rect 19525 11936 19589 11940
rect 8285 11452 8349 11456
rect 8285 11396 8289 11452
rect 8289 11396 8345 11452
rect 8345 11396 8349 11452
rect 8285 11392 8349 11396
rect 8365 11452 8429 11456
rect 8365 11396 8369 11452
rect 8369 11396 8425 11452
rect 8425 11396 8429 11452
rect 8365 11392 8429 11396
rect 8445 11452 8509 11456
rect 8445 11396 8449 11452
rect 8449 11396 8505 11452
rect 8505 11396 8509 11452
rect 8445 11392 8509 11396
rect 8525 11452 8589 11456
rect 8525 11396 8529 11452
rect 8529 11396 8585 11452
rect 8585 11396 8589 11452
rect 8525 11392 8589 11396
rect 15618 11452 15682 11456
rect 15618 11396 15622 11452
rect 15622 11396 15678 11452
rect 15678 11396 15682 11452
rect 15618 11392 15682 11396
rect 15698 11452 15762 11456
rect 15698 11396 15702 11452
rect 15702 11396 15758 11452
rect 15758 11396 15762 11452
rect 15698 11392 15762 11396
rect 15778 11452 15842 11456
rect 15778 11396 15782 11452
rect 15782 11396 15838 11452
rect 15838 11396 15842 11452
rect 15778 11392 15842 11396
rect 15858 11452 15922 11456
rect 15858 11396 15862 11452
rect 15862 11396 15918 11452
rect 15918 11396 15922 11452
rect 15858 11392 15922 11396
rect 4618 10908 4682 10912
rect 4618 10852 4622 10908
rect 4622 10852 4678 10908
rect 4678 10852 4682 10908
rect 4618 10848 4682 10852
rect 4698 10908 4762 10912
rect 4698 10852 4702 10908
rect 4702 10852 4758 10908
rect 4758 10852 4762 10908
rect 4698 10848 4762 10852
rect 4778 10908 4842 10912
rect 4778 10852 4782 10908
rect 4782 10852 4838 10908
rect 4838 10852 4842 10908
rect 4778 10848 4842 10852
rect 4858 10908 4922 10912
rect 4858 10852 4862 10908
rect 4862 10852 4918 10908
rect 4918 10852 4922 10908
rect 4858 10848 4922 10852
rect 11952 10908 12016 10912
rect 11952 10852 11956 10908
rect 11956 10852 12012 10908
rect 12012 10852 12016 10908
rect 11952 10848 12016 10852
rect 12032 10908 12096 10912
rect 12032 10852 12036 10908
rect 12036 10852 12092 10908
rect 12092 10852 12096 10908
rect 12032 10848 12096 10852
rect 12112 10908 12176 10912
rect 12112 10852 12116 10908
rect 12116 10852 12172 10908
rect 12172 10852 12176 10908
rect 12112 10848 12176 10852
rect 12192 10908 12256 10912
rect 12192 10852 12196 10908
rect 12196 10852 12252 10908
rect 12252 10852 12256 10908
rect 12192 10848 12256 10852
rect 19285 10908 19349 10912
rect 19285 10852 19289 10908
rect 19289 10852 19345 10908
rect 19345 10852 19349 10908
rect 19285 10848 19349 10852
rect 19365 10908 19429 10912
rect 19365 10852 19369 10908
rect 19369 10852 19425 10908
rect 19425 10852 19429 10908
rect 19365 10848 19429 10852
rect 19445 10908 19509 10912
rect 19445 10852 19449 10908
rect 19449 10852 19505 10908
rect 19505 10852 19509 10908
rect 19445 10848 19509 10852
rect 19525 10908 19589 10912
rect 19525 10852 19529 10908
rect 19529 10852 19585 10908
rect 19585 10852 19589 10908
rect 19525 10848 19589 10852
rect 8285 10364 8349 10368
rect 8285 10308 8289 10364
rect 8289 10308 8345 10364
rect 8345 10308 8349 10364
rect 8285 10304 8349 10308
rect 8365 10364 8429 10368
rect 8365 10308 8369 10364
rect 8369 10308 8425 10364
rect 8425 10308 8429 10364
rect 8365 10304 8429 10308
rect 8445 10364 8509 10368
rect 8445 10308 8449 10364
rect 8449 10308 8505 10364
rect 8505 10308 8509 10364
rect 8445 10304 8509 10308
rect 8525 10364 8589 10368
rect 8525 10308 8529 10364
rect 8529 10308 8585 10364
rect 8585 10308 8589 10364
rect 8525 10304 8589 10308
rect 15618 10364 15682 10368
rect 15618 10308 15622 10364
rect 15622 10308 15678 10364
rect 15678 10308 15682 10364
rect 15618 10304 15682 10308
rect 15698 10364 15762 10368
rect 15698 10308 15702 10364
rect 15702 10308 15758 10364
rect 15758 10308 15762 10364
rect 15698 10304 15762 10308
rect 15778 10364 15842 10368
rect 15778 10308 15782 10364
rect 15782 10308 15838 10364
rect 15838 10308 15842 10364
rect 15778 10304 15842 10308
rect 15858 10364 15922 10368
rect 15858 10308 15862 10364
rect 15862 10308 15918 10364
rect 15918 10308 15922 10364
rect 15858 10304 15922 10308
rect 4618 9820 4682 9824
rect 4618 9764 4622 9820
rect 4622 9764 4678 9820
rect 4678 9764 4682 9820
rect 4618 9760 4682 9764
rect 4698 9820 4762 9824
rect 4698 9764 4702 9820
rect 4702 9764 4758 9820
rect 4758 9764 4762 9820
rect 4698 9760 4762 9764
rect 4778 9820 4842 9824
rect 4778 9764 4782 9820
rect 4782 9764 4838 9820
rect 4838 9764 4842 9820
rect 4778 9760 4842 9764
rect 4858 9820 4922 9824
rect 4858 9764 4862 9820
rect 4862 9764 4918 9820
rect 4918 9764 4922 9820
rect 4858 9760 4922 9764
rect 11952 9820 12016 9824
rect 11952 9764 11956 9820
rect 11956 9764 12012 9820
rect 12012 9764 12016 9820
rect 11952 9760 12016 9764
rect 12032 9820 12096 9824
rect 12032 9764 12036 9820
rect 12036 9764 12092 9820
rect 12092 9764 12096 9820
rect 12032 9760 12096 9764
rect 12112 9820 12176 9824
rect 12112 9764 12116 9820
rect 12116 9764 12172 9820
rect 12172 9764 12176 9820
rect 12112 9760 12176 9764
rect 12192 9820 12256 9824
rect 12192 9764 12196 9820
rect 12196 9764 12252 9820
rect 12252 9764 12256 9820
rect 12192 9760 12256 9764
rect 19285 9820 19349 9824
rect 19285 9764 19289 9820
rect 19289 9764 19345 9820
rect 19345 9764 19349 9820
rect 19285 9760 19349 9764
rect 19365 9820 19429 9824
rect 19365 9764 19369 9820
rect 19369 9764 19425 9820
rect 19425 9764 19429 9820
rect 19365 9760 19429 9764
rect 19445 9820 19509 9824
rect 19445 9764 19449 9820
rect 19449 9764 19505 9820
rect 19505 9764 19509 9820
rect 19445 9760 19509 9764
rect 19525 9820 19589 9824
rect 19525 9764 19529 9820
rect 19529 9764 19585 9820
rect 19585 9764 19589 9820
rect 19525 9760 19589 9764
rect 8285 9276 8349 9280
rect 8285 9220 8289 9276
rect 8289 9220 8345 9276
rect 8345 9220 8349 9276
rect 8285 9216 8349 9220
rect 8365 9276 8429 9280
rect 8365 9220 8369 9276
rect 8369 9220 8425 9276
rect 8425 9220 8429 9276
rect 8365 9216 8429 9220
rect 8445 9276 8509 9280
rect 8445 9220 8449 9276
rect 8449 9220 8505 9276
rect 8505 9220 8509 9276
rect 8445 9216 8509 9220
rect 8525 9276 8589 9280
rect 8525 9220 8529 9276
rect 8529 9220 8585 9276
rect 8585 9220 8589 9276
rect 8525 9216 8589 9220
rect 15618 9276 15682 9280
rect 15618 9220 15622 9276
rect 15622 9220 15678 9276
rect 15678 9220 15682 9276
rect 15618 9216 15682 9220
rect 15698 9276 15762 9280
rect 15698 9220 15702 9276
rect 15702 9220 15758 9276
rect 15758 9220 15762 9276
rect 15698 9216 15762 9220
rect 15778 9276 15842 9280
rect 15778 9220 15782 9276
rect 15782 9220 15838 9276
rect 15838 9220 15842 9276
rect 15778 9216 15842 9220
rect 15858 9276 15922 9280
rect 15858 9220 15862 9276
rect 15862 9220 15918 9276
rect 15918 9220 15922 9276
rect 15858 9216 15922 9220
rect 21588 9012 21652 9076
rect 21588 8842 21652 8906
rect 4618 8732 4682 8736
rect 4618 8676 4622 8732
rect 4622 8676 4678 8732
rect 4678 8676 4682 8732
rect 4618 8672 4682 8676
rect 4698 8732 4762 8736
rect 4698 8676 4702 8732
rect 4702 8676 4758 8732
rect 4758 8676 4762 8732
rect 4698 8672 4762 8676
rect 4778 8732 4842 8736
rect 4778 8676 4782 8732
rect 4782 8676 4838 8732
rect 4838 8676 4842 8732
rect 4778 8672 4842 8676
rect 4858 8732 4922 8736
rect 4858 8676 4862 8732
rect 4862 8676 4918 8732
rect 4918 8676 4922 8732
rect 4858 8672 4922 8676
rect 11952 8732 12016 8736
rect 11952 8676 11956 8732
rect 11956 8676 12012 8732
rect 12012 8676 12016 8732
rect 11952 8672 12016 8676
rect 12032 8732 12096 8736
rect 12032 8676 12036 8732
rect 12036 8676 12092 8732
rect 12092 8676 12096 8732
rect 12032 8672 12096 8676
rect 12112 8732 12176 8736
rect 12112 8676 12116 8732
rect 12116 8676 12172 8732
rect 12172 8676 12176 8732
rect 12112 8672 12176 8676
rect 12192 8732 12256 8736
rect 12192 8676 12196 8732
rect 12196 8676 12252 8732
rect 12252 8676 12256 8732
rect 12192 8672 12256 8676
rect 19285 8732 19349 8736
rect 19285 8676 19289 8732
rect 19289 8676 19345 8732
rect 19345 8676 19349 8732
rect 19285 8672 19349 8676
rect 19365 8732 19429 8736
rect 19365 8676 19369 8732
rect 19369 8676 19425 8732
rect 19425 8676 19429 8732
rect 19365 8672 19429 8676
rect 19445 8732 19509 8736
rect 19445 8676 19449 8732
rect 19449 8676 19505 8732
rect 19505 8676 19509 8732
rect 19445 8672 19509 8676
rect 19525 8732 19589 8736
rect 19525 8676 19529 8732
rect 19529 8676 19585 8732
rect 19585 8676 19589 8732
rect 19525 8672 19589 8676
rect 8285 8188 8349 8192
rect 8285 8132 8289 8188
rect 8289 8132 8345 8188
rect 8345 8132 8349 8188
rect 8285 8128 8349 8132
rect 8365 8188 8429 8192
rect 8365 8132 8369 8188
rect 8369 8132 8425 8188
rect 8425 8132 8429 8188
rect 8365 8128 8429 8132
rect 8445 8188 8509 8192
rect 8445 8132 8449 8188
rect 8449 8132 8505 8188
rect 8505 8132 8509 8188
rect 8445 8128 8509 8132
rect 8525 8188 8589 8192
rect 8525 8132 8529 8188
rect 8529 8132 8585 8188
rect 8585 8132 8589 8188
rect 8525 8128 8589 8132
rect 15618 8188 15682 8192
rect 15618 8132 15622 8188
rect 15622 8132 15678 8188
rect 15678 8132 15682 8188
rect 15618 8128 15682 8132
rect 15698 8188 15762 8192
rect 15698 8132 15702 8188
rect 15702 8132 15758 8188
rect 15758 8132 15762 8188
rect 15698 8128 15762 8132
rect 15778 8188 15842 8192
rect 15778 8132 15782 8188
rect 15782 8132 15838 8188
rect 15838 8132 15842 8188
rect 15778 8128 15842 8132
rect 15858 8188 15922 8192
rect 15858 8132 15862 8188
rect 15862 8132 15918 8188
rect 15918 8132 15922 8188
rect 15858 8128 15922 8132
rect 4618 7644 4682 7648
rect 4618 7588 4622 7644
rect 4622 7588 4678 7644
rect 4678 7588 4682 7644
rect 4618 7584 4682 7588
rect 4698 7644 4762 7648
rect 4698 7588 4702 7644
rect 4702 7588 4758 7644
rect 4758 7588 4762 7644
rect 4698 7584 4762 7588
rect 4778 7644 4842 7648
rect 4778 7588 4782 7644
rect 4782 7588 4838 7644
rect 4838 7588 4842 7644
rect 4778 7584 4842 7588
rect 4858 7644 4922 7648
rect 4858 7588 4862 7644
rect 4862 7588 4918 7644
rect 4918 7588 4922 7644
rect 4858 7584 4922 7588
rect 11952 7644 12016 7648
rect 11952 7588 11956 7644
rect 11956 7588 12012 7644
rect 12012 7588 12016 7644
rect 11952 7584 12016 7588
rect 12032 7644 12096 7648
rect 12032 7588 12036 7644
rect 12036 7588 12092 7644
rect 12092 7588 12096 7644
rect 12032 7584 12096 7588
rect 12112 7644 12176 7648
rect 12112 7588 12116 7644
rect 12116 7588 12172 7644
rect 12172 7588 12176 7644
rect 12112 7584 12176 7588
rect 12192 7644 12256 7648
rect 12192 7588 12196 7644
rect 12196 7588 12252 7644
rect 12252 7588 12256 7644
rect 12192 7584 12256 7588
rect 19285 7644 19349 7648
rect 19285 7588 19289 7644
rect 19289 7588 19345 7644
rect 19345 7588 19349 7644
rect 19285 7584 19349 7588
rect 19365 7644 19429 7648
rect 19365 7588 19369 7644
rect 19369 7588 19425 7644
rect 19425 7588 19429 7644
rect 19365 7584 19429 7588
rect 19445 7644 19509 7648
rect 19445 7588 19449 7644
rect 19449 7588 19505 7644
rect 19505 7588 19509 7644
rect 19445 7584 19509 7588
rect 19525 7644 19589 7648
rect 19525 7588 19529 7644
rect 19529 7588 19585 7644
rect 19585 7588 19589 7644
rect 19525 7584 19589 7588
rect 8285 7100 8349 7104
rect 8285 7044 8289 7100
rect 8289 7044 8345 7100
rect 8345 7044 8349 7100
rect 8285 7040 8349 7044
rect 8365 7100 8429 7104
rect 8365 7044 8369 7100
rect 8369 7044 8425 7100
rect 8425 7044 8429 7100
rect 8365 7040 8429 7044
rect 8445 7100 8509 7104
rect 8445 7044 8449 7100
rect 8449 7044 8505 7100
rect 8505 7044 8509 7100
rect 8445 7040 8509 7044
rect 8525 7100 8589 7104
rect 8525 7044 8529 7100
rect 8529 7044 8585 7100
rect 8585 7044 8589 7100
rect 8525 7040 8589 7044
rect 15618 7100 15682 7104
rect 15618 7044 15622 7100
rect 15622 7044 15678 7100
rect 15678 7044 15682 7100
rect 15618 7040 15682 7044
rect 15698 7100 15762 7104
rect 15698 7044 15702 7100
rect 15702 7044 15758 7100
rect 15758 7044 15762 7100
rect 15698 7040 15762 7044
rect 15778 7100 15842 7104
rect 15778 7044 15782 7100
rect 15782 7044 15838 7100
rect 15838 7044 15842 7100
rect 15778 7040 15842 7044
rect 15858 7100 15922 7104
rect 15858 7044 15862 7100
rect 15862 7044 15918 7100
rect 15918 7044 15922 7100
rect 15858 7040 15922 7044
rect 4618 6556 4682 6560
rect 4618 6500 4622 6556
rect 4622 6500 4678 6556
rect 4678 6500 4682 6556
rect 4618 6496 4682 6500
rect 4698 6556 4762 6560
rect 4698 6500 4702 6556
rect 4702 6500 4758 6556
rect 4758 6500 4762 6556
rect 4698 6496 4762 6500
rect 4778 6556 4842 6560
rect 4778 6500 4782 6556
rect 4782 6500 4838 6556
rect 4838 6500 4842 6556
rect 4778 6496 4842 6500
rect 4858 6556 4922 6560
rect 4858 6500 4862 6556
rect 4862 6500 4918 6556
rect 4918 6500 4922 6556
rect 4858 6496 4922 6500
rect 11952 6556 12016 6560
rect 11952 6500 11956 6556
rect 11956 6500 12012 6556
rect 12012 6500 12016 6556
rect 11952 6496 12016 6500
rect 12032 6556 12096 6560
rect 12032 6500 12036 6556
rect 12036 6500 12092 6556
rect 12092 6500 12096 6556
rect 12032 6496 12096 6500
rect 12112 6556 12176 6560
rect 12112 6500 12116 6556
rect 12116 6500 12172 6556
rect 12172 6500 12176 6556
rect 12112 6496 12176 6500
rect 12192 6556 12256 6560
rect 12192 6500 12196 6556
rect 12196 6500 12252 6556
rect 12252 6500 12256 6556
rect 12192 6496 12256 6500
rect 19285 6556 19349 6560
rect 19285 6500 19289 6556
rect 19289 6500 19345 6556
rect 19345 6500 19349 6556
rect 19285 6496 19349 6500
rect 19365 6556 19429 6560
rect 19365 6500 19369 6556
rect 19369 6500 19425 6556
rect 19425 6500 19429 6556
rect 19365 6496 19429 6500
rect 19445 6556 19509 6560
rect 19445 6500 19449 6556
rect 19449 6500 19505 6556
rect 19505 6500 19509 6556
rect 19445 6496 19509 6500
rect 19525 6556 19589 6560
rect 19525 6500 19529 6556
rect 19529 6500 19585 6556
rect 19585 6500 19589 6556
rect 19525 6496 19589 6500
rect 8285 6012 8349 6016
rect 8285 5956 8289 6012
rect 8289 5956 8345 6012
rect 8345 5956 8349 6012
rect 8285 5952 8349 5956
rect 8365 6012 8429 6016
rect 8365 5956 8369 6012
rect 8369 5956 8425 6012
rect 8425 5956 8429 6012
rect 8365 5952 8429 5956
rect 8445 6012 8509 6016
rect 8445 5956 8449 6012
rect 8449 5956 8505 6012
rect 8505 5956 8509 6012
rect 8445 5952 8509 5956
rect 8525 6012 8589 6016
rect 8525 5956 8529 6012
rect 8529 5956 8585 6012
rect 8585 5956 8589 6012
rect 8525 5952 8589 5956
rect 15618 6012 15682 6016
rect 15618 5956 15622 6012
rect 15622 5956 15678 6012
rect 15678 5956 15682 6012
rect 15618 5952 15682 5956
rect 15698 6012 15762 6016
rect 15698 5956 15702 6012
rect 15702 5956 15758 6012
rect 15758 5956 15762 6012
rect 15698 5952 15762 5956
rect 15778 6012 15842 6016
rect 15778 5956 15782 6012
rect 15782 5956 15838 6012
rect 15838 5956 15842 6012
rect 15778 5952 15842 5956
rect 15858 6012 15922 6016
rect 15858 5956 15862 6012
rect 15862 5956 15918 6012
rect 15918 5956 15922 6012
rect 15858 5952 15922 5956
rect 4108 5748 4172 5812
rect 4618 5468 4682 5472
rect 4618 5412 4622 5468
rect 4622 5412 4678 5468
rect 4678 5412 4682 5468
rect 4618 5408 4682 5412
rect 4698 5468 4762 5472
rect 4698 5412 4702 5468
rect 4702 5412 4758 5468
rect 4758 5412 4762 5468
rect 4698 5408 4762 5412
rect 4778 5468 4842 5472
rect 4778 5412 4782 5468
rect 4782 5412 4838 5468
rect 4838 5412 4842 5468
rect 4778 5408 4842 5412
rect 4858 5468 4922 5472
rect 4858 5412 4862 5468
rect 4862 5412 4918 5468
rect 4918 5412 4922 5468
rect 4858 5408 4922 5412
rect 11952 5468 12016 5472
rect 11952 5412 11956 5468
rect 11956 5412 12012 5468
rect 12012 5412 12016 5468
rect 11952 5408 12016 5412
rect 12032 5468 12096 5472
rect 12032 5412 12036 5468
rect 12036 5412 12092 5468
rect 12092 5412 12096 5468
rect 12032 5408 12096 5412
rect 12112 5468 12176 5472
rect 12112 5412 12116 5468
rect 12116 5412 12172 5468
rect 12172 5412 12176 5468
rect 12112 5408 12176 5412
rect 12192 5468 12256 5472
rect 12192 5412 12196 5468
rect 12196 5412 12252 5468
rect 12252 5412 12256 5468
rect 12192 5408 12256 5412
rect 19285 5468 19349 5472
rect 19285 5412 19289 5468
rect 19289 5412 19345 5468
rect 19345 5412 19349 5468
rect 19285 5408 19349 5412
rect 19365 5468 19429 5472
rect 19365 5412 19369 5468
rect 19369 5412 19425 5468
rect 19425 5412 19429 5468
rect 19365 5408 19429 5412
rect 19445 5468 19509 5472
rect 19445 5412 19449 5468
rect 19449 5412 19505 5468
rect 19505 5412 19509 5468
rect 19445 5408 19509 5412
rect 19525 5468 19589 5472
rect 19525 5412 19529 5468
rect 19529 5412 19585 5468
rect 19585 5412 19589 5468
rect 19525 5408 19589 5412
rect 21588 5204 21652 5268
rect 17172 5068 17236 5132
rect 8285 4924 8349 4928
rect 8285 4868 8289 4924
rect 8289 4868 8345 4924
rect 8345 4868 8349 4924
rect 8285 4864 8349 4868
rect 8365 4924 8429 4928
rect 8365 4868 8369 4924
rect 8369 4868 8425 4924
rect 8425 4868 8429 4924
rect 8365 4864 8429 4868
rect 8445 4924 8509 4928
rect 8445 4868 8449 4924
rect 8449 4868 8505 4924
rect 8505 4868 8509 4924
rect 8445 4864 8509 4868
rect 8525 4924 8589 4928
rect 8525 4868 8529 4924
rect 8529 4868 8585 4924
rect 8585 4868 8589 4924
rect 8525 4864 8589 4868
rect 15618 4924 15682 4928
rect 15618 4868 15622 4924
rect 15622 4868 15678 4924
rect 15678 4868 15682 4924
rect 15618 4864 15682 4868
rect 15698 4924 15762 4928
rect 15698 4868 15702 4924
rect 15702 4868 15758 4924
rect 15758 4868 15762 4924
rect 15698 4864 15762 4868
rect 15778 4924 15842 4928
rect 15778 4868 15782 4924
rect 15782 4868 15838 4924
rect 15838 4868 15842 4924
rect 15778 4864 15842 4868
rect 15858 4924 15922 4928
rect 15858 4868 15862 4924
rect 15862 4868 15918 4924
rect 15918 4868 15922 4924
rect 15858 4864 15922 4868
rect 4108 4388 4172 4452
rect 15332 4388 15396 4452
rect 4618 4380 4682 4384
rect 4618 4324 4622 4380
rect 4622 4324 4678 4380
rect 4678 4324 4682 4380
rect 4618 4320 4682 4324
rect 4698 4380 4762 4384
rect 4698 4324 4702 4380
rect 4702 4324 4758 4380
rect 4758 4324 4762 4380
rect 4698 4320 4762 4324
rect 4778 4380 4842 4384
rect 4778 4324 4782 4380
rect 4782 4324 4838 4380
rect 4838 4324 4842 4380
rect 4778 4320 4842 4324
rect 4858 4380 4922 4384
rect 4858 4324 4862 4380
rect 4862 4324 4918 4380
rect 4918 4324 4922 4380
rect 4858 4320 4922 4324
rect 11952 4380 12016 4384
rect 11952 4324 11956 4380
rect 11956 4324 12012 4380
rect 12012 4324 12016 4380
rect 11952 4320 12016 4324
rect 12032 4380 12096 4384
rect 12032 4324 12036 4380
rect 12036 4324 12092 4380
rect 12092 4324 12096 4380
rect 12032 4320 12096 4324
rect 12112 4380 12176 4384
rect 12112 4324 12116 4380
rect 12116 4324 12172 4380
rect 12172 4324 12176 4380
rect 12112 4320 12176 4324
rect 12192 4380 12256 4384
rect 12192 4324 12196 4380
rect 12196 4324 12252 4380
rect 12252 4324 12256 4380
rect 12192 4320 12256 4324
rect 19285 4380 19349 4384
rect 19285 4324 19289 4380
rect 19289 4324 19345 4380
rect 19345 4324 19349 4380
rect 19285 4320 19349 4324
rect 19365 4380 19429 4384
rect 19365 4324 19369 4380
rect 19369 4324 19425 4380
rect 19425 4324 19429 4380
rect 19365 4320 19429 4324
rect 19445 4380 19509 4384
rect 19445 4324 19449 4380
rect 19449 4324 19505 4380
rect 19505 4324 19509 4380
rect 19445 4320 19509 4324
rect 19525 4380 19589 4384
rect 19525 4324 19529 4380
rect 19529 4324 19585 4380
rect 19585 4324 19589 4380
rect 19525 4320 19589 4324
rect 9628 4116 9692 4180
rect 21404 4116 21468 4180
rect 6132 3844 6196 3908
rect 9628 3980 9692 4044
rect 8285 3836 8349 3840
rect 8285 3780 8289 3836
rect 8289 3780 8345 3836
rect 8345 3780 8349 3836
rect 8285 3776 8349 3780
rect 8365 3836 8429 3840
rect 8365 3780 8369 3836
rect 8369 3780 8425 3836
rect 8425 3780 8429 3836
rect 8365 3776 8429 3780
rect 8445 3836 8509 3840
rect 8445 3780 8449 3836
rect 8449 3780 8505 3836
rect 8505 3780 8509 3836
rect 8445 3776 8509 3780
rect 8525 3836 8589 3840
rect 8525 3780 8529 3836
rect 8529 3780 8585 3836
rect 8585 3780 8589 3836
rect 8525 3776 8589 3780
rect 15618 3836 15682 3840
rect 15618 3780 15622 3836
rect 15622 3780 15678 3836
rect 15678 3780 15682 3836
rect 15618 3776 15682 3780
rect 15698 3836 15762 3840
rect 15698 3780 15702 3836
rect 15702 3780 15758 3836
rect 15758 3780 15762 3836
rect 15698 3776 15762 3780
rect 15778 3836 15842 3840
rect 15778 3780 15782 3836
rect 15782 3780 15838 3836
rect 15838 3780 15842 3836
rect 15778 3776 15842 3780
rect 15858 3836 15922 3840
rect 15858 3780 15862 3836
rect 15862 3780 15918 3836
rect 15918 3780 15922 3836
rect 15858 3776 15922 3780
rect 4618 3292 4682 3296
rect 4618 3236 4622 3292
rect 4622 3236 4678 3292
rect 4678 3236 4682 3292
rect 4618 3232 4682 3236
rect 4698 3292 4762 3296
rect 4698 3236 4702 3292
rect 4702 3236 4758 3292
rect 4758 3236 4762 3292
rect 4698 3232 4762 3236
rect 4778 3292 4842 3296
rect 4778 3236 4782 3292
rect 4782 3236 4838 3292
rect 4838 3236 4842 3292
rect 4778 3232 4842 3236
rect 4858 3292 4922 3296
rect 4858 3236 4862 3292
rect 4862 3236 4918 3292
rect 4918 3236 4922 3292
rect 4858 3232 4922 3236
rect 11952 3292 12016 3296
rect 11952 3236 11956 3292
rect 11956 3236 12012 3292
rect 12012 3236 12016 3292
rect 11952 3232 12016 3236
rect 12032 3292 12096 3296
rect 12032 3236 12036 3292
rect 12036 3236 12092 3292
rect 12092 3236 12096 3292
rect 12032 3232 12096 3236
rect 12112 3292 12176 3296
rect 12112 3236 12116 3292
rect 12116 3236 12172 3292
rect 12172 3236 12176 3292
rect 12112 3232 12176 3236
rect 12192 3292 12256 3296
rect 12192 3236 12196 3292
rect 12196 3236 12252 3292
rect 12252 3236 12256 3292
rect 12192 3232 12256 3236
rect 19285 3292 19349 3296
rect 19285 3236 19289 3292
rect 19289 3236 19345 3292
rect 19345 3236 19349 3292
rect 19285 3232 19349 3236
rect 19365 3292 19429 3296
rect 19365 3236 19369 3292
rect 19369 3236 19425 3292
rect 19425 3236 19429 3292
rect 19365 3232 19429 3236
rect 19445 3292 19509 3296
rect 19445 3236 19449 3292
rect 19449 3236 19505 3292
rect 19505 3236 19509 3292
rect 19445 3232 19509 3236
rect 19525 3292 19589 3296
rect 19525 3236 19529 3292
rect 19529 3236 19585 3292
rect 19585 3236 19589 3292
rect 19525 3232 19589 3236
rect 4108 3028 4172 3092
rect 14780 3028 14844 3092
rect 8285 2748 8349 2752
rect 8285 2692 8289 2748
rect 8289 2692 8345 2748
rect 8345 2692 8349 2748
rect 8285 2688 8349 2692
rect 8365 2748 8429 2752
rect 8365 2692 8369 2748
rect 8369 2692 8425 2748
rect 8425 2692 8429 2748
rect 8365 2688 8429 2692
rect 8445 2748 8509 2752
rect 8445 2692 8449 2748
rect 8449 2692 8505 2748
rect 8505 2692 8509 2748
rect 8445 2688 8509 2692
rect 8525 2748 8589 2752
rect 8525 2692 8529 2748
rect 8529 2692 8585 2748
rect 8585 2692 8589 2748
rect 8525 2688 8589 2692
rect 15618 2748 15682 2752
rect 15618 2692 15622 2748
rect 15622 2692 15678 2748
rect 15678 2692 15682 2748
rect 15618 2688 15682 2692
rect 15698 2748 15762 2752
rect 15698 2692 15702 2748
rect 15702 2692 15758 2748
rect 15758 2692 15762 2748
rect 15698 2688 15762 2692
rect 15778 2748 15842 2752
rect 15778 2692 15782 2748
rect 15782 2692 15838 2748
rect 15838 2692 15842 2748
rect 15778 2688 15842 2692
rect 15858 2748 15922 2752
rect 15858 2692 15862 2748
rect 15862 2692 15918 2748
rect 15918 2692 15922 2748
rect 15858 2688 15922 2692
rect 4618 2204 4682 2208
rect 4618 2148 4622 2204
rect 4622 2148 4678 2204
rect 4678 2148 4682 2204
rect 4618 2144 4682 2148
rect 4698 2204 4762 2208
rect 4698 2148 4702 2204
rect 4702 2148 4758 2204
rect 4758 2148 4762 2204
rect 4698 2144 4762 2148
rect 4778 2204 4842 2208
rect 4778 2148 4782 2204
rect 4782 2148 4838 2204
rect 4838 2148 4842 2204
rect 4778 2144 4842 2148
rect 4858 2204 4922 2208
rect 4858 2148 4862 2204
rect 4862 2148 4918 2204
rect 4918 2148 4922 2204
rect 4858 2144 4922 2148
rect 11952 2204 12016 2208
rect 11952 2148 11956 2204
rect 11956 2148 12012 2204
rect 12012 2148 12016 2204
rect 11952 2144 12016 2148
rect 12032 2204 12096 2208
rect 12032 2148 12036 2204
rect 12036 2148 12092 2204
rect 12092 2148 12096 2204
rect 12032 2144 12096 2148
rect 12112 2204 12176 2208
rect 12112 2148 12116 2204
rect 12116 2148 12172 2204
rect 12172 2148 12176 2204
rect 12112 2144 12176 2148
rect 12192 2204 12256 2208
rect 12192 2148 12196 2204
rect 12196 2148 12252 2204
rect 12252 2148 12256 2204
rect 12192 2144 12256 2148
rect 19285 2204 19349 2208
rect 19285 2148 19289 2204
rect 19289 2148 19345 2204
rect 19345 2148 19349 2204
rect 19285 2144 19349 2148
rect 19365 2204 19429 2208
rect 19365 2148 19369 2204
rect 19369 2148 19425 2204
rect 19425 2148 19429 2204
rect 19365 2144 19429 2148
rect 19445 2204 19509 2208
rect 19445 2148 19449 2204
rect 19449 2148 19505 2204
rect 19505 2148 19509 2204
rect 19445 2144 19509 2148
rect 19525 2204 19589 2208
rect 19525 2148 19529 2204
rect 19529 2148 19585 2204
rect 19585 2148 19589 2204
rect 19525 2144 19589 2148
<< metal4 >>
rect 4610 19616 4931 19632
rect 4610 19552 4618 19616
rect 4682 19552 4698 19616
rect 4762 19552 4778 19616
rect 4842 19552 4858 19616
rect 4922 19552 4931 19616
rect 4610 18528 4931 19552
rect 4610 18464 4618 18528
rect 4682 18464 4698 18528
rect 4762 18464 4778 18528
rect 4842 18464 4858 18528
rect 4922 18464 4931 18528
rect 4610 17440 4931 18464
rect 4610 17376 4618 17440
rect 4682 17376 4698 17440
rect 4762 17376 4778 17440
rect 4842 17376 4858 17440
rect 4922 17376 4931 17440
rect 4610 16352 4931 17376
rect 4610 16288 4618 16352
rect 4682 16288 4698 16352
rect 4762 16288 4778 16352
rect 4842 16288 4858 16352
rect 4922 16288 4931 16352
rect 4610 15264 4931 16288
rect 4610 15200 4618 15264
rect 4682 15200 4698 15264
rect 4762 15200 4778 15264
rect 4842 15200 4858 15264
rect 4922 15200 4931 15264
rect 4610 14176 4931 15200
rect 4610 14112 4618 14176
rect 4682 14112 4698 14176
rect 4762 14112 4778 14176
rect 4842 14112 4858 14176
rect 4922 14112 4931 14176
rect 59 13700 125 13701
rect 59 13636 60 13700
rect 124 13636 125 13700
rect 59 13635 125 13636
rect 62 13429 122 13635
rect 59 13428 125 13429
rect 59 13364 60 13428
rect 124 13364 125 13428
rect 59 13363 125 13364
rect 4610 13088 4931 14112
rect 4610 13024 4618 13088
rect 4682 13024 4698 13088
rect 4762 13024 4778 13088
rect 4842 13024 4858 13088
rect 4922 13024 4931 13088
rect 4610 12000 4931 13024
rect 8277 19072 8597 19632
rect 8277 19008 8285 19072
rect 8349 19008 8365 19072
rect 8429 19008 8445 19072
rect 8509 19008 8525 19072
rect 8589 19008 8597 19072
rect 8277 17984 8597 19008
rect 8277 17920 8285 17984
rect 8349 17920 8365 17984
rect 8429 17920 8445 17984
rect 8509 17920 8525 17984
rect 8589 17920 8597 17984
rect 8277 16896 8597 17920
rect 8277 16832 8285 16896
rect 8349 16832 8365 16896
rect 8429 16832 8445 16896
rect 8509 16832 8525 16896
rect 8589 16832 8597 16896
rect 8277 15808 8597 16832
rect 8277 15744 8285 15808
rect 8349 15744 8365 15808
rect 8429 15744 8445 15808
rect 8509 15744 8525 15808
rect 8589 15744 8597 15808
rect 8277 14720 8597 15744
rect 8277 14656 8285 14720
rect 8349 14656 8365 14720
rect 8429 14656 8445 14720
rect 8509 14656 8525 14720
rect 8589 14656 8597 14720
rect 8277 13632 8597 14656
rect 8277 13568 8285 13632
rect 8349 13568 8365 13632
rect 8429 13568 8445 13632
rect 8509 13568 8525 13632
rect 8589 13568 8597 13632
rect 6131 12884 6197 12885
rect 6131 12820 6132 12884
rect 6196 12820 6197 12884
rect 6131 12819 6197 12820
rect 4610 11936 4618 12000
rect 4682 11936 4698 12000
rect 4762 11936 4778 12000
rect 4842 11936 4858 12000
rect 4922 11936 4931 12000
rect 4610 10912 4931 11936
rect 4610 10848 4618 10912
rect 4682 10848 4698 10912
rect 4762 10848 4778 10912
rect 4842 10848 4858 10912
rect 4922 10848 4931 10912
rect 4610 9824 4931 10848
rect 4610 9760 4618 9824
rect 4682 9760 4698 9824
rect 4762 9760 4778 9824
rect 4842 9760 4858 9824
rect 4922 9760 4931 9824
rect 4610 8736 4931 9760
rect 4610 8672 4618 8736
rect 4682 8672 4698 8736
rect 4762 8672 4778 8736
rect 4842 8672 4858 8736
rect 4922 8672 4931 8736
rect 4610 7648 4931 8672
rect 4610 7584 4618 7648
rect 4682 7584 4698 7648
rect 4762 7584 4778 7648
rect 4842 7584 4858 7648
rect 4922 7584 4931 7648
rect 4610 6560 4931 7584
rect 4610 6496 4618 6560
rect 4682 6496 4698 6560
rect 4762 6496 4778 6560
rect 4842 6496 4858 6560
rect 4922 6496 4931 6560
rect 4107 5812 4173 5813
rect 4107 5748 4108 5812
rect 4172 5748 4173 5812
rect 4107 5747 4173 5748
rect 4110 5218 4170 5747
rect 4610 5472 4931 6496
rect 4610 5408 4618 5472
rect 4682 5408 4698 5472
rect 4762 5408 4778 5472
rect 4842 5408 4858 5472
rect 4922 5408 4931 5472
rect 4610 4384 4931 5408
rect 4610 4320 4618 4384
rect 4682 4320 4698 4384
rect 4762 4320 4778 4384
rect 4842 4320 4858 4384
rect 4922 4320 4931 4384
rect 4610 3296 4931 4320
rect 6134 3909 6194 12819
rect 8277 12544 8597 13568
rect 8277 12480 8285 12544
rect 8349 12480 8365 12544
rect 8429 12480 8445 12544
rect 8509 12480 8525 12544
rect 8589 12480 8597 12544
rect 8277 11456 8597 12480
rect 8277 11392 8285 11456
rect 8349 11392 8365 11456
rect 8429 11392 8445 11456
rect 8509 11392 8525 11456
rect 8589 11392 8597 11456
rect 8277 10368 8597 11392
rect 8277 10304 8285 10368
rect 8349 10304 8365 10368
rect 8429 10304 8445 10368
rect 8509 10304 8525 10368
rect 8589 10304 8597 10368
rect 8277 9280 8597 10304
rect 8277 9216 8285 9280
rect 8349 9216 8365 9280
rect 8429 9216 8445 9280
rect 8509 9216 8525 9280
rect 8589 9216 8597 9280
rect 8277 8192 8597 9216
rect 8277 8128 8285 8192
rect 8349 8128 8365 8192
rect 8429 8128 8445 8192
rect 8509 8128 8525 8192
rect 8589 8128 8597 8192
rect 8277 7104 8597 8128
rect 8277 7040 8285 7104
rect 8349 7040 8365 7104
rect 8429 7040 8445 7104
rect 8509 7040 8525 7104
rect 8589 7040 8597 7104
rect 8277 6016 8597 7040
rect 8277 5952 8285 6016
rect 8349 5952 8365 6016
rect 8429 5952 8445 6016
rect 8509 5952 8525 6016
rect 8589 5952 8597 6016
rect 8277 4928 8597 5952
rect 8277 4864 8285 4928
rect 8349 4864 8365 4928
rect 8429 4864 8445 4928
rect 8509 4864 8525 4928
rect 8589 4864 8597 4928
rect 6131 3908 6197 3909
rect 6131 3844 6132 3908
rect 6196 3844 6197 3908
rect 6131 3843 6197 3844
rect 4610 3232 4618 3296
rect 4682 3232 4698 3296
rect 4762 3232 4778 3296
rect 4842 3232 4858 3296
rect 4922 3232 4931 3296
rect 4610 2208 4931 3232
rect 4610 2144 4618 2208
rect 4682 2144 4698 2208
rect 4762 2144 4778 2208
rect 4842 2144 4858 2208
rect 4922 2144 4931 2208
rect 4610 2128 4931 2144
rect 8277 3840 8597 4864
rect 11944 19616 12264 19632
rect 11944 19552 11952 19616
rect 12016 19552 12032 19616
rect 12096 19552 12112 19616
rect 12176 19552 12192 19616
rect 12256 19552 12264 19616
rect 11944 18528 12264 19552
rect 11944 18464 11952 18528
rect 12016 18464 12032 18528
rect 12096 18464 12112 18528
rect 12176 18464 12192 18528
rect 12256 18464 12264 18528
rect 11944 17440 12264 18464
rect 11944 17376 11952 17440
rect 12016 17376 12032 17440
rect 12096 17376 12112 17440
rect 12176 17376 12192 17440
rect 12256 17376 12264 17440
rect 11944 16352 12264 17376
rect 11944 16288 11952 16352
rect 12016 16288 12032 16352
rect 12096 16288 12112 16352
rect 12176 16288 12192 16352
rect 12256 16288 12264 16352
rect 11944 15264 12264 16288
rect 11944 15200 11952 15264
rect 12016 15200 12032 15264
rect 12096 15200 12112 15264
rect 12176 15200 12192 15264
rect 12256 15200 12264 15264
rect 11944 14176 12264 15200
rect 11944 14112 11952 14176
rect 12016 14112 12032 14176
rect 12096 14112 12112 14176
rect 12176 14112 12192 14176
rect 12256 14112 12264 14176
rect 11944 13088 12264 14112
rect 11944 13024 11952 13088
rect 12016 13024 12032 13088
rect 12096 13024 12112 13088
rect 12176 13024 12192 13088
rect 12256 13024 12264 13088
rect 11944 12000 12264 13024
rect 11944 11936 11952 12000
rect 12016 11936 12032 12000
rect 12096 11936 12112 12000
rect 12176 11936 12192 12000
rect 12256 11936 12264 12000
rect 11944 10912 12264 11936
rect 11944 10848 11952 10912
rect 12016 10848 12032 10912
rect 12096 10848 12112 10912
rect 12176 10848 12192 10912
rect 12256 10848 12264 10912
rect 11944 9824 12264 10848
rect 11944 9760 11952 9824
rect 12016 9760 12032 9824
rect 12096 9760 12112 9824
rect 12176 9760 12192 9824
rect 12256 9760 12264 9824
rect 11944 8736 12264 9760
rect 11944 8672 11952 8736
rect 12016 8672 12032 8736
rect 12096 8672 12112 8736
rect 12176 8672 12192 8736
rect 12256 8672 12264 8736
rect 11944 7648 12264 8672
rect 11944 7584 11952 7648
rect 12016 7584 12032 7648
rect 12096 7584 12112 7648
rect 12176 7584 12192 7648
rect 12256 7584 12264 7648
rect 11944 6560 12264 7584
rect 11944 6496 11952 6560
rect 12016 6496 12032 6560
rect 12096 6496 12112 6560
rect 12176 6496 12192 6560
rect 12256 6496 12264 6560
rect 11944 5472 12264 6496
rect 11944 5408 11952 5472
rect 12016 5408 12032 5472
rect 12096 5408 12112 5472
rect 12176 5408 12192 5472
rect 12256 5408 12264 5472
rect 11944 4384 12264 5408
rect 15610 19072 15930 19632
rect 15610 19008 15618 19072
rect 15682 19008 15698 19072
rect 15762 19008 15778 19072
rect 15842 19008 15858 19072
rect 15922 19008 15930 19072
rect 15610 17984 15930 19008
rect 15610 17920 15618 17984
rect 15682 17920 15698 17984
rect 15762 17920 15778 17984
rect 15842 17920 15858 17984
rect 15922 17920 15930 17984
rect 15610 16896 15930 17920
rect 15610 16832 15618 16896
rect 15682 16832 15698 16896
rect 15762 16832 15778 16896
rect 15842 16832 15858 16896
rect 15922 16832 15930 16896
rect 15610 15808 15930 16832
rect 15610 15744 15618 15808
rect 15682 15744 15698 15808
rect 15762 15744 15778 15808
rect 15842 15744 15858 15808
rect 15922 15744 15930 15808
rect 15610 14720 15930 15744
rect 15610 14656 15618 14720
rect 15682 14656 15698 14720
rect 15762 14656 15778 14720
rect 15842 14656 15858 14720
rect 15922 14656 15930 14720
rect 15610 13632 15930 14656
rect 15610 13568 15618 13632
rect 15682 13568 15698 13632
rect 15762 13568 15778 13632
rect 15842 13568 15858 13632
rect 15922 13568 15930 13632
rect 15610 12544 15930 13568
rect 15610 12480 15618 12544
rect 15682 12480 15698 12544
rect 15762 12480 15778 12544
rect 15842 12480 15858 12544
rect 15922 12480 15930 12544
rect 15610 11456 15930 12480
rect 15610 11392 15618 11456
rect 15682 11392 15698 11456
rect 15762 11392 15778 11456
rect 15842 11392 15858 11456
rect 15922 11392 15930 11456
rect 15610 10368 15930 11392
rect 15610 10304 15618 10368
rect 15682 10304 15698 10368
rect 15762 10304 15778 10368
rect 15842 10304 15858 10368
rect 15922 10304 15930 10368
rect 15610 9280 15930 10304
rect 15610 9216 15618 9280
rect 15682 9216 15698 9280
rect 15762 9216 15778 9280
rect 15842 9216 15858 9280
rect 15922 9216 15930 9280
rect 15610 8192 15930 9216
rect 15610 8128 15618 8192
rect 15682 8128 15698 8192
rect 15762 8128 15778 8192
rect 15842 8128 15858 8192
rect 15922 8128 15930 8192
rect 15610 7104 15930 8128
rect 15610 7040 15618 7104
rect 15682 7040 15698 7104
rect 15762 7040 15778 7104
rect 15842 7040 15858 7104
rect 15922 7040 15930 7104
rect 15610 6016 15930 7040
rect 15610 5952 15618 6016
rect 15682 5952 15698 6016
rect 15762 5952 15778 6016
rect 15842 5952 15858 6016
rect 15922 5952 15930 6016
rect 15610 4928 15930 5952
rect 19277 19616 19597 19632
rect 19277 19552 19285 19616
rect 19349 19552 19365 19616
rect 19429 19552 19445 19616
rect 19509 19552 19525 19616
rect 19589 19552 19597 19616
rect 19277 18528 19597 19552
rect 19277 18464 19285 18528
rect 19349 18464 19365 18528
rect 19429 18464 19445 18528
rect 19509 18464 19525 18528
rect 19589 18464 19597 18528
rect 19277 17440 19597 18464
rect 19277 17376 19285 17440
rect 19349 17376 19365 17440
rect 19429 17376 19445 17440
rect 19509 17376 19525 17440
rect 19589 17376 19597 17440
rect 19277 16352 19597 17376
rect 19277 16288 19285 16352
rect 19349 16288 19365 16352
rect 19429 16288 19445 16352
rect 19509 16288 19525 16352
rect 19589 16288 19597 16352
rect 19277 15264 19597 16288
rect 19277 15200 19285 15264
rect 19349 15200 19365 15264
rect 19429 15200 19445 15264
rect 19509 15200 19525 15264
rect 19589 15200 19597 15264
rect 19277 14176 19597 15200
rect 21587 14788 21653 14789
rect 21587 14724 21588 14788
rect 21652 14724 21653 14788
rect 21587 14723 21653 14724
rect 21403 14652 21469 14653
rect 21403 14588 21404 14652
rect 21468 14650 21469 14652
rect 21590 14650 21650 14723
rect 21468 14590 21650 14650
rect 21468 14588 21469 14590
rect 21403 14587 21469 14588
rect 19277 14112 19285 14176
rect 19349 14112 19365 14176
rect 19429 14112 19445 14176
rect 19509 14112 19525 14176
rect 19589 14112 19597 14176
rect 19277 13088 19597 14112
rect 19277 13024 19285 13088
rect 19349 13024 19365 13088
rect 19429 13024 19445 13088
rect 19509 13024 19525 13088
rect 19589 13024 19597 13088
rect 19277 12000 19597 13024
rect 19277 11936 19285 12000
rect 19349 11936 19365 12000
rect 19429 11936 19445 12000
rect 19509 11936 19525 12000
rect 19589 11936 19597 12000
rect 19277 10912 19597 11936
rect 19277 10848 19285 10912
rect 19349 10848 19365 10912
rect 19429 10848 19445 10912
rect 19509 10848 19525 10912
rect 19589 10848 19597 10912
rect 19277 9824 19597 10848
rect 19277 9760 19285 9824
rect 19349 9760 19365 9824
rect 19429 9760 19445 9824
rect 19509 9760 19525 9824
rect 19589 9760 19597 9824
rect 19277 8736 19597 9760
rect 21587 9076 21653 9077
rect 21587 9012 21588 9076
rect 21652 9012 21653 9076
rect 21587 9011 21653 9012
rect 21590 8907 21650 9011
rect 21587 8906 21653 8907
rect 21587 8842 21588 8906
rect 21652 8842 21653 8906
rect 21587 8841 21653 8842
rect 19277 8672 19285 8736
rect 19349 8672 19365 8736
rect 19429 8672 19445 8736
rect 19509 8672 19525 8736
rect 19589 8672 19597 8736
rect 19277 7648 19597 8672
rect 19277 7584 19285 7648
rect 19349 7584 19365 7648
rect 19429 7584 19445 7648
rect 19509 7584 19525 7648
rect 19589 7584 19597 7648
rect 19277 6560 19597 7584
rect 19277 6496 19285 6560
rect 19349 6496 19365 6560
rect 19429 6496 19445 6560
rect 19509 6496 19525 6560
rect 19589 6496 19597 6560
rect 19277 5472 19597 6496
rect 19277 5408 19285 5472
rect 19349 5408 19365 5472
rect 19429 5408 19445 5472
rect 19509 5408 19525 5472
rect 19589 5408 19597 5472
rect 15610 4864 15618 4928
rect 15682 4864 15698 4928
rect 15762 4864 15778 4928
rect 15842 4864 15858 4928
rect 15922 4864 15930 4928
rect 11944 4320 11952 4384
rect 12016 4320 12032 4384
rect 12096 4320 12112 4384
rect 12176 4320 12192 4384
rect 12256 4320 12264 4384
rect 9627 4180 9693 4181
rect 9627 4116 9628 4180
rect 9692 4116 9693 4180
rect 9627 4115 9693 4116
rect 9630 4045 9690 4115
rect 9627 4044 9693 4045
rect 9627 3980 9628 4044
rect 9692 3980 9693 4044
rect 9627 3979 9693 3980
rect 8277 3776 8285 3840
rect 8349 3776 8365 3840
rect 8429 3776 8445 3840
rect 8509 3776 8525 3840
rect 8589 3776 8597 3840
rect 8277 2752 8597 3776
rect 8277 2688 8285 2752
rect 8349 2688 8365 2752
rect 8429 2688 8445 2752
rect 8509 2688 8525 2752
rect 8589 2688 8597 2752
rect 8277 2128 8597 2688
rect 11944 3296 12264 4320
rect 11944 3232 11952 3296
rect 12016 3232 12032 3296
rect 12096 3232 12112 3296
rect 12176 3232 12192 3296
rect 12256 3232 12264 3296
rect 11944 2208 12264 3232
rect 15610 3840 15930 4864
rect 15610 3776 15618 3840
rect 15682 3776 15698 3840
rect 15762 3776 15778 3840
rect 15842 3776 15858 3840
rect 15922 3776 15930 3840
rect 11944 2144 11952 2208
rect 12016 2144 12032 2208
rect 12096 2144 12112 2208
rect 12176 2144 12192 2208
rect 12256 2144 12264 2208
rect 11944 2128 12264 2144
rect 15610 2752 15930 3776
rect 15610 2688 15618 2752
rect 15682 2688 15698 2752
rect 15762 2688 15778 2752
rect 15842 2688 15858 2752
rect 15922 2688 15930 2752
rect 15610 2128 15930 2688
rect 19277 4384 19597 5408
rect 21587 5268 21653 5269
rect 21587 5204 21588 5268
rect 21652 5204 21653 5268
rect 21587 5203 21653 5204
rect 21590 5130 21650 5203
rect 19277 4320 19285 4384
rect 19349 4320 19365 4384
rect 19429 4320 19445 4384
rect 19509 4320 19525 4384
rect 19589 4320 19597 4384
rect 19277 3296 19597 4320
rect 21406 5070 21650 5130
rect 21406 4181 21466 5070
rect 21403 4180 21469 4181
rect 21403 4116 21404 4180
rect 21468 4116 21469 4180
rect 21403 4115 21469 4116
rect 19277 3232 19285 3296
rect 19349 3232 19365 3296
rect 19429 3232 19445 3296
rect 19509 3232 19525 3296
rect 19589 3232 19597 3296
rect 19277 2208 19597 3232
rect 19277 2144 19285 2208
rect 19349 2144 19365 2208
rect 19429 2144 19445 2208
rect 19509 2144 19525 2208
rect 19589 2144 19597 2208
rect 19277 2128 19597 2144
<< via4 >>
rect 4022 4982 4258 5218
rect 4022 4452 4258 4538
rect 4022 4388 4108 4452
rect 4108 4388 4172 4452
rect 4172 4388 4258 4452
rect 4022 4302 4258 4388
rect 4022 3092 4258 3178
rect 4022 3028 4108 3092
rect 4108 3028 4172 3092
rect 4172 3028 4258 3092
rect 4022 2942 4258 3028
rect 17086 5132 17322 5218
rect 17086 5068 17172 5132
rect 17172 5068 17236 5132
rect 17236 5068 17322 5132
rect 17086 4982 17322 5068
rect 15246 4452 15482 4538
rect 15246 4388 15332 4452
rect 15332 4388 15396 4452
rect 15396 4388 15482 4452
rect 15246 4302 15482 4388
rect 14694 3092 14930 3178
rect 14694 3028 14780 3092
rect 14780 3028 14844 3092
rect 14844 3028 14930 3092
rect 14694 2942 14930 3028
<< metal5 >>
rect 3980 5218 17364 5260
rect 3980 4982 4022 5218
rect 4258 4982 17086 5218
rect 17322 4982 17364 5218
rect 3980 4940 17364 4982
rect 3980 4538 15524 4580
rect 3980 4302 4022 4538
rect 4258 4302 15246 4538
rect 15482 4302 15524 4538
rect 3980 4260 15524 4302
rect 3980 3178 14972 3220
rect 3980 2942 4022 3178
rect 4258 2942 14694 3178
rect 14930 2942 14972 3178
rect 3980 2900 14972 2942
use scs8hd_decap_4  FILLER_1_3 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1380 0 1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_0_6 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1656 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_3  PHY_2 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1104 0 1 2720
box -38 -48 314 592
use scs8hd_decap_3  PHY_0
timestamp 1586364061
transform 1 0 1104 0 -1 2720
box -38 -48 314 592
use scs8hd_conb_1  _126_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1380 0 -1 2720
box -38 -48 314 592
use scs8hd_fill_1  FILLER_1_7 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1748 0 1 2720
box -38 -48 130 592
use scs8hd_fill_2  FILLER_0_10
timestamp 1586364061
transform 1 0 2024 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__073__B tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 2208 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_1.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 1840 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__119__B
timestamp 1586364061
transform 1 0 1840 0 1 2720
box -38 -48 222 592
use scs8hd_nor2_4  _073_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 2024 0 1 2720
box -38 -48 866 592
use scs8hd_nor2_4  _042_
timestamp 1586364061
transform 1 0 3588 0 1 2720
box -38 -48 866 592
use scs8hd_nor2_4  _072_
timestamp 1586364061
transform 1 0 2392 0 -1 2720
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__119__C
timestamp 1586364061
transform 1 0 3036 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__072__B
timestamp 1586364061
transform 1 0 3404 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__119__A
timestamp 1586364061
transform 1 0 3404 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_23
timestamp 1586364061
transform 1 0 3220 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_27
timestamp 1586364061
transform 1 0 3588 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_19
timestamp 1586364061
transform 1 0 2852 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_23
timestamp 1586364061
transform 1 0 3220 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_32
timestamp 1586364061
transform 1 0 4048 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__072__A
timestamp 1586364061
transform 1 0 3772 0 -1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_64 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 3956 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_4  FILLER_1_36
timestamp 1586364061
transform 1 0 4416 0 1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_0_37
timestamp 1586364061
transform 1 0 4508 0 -1 2720
box -38 -48 222 592
use scs8hd_inv_1  mux_right_ipin_4.tap_buf4_0_.scs8hd_inv_1 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 4232 0 -1 2720
box -38 -48 314 592
use scs8hd_fill_1  FILLER_1_40
timestamp 1586364061
transform 1 0 4784 0 1 2720
box -38 -48 130 592
use scs8hd_fill_2  FILLER_0_41
timestamp 1586364061
transform 1 0 4876 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__044__B
timestamp 1586364061
transform 1 0 4692 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__101__A
timestamp 1586364061
transform 1 0 4876 0 1 2720
box -38 -48 222 592
use scs8hd_nor2_4  _044_
timestamp 1586364061
transform 1 0 5152 0 1 2720
box -38 -48 866 592
use scs8hd_inv_8  _108_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 5244 0 -1 2720
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__108__A
timestamp 1586364061
transform 1 0 5060 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_0_54
timestamp 1586364061
transform 1 0 6072 0 -1 2720
box -38 -48 406 592
use scs8hd_fill_1  FILLER_1_43
timestamp 1586364061
transform 1 0 5060 0 1 2720
box -38 -48 130 592
use scs8hd_decap_4  FILLER_1_53
timestamp 1586364061
transform 1 0 5980 0 1 2720
box -38 -48 406 592
use scs8hd_fill_1  FILLER_1_60
timestamp 1586364061
transform 1 0 6624 0 1 2720
box -38 -48 130 592
use scs8hd_fill_1  FILLER_1_57
timestamp 1586364061
transform 1 0 6348 0 1 2720
box -38 -48 130 592
use scs8hd_fill_2  FILLER_0_60
timestamp 1586364061
transform 1 0 6624 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__077__A
timestamp 1586364061
transform 1 0 6440 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__077__B
timestamp 1586364061
transform 1 0 6440 0 1 2720
box -38 -48 222 592
use scs8hd_decap_3  FILLER_1_62
timestamp 1586364061
transform 1 0 6808 0 1 2720
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_70
timestamp 1586364061
transform 1 0 6716 0 1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_65
timestamp 1586364061
transform 1 0 6808 0 -1 2720
box -38 -48 130 592
use scs8hd_buf_2  _149_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 7084 0 1 2720
box -38 -48 406 592
use scs8hd_conb_1  _130_
timestamp 1586364061
transform 1 0 6900 0 -1 2720
box -38 -48 314 592
use scs8hd_fill_2  FILLER_1_69
timestamp 1586364061
transform 1 0 7452 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_66
timestamp 1586364061
transform 1 0 7176 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__042__B
timestamp 1586364061
transform 1 0 7360 0 -1 2720
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_right_ipin_4.LATCH_4_.latch tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 8188 0 1 2720
box -38 -48 1050 592
use scs8hd_lpflow_inputisolatch_1  mem_right_ipin_4.LATCH_5_.latch
timestamp 1586364061
transform 1 0 7912 0 -1 2720
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA__149__A
timestamp 1586364061
transform 1 0 7636 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_4.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 7728 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_4.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 8004 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_70
timestamp 1586364061
transform 1 0 7544 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_73
timestamp 1586364061
transform 1 0 7820 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_88
timestamp 1586364061
transform 1 0 9200 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_89
timestamp 1586364061
transform 1 0 9292 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_85
timestamp 1586364061
transform 1 0 8924 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_4.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 9108 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_96
timestamp 1586364061
transform 1 0 9936 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_92
timestamp 1586364061
transform 1 0 9568 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_4.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 9752 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_4.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 9384 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_4.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9476 0 -1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_66
timestamp 1586364061
transform 1 0 9660 0 -1 2720
box -38 -48 130 592
use scs8hd_ebufn_2  mux_right_ipin_4.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 9752 0 -1 2720
box -38 -48 866 592
use scs8hd_or3_4  _115_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 10764 0 1 2720
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__115__C
timestamp 1586364061
transform 1 0 10580 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__115__A
timestamp 1586364061
transform 1 0 10764 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__111__C
timestamp 1586364061
transform 1 0 11224 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_4.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10120 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_103
timestamp 1586364061
transform 1 0 10580 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_3  FILLER_0_107
timestamp 1586364061
transform 1 0 10948 0 -1 2720
box -38 -48 314 592
use scs8hd_decap_3  FILLER_1_100
timestamp 1586364061
transform 1 0 10304 0 1 2720
box -38 -48 314 592
use scs8hd_fill_2  FILLER_1_114
timestamp 1586364061
transform 1 0 11592 0 1 2720
box -38 -48 222 592
use scs8hd_buf_2  _143_
timestamp 1586364061
transform 1 0 11408 0 -1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_1_118
timestamp 1586364061
transform 1 0 11960 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_120
timestamp 1586364061
transform 1 0 12144 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_116
timestamp 1586364061
transform 1 0 11776 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__111__B
timestamp 1586364061
transform 1 0 12144 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__143__A
timestamp 1586364061
transform 1 0 11960 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__111__A
timestamp 1586364061
transform 1 0 11776 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_123
timestamp 1586364061
transform 1 0 12420 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 12328 0 -1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_71
timestamp 1586364061
transform 1 0 12328 0 1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_67
timestamp 1586364061
transform 1 0 12512 0 -1 2720
box -38 -48 130 592
use scs8hd_fill_2  FILLER_1_127
timestamp 1586364061
transform 1 0 12788 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_128
timestamp 1586364061
transform 1 0 12880 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__100__A
timestamp 1586364061
transform 1 0 13064 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__100__B
timestamp 1586364061
transform 1 0 12604 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__100__C
timestamp 1586364061
transform 1 0 12972 0 1 2720
box -38 -48 222 592
use scs8hd_inv_1  mux_right_ipin_0.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 12604 0 -1 2720
box -38 -48 314 592
use scs8hd_fill_2  FILLER_0_132
timestamp 1586364061
transform 1 0 13248 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_1.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 13432 0 -1 2720
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_left_ipin_1.LATCH_1_.latch
timestamp 1586364061
transform 1 0 13616 0 -1 2720
box -38 -48 1050 592
use scs8hd_nor3_4  _099_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 13156 0 1 2720
box -38 -48 1234 592
use scs8hd_diode_2  ANTENNA__099__B
timestamp 1586364061
transform 1 0 14536 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__099__C
timestamp 1586364061
transform 1 0 14904 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_1.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 14812 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_147
timestamp 1586364061
transform 1 0 14628 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_151
timestamp 1586364061
transform 1 0 14996 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_144
timestamp 1586364061
transform 1 0 14352 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_148
timestamp 1586364061
transform 1 0 14720 0 1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_1_152
timestamp 1586364061
transform 1 0 15088 0 1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_1_158
timestamp 1586364061
transform 1 0 15640 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_159
timestamp 1586364061
transform 1 0 15732 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_0.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 15180 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 15456 0 1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_68
timestamp 1586364061
transform 1 0 15364 0 -1 2720
box -38 -48 130 592
use scs8hd_inv_1  mux_right_ipin_0.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 15456 0 -1 2720
box -38 -48 314 592
use scs8hd_fill_2  FILLER_0_163
timestamp 1586364061
transform 1 0 16100 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 15824 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_0.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 16284 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 15916 0 -1 2720
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_ipin_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 16008 0 1 2720
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  mem_right_ipin_0.LATCH_5_.latch
timestamp 1586364061
transform 1 0 16468 0 -1 2720
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 17020 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__109__A
timestamp 1586364061
transform 1 0 17388 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_178
timestamp 1586364061
transform 1 0 17480 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_171
timestamp 1586364061
transform 1 0 16836 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_175
timestamp 1586364061
transform 1 0 17204 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_179
timestamp 1586364061
transform 1 0 17572 0 1 2720
box -38 -48 222 592
use scs8hd_inv_8  _103_
timestamp 1586364061
transform 1 0 18032 0 1 2720
box -38 -48 866 592
use scs8hd_ebufn_2  mux_right_ipin_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18308 0 -1 2720
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_69
timestamp 1586364061
transform 1 0 18216 0 -1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_72
timestamp 1586364061
transform 1 0 17940 0 1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__103__A
timestamp 1586364061
transform 1 0 17756 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 18032 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 17664 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_182
timestamp 1586364061
transform 1 0 17848 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_193
timestamp 1586364061
transform 1 0 18860 0 1 2720
box -38 -48 222 592
use scs8hd_inv_1  mux_right_ipin_0.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 19596 0 1 2720
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 20056 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__084__B
timestamp 1586364061
transform 1 0 19044 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__084__A
timestamp 1586364061
transform 1 0 19412 0 1 2720
box -38 -48 222 592
use scs8hd_decap_12  FILLER_0_196 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 19136 0 -1 2720
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_1_197
timestamp 1586364061
transform 1 0 19228 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_204
timestamp 1586364061
transform 1 0 19872 0 1 2720
box -38 -48 222 592
use scs8hd_decap_3  PHY_1
timestamp 1586364061
transform -1 0 20884 0 -1 2720
box -38 -48 314 592
use scs8hd_decap_3  PHY_3
timestamp 1586364061
transform -1 0 20884 0 1 2720
box -38 -48 314 592
use scs8hd_decap_4  FILLER_0_208
timestamp 1586364061
transform 1 0 20240 0 -1 2720
box -38 -48 406 592
use scs8hd_decap_4  FILLER_1_208
timestamp 1586364061
transform 1 0 20240 0 1 2720
box -38 -48 406 592
use scs8hd_conb_1  _125_
timestamp 1586364061
transform 1 0 1380 0 -1 3808
box -38 -48 314 592
use scs8hd_decap_3  PHY_4
timestamp 1586364061
transform 1 0 1104 0 -1 3808
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__121__A
timestamp 1586364061
transform 1 0 2024 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_2_6
timestamp 1586364061
transform 1 0 1656 0 -1 3808
box -38 -48 406 592
use scs8hd_fill_2  FILLER_2_12
timestamp 1586364061
transform 1 0 2208 0 -1 3808
box -38 -48 222 592
use scs8hd_or3_4  _119_
timestamp 1586364061
transform 1 0 2392 0 -1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__121__C
timestamp 1586364061
transform 1 0 3404 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_23
timestamp 1586364061
transform 1 0 3220 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_27
timestamp 1586364061
transform 1 0 3588 0 -1 3808
box -38 -48 222 592
use scs8hd_inv_8  _101_
timestamp 1586364061
transform 1 0 4876 0 -1 3808
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_73
timestamp 1586364061
transform 1 0 3956 0 -1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__042__A
timestamp 1586364061
transform 1 0 3772 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__073__A
timestamp 1586364061
transform 1 0 4232 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__046__A
timestamp 1586364061
transform 1 0 4692 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_32
timestamp 1586364061
transform 1 0 4048 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_3  FILLER_2_36
timestamp 1586364061
transform 1 0 4416 0 -1 3808
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__044__A
timestamp 1586364061
transform 1 0 5888 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_50
timestamp 1586364061
transform 1 0 5704 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_54
timestamp 1586364061
transform 1 0 6072 0 -1 3808
box -38 -48 222 592
use scs8hd_nor2_4  _077_
timestamp 1586364061
transform 1 0 6440 0 -1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__076__A
timestamp 1586364061
transform 1 0 6256 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__046__B
timestamp 1586364061
transform 1 0 7452 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_67
timestamp 1586364061
transform 1 0 7268 0 -1 3808
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_ipin_4.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 8004 0 -1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_4.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 7820 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_71
timestamp 1586364061
transform 1 0 7636 0 -1 3808
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_ipin_4.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9660 0 -1 3808
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_74
timestamp 1586364061
transform 1 0 9568 0 -1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_4.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 9016 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_4.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 9384 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_84
timestamp 1586364061
transform 1 0 8832 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_88
timestamp 1586364061
transform 1 0 9200 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__115__B
timestamp 1586364061
transform 1 0 10764 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_4.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11132 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_3  FILLER_2_102
timestamp 1586364061
transform 1 0 10488 0 -1 3808
box -38 -48 314 592
use scs8hd_fill_2  FILLER_2_107
timestamp 1586364061
transform 1 0 10948 0 -1 3808
box -38 -48 222 592
use scs8hd_or3_4  _111_
timestamp 1586364061
transform 1 0 11408 0 -1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__063__B
timestamp 1586364061
transform 1 0 12512 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_1  FILLER_2_111
timestamp 1586364061
transform 1 0 11316 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_3  FILLER_2_121
timestamp 1586364061
transform 1 0 12236 0 -1 3808
box -38 -48 314 592
use scs8hd_nor3_4  _100_
timestamp 1586364061
transform 1 0 13248 0 -1 3808
box -38 -48 1234 592
use scs8hd_diode_2  ANTENNA__099__A
timestamp 1586364061
transform 1 0 13064 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_2_126
timestamp 1586364061
transform 1 0 12696 0 -1 3808
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_1.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 14628 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14996 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_145
timestamp 1586364061
transform 1 0 14444 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_149
timestamp 1586364061
transform 1 0 14812 0 -1 3808
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_ipin_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15640 0 -1 3808
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_75
timestamp 1586364061
transform 1 0 15180 0 -1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 15456 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_154
timestamp 1586364061
transform 1 0 15272 0 -1 3808
box -38 -48 222 592
use scs8hd_inv_8  _109_
timestamp 1586364061
transform 1 0 17204 0 -1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 16652 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_167
timestamp 1586364061
transform 1 0 16468 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_2_171
timestamp 1586364061
transform 1 0 16836 0 -1 3808
box -38 -48 406 592
use scs8hd_nor2_4  _084_
timestamp 1586364061
transform 1 0 18768 0 -1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_0.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 18216 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 18584 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_184
timestamp 1586364061
transform 1 0 18032 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_188
timestamp 1586364061
transform 1 0 18400 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_8  FILLER_2_201 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 19596 0 -1 3808
box -38 -48 774 592
use scs8hd_decap_3  PHY_5
timestamp 1586364061
transform -1 0 20884 0 -1 3808
box -38 -48 314 592
use scs8hd_decap_3  FILLER_2_209
timestamp 1586364061
transform 1 0 20332 0 -1 3808
box -38 -48 314 592
use scs8hd_or3_4  _121_
timestamp 1586364061
transform 1 0 2024 0 1 3808
box -38 -48 866 592
use scs8hd_decap_3  PHY_6
timestamp 1586364061
transform 1 0 1104 0 1 3808
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__123__A
timestamp 1586364061
transform 1 0 1840 0 1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_3_3
timestamp 1586364061
transform 1 0 1380 0 1 3808
box -38 -48 406 592
use scs8hd_fill_1  FILLER_3_7
timestamp 1586364061
transform 1 0 1748 0 1 3808
box -38 -48 130 592
use scs8hd_nor2_4  _043_
timestamp 1586364061
transform 1 0 3588 0 1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__123__C
timestamp 1586364061
transform 1 0 3036 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__123__B
timestamp 1586364061
transform 1 0 3404 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_19
timestamp 1586364061
transform 1 0 2852 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_23
timestamp 1586364061
transform 1 0 3220 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__074__A
timestamp 1586364061
transform 1 0 4600 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_36
timestamp 1586364061
transform 1 0 4416 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_40
timestamp 1586364061
transform 1 0 4784 0 1 3808
box -38 -48 222 592
use scs8hd_nor2_4  _074_
timestamp 1586364061
transform 1 0 5152 0 1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__076__B
timestamp 1586364061
transform 1 0 6164 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__074__B
timestamp 1586364061
transform 1 0 4968 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_53
timestamp 1586364061
transform 1 0 5980 0 1 3808
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_right_ipin_4.LATCH_0_.latch
timestamp 1586364061
transform 1 0 7084 0 1 3808
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_76
timestamp 1586364061
transform 1 0 6716 0 1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_4.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 6532 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_57
timestamp 1586364061
transform 1 0 6348 0 1 3808
box -38 -48 222 592
use scs8hd_decap_3  FILLER_3_62
timestamp 1586364061
transform 1 0 6808 0 1 3808
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__043__B
timestamp 1586364061
transform 1 0 8280 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_4.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 8648 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_76
timestamp 1586364061
transform 1 0 8096 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_80
timestamp 1586364061
transform 1 0 8464 0 1 3808
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_right_ipin_4.LATCH_3_.latch
timestamp 1586364061
transform 1 0 9568 0 1 3808
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_4.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 9384 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_4.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 9016 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_84
timestamp 1586364061
transform 1 0 8832 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_88
timestamp 1586364061
transform 1 0 9200 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__040__B
timestamp 1586364061
transform 1 0 11132 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_4.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 10764 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_103
timestamp 1586364061
transform 1 0 10580 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_107
timestamp 1586364061
transform 1 0 10948 0 1 3808
box -38 -48 222 592
use scs8hd_or2_4  _063_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 12512 0 1 3808
box -38 -48 682 592
use scs8hd_inv_1  mux_right_ipin_7.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 11316 0 1 3808
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_77
timestamp 1586364061
transform 1 0 12328 0 1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__040__A
timestamp 1586364061
transform 1 0 11960 0 1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_3_114
timestamp 1586364061
transform 1 0 11592 0 1 3808
box -38 -48 406 592
use scs8hd_fill_2  FILLER_3_120
timestamp 1586364061
transform 1 0 12144 0 1 3808
box -38 -48 222 592
use scs8hd_fill_1  FILLER_3_123
timestamp 1586364061
transform 1 0 12420 0 1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__063__A
timestamp 1586364061
transform 1 0 13340 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_1.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 13708 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_131
timestamp 1586364061
transform 1 0 13156 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_135
timestamp 1586364061
transform 1 0 13524 0 1 3808
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_left_ipin_1.LATCH_0_.latch
timestamp 1586364061
transform 1 0 13892 0 1 3808
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 15088 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_150
timestamp 1586364061
transform 1 0 14904 0 1 3808
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_ipin_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15640 0 1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 15456 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_154
timestamp 1586364061
transform 1 0 15272 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_0.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 16836 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_0.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 17204 0 1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_3_167
timestamp 1586364061
transform 1 0 16468 0 1 3808
box -38 -48 406 592
use scs8hd_fill_2  FILLER_3_173
timestamp 1586364061
transform 1 0 17020 0 1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_3_177
timestamp 1586364061
transform 1 0 17388 0 1 3808
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_right_ipin_0.LATCH_4_.latch
timestamp 1586364061
transform 1 0 18032 0 1 3808
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_78
timestamp 1586364061
transform 1 0 17940 0 1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_0.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 17756 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 19228 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_195
timestamp 1586364061
transform 1 0 19044 0 1 3808
box -38 -48 222 592
use scs8hd_decap_12  FILLER_3_199
timestamp 1586364061
transform 1 0 19412 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_3  PHY_7
timestamp 1586364061
transform -1 0 20884 0 1 3808
box -38 -48 314 592
use scs8hd_fill_1  FILLER_3_211
timestamp 1586364061
transform 1 0 20516 0 1 3808
box -38 -48 130 592
use scs8hd_inv_1  mux_left_ipin_1.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1380 0 -1 4896
box -38 -48 314 592
use scs8hd_decap_3  PHY_8
timestamp 1586364061
transform 1 0 1104 0 -1 4896
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__121__B
timestamp 1586364061
transform 1 0 2024 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_4_6
timestamp 1586364061
transform 1 0 1656 0 -1 4896
box -38 -48 406 592
use scs8hd_fill_2  FILLER_4_12
timestamp 1586364061
transform 1 0 2208 0 -1 4896
box -38 -48 222 592
use scs8hd_or3_4  _123_
timestamp 1586364061
transform 1 0 2392 0 -1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__071__A
timestamp 1586364061
transform 1 0 3404 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_23
timestamp 1586364061
transform 1 0 3220 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_27
timestamp 1586364061
transform 1 0 3588 0 -1 4896
box -38 -48 222 592
use scs8hd_nor2_4  _046_
timestamp 1586364061
transform 1 0 4876 0 -1 4896
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_79
timestamp 1586364061
transform 1 0 3956 0 -1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__048__A
timestamp 1586364061
transform 1 0 4324 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__048__B
timestamp 1586364061
transform 1 0 4692 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__043__A
timestamp 1586364061
transform 1 0 3772 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_3  FILLER_4_32
timestamp 1586364061
transform 1 0 4048 0 -1 4896
box -38 -48 314 592
use scs8hd_fill_2  FILLER_4_37
timestamp 1586364061
transform 1 0 4508 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__092__B
timestamp 1586364061
transform 1 0 5888 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_50
timestamp 1586364061
transform 1 0 5704 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_54
timestamp 1586364061
transform 1 0 6072 0 -1 4896
box -38 -48 222 592
use scs8hd_nor2_4  _076_
timestamp 1586364061
transform 1 0 6440 0 -1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_4.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 7452 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__092__C
timestamp 1586364061
transform 1 0 6256 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_67
timestamp 1586364061
transform 1 0 7268 0 -1 4896
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_ipin_4.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 8004 0 -1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_4.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 7820 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_71
timestamp 1586364061
transform 1 0 7636 0 -1 4896
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_ipin_4.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9660 0 -1 4896
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_80
timestamp 1586364061
transform 1 0 9568 0 -1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_4.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 9108 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_3  FILLER_4_84
timestamp 1586364061
transform 1 0 8832 0 -1 4896
box -38 -48 314 592
use scs8hd_decap_3  FILLER_4_89
timestamp 1586364061
transform 1 0 9292 0 -1 4896
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__117__A
timestamp 1586364061
transform 1 0 10764 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_3  FILLER_4_102
timestamp 1586364061
transform 1 0 10488 0 -1 4896
box -38 -48 314 592
use scs8hd_decap_4  FILLER_4_107
timestamp 1586364061
transform 1 0 10948 0 -1 4896
box -38 -48 406 592
use scs8hd_or3_4  _040_
timestamp 1586364061
transform 1 0 11960 0 -1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_7.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 11316 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__040__C
timestamp 1586364061
transform 1 0 11776 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_3  FILLER_4_113
timestamp 1586364061
transform 1 0 11500 0 -1 4896
box -38 -48 314 592
use scs8hd_inv_8  _110_
timestamp 1586364061
transform 1 0 13616 0 -1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__110__A
timestamp 1586364061
transform 1 0 13432 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_4.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 12972 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_127
timestamp 1586364061
transform 1 0 12788 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_3  FILLER_4_131
timestamp 1586364061
transform 1 0 13156 0 -1 4896
box -38 -48 314 592
use scs8hd_decap_8  FILLER_4_145
timestamp 1586364061
transform 1 0 14444 0 -1 4896
box -38 -48 774 592
use scs8hd_ebufn_2  mux_left_ipin_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15272 0 -1 4896
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_81
timestamp 1586364061
transform 1 0 15180 0 -1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_0.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 16284 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_163
timestamp 1586364061
transform 1 0 16100 0 -1 4896
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_right_ipin_0.LATCH_3_.latch
timestamp 1586364061
transform 1 0 16836 0 -1 4896
box -38 -48 1050 592
use scs8hd_decap_4  FILLER_4_167
timestamp 1586364061
transform 1 0 16468 0 -1 4896
box -38 -48 406 592
use scs8hd_ebufn_2  mux_right_ipin_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18584 0 -1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 18032 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 18400 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_182
timestamp 1586364061
transform 1 0 17848 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_186
timestamp 1586364061
transform 1 0 18216 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__085__C
timestamp 1586364061
transform 1 0 19596 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_199
timestamp 1586364061
transform 1 0 19412 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_8  FILLER_4_203
timestamp 1586364061
transform 1 0 19780 0 -1 4896
box -38 -48 774 592
use scs8hd_decap_3  PHY_9
timestamp 1586364061
transform -1 0 20884 0 -1 4896
box -38 -48 314 592
use scs8hd_fill_1  FILLER_4_211
timestamp 1586364061
transform 1 0 20516 0 -1 4896
box -38 -48 130 592
use scs8hd_inv_1  mux_right_ipin_4.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1564 0 1 4896
box -38 -48 314 592
use scs8hd_decap_3  PHY_10
timestamp 1586364061
transform 1 0 1104 0 1 4896
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_4.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 2024 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_3
timestamp 1586364061
transform 1 0 1380 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_8
timestamp 1586364061
transform 1 0 1840 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_12
timestamp 1586364061
transform 1 0 2208 0 1 4896
box -38 -48 222 592
use scs8hd_or3_4  _041_
timestamp 1586364061
transform 1 0 3588 0 1 4896
box -38 -48 866 592
use scs8hd_inv_1  mux_left_ipin_1.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 2576 0 1 4896
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__071__B
timestamp 1586364061
transform 1 0 2392 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__041__B
timestamp 1586364061
transform 1 0 3404 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_1.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 3036 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_19
timestamp 1586364061
transform 1 0 2852 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_23
timestamp 1586364061
transform 1 0 3220 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__055__A
timestamp 1586364061
transform 1 0 4600 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_36
timestamp 1586364061
transform 1 0 4416 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_40
timestamp 1586364061
transform 1 0 4784 0 1 4896
box -38 -48 222 592
use scs8hd_or3_4  _055_
timestamp 1586364061
transform 1 0 5152 0 1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__092__A
timestamp 1586364061
transform 1 0 6164 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__055__B
timestamp 1586364061
transform 1 0 4968 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_53
timestamp 1586364061
transform 1 0 5980 0 1 4896
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_right_ipin_4.LATCH_1_.latch
timestamp 1586364061
transform 1 0 7360 0 1 4896
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_82
timestamp 1586364061
transform 1 0 6716 0 1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_4.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 7176 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__092__D
timestamp 1586364061
transform 1 0 6532 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_57
timestamp 1586364061
transform 1 0 6348 0 1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_5_62
timestamp 1586364061
transform 1 0 6808 0 1 4896
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_4.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 8556 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_79
timestamp 1586364061
transform 1 0 8372 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_83
timestamp 1586364061
transform 1 0 8740 0 1 4896
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_ipin_4.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9108 0 1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_4.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 8924 0 1 4896
box -38 -48 222 592
use scs8hd_decap_3  FILLER_5_96
timestamp 1586364061
transform 1 0 9936 0 1 4896
box -38 -48 314 592
use scs8hd_or3_4  _117_
timestamp 1586364061
transform 1 0 10764 0 1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__117__B
timestamp 1586364061
transform 1 0 10580 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__117__C
timestamp 1586364061
transform 1 0 10212 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_101
timestamp 1586364061
transform 1 0 10396 0 1 4896
box -38 -48 222 592
use scs8hd_or3_4  _112_
timestamp 1586364061
transform 1 0 12420 0 1 4896
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_83
timestamp 1586364061
transform 1 0 12328 0 1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__112__B
timestamp 1586364061
transform 1 0 12144 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__105__A
timestamp 1586364061
transform 1 0 11776 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_114
timestamp 1586364061
transform 1 0 11592 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_118
timestamp 1586364061
transform 1 0 11960 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__102__A
timestamp 1586364061
transform 1 0 13800 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__106__A
timestamp 1586364061
transform 1 0 13432 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_132
timestamp 1586364061
transform 1 0 13248 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_136
timestamp 1586364061
transform 1 0 13616 0 1 4896
box -38 -48 222 592
use scs8hd_inv_8  _102_
timestamp 1586364061
transform 1 0 13984 0 1 4896
box -38 -48 866 592
use scs8hd_decap_4  FILLER_5_149
timestamp 1586364061
transform 1 0 14812 0 1 4896
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_right_ipin_0.LATCH_1_.latch
timestamp 1586364061
transform 1 0 15732 0 1 4896
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_0.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 15548 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 15180 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_155
timestamp 1586364061
transform 1 0 15364 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 17480 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 16928 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_170
timestamp 1586364061
transform 1 0 16744 0 1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_5_174
timestamp 1586364061
transform 1 0 17112 0 1 4896
box -38 -48 406 592
use scs8hd_ebufn_2  mux_right_ipin_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18032 0 1 4896
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_84
timestamp 1586364061
transform 1 0 17940 0 1 4896
box -38 -48 130 592
use scs8hd_decap_3  FILLER_5_180
timestamp 1586364061
transform 1 0 17664 0 1 4896
box -38 -48 314 592
use scs8hd_fill_2  FILLER_5_193
timestamp 1586364061
transform 1 0 18860 0 1 4896
box -38 -48 222 592
use scs8hd_inv_1  mux_right_ipin_5.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 19596 0 1 4896
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__085__A
timestamp 1586364061
transform 1 0 19044 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_5.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 20056 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__085__B
timestamp 1586364061
transform 1 0 19412 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_197
timestamp 1586364061
transform 1 0 19228 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_204
timestamp 1586364061
transform 1 0 19872 0 1 4896
box -38 -48 222 592
use scs8hd_decap_3  PHY_11
timestamp 1586364061
transform -1 0 20884 0 1 4896
box -38 -48 314 592
use scs8hd_decap_4  FILLER_5_208
timestamp 1586364061
transform 1 0 20240 0 1 4896
box -38 -48 406 592
use scs8hd_decap_4  FILLER_7_3
timestamp 1586364061
transform 1 0 1380 0 1 5984
box -38 -48 406 592
use scs8hd_fill_2  FILLER_6_6
timestamp 1586364061
transform 1 0 1656 0 -1 5984
box -38 -48 222 592
use scs8hd_decap_3  PHY_14
timestamp 1586364061
transform 1 0 1104 0 1 5984
box -38 -48 314 592
use scs8hd_decap_3  PHY_12
timestamp 1586364061
transform 1 0 1104 0 -1 5984
box -38 -48 314 592
use scs8hd_inv_1  mux_right_ipin_2.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1380 0 -1 5984
box -38 -48 314 592
use scs8hd_fill_1  FILLER_7_7
timestamp 1586364061
transform 1 0 1748 0 1 5984
box -38 -48 130 592
use scs8hd_fill_2  FILLER_6_10
timestamp 1586364061
transform 1 0 2024 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__071__C
timestamp 1586364061
transform 1 0 2208 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_2.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 1840 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__062__B
timestamp 1586364061
transform 1 0 1840 0 1 5984
box -38 -48 222 592
use scs8hd_or3_4  _062_
timestamp 1586364061
transform 1 0 2024 0 1 5984
box -38 -48 866 592
use scs8hd_nor2_4  _047_
timestamp 1586364061
transform 1 0 3588 0 1 5984
box -38 -48 866 592
use scs8hd_or3_4  _071_
timestamp 1586364061
transform 1 0 2392 0 -1 5984
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__062__A
timestamp 1586364061
transform 1 0 3036 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__041__A
timestamp 1586364061
transform 1 0 3588 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__062__C
timestamp 1586364061
transform 1 0 3404 0 1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_6_23
timestamp 1586364061
transform 1 0 3220 0 -1 5984
box -38 -48 406 592
use scs8hd_fill_2  FILLER_7_19
timestamp 1586364061
transform 1 0 2852 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_23
timestamp 1586364061
transform 1 0 3220 0 1 5984
box -38 -48 222 592
use scs8hd_or3_4  _048_
timestamp 1586364061
transform 1 0 4324 0 -1 5984
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_85
timestamp 1586364061
transform 1 0 3956 0 -1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__097__B
timestamp 1586364061
transform 1 0 4600 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_29
timestamp 1586364061
transform 1 0 3772 0 -1 5984
box -38 -48 222 592
use scs8hd_decap_3  FILLER_6_32
timestamp 1586364061
transform 1 0 4048 0 -1 5984
box -38 -48 314 592
use scs8hd_fill_2  FILLER_7_36
timestamp 1586364061
transform 1 0 4416 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_40
timestamp 1586364061
transform 1 0 4784 0 1 5984
box -38 -48 222 592
use scs8hd_or4_4  _092_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 5888 0 -1 5984
box -38 -48 866 592
use scs8hd_inv_8  _104_
timestamp 1586364061
transform 1 0 5152 0 1 5984
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__104__A
timestamp 1586364061
transform 1 0 4968 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__055__C
timestamp 1586364061
transform 1 0 5336 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__075__A
timestamp 1586364061
transform 1 0 6164 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__097__A
timestamp 1586364061
transform 1 0 5704 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_44
timestamp 1586364061
transform 1 0 5152 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_48
timestamp 1586364061
transform 1 0 5520 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_53
timestamp 1586364061
transform 1 0 5980 0 1 5984
box -38 -48 222 592
use scs8hd_nor2_4  _075_
timestamp 1586364061
transform 1 0 6808 0 1 5984
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  mem_right_ipin_4.LATCH_2_.latch
timestamp 1586364061
transform 1 0 7452 0 -1 5984
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_88
timestamp 1586364061
transform 1 0 6716 0 1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_2.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 6532 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__075__B
timestamp 1586364061
transform 1 0 6900 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_2.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 7268 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_61
timestamp 1586364061
transform 1 0 6716 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_65
timestamp 1586364061
transform 1 0 7084 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_57
timestamp 1586364061
transform 1 0 6348 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_7.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 8556 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_4.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 8004 0 1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_6_80
timestamp 1586364061
transform 1 0 8464 0 -1 5984
box -38 -48 406 592
use scs8hd_decap_4  FILLER_7_71
timestamp 1586364061
transform 1 0 7636 0 1 5984
box -38 -48 406 592
use scs8hd_decap_4  FILLER_7_77
timestamp 1586364061
transform 1 0 8188 0 1 5984
box -38 -48 406 592
use scs8hd_fill_1  FILLER_7_83
timestamp 1586364061
transform 1 0 8740 0 1 5984
box -38 -48 130 592
use scs8hd_ebufn_2  mux_right_ipin_4.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9660 0 -1 5984
box -38 -48 866 592
use scs8hd_ebufn_2  mux_right_ipin_4.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 8832 0 1 5984
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_86
timestamp 1586364061
transform 1 0 9568 0 -1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__113__A
timestamp 1586364061
transform 1 0 9936 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_4.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 8832 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_4.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9200 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_86
timestamp 1586364061
transform 1 0 9016 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_90
timestamp 1586364061
transform 1 0 9384 0 -1 5984
box -38 -48 222 592
use scs8hd_decap_3  FILLER_7_93
timestamp 1586364061
transform 1 0 9660 0 1 5984
box -38 -48 314 592
use scs8hd_ebufn_2  mux_right_ipin_4.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10396 0 1 5984
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__113__B
timestamp 1586364061
transform 1 0 10672 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_4.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11040 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_102
timestamp 1586364061
transform 1 0 10488 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_106
timestamp 1586364061
transform 1 0 10856 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_1  FILLER_6_110
timestamp 1586364061
transform 1 0 11224 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_3  FILLER_7_98
timestamp 1586364061
transform 1 0 10120 0 1 5984
box -38 -48 314 592
use scs8hd_fill_2  FILLER_7_110
timestamp 1586364061
transform 1 0 11224 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_114
timestamp 1586364061
transform 1 0 11592 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_7.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 11776 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__113__C
timestamp 1586364061
transform 1 0 11408 0 1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_7_123
timestamp 1586364061
transform 1 0 12420 0 1 5984
box -38 -48 406 592
use scs8hd_fill_2  FILLER_7_118
timestamp 1586364061
transform 1 0 11960 0 1 5984
box -38 -48 222 592
use scs8hd_decap_3  FILLER_6_120
timestamp 1586364061
transform 1 0 12144 0 -1 5984
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_7.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 12144 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__112__A
timestamp 1586364061
transform 1 0 12420 0 -1 5984
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_89
timestamp 1586364061
transform 1 0 12328 0 1 5984
box -38 -48 130 592
use scs8hd_inv_8  _105_
timestamp 1586364061
transform 1 0 11316 0 -1 5984
box -38 -48 866 592
use scs8hd_inv_8  _106_
timestamp 1586364061
transform 1 0 13156 0 -1 5984
box -38 -48 866 592
use scs8hd_inv_8  _107_
timestamp 1586364061
transform 1 0 13340 0 1 5984
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__107__A
timestamp 1586364061
transform 1 0 13156 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__078__A
timestamp 1586364061
transform 1 0 12788 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__112__C
timestamp 1586364061
transform 1 0 12788 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_125
timestamp 1586364061
transform 1 0 12604 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_129
timestamp 1586364061
transform 1 0 12972 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_129
timestamp 1586364061
transform 1 0 12972 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__078__C
timestamp 1586364061
transform 1 0 14352 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__078__B
timestamp 1586364061
transform 1 0 14168 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_0.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 14996 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_140
timestamp 1586364061
transform 1 0 13984 0 -1 5984
box -38 -48 222 592
use scs8hd_decap_8  FILLER_6_144
timestamp 1586364061
transform 1 0 14352 0 -1 5984
box -38 -48 774 592
use scs8hd_fill_1  FILLER_6_152
timestamp 1586364061
transform 1 0 15088 0 -1 5984
box -38 -48 130 592
use scs8hd_fill_2  FILLER_7_142
timestamp 1586364061
transform 1 0 14168 0 1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_7_146
timestamp 1586364061
transform 1 0 14536 0 1 5984
box -38 -48 406 592
use scs8hd_fill_1  FILLER_7_150
timestamp 1586364061
transform 1 0 14904 0 1 5984
box -38 -48 130 592
use scs8hd_nor2_4  _081_
timestamp 1586364061
transform 1 0 15548 0 1 5984
box -38 -48 866 592
use scs8hd_ebufn_2  mux_right_ipin_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15916 0 -1 5984
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_87
timestamp 1586364061
transform 1 0 15180 0 -1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__081__B
timestamp 1586364061
transform 1 0 15364 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__081__A
timestamp 1586364061
transform 1 0 15548 0 -1 5984
box -38 -48 222 592
use scs8hd_decap_3  FILLER_6_154
timestamp 1586364061
transform 1 0 15272 0 -1 5984
box -38 -48 314 592
use scs8hd_fill_2  FILLER_6_159
timestamp 1586364061
transform 1 0 15732 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_153
timestamp 1586364061
transform 1 0 15180 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_166
timestamp 1586364061
transform 1 0 16376 0 1 5984
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_ipin_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 17480 0 -1 5984
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_0.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 17572 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_0.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 16560 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 17204 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 17296 0 -1 5984
box -38 -48 222 592
use scs8hd_decap_6  FILLER_6_170 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 16744 0 -1 5984
box -38 -48 590 592
use scs8hd_decap_4  FILLER_7_170
timestamp 1586364061
transform 1 0 16744 0 1 5984
box -38 -48 406 592
use scs8hd_fill_1  FILLER_7_174
timestamp 1586364061
transform 1 0 17112 0 1 5984
box -38 -48 130 592
use scs8hd_fill_2  FILLER_7_177
timestamp 1586364061
transform 1 0 17388 0 1 5984
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_ipin_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18032 0 1 5984
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_90
timestamp 1586364061
transform 1 0 17940 0 1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 18492 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_187
timestamp 1586364061
transform 1 0 18308 0 -1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_6_191
timestamp 1586364061
transform 1 0 18676 0 -1 5984
box -38 -48 406 592
use scs8hd_fill_2  FILLER_7_181
timestamp 1586364061
transform 1 0 17756 0 1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_7_193
timestamp 1586364061
transform 1 0 18860 0 1 5984
box -38 -48 406 592
use scs8hd_or3_4  _085_
timestamp 1586364061
transform 1 0 19044 0 -1 5984
box -38 -48 866 592
use scs8hd_inv_1  mux_right_ipin_5.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 19596 0 1 5984
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__140__A
timestamp 1586364061
transform 1 0 19320 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_5.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 20056 0 1 5984
box -38 -48 222 592
use scs8hd_decap_8  FILLER_6_204
timestamp 1586364061
transform 1 0 19872 0 -1 5984
box -38 -48 774 592
use scs8hd_fill_1  FILLER_7_197
timestamp 1586364061
transform 1 0 19228 0 1 5984
box -38 -48 130 592
use scs8hd_fill_1  FILLER_7_200
timestamp 1586364061
transform 1 0 19504 0 1 5984
box -38 -48 130 592
use scs8hd_fill_2  FILLER_7_204
timestamp 1586364061
transform 1 0 19872 0 1 5984
box -38 -48 222 592
use scs8hd_decap_3  PHY_13
timestamp 1586364061
transform -1 0 20884 0 -1 5984
box -38 -48 314 592
use scs8hd_decap_3  PHY_15
timestamp 1586364061
transform -1 0 20884 0 1 5984
box -38 -48 314 592
use scs8hd_decap_4  FILLER_7_208
timestamp 1586364061
transform 1 0 20240 0 1 5984
box -38 -48 406 592
use scs8hd_inv_1  mux_right_ipin_4.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1380 0 -1 7072
box -38 -48 314 592
use scs8hd_decap_3  PHY_16
timestamp 1586364061
transform 1 0 1104 0 -1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_4.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 1840 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__061__B
timestamp 1586364061
transform 1 0 2208 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_6
timestamp 1586364061
transform 1 0 1656 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_10
timestamp 1586364061
transform 1 0 2024 0 -1 7072
box -38 -48 222 592
use scs8hd_nor2_4  _045_
timestamp 1586364061
transform 1 0 2392 0 -1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__057__A
timestamp 1586364061
transform 1 0 3588 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_8_23
timestamp 1586364061
transform 1 0 3220 0 -1 7072
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_91
timestamp 1586364061
transform 1 0 3956 0 -1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__047__A
timestamp 1586364061
transform 1 0 4232 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__048__C
timestamp 1586364061
transform 1 0 4600 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_29
timestamp 1586364061
transform 1 0 3772 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_32
timestamp 1586364061
transform 1 0 4048 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_36
timestamp 1586364061
transform 1 0 4416 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_40
timestamp 1586364061
transform 1 0 4784 0 -1 7072
box -38 -48 222 592
use scs8hd_nor2_4  _097_
timestamp 1586364061
transform 1 0 4968 0 -1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_4.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 5980 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_51
timestamp 1586364061
transform 1 0 5796 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_8_55
timestamp 1586364061
transform 1 0 6164 0 -1 7072
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_right_ipin_2.LATCH_0_.latch
timestamp 1586364061
transform 1 0 6532 0 -1 7072
box -38 -48 1050 592
use scs8hd_inv_1  mux_right_ipin_7.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 8556 0 -1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 7820 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_3  FILLER_8_70
timestamp 1586364061
transform 1 0 7544 0 -1 7072
box -38 -48 314 592
use scs8hd_decap_6  FILLER_8_75
timestamp 1586364061
transform 1 0 8004 0 -1 7072
box -38 -48 590 592
use scs8hd_or3_4  _113_
timestamp 1586364061
transform 1 0 9936 0 -1 7072
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_92
timestamp 1586364061
transform 1 0 9568 0 -1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_4.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9384 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_4.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9016 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_84
timestamp 1586364061
transform 1 0 8832 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_88
timestamp 1586364061
transform 1 0 9200 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_3  FILLER_8_93
timestamp 1586364061
transform 1 0 9660 0 -1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_4.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10948 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_105
timestamp 1586364061
transform 1 0 10764 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_8_109
timestamp 1586364061
transform 1 0 11132 0 -1 7072
box -38 -48 406 592
use scs8hd_ebufn_2  mux_right_ipin_7.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 11500 0 -1 7072
box -38 -48 866 592
use scs8hd_decap_8  FILLER_8_122
timestamp 1586364061
transform 1 0 12328 0 -1 7072
box -38 -48 774 592
use scs8hd_or3_4  _078_
timestamp 1586364061
transform 1 0 13616 0 -1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_7.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 13248 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_130
timestamp 1586364061
transform 1 0 13064 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_134
timestamp 1586364061
transform 1 0 13432 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_8  FILLER_8_145
timestamp 1586364061
transform 1 0 14444 0 -1 7072
box -38 -48 774 592
use scs8hd_lpflow_inputisolatch_1  mem_right_ipin_0.LATCH_0_.latch
timestamp 1586364061
transform 1 0 15824 0 -1 7072
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_93
timestamp 1586364061
transform 1 0 15180 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_6  FILLER_8_154
timestamp 1586364061
transform 1 0 15272 0 -1 7072
box -38 -48 590 592
use scs8hd_lpflow_inputisolatch_1  mem_right_ipin_0.LATCH_2_.latch
timestamp 1586364061
transform 1 0 17572 0 -1 7072
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_0.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 17388 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 17020 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_171
timestamp 1586364061
transform 1 0 16836 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_175
timestamp 1586364061
transform 1 0 17204 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_8  FILLER_8_190
timestamp 1586364061
transform 1 0 18584 0 -1 7072
box -38 -48 774 592
use scs8hd_buf_2  _140_
timestamp 1586364061
transform 1 0 19320 0 -1 7072
box -38 -48 406 592
use scs8hd_decap_8  FILLER_8_202
timestamp 1586364061
transform 1 0 19688 0 -1 7072
box -38 -48 774 592
use scs8hd_decap_3  PHY_17
timestamp 1586364061
transform -1 0 20884 0 -1 7072
box -38 -48 314 592
use scs8hd_fill_2  FILLER_8_210
timestamp 1586364061
transform 1 0 20424 0 -1 7072
box -38 -48 222 592
use scs8hd_nor2_4  _061_
timestamp 1586364061
transform 1 0 2024 0 1 7072
box -38 -48 866 592
use scs8hd_decap_3  PHY_18
timestamp 1586364061
transform 1 0 1104 0 1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_2.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 1840 0 1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_9_3
timestamp 1586364061
transform 1 0 1380 0 1 7072
box -38 -48 406 592
use scs8hd_fill_1  FILLER_9_7
timestamp 1586364061
transform 1 0 1748 0 1 7072
box -38 -48 130 592
use scs8hd_nor2_4  _057_
timestamp 1586364061
transform 1 0 3588 0 1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 3036 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__057__B
timestamp 1586364061
transform 1 0 3404 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_19
timestamp 1586364061
transform 1 0 2852 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_23
timestamp 1586364061
transform 1 0 3220 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__095__A
timestamp 1586364061
transform 1 0 4600 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_36
timestamp 1586364061
transform 1 0 4416 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_40
timestamp 1586364061
transform 1 0 4784 0 1 7072
box -38 -48 222 592
use scs8hd_nor2_4  _095_
timestamp 1586364061
transform 1 0 5152 0 1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_2.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 6164 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__095__B
timestamp 1586364061
transform 1 0 4968 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_53
timestamp 1586364061
transform 1 0 5980 0 1 7072
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_right_ipin_2.LATCH_4_.latch
timestamp 1586364061
transform 1 0 6900 0 1 7072
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_94
timestamp 1586364061
transform 1 0 6716 0 1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_7.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 6532 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_57
timestamp 1586364061
transform 1 0 6348 0 1 7072
box -38 -48 222 592
use scs8hd_fill_1  FILLER_9_62
timestamp 1586364061
transform 1 0 6808 0 1 7072
box -38 -48 130 592
use scs8hd_ebufn_2  mux_right_ipin_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 8648 0 1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 8096 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 8464 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_74
timestamp 1586364061
transform 1 0 7912 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_78
timestamp 1586364061
transform 1 0 8280 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_2.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9660 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_91
timestamp 1586364061
transform 1 0 9476 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_95
timestamp 1586364061
transform 1 0 9844 0 1 7072
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_ipin_2.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10212 0 1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_7.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 11224 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_2.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10028 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_108
timestamp 1586364061
transform 1 0 11040 0 1 7072
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_95
timestamp 1586364061
transform 1 0 12328 0 1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_7.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 11592 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_112
timestamp 1586364061
transform 1 0 11408 0 1 7072
box -38 -48 222 592
use scs8hd_decap_6  FILLER_9_116
timestamp 1586364061
transform 1 0 11776 0 1 7072
box -38 -48 590 592
use scs8hd_fill_2  FILLER_9_123
timestamp 1586364061
transform 1 0 12420 0 1 7072
box -38 -48 222 592
use scs8hd_buf_2  _142_
timestamp 1586364061
transform 1 0 12604 0 1 7072
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_right_ipin_7.LATCH_5_.latch
timestamp 1586364061
transform 1 0 13708 0 1 7072
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA__142__A
timestamp 1586364061
transform 1 0 13156 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_7.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 13524 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_129
timestamp 1586364061
transform 1 0 12972 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_133
timestamp 1586364061
transform 1 0 13340 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_7.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 14904 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_148
timestamp 1586364061
transform 1 0 14720 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_152
timestamp 1586364061
transform 1 0 15088 0 1 7072
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_ipin_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 16376 0 1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__082__B
timestamp 1586364061
transform 1 0 15732 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__082__A
timestamp 1586364061
transform 1 0 16100 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_7.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 15272 0 1 7072
box -38 -48 222 592
use scs8hd_decap_3  FILLER_9_156
timestamp 1586364061
transform 1 0 15456 0 1 7072
box -38 -48 314 592
use scs8hd_fill_2  FILLER_9_161
timestamp 1586364061
transform 1 0 15916 0 1 7072
box -38 -48 222 592
use scs8hd_fill_1  FILLER_9_165
timestamp 1586364061
transform 1 0 16284 0 1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 17388 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_175
timestamp 1586364061
transform 1 0 17204 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_179
timestamp 1586364061
transform 1 0 17572 0 1 7072
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_ipin_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18032 0 1 7072
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_96
timestamp 1586364061
transform 1 0 17940 0 1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 17756 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_193
timestamp 1586364061
transform 1 0 18860 0 1 7072
box -38 -48 222 592
use scs8hd_inv_1  mux_right_ipin_5.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 19596 0 1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_5.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 20056 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__093__B
timestamp 1586364061
transform 1 0 19044 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__093__A
timestamp 1586364061
transform 1 0 19412 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_197
timestamp 1586364061
transform 1 0 19228 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_204
timestamp 1586364061
transform 1 0 19872 0 1 7072
box -38 -48 222 592
use scs8hd_decap_3  PHY_19
timestamp 1586364061
transform -1 0 20884 0 1 7072
box -38 -48 314 592
use scs8hd_decap_4  FILLER_9_208
timestamp 1586364061
transform 1 0 20240 0 1 7072
box -38 -48 406 592
use scs8hd_inv_1  mux_right_ipin_2.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1932 0 -1 8160
box -38 -48 314 592
use scs8hd_decap_3  PHY_20
timestamp 1586364061
transform 1 0 1104 0 -1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__045__B
timestamp 1586364061
transform 1 0 1748 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_10_3
timestamp 1586364061
transform 1 0 1380 0 -1 8160
box -38 -48 406 592
use scs8hd_fill_2  FILLER_10_12
timestamp 1586364061
transform 1 0 2208 0 -1 8160
box -38 -48 222 592
use scs8hd_inv_1  mux_right_ipin_0.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 2944 0 -1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__058__A
timestamp 1586364061
transform 1 0 3404 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__045__A
timestamp 1586364061
transform 1 0 2392 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__061__A
timestamp 1586364061
transform 1 0 2760 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_16
timestamp 1586364061
transform 1 0 2576 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_23
timestamp 1586364061
transform 1 0 3220 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_27
timestamp 1586364061
transform 1 0 3588 0 -1 8160
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_ipin_2.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 4876 0 -1 8160
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_97
timestamp 1586364061
transform 1 0 3956 0 -1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__041__C
timestamp 1586364061
transform 1 0 3772 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__047__B
timestamp 1586364061
transform 1 0 4232 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_2.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 4692 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_32
timestamp 1586364061
transform 1 0 4048 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_3  FILLER_10_36
timestamp 1586364061
transform 1 0 4416 0 -1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_2.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 5888 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_50
timestamp 1586364061
transform 1 0 5704 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_8  FILLER_10_54
timestamp 1586364061
transform 1 0 6072 0 -1 8160
box -38 -48 774 592
use scs8hd_inv_1  mux_right_ipin_7.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 6808 0 -1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_2.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 7268 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_65
timestamp 1586364061
transform 1 0 7084 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_69
timestamp 1586364061
transform 1 0 7452 0 -1 8160
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_ipin_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 7820 0 -1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 7636 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_82
timestamp 1586364061
transform 1 0 8648 0 -1 8160
box -38 -48 222 592
use scs8hd_conb_1  _133_
timestamp 1586364061
transform 1 0 9844 0 -1 8160
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_98
timestamp 1586364061
transform 1 0 9568 0 -1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_2.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 9200 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 8832 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_86
timestamp 1586364061
transform 1 0 9016 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_90
timestamp 1586364061
transform 1 0 9384 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_93
timestamp 1586364061
transform 1 0 9660 0 -1 8160
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_right_ipin_7.LATCH_1_.latch
timestamp 1586364061
transform 1 0 10856 0 -1 8160
box -38 -48 1050 592
use scs8hd_decap_8  FILLER_10_98
timestamp 1586364061
transform 1 0 10120 0 -1 8160
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_7.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 12420 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_6  FILLER_10_117
timestamp 1586364061
transform 1 0 11868 0 -1 8160
box -38 -48 590 592
use scs8hd_lpflow_inputisolatch_1  mem_right_ipin_7.LATCH_3_.latch
timestamp 1586364061
transform 1 0 13248 0 -1 8160
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_7.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 12788 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_125
timestamp 1586364061
transform 1 0 12604 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_3  FILLER_10_129
timestamp 1586364061
transform 1 0 12972 0 -1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_7.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 14444 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_143
timestamp 1586364061
transform 1 0 14260 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_6  FILLER_10_147
timestamp 1586364061
transform 1 0 14628 0 -1 8160
box -38 -48 590 592
use scs8hd_nor2_4  _082_
timestamp 1586364061
transform 1 0 15732 0 -1 8160
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_99
timestamp 1586364061
transform 1 0 15180 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_4  FILLER_10_154
timestamp 1586364061
transform 1 0 15272 0 -1 8160
box -38 -48 406 592
use scs8hd_fill_1  FILLER_10_158
timestamp 1586364061
transform 1 0 15640 0 -1 8160
box -38 -48 130 592
use scs8hd_ebufn_2  mux_right_ipin_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 17296 0 -1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 16744 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 17112 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_168
timestamp 1586364061
transform 1 0 16560 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_172
timestamp 1586364061
transform 1 0 16928 0 -1 8160
box -38 -48 222 592
use scs8hd_nor2_4  _093_
timestamp 1586364061
transform 1 0 18860 0 -1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_5.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 18308 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 18676 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_185
timestamp 1586364061
transform 1 0 18124 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_189
timestamp 1586364061
transform 1 0 18492 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_8  FILLER_10_202
timestamp 1586364061
transform 1 0 19688 0 -1 8160
box -38 -48 774 592
use scs8hd_decap_3  PHY_21
timestamp 1586364061
transform -1 0 20884 0 -1 8160
box -38 -48 314 592
use scs8hd_fill_2  FILLER_10_210
timestamp 1586364061
transform 1 0 20424 0 -1 8160
box -38 -48 222 592
use scs8hd_inv_1  mux_right_ipin_2.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 2024 0 1 8160
box -38 -48 314 592
use scs8hd_decap_3  PHY_22
timestamp 1586364061
transform 1 0 1104 0 1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_2.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 1840 0 1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_11_3
timestamp 1586364061
transform 1 0 1380 0 1 8160
box -38 -48 406 592
use scs8hd_fill_1  FILLER_11_7
timestamp 1586364061
transform 1 0 1748 0 1 8160
box -38 -48 130 592
use scs8hd_fill_2  FILLER_11_13
timestamp 1586364061
transform 1 0 2300 0 1 8160
box -38 -48 222 592
use scs8hd_nor2_4  _058_
timestamp 1586364061
transform 1 0 3036 0 1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_2.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 2484 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__058__B
timestamp 1586364061
transform 1 0 2852 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_17
timestamp 1586364061
transform 1 0 2668 0 1 8160
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_right_ipin_2.LATCH_5_.latch
timestamp 1586364061
transform 1 0 4600 0 1 8160
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_2.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 4416 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_2.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 4048 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_30
timestamp 1586364061
transform 1 0 3864 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_34
timestamp 1586364061
transform 1 0 4232 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__094__B
timestamp 1586364061
transform 1 0 5796 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__094__A
timestamp 1586364061
transform 1 0 6164 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_49
timestamp 1586364061
transform 1 0 5612 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_53
timestamp 1586364061
transform 1 0 5980 0 1 8160
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_100
timestamp 1586364061
transform 1 0 6716 0 1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_2.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 6992 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_2.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 7360 0 1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_11_57
timestamp 1586364061
transform 1 0 6348 0 1 8160
box -38 -48 406 592
use scs8hd_fill_2  FILLER_11_62
timestamp 1586364061
transform 1 0 6808 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_66
timestamp 1586364061
transform 1 0 7176 0 1 8160
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_ipin_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 7636 0 1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_6.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 8648 0 1 8160
box -38 -48 222 592
use scs8hd_fill_1  FILLER_11_70
timestamp 1586364061
transform 1 0 7544 0 1 8160
box -38 -48 130 592
use scs8hd_fill_2  FILLER_11_80
timestamp 1586364061
transform 1 0 8464 0 1 8160
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_right_ipin_2.LATCH_3_.latch
timestamp 1586364061
transform 1 0 9200 0 1 8160
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_2.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 9016 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_84
timestamp 1586364061
transform 1 0 8832 0 1 8160
box -38 -48 222 592
use scs8hd_or2_4  _064_
timestamp 1586364061
transform 1 0 10948 0 1 8160
box -38 -48 682 592
use scs8hd_diode_2  ANTENNA__138__A
timestamp 1586364061
transform 1 0 10396 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__064__B
timestamp 1586364061
transform 1 0 10764 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_99
timestamp 1586364061
transform 1 0 10212 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_103
timestamp 1586364061
transform 1 0 10580 0 1 8160
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_ipin_7.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12420 0 1 8160
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_101
timestamp 1586364061
transform 1 0 12328 0 1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__064__A
timestamp 1586364061
transform 1 0 11776 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_7.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 12144 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_114
timestamp 1586364061
transform 1 0 11592 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_118
timestamp 1586364061
transform 1 0 11960 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_7.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 13616 0 1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_11_132
timestamp 1586364061
transform 1 0 13248 0 1 8160
box -38 -48 406 592
use scs8hd_decap_4  FILLER_11_138
timestamp 1586364061
transform 1 0 13800 0 1 8160
box -38 -48 406 592
use scs8hd_ebufn_2  mux_right_ipin_7.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 14352 0 1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_7.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14168 0 1 8160
box -38 -48 222 592
use scs8hd_nor2_4  _080_
timestamp 1586364061
transform 1 0 15916 0 1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__139__A
timestamp 1586364061
transform 1 0 15456 0 1 8160
box -38 -48 222 592
use scs8hd_decap_3  FILLER_11_153
timestamp 1586364061
transform 1 0 15180 0 1 8160
box -38 -48 314 592
use scs8hd_decap_3  FILLER_11_158
timestamp 1586364061
transform 1 0 15640 0 1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_5.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 16928 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_5.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 17296 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_170
timestamp 1586364061
transform 1 0 16744 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_174
timestamp 1586364061
transform 1 0 17112 0 1 8160
box -38 -48 222 592
use scs8hd_decap_3  FILLER_11_178
timestamp 1586364061
transform 1 0 17480 0 1 8160
box -38 -48 314 592
use scs8hd_ebufn_2  mux_right_ipin_5.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18124 0 1 8160
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_102
timestamp 1586364061
transform 1 0 17940 0 1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_5.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 17756 0 1 8160
box -38 -48 222 592
use scs8hd_fill_1  FILLER_11_184
timestamp 1586364061
transform 1 0 18032 0 1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_5.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 19136 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_5.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 19504 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_194
timestamp 1586364061
transform 1 0 18952 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_198
timestamp 1586364061
transform 1 0 19320 0 1 8160
box -38 -48 222 592
use scs8hd_decap_8  FILLER_11_202
timestamp 1586364061
transform 1 0 19688 0 1 8160
box -38 -48 774 592
use scs8hd_decap_3  PHY_23
timestamp 1586364061
transform -1 0 20884 0 1 8160
box -38 -48 314 592
use scs8hd_fill_2  FILLER_11_210
timestamp 1586364061
transform 1 0 20424 0 1 8160
box -38 -48 222 592
use scs8hd_inv_1  mux_right_ipin_2.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1932 0 -1 9248
box -38 -48 314 592
use scs8hd_decap_3  PHY_24
timestamp 1586364061
transform 1 0 1104 0 -1 9248
box -38 -48 314 592
use scs8hd_decap_6  FILLER_12_3
timestamp 1586364061
transform 1 0 1380 0 -1 9248
box -38 -48 590 592
use scs8hd_decap_6  FILLER_12_12
timestamp 1586364061
transform 1 0 2208 0 -1 9248
box -38 -48 590 592
use scs8hd_inv_1  mux_right_ipin_2.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 2944 0 -1 9248
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__056__B
timestamp 1586364061
transform 1 0 3588 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_2.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 2760 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_12_23
timestamp 1586364061
transform 1 0 3220 0 -1 9248
box -38 -48 406 592
use scs8hd_conb_1  _128_
timestamp 1586364061
transform 1 0 4140 0 -1 9248
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_103
timestamp 1586364061
transform 1 0 3956 0 -1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__059__A
timestamp 1586364061
transform 1 0 4600 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_29
timestamp 1586364061
transform 1 0 3772 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_1  FILLER_12_32
timestamp 1586364061
transform 1 0 4048 0 -1 9248
box -38 -48 130 592
use scs8hd_fill_2  FILLER_12_36
timestamp 1586364061
transform 1 0 4416 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_40
timestamp 1586364061
transform 1 0 4784 0 -1 9248
box -38 -48 222 592
use scs8hd_nor2_4  _094_
timestamp 1586364061
transform 1 0 5152 0 -1 9248
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_2.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 4968 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_2.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 6164 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_53
timestamp 1586364061
transform 1 0 5980 0 -1 9248
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_right_ipin_2.LATCH_1_.latch
timestamp 1586364061
transform 1 0 6716 0 -1 9248
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_2.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 6532 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_57
timestamp 1586364061
transform 1 0 6348 0 -1 9248
box -38 -48 222 592
use scs8hd_inv_1  mux_right_ipin_6.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 8556 0 -1 9248
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_2.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 7912 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 8280 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_72
timestamp 1586364061
transform 1 0 7728 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_76
timestamp 1586364061
transform 1 0 8096 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_1  FILLER_12_80
timestamp 1586364061
transform 1 0 8464 0 -1 9248
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_104
timestamp 1586364061
transform 1 0 9568 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_8  FILLER_12_84
timestamp 1586364061
transform 1 0 8832 0 -1 9248
box -38 -48 774 592
use scs8hd_decap_4  FILLER_12_93
timestamp 1586364061
transform 1 0 9660 0 -1 9248
box -38 -48 406 592
use scs8hd_buf_2  _138_
timestamp 1586364061
transform 1 0 10028 0 -1 9248
box -38 -48 406 592
use scs8hd_ebufn_2  mux_right_ipin_7.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 11132 0 -1 9248
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_7.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 10580 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_7.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10948 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_101
timestamp 1586364061
transform 1 0 10396 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_105
timestamp 1586364061
transform 1 0 10764 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_6  FILLER_12_118
timestamp 1586364061
transform 1 0 11960 0 -1 9248
box -38 -48 590 592
use scs8hd_fill_1  FILLER_12_124
timestamp 1586364061
transform 1 0 12512 0 -1 9248
box -38 -48 130 592
use scs8hd_ebufn_2  mux_right_ipin_7.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 13616 0 -1 9248
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_7.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 12604 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_7.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 13432 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_6  FILLER_12_127
timestamp 1586364061
transform 1 0 12788 0 -1 9248
box -38 -48 590 592
use scs8hd_fill_1  FILLER_12_133
timestamp 1586364061
transform 1 0 13340 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_8  FILLER_12_145
timestamp 1586364061
transform 1 0 14444 0 -1 9248
box -38 -48 774 592
use scs8hd_buf_2  _139_
timestamp 1586364061
transform 1 0 15456 0 -1 9248
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_105
timestamp 1586364061
transform 1 0 15180 0 -1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__080__B
timestamp 1586364061
transform 1 0 16008 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__080__A
timestamp 1586364061
transform 1 0 16376 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_154
timestamp 1586364061
transform 1 0 15272 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_160
timestamp 1586364061
transform 1 0 15824 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_164
timestamp 1586364061
transform 1 0 16192 0 -1 9248
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_right_ipin_5.LATCH_0_.latch
timestamp 1586364061
transform 1 0 16560 0 -1 9248
box -38 -48 1050 592
use scs8hd_decap_4  FILLER_12_179
timestamp 1586364061
transform 1 0 17572 0 -1 9248
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_right_ipin_5.LATCH_2_.latch
timestamp 1586364061
transform 1 0 18308 0 -1 9248
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_5.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 18032 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_1  FILLER_12_183
timestamp 1586364061
transform 1 0 17940 0 -1 9248
box -38 -48 130 592
use scs8hd_fill_1  FILLER_12_186
timestamp 1586364061
transform 1 0 18216 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_12  FILLER_12_198
timestamp 1586364061
transform 1 0 19320 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_3  PHY_25
timestamp 1586364061
transform -1 0 20884 0 -1 9248
box -38 -48 314 592
use scs8hd_fill_2  FILLER_12_210
timestamp 1586364061
transform 1 0 20424 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_3
timestamp 1586364061
transform 1 0 1380 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__134__A
timestamp 1586364061
transform 1 0 1564 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_3  PHY_28
timestamp 1586364061
transform 1 0 1104 0 -1 10336
box -38 -48 314 592
use scs8hd_decap_3  PHY_26
timestamp 1586364061
transform 1 0 1104 0 1 9248
box -38 -48 314 592
use scs8hd_buf_2  _141_
timestamp 1586364061
transform 1 0 1380 0 1 9248
box -38 -48 406 592
use scs8hd_fill_2  FILLER_14_7
timestamp 1586364061
transform 1 0 1748 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_11
timestamp 1586364061
transform 1 0 2116 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_7
timestamp 1586364061
transform 1 0 1748 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_7.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 2300 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__141__A
timestamp 1586364061
transform 1 0 1932 0 1 9248
box -38 -48 222 592
use scs8hd_inv_1  mux_right_ipin_7.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1932 0 -1 10336
box -38 -48 314 592
use scs8hd_decap_8  FILLER_14_12
timestamp 1586364061
transform 1 0 2208 0 -1 10336
box -38 -48 774 592
use scs8hd_fill_2  FILLER_13_19
timestamp 1586364061
transform 1 0 2852 0 1 9248
box -38 -48 222 592
use scs8hd_fill_1  FILLER_13_15
timestamp 1586364061
transform 1 0 2484 0 1 9248
box -38 -48 130 592
use scs8hd_inv_1  mux_right_ipin_7.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 2576 0 1 9248
box -38 -48 314 592
use scs8hd_inv_1  mux_right_ipin_7.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 2944 0 -1 10336
box -38 -48 314 592
use scs8hd_decap_4  FILLER_14_23
timestamp 1586364061
transform 1 0 3220 0 -1 10336
box -38 -48 406 592
use scs8hd_fill_2  FILLER_13_23
timestamp 1586364061
transform 1 0 3220 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__060__B
timestamp 1586364061
transform 1 0 3588 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_7.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 3404 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_7.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 3036 0 1 9248
box -38 -48 222 592
use scs8hd_nor2_4  _056_
timestamp 1586364061
transform 1 0 3588 0 1 9248
box -38 -48 866 592
use scs8hd_nor2_4  _059_
timestamp 1586364061
transform 1 0 4324 0 -1 10336
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_109
timestamp 1586364061
transform 1 0 3956 0 -1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__059__B
timestamp 1586364061
transform 1 0 4600 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_36
timestamp 1586364061
transform 1 0 4416 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_40
timestamp 1586364061
transform 1 0 4784 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_29
timestamp 1586364061
transform 1 0 3772 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_3  FILLER_14_32
timestamp 1586364061
transform 1 0 4048 0 -1 10336
box -38 -48 314 592
use scs8hd_ebufn_2  mux_right_ipin_2.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 5152 0 1 9248
box -38 -48 866 592
use scs8hd_ebufn_2  mux_right_ipin_2.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 5888 0 -1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__056__A
timestamp 1586364061
transform 1 0 4968 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__098__A
timestamp 1586364061
transform 1 0 5336 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__070__A
timestamp 1586364061
transform 1 0 5704 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_2.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 6164 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_53
timestamp 1586364061
transform 1 0 5980 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_44
timestamp 1586364061
transform 1 0 5152 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_48
timestamp 1586364061
transform 1 0 5520 0 -1 10336
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_right_ipin_2.LATCH_2_.latch
timestamp 1586364061
transform 1 0 6808 0 1 9248
box -38 -48 1050 592
use scs8hd_ebufn_2  mux_right_ipin_2.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 7452 0 -1 10336
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_106
timestamp 1586364061
transform 1 0 6716 0 1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_2.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 6532 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_2.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 6900 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 7268 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_57
timestamp 1586364061
transform 1 0 6348 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_61
timestamp 1586364061
transform 1 0 6716 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_65
timestamp 1586364061
transform 1 0 7084 0 -1 10336
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_ipin_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 8556 0 1 9248
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 8372 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_2.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 8004 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 8556 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_73
timestamp 1586364061
transform 1 0 7820 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_77
timestamp 1586364061
transform 1 0 8188 0 1 9248
box -38 -48 222 592
use scs8hd_decap_3  FILLER_14_78
timestamp 1586364061
transform 1 0 8280 0 -1 10336
box -38 -48 314 592
use scs8hd_decap_8  FILLER_14_83
timestamp 1586364061
transform 1 0 8740 0 -1 10336
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_110
timestamp 1586364061
transform 1 0 9568 0 -1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_3.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 9844 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_7.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9660 0 1 9248
box -38 -48 222 592
use scs8hd_decap_3  FILLER_13_90
timestamp 1586364061
transform 1 0 9384 0 1 9248
box -38 -48 314 592
use scs8hd_fill_2  FILLER_13_95
timestamp 1586364061
transform 1 0 9844 0 1 9248
box -38 -48 222 592
use scs8hd_fill_1  FILLER_14_91
timestamp 1586364061
transform 1 0 9476 0 -1 10336
box -38 -48 130 592
use scs8hd_fill_2  FILLER_14_93
timestamp 1586364061
transform 1 0 9660 0 -1 10336
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_right_ipin_7.LATCH_0_.latch
timestamp 1586364061
transform 1 0 10488 0 1 9248
box -38 -48 1050 592
use scs8hd_inv_1  mux_right_ipin_6.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 10028 0 -1 10336
box -38 -48 314 592
use scs8hd_ebufn_2  mux_right_ipin_7.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 11040 0 -1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_6.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 10028 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_7.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 10488 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_3.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10856 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_3  FILLER_13_99
timestamp 1586364061
transform 1 0 10212 0 1 9248
box -38 -48 314 592
use scs8hd_fill_2  FILLER_14_100
timestamp 1586364061
transform 1 0 10304 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_104
timestamp 1586364061
transform 1 0 10672 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_113
timestamp 1586364061
transform 1 0 11500 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_117
timestamp 1586364061
transform 1 0 11868 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_3  FILLER_13_117
timestamp 1586364061
transform 1 0 11868 0 1 9248
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_7.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 11684 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_121
timestamp 1586364061
transform 1 0 12236 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_3.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 12052 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_7.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 12144 0 1 9248
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_107
timestamp 1586364061
transform 1 0 12328 0 1 9248
box -38 -48 130 592
use scs8hd_fill_2  FILLER_13_123
timestamp 1586364061
transform 1 0 12420 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_7.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 12420 0 -1 10336
box -38 -48 222 592
use scs8hd_buf_2  _136_
timestamp 1586364061
transform 1 0 12604 0 1 9248
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_right_ipin_7.LATCH_2_.latch
timestamp 1586364061
transform 1 0 12604 0 -1 10336
box -38 -48 1050 592
use scs8hd_lpflow_inputisolatch_1  mem_right_ipin_7.LATCH_4_.latch
timestamp 1586364061
transform 1 0 13708 0 1 9248
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA__136__A
timestamp 1586364061
transform 1 0 13156 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_7.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 13524 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_7.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 13800 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_129
timestamp 1586364061
transform 1 0 12972 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_133
timestamp 1586364061
transform 1 0 13340 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_136
timestamp 1586364061
transform 1 0 13616 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_7.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14260 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_6  FILLER_13_148
timestamp 1586364061
transform 1 0 14720 0 1 9248
box -38 -48 590 592
use scs8hd_decap_3  FILLER_14_140
timestamp 1586364061
transform 1 0 13984 0 -1 10336
box -38 -48 314 592
use scs8hd_decap_8  FILLER_14_145
timestamp 1586364061
transform 1 0 14444 0 -1 10336
box -38 -48 774 592
use scs8hd_fill_2  FILLER_14_158
timestamp 1586364061
transform 1 0 15640 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_13_156
timestamp 1586364061
transform 1 0 15456 0 1 9248
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__135__A
timestamp 1586364061
transform 1 0 15272 0 1 9248
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_111
timestamp 1586364061
transform 1 0 15180 0 -1 10336
box -38 -48 130 592
use scs8hd_buf_2  _135_
timestamp 1586364061
transform 1 0 15272 0 -1 10336
box -38 -48 406 592
use scs8hd_fill_2  FILLER_14_162
timestamp 1586364061
transform 1 0 16008 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_162
timestamp 1586364061
transform 1 0 16008 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_5.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 16192 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_5.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 15824 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_5.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 15824 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_5.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 16192 0 1 9248
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_ipin_5.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 16376 0 1 9248
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  mem_right_ipin_5.LATCH_3_.latch
timestamp 1586364061
transform 1 0 16376 0 -1 10336
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_5.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 17388 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_175
timestamp 1586364061
transform 1 0 17204 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_179
timestamp 1586364061
transform 1 0 17572 0 1 9248
box -38 -48 222 592
use scs8hd_decap_8  FILLER_14_177
timestamp 1586364061
transform 1 0 17388 0 -1 10336
box -38 -48 774 592
use scs8hd_ebufn_2  mux_right_ipin_5.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18032 0 1 9248
box -38 -48 866 592
use scs8hd_ebufn_2  mux_right_ipin_5.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18308 0 -1 10336
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_108
timestamp 1586364061
transform 1 0 17940 0 1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_5.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 17756 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_193
timestamp 1586364061
transform 1 0 18860 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_185
timestamp 1586364061
transform 1 0 18124 0 -1 10336
box -38 -48 222 592
use scs8hd_conb_1  _131_
timestamp 1586364061
transform 1 0 19596 0 1 9248
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_5.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 19044 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_5.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 19412 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_5.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 19320 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_197
timestamp 1586364061
transform 1 0 19228 0 1 9248
box -38 -48 222 592
use scs8hd_decap_8  FILLER_13_204
timestamp 1586364061
transform 1 0 19872 0 1 9248
box -38 -48 774 592
use scs8hd_fill_2  FILLER_14_196
timestamp 1586364061
transform 1 0 19136 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_12  FILLER_14_200
timestamp 1586364061
transform 1 0 19504 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_3  PHY_27
timestamp 1586364061
transform -1 0 20884 0 1 9248
box -38 -48 314 592
use scs8hd_decap_3  PHY_29
timestamp 1586364061
transform -1 0 20884 0 -1 10336
box -38 -48 314 592
use scs8hd_inv_1  mux_right_ipin_2.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1564 0 1 10336
box -38 -48 314 592
use scs8hd_decap_3  PHY_30
timestamp 1586364061
transform 1 0 1104 0 1 10336
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_2.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 2024 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_3
timestamp 1586364061
transform 1 0 1380 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_8
timestamp 1586364061
transform 1 0 1840 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_12
timestamp 1586364061
transform 1 0 2208 0 1 10336
box -38 -48 222 592
use scs8hd_nor2_4  _060_
timestamp 1586364061
transform 1 0 3588 0 1 10336
box -38 -48 866 592
use scs8hd_inv_1  mux_right_ipin_2.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 2576 0 1 10336
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_2.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 3036 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_3.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 3404 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__060__A
timestamp 1586364061
transform 1 0 2392 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_19
timestamp 1586364061
transform 1 0 2852 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_23
timestamp 1586364061
transform 1 0 3220 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__070__B
timestamp 1586364061
transform 1 0 4600 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_36
timestamp 1586364061
transform 1 0 4416 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_40
timestamp 1586364061
transform 1 0 4784 0 1 10336
box -38 -48 222 592
use scs8hd_nor2_4  _098_
timestamp 1586364061
transform 1 0 5152 0 1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__098__B
timestamp 1586364061
transform 1 0 4968 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__096__B
timestamp 1586364061
transform 1 0 6164 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_53
timestamp 1586364061
transform 1 0 5980 0 1 10336
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_112
timestamp 1586364061
transform 1 0 6716 0 1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__096__A
timestamp 1586364061
transform 1 0 6532 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 7268 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_57
timestamp 1586364061
transform 1 0 6348 0 1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_15_62
timestamp 1586364061
transform 1 0 6808 0 1 10336
box -38 -48 406 592
use scs8hd_fill_1  FILLER_15_66
timestamp 1586364061
transform 1 0 7176 0 1 10336
box -38 -48 130 592
use scs8hd_decap_3  FILLER_15_69
timestamp 1586364061
transform 1 0 7452 0 1 10336
box -38 -48 314 592
use scs8hd_ebufn_2  mux_left_ipin_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 7728 0 1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 8740 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_81
timestamp 1586364061
transform 1 0 8556 0 1 10336
box -38 -48 222 592
use scs8hd_inv_1  mux_left_ipin_0.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 9292 0 1 10336
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 9752 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_3.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9108 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_85
timestamp 1586364061
transform 1 0 8924 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_92
timestamp 1586364061
transform 1 0 9568 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_96
timestamp 1586364061
transform 1 0 9936 0 1 10336
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_ipin_3.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10488 0 1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_3.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 10120 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_100
timestamp 1586364061
transform 1 0 10304 0 1 10336
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_113
timestamp 1586364061
transform 1 0 12328 0 1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_3.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 11500 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_7.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 12144 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_111
timestamp 1586364061
transform 1 0 11316 0 1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_15_115
timestamp 1586364061
transform 1 0 11684 0 1 10336
box -38 -48 406 592
use scs8hd_fill_1  FILLER_15_119
timestamp 1586364061
transform 1 0 12052 0 1 10336
box -38 -48 130 592
use scs8hd_decap_3  FILLER_15_123
timestamp 1586364061
transform 1 0 12420 0 1 10336
box -38 -48 314 592
use scs8hd_ebufn_2  mux_right_ipin_7.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12696 0 1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_7.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 13708 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_135
timestamp 1586364061
transform 1 0 13524 0 1 10336
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_ipin_7.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 14260 0 1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_7.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 14076 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_139
timestamp 1586364061
transform 1 0 13892 0 1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_15_152
timestamp 1586364061
transform 1 0 15088 0 1 10336
box -38 -48 406 592
use scs8hd_ebufn_2  mux_right_ipin_5.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 16376 0 1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_5.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 15548 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_5.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 16192 0 1 10336
box -38 -48 222 592
use scs8hd_fill_1  FILLER_15_156
timestamp 1586364061
transform 1 0 15456 0 1 10336
box -38 -48 130 592
use scs8hd_decap_4  FILLER_15_159
timestamp 1586364061
transform 1 0 15732 0 1 10336
box -38 -48 406 592
use scs8hd_fill_1  FILLER_15_163
timestamp 1586364061
transform 1 0 16100 0 1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_5.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 17388 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_175
timestamp 1586364061
transform 1 0 17204 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_179
timestamp 1586364061
transform 1 0 17572 0 1 10336
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_ipin_5.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18492 0 1 10336
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_114
timestamp 1586364061
transform 1 0 17940 0 1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_5.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 18308 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_5.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 17756 0 1 10336
box -38 -48 222 592
use scs8hd_decap_3  FILLER_15_184
timestamp 1586364061
transform 1 0 18032 0 1 10336
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_5.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 19504 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_5.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 19872 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_198
timestamp 1586364061
transform 1 0 19320 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_202
timestamp 1586364061
transform 1 0 19688 0 1 10336
box -38 -48 222 592
use scs8hd_decap_6  FILLER_15_206
timestamp 1586364061
transform 1 0 20056 0 1 10336
box -38 -48 590 592
use scs8hd_decap_3  PHY_31
timestamp 1586364061
transform -1 0 20884 0 1 10336
box -38 -48 314 592
use scs8hd_buf_2  _134_
timestamp 1586364061
transform 1 0 1380 0 -1 11424
box -38 -48 406 592
use scs8hd_decap_3  PHY_32
timestamp 1586364061
transform 1 0 1104 0 -1 11424
box -38 -48 314 592
use scs8hd_decap_12  FILLER_16_7
timestamp 1586364061
transform 1 0 1748 0 -1 11424
box -38 -48 1142 592
use scs8hd_inv_1  mux_right_ipin_3.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 2944 0 -1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__069__B
timestamp 1586364061
transform 1 0 3588 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_1  FILLER_16_19
timestamp 1586364061
transform 1 0 2852 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_4  FILLER_16_23
timestamp 1586364061
transform 1 0 3220 0 -1 11424
box -38 -48 406 592
use scs8hd_nor2_4  _070_
timestamp 1586364061
transform 1 0 4140 0 -1 11424
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_115
timestamp 1586364061
transform 1 0 3956 0 -1 11424
box -38 -48 130 592
use scs8hd_fill_2  FILLER_16_29
timestamp 1586364061
transform 1 0 3772 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_1  FILLER_16_32
timestamp 1586364061
transform 1 0 4048 0 -1 11424
box -38 -48 130 592
use scs8hd_nor2_4  _096_
timestamp 1586364061
transform 1 0 5704 0 -1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__122__B
timestamp 1586364061
transform 1 0 5152 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__090__A
timestamp 1586364061
transform 1 0 5520 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_42
timestamp 1586364061
transform 1 0 4968 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_46
timestamp 1586364061
transform 1 0 5336 0 -1 11424
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_ipin_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 7268 0 -1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_0.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 6716 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_0.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 7084 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_59
timestamp 1586364061
transform 1 0 6532 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_63
timestamp 1586364061
transform 1 0 6900 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 8280 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 8648 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_76
timestamp 1586364061
transform 1 0 8096 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_80
timestamp 1586364061
transform 1 0 8464 0 -1 11424
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_right_ipin_3.LATCH_0_.latch
timestamp 1586364061
transform 1 0 9752 0 -1 11424
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_116
timestamp 1586364061
transform 1 0 9568 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_8  FILLER_16_84
timestamp 1586364061
transform 1 0 8832 0 -1 11424
box -38 -48 774 592
use scs8hd_fill_1  FILLER_16_93
timestamp 1586364061
transform 1 0 9660 0 -1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_3.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11224 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_16_105
timestamp 1586364061
transform 1 0 10764 0 -1 11424
box -38 -48 406 592
use scs8hd_fill_1  FILLER_16_109
timestamp 1586364061
transform 1 0 11132 0 -1 11424
box -38 -48 130 592
use scs8hd_ebufn_2  mux_right_ipin_3.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 11500 0 -1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_7.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 12512 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_1  FILLER_16_112
timestamp 1586364061
transform 1 0 11408 0 -1 11424
box -38 -48 130 592
use scs8hd_fill_2  FILLER_16_122
timestamp 1586364061
transform 1 0 12328 0 -1 11424
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_ipin_7.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 13248 0 -1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_6.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 12880 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_126
timestamp 1586364061
transform 1 0 12696 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_130
timestamp 1586364061
transform 1 0 13064 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14812 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_6.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14260 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_141
timestamp 1586364061
transform 1 0 14076 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_16_145
timestamp 1586364061
transform 1 0 14444 0 -1 11424
box -38 -48 406 592
use scs8hd_fill_2  FILLER_16_151
timestamp 1586364061
transform 1 0 14996 0 -1 11424
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_right_ipin_5.LATCH_1_.latch
timestamp 1586364061
transform 1 0 15548 0 -1 11424
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_117
timestamp 1586364061
transform 1 0 15180 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_3  FILLER_16_154
timestamp 1586364061
transform 1 0 15272 0 -1 11424
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_right_ipin_5.LATCH_4_.latch
timestamp 1586364061
transform 1 0 17296 0 -1 11424
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 16744 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_5.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 17112 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_168
timestamp 1586364061
transform 1 0 16560 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_172
timestamp 1586364061
transform 1 0 16928 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_5.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 18584 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_3  FILLER_16_187
timestamp 1586364061
transform 1 0 18308 0 -1 11424
box -38 -48 314 592
use scs8hd_decap_3  FILLER_16_192
timestamp 1586364061
transform 1 0 18768 0 -1 11424
box -38 -48 314 592
use scs8hd_ebufn_2  mux_right_ipin_5.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 19044 0 -1 11424
box -38 -48 866 592
use scs8hd_decap_8  FILLER_16_204
timestamp 1586364061
transform 1 0 19872 0 -1 11424
box -38 -48 774 592
use scs8hd_decap_3  PHY_33
timestamp 1586364061
transform -1 0 20884 0 -1 11424
box -38 -48 314 592
use scs8hd_inv_1  mux_left_ipin_0.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1564 0 1 11424
box -38 -48 314 592
use scs8hd_decap_3  PHY_34
timestamp 1586364061
transform 1 0 1104 0 1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 2024 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_3
timestamp 1586364061
transform 1 0 1380 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_8
timestamp 1586364061
transform 1 0 1840 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_12
timestamp 1586364061
transform 1 0 2208 0 1 11424
box -38 -48 222 592
use scs8hd_nor2_4  _069_
timestamp 1586364061
transform 1 0 3588 0 1 11424
box -38 -48 866 592
use scs8hd_inv_1  mux_right_ipin_3.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 2576 0 1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_3.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 3036 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_3.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 3404 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 2392 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_19
timestamp 1586364061
transform 1 0 2852 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_23
timestamp 1586364061
transform 1 0 3220 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__122__A
timestamp 1586364061
transform 1 0 4600 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_36
timestamp 1586364061
transform 1 0 4416 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_40
timestamp 1586364061
transform 1 0 4784 0 1 11424
box -38 -48 222 592
use scs8hd_nor2_4  _090_
timestamp 1586364061
transform 1 0 5152 0 1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_0.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 6164 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__090__B
timestamp 1586364061
transform 1 0 4968 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_53
timestamp 1586364061
transform 1 0 5980 0 1 11424
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_left_ipin_0.LATCH_1_.latch
timestamp 1586364061
transform 1 0 6808 0 1 11424
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_118
timestamp 1586364061
transform 1 0 6716 0 1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_0.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 6532 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_57
timestamp 1586364061
transform 1 0 6348 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 8004 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_3.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 8556 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_73
timestamp 1586364061
transform 1 0 7820 0 1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_17_77
timestamp 1586364061
transform 1 0 8188 0 1 11424
box -38 -48 406 592
use scs8hd_fill_2  FILLER_17_83
timestamp 1586364061
transform 1 0 8740 0 1 11424
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_right_ipin_3.LATCH_1_.latch
timestamp 1586364061
transform 1 0 9476 0 1 11424
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_3.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 9292 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 8924 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_87
timestamp 1586364061
transform 1 0 9108 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_3.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 11132 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10672 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_102
timestamp 1586364061
transform 1 0 10488 0 1 11424
box -38 -48 222 592
use scs8hd_decap_3  FILLER_17_106
timestamp 1586364061
transform 1 0 10856 0 1 11424
box -38 -48 314 592
use scs8hd_inv_1  mux_right_ipin_5.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 11316 0 1 11424
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_119
timestamp 1586364061
transform 1 0 12328 0 1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_5.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 11776 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_114
timestamp 1586364061
transform 1 0 11592 0 1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_17_118
timestamp 1586364061
transform 1 0 11960 0 1 11424
box -38 -48 406 592
use scs8hd_decap_3  FILLER_17_123
timestamp 1586364061
transform 1 0 12420 0 1 11424
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_right_ipin_6.LATCH_1_.latch
timestamp 1586364061
transform 1 0 12880 0 1 11424
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_6.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 12696 0 1 11424
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_ipin_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 14812 0 1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 14628 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_6.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 14076 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_139
timestamp 1586364061
transform 1 0 13892 0 1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_17_143
timestamp 1586364061
transform 1 0 14260 0 1 11424
box -38 -48 406 592
use scs8hd_ebufn_2  mux_right_ipin_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 16376 0 1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 16192 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_6.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 15824 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_158
timestamp 1586364061
transform 1 0 15640 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_162
timestamp 1586364061
transform 1 0 16008 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_5.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 17388 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_175
timestamp 1586364061
transform 1 0 17204 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_179
timestamp 1586364061
transform 1 0 17572 0 1 11424
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_ipin_5.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18584 0 1 11424
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_120
timestamp 1586364061
transform 1 0 17940 0 1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_5.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 18400 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_5.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 17756 0 1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_17_184
timestamp 1586364061
transform 1 0 18032 0 1 11424
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_5.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 19596 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_5.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 19964 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_199
timestamp 1586364061
transform 1 0 19412 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_203
timestamp 1586364061
transform 1 0 19780 0 1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_17_207
timestamp 1586364061
transform 1 0 20148 0 1 11424
box -38 -48 406 592
use scs8hd_decap_3  PHY_35
timestamp 1586364061
transform -1 0 20884 0 1 11424
box -38 -48 314 592
use scs8hd_fill_1  FILLER_17_211
timestamp 1586364061
transform 1 0 20516 0 1 11424
box -38 -48 130 592
use scs8hd_inv_1  mux_left_ipin_0.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1932 0 -1 12512
box -38 -48 314 592
use scs8hd_decap_3  PHY_36
timestamp 1586364061
transform 1 0 1104 0 -1 12512
box -38 -48 314 592
use scs8hd_decap_6  FILLER_18_3
timestamp 1586364061
transform 1 0 1380 0 -1 12512
box -38 -48 590 592
use scs8hd_decap_8  FILLER_18_12
timestamp 1586364061
transform 1 0 2208 0 -1 12512
box -38 -48 774 592
use scs8hd_inv_1  mux_right_ipin_3.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 2944 0 -1 12512
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__069__A
timestamp 1586364061
transform 1 0 3588 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_18_23
timestamp 1586364061
transform 1 0 3220 0 -1 12512
box -38 -48 406 592
use scs8hd_nor2_4  _122_
timestamp 1586364061
transform 1 0 4600 0 -1 12512
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_121
timestamp 1586364061
transform 1 0 3956 0 -1 12512
box -38 -48 130 592
use scs8hd_fill_2  FILLER_18_29
timestamp 1586364061
transform 1 0 3772 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_6  FILLER_18_32
timestamp 1586364061
transform 1 0 4048 0 -1 12512
box -38 -48 590 592
use scs8hd_lpflow_inputisolatch_1  mem_left_ipin_0.LATCH_0_.latch
timestamp 1586364061
transform 1 0 6164 0 -1 12512
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA__039__A
timestamp 1586364061
transform 1 0 5612 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 5980 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_47
timestamp 1586364061
transform 1 0 5428 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_51
timestamp 1586364061
transform 1 0 5796 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 7360 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_66
timestamp 1586364061
transform 1 0 7176 0 -1 12512
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_ipin_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 7912 0 -1 12512
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 7728 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_70
timestamp 1586364061
transform 1 0 7544 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_83
timestamp 1586364061
transform 1 0 8740 0 -1 12512
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_ipin_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9660 0 -1 12512
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_122
timestamp 1586364061
transform 1 0 9568 0 -1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 8924 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_18_87
timestamp 1586364061
transform 1 0 9108 0 -1 12512
box -38 -48 406 592
use scs8hd_fill_1  FILLER_18_91
timestamp 1586364061
transform 1 0 9476 0 -1 12512
box -38 -48 130 592
use scs8hd_ebufn_2  mux_right_ipin_3.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 11224 0 -1 12512
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_3.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10672 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_102
timestamp 1586364061
transform 1 0 10488 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_18_106
timestamp 1586364061
transform 1 0 10856 0 -1 12512
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_6.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 12236 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_119
timestamp 1586364061
transform 1 0 12052 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_3  FILLER_18_123
timestamp 1586364061
transform 1 0 12420 0 -1 12512
box -38 -48 314 592
use scs8hd_ebufn_2  mux_right_ipin_6.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 13616 0 -1 12512
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_6.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 12696 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_6.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 13432 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_6  FILLER_18_128
timestamp 1586364061
transform 1 0 12880 0 -1 12512
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_6.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14996 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_6.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14628 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_145
timestamp 1586364061
transform 1 0 14444 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_149
timestamp 1586364061
transform 1 0 14812 0 -1 12512
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_ipin_6.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15272 0 -1 12512
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_123
timestamp 1586364061
transform 1 0 15180 0 -1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_1.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 16284 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_163
timestamp 1586364061
transform 1 0 16100 0 -1 12512
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_right_ipin_5.LATCH_5_.latch
timestamp 1586364061
transform 1 0 17112 0 -1 12512
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_1.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 16652 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_167
timestamp 1586364061
transform 1 0 16468 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_3  FILLER_18_171
timestamp 1586364061
transform 1 0 16836 0 -1 12512
box -38 -48 314 592
use scs8hd_ebufn_2  mux_right_ipin_5.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18860 0 -1 12512
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 18308 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 18676 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_185
timestamp 1586364061
transform 1 0 18124 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_189
timestamp 1586364061
transform 1 0 18492 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_8  FILLER_18_202
timestamp 1586364061
transform 1 0 19688 0 -1 12512
box -38 -48 774 592
use scs8hd_decap_3  PHY_37
timestamp 1586364061
transform -1 0 20884 0 -1 12512
box -38 -48 314 592
use scs8hd_fill_2  FILLER_18_210
timestamp 1586364061
transform 1 0 20424 0 -1 12512
box -38 -48 222 592
use scs8hd_inv_1  mux_right_ipin_4.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 2116 0 1 12512
box -38 -48 314 592
use scs8hd_decap_3  PHY_38
timestamp 1586364061
transform 1 0 1104 0 1 12512
box -38 -48 314 592
use scs8hd_decap_3  PHY_40
timestamp 1586364061
transform 1 0 1104 0 -1 13600
box -38 -48 314 592
use scs8hd_decap_8  FILLER_19_3
timestamp 1586364061
transform 1 0 1380 0 1 12512
box -38 -48 774 592
use scs8hd_decap_12  FILLER_20_3
timestamp 1586364061
transform 1 0 1380 0 -1 13600
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_20_19
timestamp 1586364061
transform 1 0 2852 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_4  FILLER_20_15
timestamp 1586364061
transform 1 0 2484 0 -1 13600
box -38 -48 406 592
use scs8hd_fill_2  FILLER_19_18
timestamp 1586364061
transform 1 0 2760 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_14
timestamp 1586364061
transform 1 0 2392 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_4.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 2944 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_4.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 2576 0 1 12512
box -38 -48 222 592
use scs8hd_inv_1  mux_right_ipin_4.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 2944 0 -1 13600
box -38 -48 314 592
use scs8hd_fill_2  FILLER_19_25
timestamp 1586364061
transform 1 0 3404 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_3.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 3588 0 1 12512
box -38 -48 222 592
use scs8hd_inv_1  mux_right_ipin_3.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 3128 0 1 12512
box -38 -48 314 592
use scs8hd_decap_8  FILLER_20_23
timestamp 1586364061
transform 1 0 3220 0 -1 13600
box -38 -48 774 592
use scs8hd_nor2_4  _120_
timestamp 1586364061
transform 1 0 4784 0 -1 13600
box -38 -48 866 592
use scs8hd_inv_1  mux_left_ipin_0.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 4140 0 1 12512
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_127
timestamp 1586364061
transform 1 0 3956 0 -1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 4600 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__120__B
timestamp 1586364061
transform 1 0 3956 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_29
timestamp 1586364061
transform 1 0 3772 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_36
timestamp 1586364061
transform 1 0 4416 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_40
timestamp 1586364061
transform 1 0 4784 0 1 12512
box -38 -48 222 592
use scs8hd_decap_8  FILLER_20_32
timestamp 1586364061
transform 1 0 4048 0 -1 13600
box -38 -48 774 592
use scs8hd_nor2_4  _039_
timestamp 1586364061
transform 1 0 5152 0 1 12512
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__120__A
timestamp 1586364061
transform 1 0 4968 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__116__A
timestamp 1586364061
transform 1 0 5796 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__116__B
timestamp 1586364061
transform 1 0 6164 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__039__B
timestamp 1586364061
transform 1 0 6164 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_53
timestamp 1586364061
transform 1 0 5980 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_49
timestamp 1586364061
transform 1 0 5612 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_53
timestamp 1586364061
transform 1 0 5980 0 -1 13600
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_ipin_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 6348 0 -1 13600
box -38 -48 866 592
use scs8hd_ebufn_2  mux_left_ipin_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 6992 0 1 12512
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_124
timestamp 1586364061
transform 1 0 6716 0 1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 6532 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_0.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 7360 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_57
timestamp 1586364061
transform 1 0 6348 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_62
timestamp 1586364061
transform 1 0 6808 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_66
timestamp 1586364061
transform 1 0 7176 0 -1 13600
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_ipin_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 8740 0 1 12512
box -38 -48 866 592
use scs8hd_ebufn_2  mux_left_ipin_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 7912 0 -1 13600
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 8004 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 8556 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 7728 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_73
timestamp 1586364061
transform 1 0 7820 0 1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_19_77
timestamp 1586364061
transform 1 0 8188 0 1 12512
box -38 -48 406 592
use scs8hd_fill_2  FILLER_20_70
timestamp 1586364061
transform 1 0 7544 0 -1 13600
box -38 -48 222 592
use scs8hd_decap_8  FILLER_20_83
timestamp 1586364061
transform 1 0 8740 0 -1 13600
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_128
timestamp 1586364061
transform 1 0 9568 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_6  FILLER_19_92
timestamp 1586364061
transform 1 0 9568 0 1 12512
box -38 -48 590 592
use scs8hd_fill_1  FILLER_20_91
timestamp 1586364061
transform 1 0 9476 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_6  FILLER_20_93
timestamp 1586364061
transform 1 0 9660 0 -1 13600
box -38 -48 590 592
use scs8hd_ebufn_2  mux_right_ipin_3.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10304 0 1 12512
box -38 -48 866 592
use scs8hd_ebufn_2  mux_right_ipin_3.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10488 0 -1 13600
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_3.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10120 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_3.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10304 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_109
timestamp 1586364061
transform 1 0 11132 0 1 12512
box -38 -48 222 592
use scs8hd_fill_1  FILLER_20_99
timestamp 1586364061
transform 1 0 10212 0 -1 13600
box -38 -48 130 592
use scs8hd_fill_2  FILLER_20_115
timestamp 1586364061
transform 1 0 11684 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_111
timestamp 1586364061
transform 1 0 11316 0 -1 13600
box -38 -48 222 592
use scs8hd_decap_3  FILLER_19_113
timestamp 1586364061
transform 1 0 11500 0 1 12512
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11868 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_6.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 11776 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 11500 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_3.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 11316 0 1 12512
box -38 -48 222 592
use scs8hd_decap_3  FILLER_19_123
timestamp 1586364061
transform 1 0 12420 0 1 12512
box -38 -48 314 592
use scs8hd_fill_2  FILLER_19_118
timestamp 1586364061
transform 1 0 11960 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_6.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 12144 0 1 12512
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_125
timestamp 1586364061
transform 1 0 12328 0 1 12512
box -38 -48 130 592
use scs8hd_ebufn_2  mux_right_ipin_6.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12052 0 -1 13600
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  mem_right_ipin_6.LATCH_0_.latch
timestamp 1586364061
transform 1 0 12696 0 1 12512
box -38 -48 1050 592
use scs8hd_ebufn_2  mux_right_ipin_6.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 13616 0 -1 13600
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_6.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 13340 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_137
timestamp 1586364061
transform 1 0 13708 0 1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_20_128
timestamp 1586364061
transform 1 0 12880 0 -1 13600
box -38 -48 406 592
use scs8hd_fill_1  FILLER_20_132
timestamp 1586364061
transform 1 0 13248 0 -1 13600
box -38 -48 130 592
use scs8hd_fill_1  FILLER_20_135
timestamp 1586364061
transform 1 0 13524 0 -1 13600
box -38 -48 130 592
use scs8hd_ebufn_2  mux_right_ipin_6.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 14444 0 1 12512
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_6.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 14260 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_6.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 13892 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_141
timestamp 1586364061
transform 1 0 14076 0 1 12512
box -38 -48 222 592
use scs8hd_decap_8  FILLER_20_145
timestamp 1586364061
transform 1 0 14444 0 -1 13600
box -38 -48 774 592
use scs8hd_decap_6  FILLER_20_157
timestamp 1586364061
transform 1 0 15548 0 -1 13600
box -38 -48 590 592
use scs8hd_decap_3  FILLER_19_158
timestamp 1586364061
transform 1 0 15640 0 1 12512
box -38 -48 314 592
use scs8hd_fill_2  FILLER_19_154
timestamp 1586364061
transform 1 0 15272 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_5.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 15456 0 1 12512
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_129
timestamp 1586364061
transform 1 0 15180 0 -1 13600
box -38 -48 130 592
use scs8hd_inv_1  mux_right_ipin_5.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 15272 0 -1 13600
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_1.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 16100 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_1.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 15916 0 1 12512
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_right_ipin_1.LATCH_1_.latch
timestamp 1586364061
transform 1 0 16100 0 1 12512
box -38 -48 1050 592
use scs8hd_lpflow_inputisolatch_1  mem_right_ipin_1.LATCH_0_.latch
timestamp 1586364061
transform 1 0 16284 0 -1 13600
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_1.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 17480 0 -1 13600
box -38 -48 222 592
use scs8hd_decap_6  FILLER_19_174
timestamp 1586364061
transform 1 0 17112 0 1 12512
box -38 -48 590 592
use scs8hd_fill_2  FILLER_20_176
timestamp 1586364061
transform 1 0 17296 0 -1 13600
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_ipin_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18216 0 -1 13600
box -38 -48 866 592
use scs8hd_ebufn_2  mux_right_ipin_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18492 0 1 12512
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_126
timestamp 1586364061
transform 1 0 17940 0 1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 18308 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 17756 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 18032 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_1  FILLER_19_180
timestamp 1586364061
transform 1 0 17664 0 1 12512
box -38 -48 130 592
use scs8hd_decap_3  FILLER_19_184
timestamp 1586364061
transform 1 0 18032 0 1 12512
box -38 -48 314 592
use scs8hd_decap_4  FILLER_20_180
timestamp 1586364061
transform 1 0 17664 0 -1 13600
box -38 -48 406 592
use scs8hd_decap_12  FILLER_19_198
timestamp 1586364061
transform 1 0 19320 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_195
timestamp 1586364061
transform 1 0 19044 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_20_207
timestamp 1586364061
transform 1 0 20148 0 -1 13600
box -38 -48 406 592
use scs8hd_decap_3  PHY_39
timestamp 1586364061
transform -1 0 20884 0 1 12512
box -38 -48 314 592
use scs8hd_decap_3  PHY_41
timestamp 1586364061
transform -1 0 20884 0 -1 13600
box -38 -48 314 592
use scs8hd_fill_2  FILLER_19_210
timestamp 1586364061
transform 1 0 20424 0 1 12512
box -38 -48 222 592
use scs8hd_fill_1  FILLER_20_211
timestamp 1586364061
transform 1 0 20516 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_3  PHY_42
timestamp 1586364061
transform 1 0 1104 0 1 13600
box -38 -48 314 592
use scs8hd_decap_12  FILLER_21_3
timestamp 1586364061
transform 1 0 1380 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_21_15
timestamp 1586364061
transform 1 0 2484 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_21_27
timestamp 1586364061
transform 1 0 3588 0 1 13600
box -38 -48 590 592
use scs8hd_inv_1  mux_left_ipin_0.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 4140 0 1 13600
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_4.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 4600 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_36
timestamp 1586364061
transform 1 0 4416 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_40
timestamp 1586364061
transform 1 0 4784 0 1 13600
box -38 -48 222 592
use scs8hd_nor2_4  _118_
timestamp 1586364061
transform 1 0 5152 0 1 13600
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 4968 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_0.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 6164 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_53
timestamp 1586364061
transform 1 0 5980 0 1 13600
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_left_ipin_0.LATCH_2_.latch
timestamp 1586364061
transform 1 0 6808 0 1 13600
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_130
timestamp 1586364061
transform 1 0 6716 0 1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_0.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 6532 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_57
timestamp 1586364061
transform 1 0 6348 0 1 13600
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_left_ipin_0.LATCH_3_.latch
timestamp 1586364061
transform 1 0 8740 0 1 13600
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_0.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 8556 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_0.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 8004 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_73
timestamp 1586364061
transform 1 0 7820 0 1 13600
box -38 -48 222 592
use scs8hd_decap_4  FILLER_21_77
timestamp 1586364061
transform 1 0 8188 0 1 13600
box -38 -48 406 592
use scs8hd_decap_3  FILLER_21_94
timestamp 1586364061
transform 1 0 9752 0 1 13600
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_right_ipin_3.LATCH_2_.latch
timestamp 1586364061
transform 1 0 10488 0 1 13600
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_6.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 10028 0 1 13600
box -38 -48 222 592
use scs8hd_decap_3  FILLER_21_99
timestamp 1586364061
transform 1 0 10212 0 1 13600
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_right_ipin_6.LATCH_2_.latch
timestamp 1586364061
transform 1 0 12420 0 1 13600
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_131
timestamp 1586364061
transform 1 0 12328 0 1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_6.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 12144 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_3.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 11684 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_113
timestamp 1586364061
transform 1 0 11500 0 1 13600
box -38 -48 222 592
use scs8hd_decap_3  FILLER_21_117
timestamp 1586364061
transform 1 0 11868 0 1 13600
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_6.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 13616 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_134
timestamp 1586364061
transform 1 0 13432 0 1 13600
box -38 -48 222 592
use scs8hd_decap_3  FILLER_21_138
timestamp 1586364061
transform 1 0 13800 0 1 13600
box -38 -48 314 592
use scs8hd_ebufn_2  mux_right_ipin_6.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 14260 0 1 13600
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_6.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 14076 0 1 13600
box -38 -48 222 592
use scs8hd_decap_6  FILLER_21_152
timestamp 1586364061
transform 1 0 15088 0 1 13600
box -38 -48 590 592
use scs8hd_lpflow_inputisolatch_1  mem_right_ipin_1.LATCH_2_.latch
timestamp 1586364061
transform 1 0 16192 0 1 13600
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA__148__A
timestamp 1586364061
transform 1 0 15640 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_1.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 16008 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_160
timestamp 1586364061
transform 1 0 15824 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_1.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 17388 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_175
timestamp 1586364061
transform 1 0 17204 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_179
timestamp 1586364061
transform 1 0 17572 0 1 13600
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_ipin_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18032 0 1 13600
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_132
timestamp 1586364061
transform 1 0 17940 0 1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 17756 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_193
timestamp 1586364061
transform 1 0 18860 0 1 13600
box -38 -48 222 592
use scs8hd_inv_1  mux_right_ipin_5.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 19596 0 1 13600
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 19044 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 19412 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_5.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 20056 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_197
timestamp 1586364061
transform 1 0 19228 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_204
timestamp 1586364061
transform 1 0 19872 0 1 13600
box -38 -48 222 592
use scs8hd_decap_3  PHY_43
timestamp 1586364061
transform -1 0 20884 0 1 13600
box -38 -48 314 592
use scs8hd_decap_4  FILLER_21_208
timestamp 1586364061
transform 1 0 20240 0 1 13600
box -38 -48 406 592
use scs8hd_decap_3  PHY_44
timestamp 1586364061
transform 1 0 1104 0 -1 14688
box -38 -48 314 592
use scs8hd_decap_12  FILLER_22_3
timestamp 1586364061
transform 1 0 1380 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_15
timestamp 1586364061
transform 1 0 2484 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_22_27
timestamp 1586364061
transform 1 0 3588 0 -1 14688
box -38 -48 406 592
use scs8hd_inv_1  mux_right_ipin_4.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 4324 0 -1 14688
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_133
timestamp 1586364061
transform 1 0 3956 0 -1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__118__B
timestamp 1586364061
transform 1 0 4784 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_3  FILLER_22_32
timestamp 1586364061
transform 1 0 4048 0 -1 14688
box -38 -48 314 592
use scs8hd_fill_2  FILLER_22_38
timestamp 1586364061
transform 1 0 4600 0 -1 14688
box -38 -48 222 592
use scs8hd_nor2_4  _116_
timestamp 1586364061
transform 1 0 5336 0 -1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__118__A
timestamp 1586364061
transform 1 0 5152 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_42
timestamp 1586364061
transform 1 0 4968 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_8  FILLER_22_55
timestamp 1586364061
transform 1 0 6164 0 -1 14688
box -38 -48 774 592
use scs8hd_lpflow_inputisolatch_1  mem_left_ipin_0.LATCH_4_.latch
timestamp 1586364061
transform 1 0 6900 0 -1 14688
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_0.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 8740 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_8  FILLER_22_74
timestamp 1586364061
transform 1 0 7912 0 -1 14688
box -38 -48 774 592
use scs8hd_fill_1  FILLER_22_82
timestamp 1586364061
transform 1 0 8648 0 -1 14688
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_134
timestamp 1586364061
transform 1 0 9568 0 -1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_3.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 9844 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_3.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9108 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_85
timestamp 1586364061
transform 1 0 8924 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_3  FILLER_22_89
timestamp 1586364061
transform 1 0 9292 0 -1 14688
box -38 -48 314 592
use scs8hd_fill_2  FILLER_22_93
timestamp 1586364061
transform 1 0 9660 0 -1 14688
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_ipin_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 11040 0 -1 14688
box -38 -48 866 592
use scs8hd_inv_1  mux_right_ipin_6.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 10028 0 -1 14688
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_3.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 10488 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_3.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 10856 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_100
timestamp 1586364061
transform 1 0 10304 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_104
timestamp 1586364061
transform 1 0 10672 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_6.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 12420 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_6  FILLER_22_117
timestamp 1586364061
transform 1 0 11868 0 -1 14688
box -38 -48 590 592
use scs8hd_ebufn_2  mux_right_ipin_6.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 13340 0 -1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_6.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 13156 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_6.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 12788 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_125
timestamp 1586364061
transform 1 0 12604 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_129
timestamp 1586364061
transform 1 0 12972 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_6.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14352 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_6.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14996 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_142
timestamp 1586364061
transform 1 0 14168 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_22_146
timestamp 1586364061
transform 1 0 14536 0 -1 14688
box -38 -48 406 592
use scs8hd_fill_1  FILLER_22_150
timestamp 1586364061
transform 1 0 14904 0 -1 14688
box -38 -48 130 592
use scs8hd_buf_2  _148_
timestamp 1586364061
transform 1 0 15640 0 -1 14688
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_135
timestamp 1586364061
transform 1 0 15180 0 -1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_1.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 16192 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_6.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 15456 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_154
timestamp 1586364061
transform 1 0 15272 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_162
timestamp 1586364061
transform 1 0 16008 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_22_166
timestamp 1586364061
transform 1 0 16376 0 -1 14688
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_right_ipin_1.LATCH_3_.latch
timestamp 1586364061
transform 1 0 16744 0 -1 14688
box -38 -48 1050 592
use scs8hd_ebufn_2  mux_right_ipin_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18492 0 -1 14688
box -38 -48 866 592
use scs8hd_decap_8  FILLER_22_181
timestamp 1586364061
transform 1 0 17756 0 -1 14688
box -38 -48 774 592
use scs8hd_decap_12  FILLER_22_198
timestamp 1586364061
transform 1 0 19320 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_3  PHY_45
timestamp 1586364061
transform -1 0 20884 0 -1 14688
box -38 -48 314 592
use scs8hd_fill_2  FILLER_22_210
timestamp 1586364061
transform 1 0 20424 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_3  PHY_46
timestamp 1586364061
transform 1 0 1104 0 1 14688
box -38 -48 314 592
use scs8hd_decap_12  FILLER_23_3
timestamp 1586364061
transform 1 0 1380 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_15
timestamp 1586364061
transform 1 0 2484 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_27
timestamp 1586364061
transform 1 0 3588 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_23_39
timestamp 1586364061
transform 1 0 4692 0 1 14688
box -38 -48 774 592
use scs8hd_inv_1  mux_left_ipin_0.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 5704 0 1 14688
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 6164 0 1 14688
box -38 -48 222 592
use scs8hd_decap_3  FILLER_23_47
timestamp 1586364061
transform 1 0 5428 0 1 14688
box -38 -48 314 592
use scs8hd_fill_2  FILLER_23_53
timestamp 1586364061
transform 1 0 5980 0 1 14688
box -38 -48 222 592
use scs8hd_nor2_4  _114_
timestamp 1586364061
transform 1 0 6808 0 1 14688
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_136
timestamp 1586364061
transform 1 0 6716 0 1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__114__A
timestamp 1586364061
transform 1 0 6532 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_57
timestamp 1586364061
transform 1 0 6348 0 1 14688
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_ipin_3.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 8464 0 1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_0.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 7820 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_0.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 8188 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_71
timestamp 1586364061
transform 1 0 7636 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_75
timestamp 1586364061
transform 1 0 8004 0 1 14688
box -38 -48 222 592
use scs8hd_fill_1  FILLER_23_79
timestamp 1586364061
transform 1 0 8372 0 1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_3.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 9752 0 1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_23_89
timestamp 1586364061
transform 1 0 9292 0 1 14688
box -38 -48 406 592
use scs8hd_fill_1  FILLER_23_93
timestamp 1586364061
transform 1 0 9660 0 1 14688
box -38 -48 130 592
use scs8hd_fill_1  FILLER_23_96
timestamp 1586364061
transform 1 0 9936 0 1 14688
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  mem_right_ipin_3.LATCH_3_.latch
timestamp 1586364061
transform 1 0 10028 0 1 14688
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_3.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 11224 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_108
timestamp 1586364061
transform 1 0 11040 0 1 14688
box -38 -48 222 592
use scs8hd_inv_1  mux_right_ipin_6.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 12420 0 1 14688
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_137
timestamp 1586364061
transform 1 0 12328 0 1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_3.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 11592 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_3.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11960 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_112
timestamp 1586364061
transform 1 0 11408 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_116
timestamp 1586364061
transform 1 0 11776 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_120
timestamp 1586364061
transform 1 0 12144 0 1 14688
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_right_ipin_6.LATCH_4_.latch
timestamp 1586364061
transform 1 0 13432 0 1 14688
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_6.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 12880 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_6.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 13248 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_126
timestamp 1586364061
transform 1 0 12696 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_130
timestamp 1586364061
transform 1 0 13064 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_6.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 14996 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_6.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 14628 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_145
timestamp 1586364061
transform 1 0 14444 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_149
timestamp 1586364061
transform 1 0 14812 0 1 14688
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_ipin_6.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15180 0 1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_1.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 16284 0 1 14688
box -38 -48 222 592
use scs8hd_decap_3  FILLER_23_162
timestamp 1586364061
transform 1 0 16008 0 1 14688
box -38 -48 314 592
use scs8hd_buf_2  _147_
timestamp 1586364061
transform 1 0 16836 0 1 14688
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__147__A
timestamp 1586364061
transform 1 0 17388 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_1.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 16652 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_167
timestamp 1586364061
transform 1 0 16468 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_175
timestamp 1586364061
transform 1 0 17204 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_179
timestamp 1586364061
transform 1 0 17572 0 1 14688
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_ipin_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18400 0 1 14688
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_138
timestamp 1586364061
transform 1 0 17940 0 1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_1.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 18216 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 17756 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_184
timestamp 1586364061
transform 1 0 18032 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_1.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 19412 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 19780 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_197
timestamp 1586364061
transform 1 0 19228 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_201
timestamp 1586364061
transform 1 0 19596 0 1 14688
box -38 -48 222 592
use scs8hd_decap_6  FILLER_23_205
timestamp 1586364061
transform 1 0 19964 0 1 14688
box -38 -48 590 592
use scs8hd_decap_3  PHY_47
timestamp 1586364061
transform -1 0 20884 0 1 14688
box -38 -48 314 592
use scs8hd_fill_1  FILLER_23_211
timestamp 1586364061
transform 1 0 20516 0 1 14688
box -38 -48 130 592
use scs8hd_decap_3  PHY_48
timestamp 1586364061
transform 1 0 1104 0 -1 15776
box -38 -48 314 592
use scs8hd_decap_12  FILLER_24_3
timestamp 1586364061
transform 1 0 1380 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_15
timestamp 1586364061
transform 1 0 2484 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_24_27
timestamp 1586364061
transform 1 0 3588 0 -1 15776
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_139
timestamp 1586364061
transform 1 0 3956 0 -1 15776
box -38 -48 130 592
use scs8hd_decap_12  FILLER_24_32
timestamp 1586364061
transform 1 0 4048 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_44
timestamp 1586364061
transform 1 0 5152 0 -1 15776
box -38 -48 1142 592
use scs8hd_conb_1  _124_
timestamp 1586364061
transform 1 0 6256 0 -1 15776
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_left_ipin_0.LATCH_5_.latch
timestamp 1586364061
transform 1 0 7268 0 -1 15776
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA__114__B
timestamp 1586364061
transform 1 0 6808 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_3  FILLER_24_59
timestamp 1586364061
transform 1 0 6532 0 -1 15776
box -38 -48 314 592
use scs8hd_decap_3  FILLER_24_64
timestamp 1586364061
transform 1 0 6992 0 -1 15776
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 8464 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_78
timestamp 1586364061
transform 1 0 8280 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_82
timestamp 1586364061
transform 1 0 8648 0 -1 15776
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_right_ipin_3.LATCH_4_.latch
timestamp 1586364061
transform 1 0 9752 0 -1 15776
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_140
timestamp 1586364061
transform 1 0 9568 0 -1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__068__A
timestamp 1586364061
transform 1 0 9384 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_3.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 8832 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_24_86
timestamp 1586364061
transform 1 0 9016 0 -1 15776
box -38 -48 406 592
use scs8hd_fill_1  FILLER_24_93
timestamp 1586364061
transform 1 0 9660 0 -1 15776
box -38 -48 130 592
use scs8hd_decap_8  FILLER_24_105
timestamp 1586364061
transform 1 0 10764 0 -1 15776
box -38 -48 774 592
use scs8hd_ebufn_2  mux_right_ipin_3.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 11500 0 -1 15776
box -38 -48 866 592
use scs8hd_decap_8  FILLER_24_122
timestamp 1586364061
transform 1 0 12328 0 -1 15776
box -38 -48 774 592
use scs8hd_lpflow_inputisolatch_1  mem_right_ipin_6.LATCH_3_.latch
timestamp 1586364061
transform 1 0 13432 0 -1 15776
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA__089__B
timestamp 1586364061
transform 1 0 13156 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_1  FILLER_24_130
timestamp 1586364061
transform 1 0 13064 0 -1 15776
box -38 -48 130 592
use scs8hd_fill_1  FILLER_24_133
timestamp 1586364061
transform 1 0 13340 0 -1 15776
box -38 -48 130 592
use scs8hd_decap_8  FILLER_24_145
timestamp 1586364061
transform 1 0 14444 0 -1 15776
box -38 -48 774 592
use scs8hd_inv_1  mux_right_ipin_6.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 15272 0 -1 15776
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_141
timestamp 1586364061
transform 1 0 15180 0 -1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__079__A
timestamp 1586364061
transform 1 0 15916 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_24_157
timestamp 1586364061
transform 1 0 15548 0 -1 15776
box -38 -48 406 592
use scs8hd_decap_6  FILLER_24_163
timestamp 1586364061
transform 1 0 16100 0 -1 15776
box -38 -48 590 592
use scs8hd_lpflow_inputisolatch_1  mem_right_ipin_1.LATCH_5_.latch
timestamp 1586364061
transform 1 0 16744 0 -1 15776
box -38 -48 1050 592
use scs8hd_fill_1  FILLER_24_169
timestamp 1586364061
transform 1 0 16652 0 -1 15776
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  mem_right_ipin_1.LATCH_4_.latch
timestamp 1586364061
transform 1 0 18492 0 -1 15776
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_1.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 18032 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_3  FILLER_24_181
timestamp 1586364061
transform 1 0 17756 0 -1 15776
box -38 -48 314 592
use scs8hd_decap_3  FILLER_24_186
timestamp 1586364061
transform 1 0 18216 0 -1 15776
box -38 -48 314 592
use scs8hd_decap_12  FILLER_24_200
timestamp 1586364061
transform 1 0 19504 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_3  PHY_49
timestamp 1586364061
transform -1 0 20884 0 -1 15776
box -38 -48 314 592
use scs8hd_buf_2  _151_
timestamp 1586364061
transform 1 0 1380 0 1 15776
box -38 -48 406 592
use scs8hd_decap_3  PHY_50
timestamp 1586364061
transform 1 0 1104 0 1 15776
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__151__A
timestamp 1586364061
transform 1 0 1932 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_7
timestamp 1586364061
transform 1 0 1748 0 1 15776
box -38 -48 222 592
use scs8hd_decap_12  FILLER_25_11
timestamp 1586364061
transform 1 0 2116 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_23
timestamp 1586364061
transform 1 0 3220 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_35
timestamp 1586364061
transform 1 0 4324 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_47
timestamp 1586364061
transform 1 0 5428 0 1 15776
box -38 -48 1142 592
use scs8hd_inv_1  mux_right_ipin_4.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 6900 0 1 15776
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_142
timestamp 1586364061
transform 1 0 6716 0 1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_4.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 7360 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_59
timestamp 1586364061
transform 1 0 6532 0 1 15776
box -38 -48 222 592
use scs8hd_fill_1  FILLER_25_62
timestamp 1586364061
transform 1 0 6808 0 1 15776
box -38 -48 130 592
use scs8hd_fill_2  FILLER_25_66
timestamp 1586364061
transform 1 0 7176 0 1 15776
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_ipin_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 7912 0 1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__066__B
timestamp 1586364061
transform 1 0 7728 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_70
timestamp 1586364061
transform 1 0 7544 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_83
timestamp 1586364061
transform 1 0 8740 0 1 15776
box -38 -48 222 592
use scs8hd_inv_1  mux_right_ipin_3.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 9568 0 1 15776
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__068__B
timestamp 1586364061
transform 1 0 9384 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__066__A
timestamp 1586364061
transform 1 0 8924 0 1 15776
box -38 -48 222 592
use scs8hd_decap_3  FILLER_25_87
timestamp 1586364061
transform 1 0 9108 0 1 15776
box -38 -48 314 592
use scs8hd_fill_2  FILLER_25_95
timestamp 1586364061
transform 1 0 9844 0 1 15776
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_right_ipin_3.LATCH_5_.latch
timestamp 1586364061
transform 1 0 10580 0 1 15776
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_3.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 10028 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_3.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 10396 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_99
timestamp 1586364061
transform 1 0 10212 0 1 15776
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_143
timestamp 1586364061
transform 1 0 12328 0 1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_3.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11776 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_3.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 12144 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_114
timestamp 1586364061
transform 1 0 11592 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_118
timestamp 1586364061
transform 1 0 11960 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_123
timestamp 1586364061
transform 1 0 12420 0 1 15776
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_right_ipin_6.LATCH_5_.latch
timestamp 1586364061
transform 1 0 13156 0 1 15776
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_6.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 12972 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__089__A
timestamp 1586364061
transform 1 0 12604 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_127
timestamp 1586364061
transform 1 0 12788 0 1 15776
box -38 -48 222 592
use scs8hd_conb_1  _132_
timestamp 1586364061
transform 1 0 14904 0 1 15776
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__087__A
timestamp 1586364061
transform 1 0 14720 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_6.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 14352 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_142
timestamp 1586364061
transform 1 0 14168 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_146
timestamp 1586364061
transform 1 0 14536 0 1 15776
box -38 -48 222 592
use scs8hd_nor2_4  _079_
timestamp 1586364061
transform 1 0 15916 0 1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__079__B
timestamp 1586364061
transform 1 0 15732 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__087__B
timestamp 1586364061
transform 1 0 15364 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_153
timestamp 1586364061
transform 1 0 15180 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_157
timestamp 1586364061
transform 1 0 15548 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 17388 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 17020 0 1 15776
box -38 -48 222 592
use scs8hd_decap_3  FILLER_25_170
timestamp 1586364061
transform 1 0 16744 0 1 15776
box -38 -48 314 592
use scs8hd_fill_2  FILLER_25_175
timestamp 1586364061
transform 1 0 17204 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_179
timestamp 1586364061
transform 1 0 17572 0 1 15776
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_ipin_1.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18032 0 1 15776
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_144
timestamp 1586364061
transform 1 0 17940 0 1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_1.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 17756 0 1 15776
box -38 -48 222 592
use scs8hd_decap_6  FILLER_25_193
timestamp 1586364061
transform 1 0 18860 0 1 15776
box -38 -48 590 592
use scs8hd_inv_1  mux_right_ipin_1.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 19596 0 1 15776
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__144__A
timestamp 1586364061
transform 1 0 19412 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_1.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 20056 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_204
timestamp 1586364061
transform 1 0 19872 0 1 15776
box -38 -48 222 592
use scs8hd_decap_3  PHY_51
timestamp 1586364061
transform -1 0 20884 0 1 15776
box -38 -48 314 592
use scs8hd_decap_4  FILLER_25_208
timestamp 1586364061
transform 1 0 20240 0 1 15776
box -38 -48 406 592
use scs8hd_decap_3  PHY_52
timestamp 1586364061
transform 1 0 1104 0 -1 16864
box -38 -48 314 592
use scs8hd_decap_3  PHY_54
timestamp 1586364061
transform 1 0 1104 0 1 16864
box -38 -48 314 592
use scs8hd_decap_12  FILLER_26_3
timestamp 1586364061
transform 1 0 1380 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_3
timestamp 1586364061
transform 1 0 1380 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_26_15
timestamp 1586364061
transform 1 0 2484 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_26_27
timestamp 1586364061
transform 1 0 3588 0 -1 16864
box -38 -48 406 592
use scs8hd_decap_12  FILLER_27_15
timestamp 1586364061
transform 1 0 2484 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_27
timestamp 1586364061
transform 1 0 3588 0 1 16864
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_145
timestamp 1586364061
transform 1 0 3956 0 -1 16864
box -38 -48 130 592
use scs8hd_decap_12  FILLER_26_32
timestamp 1586364061
transform 1 0 4048 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_39
timestamp 1586364061
transform 1 0 4692 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_26_44
timestamp 1586364061
transform 1 0 5152 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_27_51
timestamp 1586364061
transform 1 0 5796 0 1 16864
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_148
timestamp 1586364061
transform 1 0 6716 0 1 16864
box -38 -48 130 592
use scs8hd_decap_12  FILLER_26_56
timestamp 1586364061
transform 1 0 6256 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_26_68
timestamp 1586364061
transform 1 0 7360 0 -1 16864
box -38 -48 406 592
use scs8hd_fill_2  FILLER_27_59
timestamp 1586364061
transform 1 0 6532 0 1 16864
box -38 -48 222 592
use scs8hd_decap_12  FILLER_27_62
timestamp 1586364061
transform 1 0 6808 0 1 16864
box -38 -48 1142 592
use scs8hd_nor2_4  _066_
timestamp 1586364061
transform 1 0 8004 0 -1 16864
box -38 -48 866 592
use scs8hd_inv_1  mux_left_ipin_0.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 8372 0 1 16864
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 7820 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_1  FILLER_26_72
timestamp 1586364061
transform 1 0 7728 0 -1 16864
box -38 -48 130 592
use scs8hd_decap_4  FILLER_27_74
timestamp 1586364061
transform 1 0 7912 0 1 16864
box -38 -48 406 592
use scs8hd_fill_1  FILLER_27_78
timestamp 1586364061
transform 1 0 8280 0 1 16864
box -38 -48 130 592
use scs8hd_fill_2  FILLER_27_82
timestamp 1586364061
transform 1 0 8648 0 1 16864
box -38 -48 222 592
use scs8hd_nor2_4  _067_
timestamp 1586364061
transform 1 0 9384 0 1 16864
box -38 -48 866 592
use scs8hd_nor2_4  _068_
timestamp 1586364061
transform 1 0 9660 0 -1 16864
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_146
timestamp 1586364061
transform 1 0 9568 0 -1 16864
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__067__B
timestamp 1586364061
transform 1 0 9200 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__067__A
timestamp 1586364061
transform 1 0 9384 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 8832 0 1 16864
box -38 -48 222 592
use scs8hd_decap_6  FILLER_26_84
timestamp 1586364061
transform 1 0 8832 0 -1 16864
box -38 -48 590 592
use scs8hd_fill_2  FILLER_27_86
timestamp 1586364061
transform 1 0 9016 0 1 16864
box -38 -48 222 592
use scs8hd_conb_1  _129_
timestamp 1586364061
transform 1 0 11040 0 1 16864
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__065__B
timestamp 1586364061
transform 1 0 10396 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__065__A
timestamp 1586364061
transform 1 0 10764 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_3.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 10672 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_102
timestamp 1586364061
transform 1 0 10488 0 -1 16864
box -38 -48 222 592
use scs8hd_decap_8  FILLER_26_106
timestamp 1586364061
transform 1 0 10856 0 -1 16864
box -38 -48 774 592
use scs8hd_fill_2  FILLER_27_99
timestamp 1586364061
transform 1 0 10212 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_103
timestamp 1586364061
transform 1 0 10580 0 1 16864
box -38 -48 222 592
use scs8hd_fill_1  FILLER_27_107
timestamp 1586364061
transform 1 0 10948 0 1 16864
box -38 -48 130 592
use scs8hd_nor2_4  _091_
timestamp 1586364061
transform 1 0 12420 0 1 16864
box -38 -48 866 592
use scs8hd_ebufn_2  mux_right_ipin_3.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 11592 0 -1 16864
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_149
timestamp 1586364061
transform 1 0 12328 0 1 16864
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__091__B
timestamp 1586364061
transform 1 0 12144 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_123
timestamp 1586364061
transform 1 0 12420 0 -1 16864
box -38 -48 222 592
use scs8hd_decap_8  FILLER_27_111
timestamp 1586364061
transform 1 0 11316 0 1 16864
box -38 -48 774 592
use scs8hd_fill_1  FILLER_27_119
timestamp 1586364061
transform 1 0 12052 0 1 16864
box -38 -48 130 592
use scs8hd_nor2_4  _089_
timestamp 1586364061
transform 1 0 13156 0 -1 16864
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__088__B
timestamp 1586364061
transform 1 0 13432 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__088__A
timestamp 1586364061
transform 1 0 12604 0 -1 16864
box -38 -48 222 592
use scs8hd_decap_4  FILLER_26_127
timestamp 1586364061
transform 1 0 12788 0 -1 16864
box -38 -48 406 592
use scs8hd_fill_2  FILLER_27_132
timestamp 1586364061
transform 1 0 13248 0 1 16864
box -38 -48 222 592
use scs8hd_decap_4  FILLER_27_136
timestamp 1586364061
transform 1 0 13616 0 1 16864
box -38 -48 406 592
use scs8hd_fill_1  FILLER_27_140
timestamp 1586364061
transform 1 0 13984 0 1 16864
box -38 -48 130 592
use scs8hd_fill_2  FILLER_26_145
timestamp 1586364061
transform 1 0 14444 0 -1 16864
box -38 -48 222 592
use scs8hd_decap_3  FILLER_26_140
timestamp 1586364061
transform 1 0 13984 0 -1 16864
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_6.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14260 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_6.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 14076 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_152
timestamp 1586364061
transform 1 0 15088 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_149
timestamp 1586364061
transform 1 0 14812 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_6.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 14628 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__083__A
timestamp 1586364061
transform 1 0 14996 0 -1 16864
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_ipin_6.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 14260 0 1 16864
box -38 -48 866 592
use scs8hd_nor2_4  _049_
timestamp 1586364061
transform 1 0 15824 0 1 16864
box -38 -48 866 592
use scs8hd_nor2_4  _087_
timestamp 1586364061
transform 1 0 15272 0 -1 16864
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_147
timestamp 1586364061
transform 1 0 15180 0 -1 16864
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__049__B
timestamp 1586364061
transform 1 0 15640 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__083__B
timestamp 1586364061
transform 1 0 15272 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__049__A
timestamp 1586364061
transform 1 0 16284 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_163
timestamp 1586364061
transform 1 0 16100 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_156
timestamp 1586364061
transform 1 0 15456 0 1 16864
box -38 -48 222 592
use scs8hd_conb_1  _127_
timestamp 1586364061
transform 1 0 16836 0 -1 16864
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__053__B
timestamp 1586364061
transform 1 0 16836 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__053__A
timestamp 1586364061
transform 1 0 17204 0 1 16864
box -38 -48 222 592
use scs8hd_decap_4  FILLER_26_167
timestamp 1586364061
transform 1 0 16468 0 -1 16864
box -38 -48 406 592
use scs8hd_decap_8  FILLER_26_174
timestamp 1586364061
transform 1 0 17112 0 -1 16864
box -38 -48 774 592
use scs8hd_fill_2  FILLER_27_169
timestamp 1586364061
transform 1 0 16652 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_173
timestamp 1586364061
transform 1 0 17020 0 1 16864
box -38 -48 222 592
use scs8hd_decap_4  FILLER_27_177
timestamp 1586364061
transform 1 0 17388 0 1 16864
box -38 -48 406 592
use scs8hd_nor2_4  _052_
timestamp 1586364061
transform 1 0 18032 0 1 16864
box -38 -48 866 592
use scs8hd_ebufn_2  mux_right_ipin_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 17848 0 -1 16864
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_150
timestamp 1586364061
transform 1 0 17940 0 1 16864
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__052__B
timestamp 1586364061
transform 1 0 17756 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__050__A
timestamp 1586364061
transform 1 0 18860 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_191
timestamp 1586364061
transform 1 0 18676 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_193
timestamp 1586364061
transform 1 0 18860 0 1 16864
box -38 -48 222 592
use scs8hd_buf_2  _144_
timestamp 1586364061
transform 1 0 19412 0 -1 16864
box -38 -48 406 592
use scs8hd_inv_1  mux_right_ipin_1.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 19596 0 1 16864
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_1.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 20056 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__050__B
timestamp 1586364061
transform 1 0 19044 0 1 16864
box -38 -48 222 592
use scs8hd_decap_4  FILLER_26_195
timestamp 1586364061
transform 1 0 19044 0 -1 16864
box -38 -48 406 592
use scs8hd_decap_8  FILLER_26_203
timestamp 1586364061
transform 1 0 19780 0 -1 16864
box -38 -48 774 592
use scs8hd_decap_4  FILLER_27_197
timestamp 1586364061
transform 1 0 19228 0 1 16864
box -38 -48 406 592
use scs8hd_fill_2  FILLER_27_204
timestamp 1586364061
transform 1 0 19872 0 1 16864
box -38 -48 222 592
use scs8hd_decap_3  PHY_53
timestamp 1586364061
transform -1 0 20884 0 -1 16864
box -38 -48 314 592
use scs8hd_decap_3  PHY_55
timestamp 1586364061
transform -1 0 20884 0 1 16864
box -38 -48 314 592
use scs8hd_fill_1  FILLER_26_211
timestamp 1586364061
transform 1 0 20516 0 -1 16864
box -38 -48 130 592
use scs8hd_decap_4  FILLER_27_208
timestamp 1586364061
transform 1 0 20240 0 1 16864
box -38 -48 406 592
use scs8hd_decap_3  PHY_56
timestamp 1586364061
transform 1 0 1104 0 -1 17952
box -38 -48 314 592
use scs8hd_decap_12  FILLER_28_3
timestamp 1586364061
transform 1 0 1380 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_15
timestamp 1586364061
transform 1 0 2484 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_28_27
timestamp 1586364061
transform 1 0 3588 0 -1 17952
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_151
timestamp 1586364061
transform 1 0 3956 0 -1 17952
box -38 -48 130 592
use scs8hd_decap_12  FILLER_28_32
timestamp 1586364061
transform 1 0 4048 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_44
timestamp 1586364061
transform 1 0 5152 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_56
timestamp 1586364061
transform 1 0 6256 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_68
timestamp 1586364061
transform 1 0 7360 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_80
timestamp 1586364061
transform 1 0 8464 0 -1 17952
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_152
timestamp 1586364061
transform 1 0 9568 0 -1 17952
box -38 -48 130 592
use scs8hd_decap_6  FILLER_28_93
timestamp 1586364061
transform 1 0 9660 0 -1 17952
box -38 -48 590 592
use scs8hd_nor2_4  _065_
timestamp 1586364061
transform 1 0 10212 0 -1 17952
box -38 -48 866 592
use scs8hd_decap_12  FILLER_28_108
timestamp 1586364061
transform 1 0 11040 0 -1 17952
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA__091__A
timestamp 1586364061
transform 1 0 12420 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_3  FILLER_28_120
timestamp 1586364061
transform 1 0 12144 0 -1 17952
box -38 -48 314 592
use scs8hd_nor2_4  _088_
timestamp 1586364061
transform 1 0 12604 0 -1 17952
box -38 -48 866 592
use scs8hd_decap_8  FILLER_28_134
timestamp 1586364061
transform 1 0 13432 0 -1 17952
box -38 -48 774 592
use scs8hd_inv_1  mux_right_ipin_6.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 14168 0 -1 17952
box -38 -48 314 592
use scs8hd_decap_8  FILLER_28_145
timestamp 1586364061
transform 1 0 14444 0 -1 17952
box -38 -48 774 592
use scs8hd_nor2_4  _083_
timestamp 1586364061
transform 1 0 15272 0 -1 17952
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_153
timestamp 1586364061
transform 1 0 15180 0 -1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__051__A
timestamp 1586364061
transform 1 0 16284 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_163
timestamp 1586364061
transform 1 0 16100 0 -1 17952
box -38 -48 222 592
use scs8hd_nor2_4  _053_
timestamp 1586364061
transform 1 0 16836 0 -1 17952
box -38 -48 866 592
use scs8hd_decap_4  FILLER_28_167
timestamp 1586364061
transform 1 0 16468 0 -1 17952
box -38 -48 406 592
use scs8hd_nor2_4  _050_
timestamp 1586364061
transform 1 0 18400 0 -1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__052__A
timestamp 1586364061
transform 1 0 18032 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_4  FILLER_28_180
timestamp 1586364061
transform 1 0 17664 0 -1 17952
box -38 -48 406 592
use scs8hd_fill_2  FILLER_28_186
timestamp 1586364061
transform 1 0 18216 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_12  FILLER_28_197
timestamp 1586364061
transform 1 0 19228 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_3  PHY_57
timestamp 1586364061
transform -1 0 20884 0 -1 17952
box -38 -48 314 592
use scs8hd_decap_3  FILLER_28_209
timestamp 1586364061
transform 1 0 20332 0 -1 17952
box -38 -48 314 592
use scs8hd_buf_2  _146_
timestamp 1586364061
transform 1 0 1380 0 1 17952
box -38 -48 406 592
use scs8hd_decap_3  PHY_58
timestamp 1586364061
transform 1 0 1104 0 1 17952
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__146__A
timestamp 1586364061
transform 1 0 1932 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_7
timestamp 1586364061
transform 1 0 1748 0 1 17952
box -38 -48 222 592
use scs8hd_decap_12  FILLER_29_11
timestamp 1586364061
transform 1 0 2116 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_23
timestamp 1586364061
transform 1 0 3220 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_35
timestamp 1586364061
transform 1 0 4324 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_47
timestamp 1586364061
transform 1 0 5428 0 1 17952
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_154
timestamp 1586364061
transform 1 0 6716 0 1 17952
box -38 -48 130 592
use scs8hd_fill_2  FILLER_29_59
timestamp 1586364061
transform 1 0 6532 0 1 17952
box -38 -48 222 592
use scs8hd_decap_12  FILLER_29_62
timestamp 1586364061
transform 1 0 6808 0 1 17952
box -38 -48 1142 592
use scs8hd_buf_2  _137_
timestamp 1586364061
transform 1 0 7912 0 1 17952
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__137__A
timestamp 1586364061
transform 1 0 8464 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_78
timestamp 1586364061
transform 1 0 8280 0 1 17952
box -38 -48 222 592
use scs8hd_decap_12  FILLER_29_82
timestamp 1586364061
transform 1 0 8648 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_29_94
timestamp 1586364061
transform 1 0 9752 0 1 17952
box -38 -48 590 592
use scs8hd_inv_1  mux_right_ipin_3.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 10396 0 1 17952
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_3.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 10856 0 1 17952
box -38 -48 222 592
use scs8hd_fill_1  FILLER_29_100
timestamp 1586364061
transform 1 0 10304 0 1 17952
box -38 -48 130 592
use scs8hd_fill_2  FILLER_29_104
timestamp 1586364061
transform 1 0 10672 0 1 17952
box -38 -48 222 592
use scs8hd_decap_8  FILLER_29_108
timestamp 1586364061
transform 1 0 11040 0 1 17952
box -38 -48 774 592
use scs8hd_nor2_4  _086_
timestamp 1586364061
transform 1 0 12512 0 1 17952
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_155
timestamp 1586364061
transform 1 0 12328 0 1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__086__B
timestamp 1586364061
transform 1 0 12144 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_3.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 11776 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_118
timestamp 1586364061
transform 1 0 11960 0 1 17952
box -38 -48 222 592
use scs8hd_fill_1  FILLER_29_123
timestamp 1586364061
transform 1 0 12420 0 1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 13524 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_133
timestamp 1586364061
transform 1 0 13340 0 1 17952
box -38 -48 222 592
use scs8hd_decap_4  FILLER_29_137
timestamp 1586364061
transform 1 0 13708 0 1 17952
box -38 -48 406 592
use scs8hd_buf_2  _150_
timestamp 1586364061
transform 1 0 14352 0 1 17952
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__150__A
timestamp 1586364061
transform 1 0 14904 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_7.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 14168 0 1 17952
box -38 -48 222 592
use scs8hd_fill_1  FILLER_29_141
timestamp 1586364061
transform 1 0 14076 0 1 17952
box -38 -48 130 592
use scs8hd_fill_2  FILLER_29_148
timestamp 1586364061
transform 1 0 14720 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_152
timestamp 1586364061
transform 1 0 15088 0 1 17952
box -38 -48 222 592
use scs8hd_nor2_4  _054_
timestamp 1586364061
transform 1 0 15456 0 1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__054__B
timestamp 1586364061
transform 1 0 15272 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_165
timestamp 1586364061
transform 1 0 16284 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_1.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 17572 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__051__B
timestamp 1586364061
transform 1 0 16468 0 1 17952
box -38 -48 222 592
use scs8hd_decap_8  FILLER_29_169
timestamp 1586364061
transform 1 0 16652 0 1 17952
box -38 -48 774 592
use scs8hd_fill_2  FILLER_29_177
timestamp 1586364061
transform 1 0 17388 0 1 17952
box -38 -48 222 592
use scs8hd_buf_2  _145_
timestamp 1586364061
transform 1 0 18032 0 1 17952
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_156
timestamp 1586364061
transform 1 0 17940 0 1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__145__A
timestamp 1586364061
transform 1 0 18584 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_181
timestamp 1586364061
transform 1 0 17756 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_188
timestamp 1586364061
transform 1 0 18400 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_192
timestamp 1586364061
transform 1 0 18768 0 1 17952
box -38 -48 222 592
use scs8hd_inv_1  mux_right_ipin_1.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 19136 0 1 17952
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_1.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 19596 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_1.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 18952 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_1.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 19964 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_199
timestamp 1586364061
transform 1 0 19412 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_203
timestamp 1586364061
transform 1 0 19780 0 1 17952
box -38 -48 222 592
use scs8hd_decap_4  FILLER_29_207
timestamp 1586364061
transform 1 0 20148 0 1 17952
box -38 -48 406 592
use scs8hd_decap_3  PHY_59
timestamp 1586364061
transform -1 0 20884 0 1 17952
box -38 -48 314 592
use scs8hd_fill_1  FILLER_29_211
timestamp 1586364061
transform 1 0 20516 0 1 17952
box -38 -48 130 592
use scs8hd_decap_3  PHY_60
timestamp 1586364061
transform 1 0 1104 0 -1 19040
box -38 -48 314 592
use scs8hd_decap_12  FILLER_30_3
timestamp 1586364061
transform 1 0 1380 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_15
timestamp 1586364061
transform 1 0 2484 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_30_27
timestamp 1586364061
transform 1 0 3588 0 -1 19040
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_157
timestamp 1586364061
transform 1 0 3956 0 -1 19040
box -38 -48 130 592
use scs8hd_decap_12  FILLER_30_32
timestamp 1586364061
transform 1 0 4048 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_44
timestamp 1586364061
transform 1 0 5152 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_56
timestamp 1586364061
transform 1 0 6256 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_68
timestamp 1586364061
transform 1 0 7360 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_80
timestamp 1586364061
transform 1 0 8464 0 -1 19040
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_158
timestamp 1586364061
transform 1 0 9568 0 -1 19040
box -38 -48 130 592
use scs8hd_decap_12  FILLER_30_93
timestamp 1586364061
transform 1 0 9660 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_105
timestamp 1586364061
transform 1 0 10764 0 -1 19040
box -38 -48 1142 592
use scs8hd_inv_1  mux_right_ipin_3.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 12144 0 -1 19040
box -38 -48 314 592
use scs8hd_decap_3  FILLER_30_117
timestamp 1586364061
transform 1 0 11868 0 -1 19040
box -38 -48 314 592
use scs8hd_fill_2  FILLER_30_123
timestamp 1586364061
transform 1 0 12420 0 -1 19040
box -38 -48 222 592
use scs8hd_inv_1  mux_right_ipin_0.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 13156 0 -1 19040
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__086__A
timestamp 1586364061
transform 1 0 12604 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_4  FILLER_30_127
timestamp 1586364061
transform 1 0 12788 0 -1 19040
box -38 -48 406 592
use scs8hd_decap_8  FILLER_30_134
timestamp 1586364061
transform 1 0 13432 0 -1 19040
box -38 -48 774 592
use scs8hd_inv_1  mux_right_ipin_7.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 14168 0 -1 19040
box -38 -48 314 592
use scs8hd_decap_8  FILLER_30_145
timestamp 1586364061
transform 1 0 14444 0 -1 19040
box -38 -48 774 592
use scs8hd_nor2_4  _051_
timestamp 1586364061
transform 1 0 15732 0 -1 19040
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_159
timestamp 1586364061
transform 1 0 15180 0 -1 19040
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__054__A
timestamp 1586364061
transform 1 0 15456 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_154
timestamp 1586364061
transform 1 0 15272 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_1  FILLER_30_158
timestamp 1586364061
transform 1 0 15640 0 -1 19040
box -38 -48 130 592
use scs8hd_inv_1  mux_right_ipin_1.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 17572 0 -1 19040
box -38 -48 314 592
use scs8hd_decap_8  FILLER_30_168
timestamp 1586364061
transform 1 0 16560 0 -1 19040
box -38 -48 774 592
use scs8hd_decap_3  FILLER_30_176
timestamp 1586364061
transform 1 0 17296 0 -1 19040
box -38 -48 314 592
use scs8hd_inv_1  mux_right_ipin_1.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 18584 0 -1 19040
box -38 -48 314 592
use scs8hd_decap_8  FILLER_30_182
timestamp 1586364061
transform 1 0 17848 0 -1 19040
box -38 -48 774 592
use scs8hd_decap_8  FILLER_30_193
timestamp 1586364061
transform 1 0 18860 0 -1 19040
box -38 -48 774 592
use scs8hd_inv_1  mux_right_ipin_1.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 19596 0 -1 19040
box -38 -48 314 592
use scs8hd_decap_8  FILLER_30_204
timestamp 1586364061
transform 1 0 19872 0 -1 19040
box -38 -48 774 592
use scs8hd_decap_3  PHY_61
timestamp 1586364061
transform -1 0 20884 0 -1 19040
box -38 -48 314 592
use scs8hd_decap_3  PHY_62
timestamp 1586364061
transform 1 0 1104 0 1 19040
box -38 -48 314 592
use scs8hd_decap_12  FILLER_31_3
timestamp 1586364061
transform 1 0 1380 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_15
timestamp 1586364061
transform 1 0 2484 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_31_27
timestamp 1586364061
transform 1 0 3588 0 1 19040
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_160
timestamp 1586364061
transform 1 0 3956 0 1 19040
box -38 -48 130 592
use scs8hd_decap_12  FILLER_31_32
timestamp 1586364061
transform 1 0 4048 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_44
timestamp 1586364061
transform 1 0 5152 0 1 19040
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_161
timestamp 1586364061
transform 1 0 6808 0 1 19040
box -38 -48 130 592
use scs8hd_decap_6  FILLER_31_56
timestamp 1586364061
transform 1 0 6256 0 1 19040
box -38 -48 590 592
use scs8hd_decap_12  FILLER_31_63
timestamp 1586364061
transform 1 0 6900 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_75
timestamp 1586364061
transform 1 0 8004 0 1 19040
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_162
timestamp 1586364061
transform 1 0 9660 0 1 19040
box -38 -48 130 592
use scs8hd_decap_6  FILLER_31_87
timestamp 1586364061
transform 1 0 9108 0 1 19040
box -38 -48 590 592
use scs8hd_decap_12  FILLER_31_94
timestamp 1586364061
transform 1 0 9752 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_106
timestamp 1586364061
transform 1 0 10856 0 1 19040
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_163
timestamp 1586364061
transform 1 0 12512 0 1 19040
box -38 -48 130 592
use scs8hd_decap_6  FILLER_31_118
timestamp 1586364061
transform 1 0 11960 0 1 19040
box -38 -48 590 592
use scs8hd_inv_1  mux_right_ipin_0.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 13340 0 1 19040
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 13800 0 1 19040
box -38 -48 222 592
use scs8hd_decap_8  FILLER_31_125
timestamp 1586364061
transform 1 0 12604 0 1 19040
box -38 -48 774 592
use scs8hd_fill_2  FILLER_31_136
timestamp 1586364061
transform 1 0 13616 0 1 19040
box -38 -48 222 592
use scs8hd_inv_1  mux_right_ipin_0.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 14352 0 1 19040
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 14812 0 1 19040
box -38 -48 222 592
use scs8hd_decap_4  FILLER_31_140
timestamp 1586364061
transform 1 0 13984 0 1 19040
box -38 -48 406 592
use scs8hd_fill_2  FILLER_31_147
timestamp 1586364061
transform 1 0 14628 0 1 19040
box -38 -48 222 592
use scs8hd_decap_4  FILLER_31_151
timestamp 1586364061
transform 1 0 14996 0 1 19040
box -38 -48 406 592
use scs8hd_inv_1  mux_right_ipin_6.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 15456 0 1 19040
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_164
timestamp 1586364061
transform 1 0 15364 0 1 19040
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_6.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 15916 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_159
timestamp 1586364061
transform 1 0 15732 0 1 19040
box -38 -48 222 592
use scs8hd_decap_12  FILLER_31_163
timestamp 1586364061
transform 1 0 16100 0 1 19040
box -38 -48 1142 592
use scs8hd_inv_1  mux_right_ipin_5.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 17204 0 1 19040
box -38 -48 314 592
use scs8hd_fill_2  FILLER_31_178
timestamp 1586364061
transform 1 0 17480 0 1 19040
box -38 -48 222 592
use scs8hd_inv_1  mux_right_ipin_1.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 18308 0 1 19040
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_165
timestamp 1586364061
transform 1 0 18216 0 1 19040
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_5.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 17664 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_1.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 18768 0 1 19040
box -38 -48 222 592
use scs8hd_decap_4  FILLER_31_182
timestamp 1586364061
transform 1 0 17848 0 1 19040
box -38 -48 406 592
use scs8hd_fill_2  FILLER_31_190
timestamp 1586364061
transform 1 0 18584 0 1 19040
box -38 -48 222 592
use scs8hd_inv_1  mux_left_ipin_1.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 19320 0 1 19040
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_1.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 19780 0 1 19040
box -38 -48 222 592
use scs8hd_decap_4  FILLER_31_194
timestamp 1586364061
transform 1 0 18952 0 1 19040
box -38 -48 406 592
use scs8hd_fill_2  FILLER_31_201
timestamp 1586364061
transform 1 0 19596 0 1 19040
box -38 -48 222 592
use scs8hd_decap_6  FILLER_31_205
timestamp 1586364061
transform 1 0 19964 0 1 19040
box -38 -48 590 592
use scs8hd_decap_3  PHY_63
timestamp 1586364061
transform -1 0 20884 0 1 19040
box -38 -48 314 592
use scs8hd_fill_1  FILLER_31_211
timestamp 1586364061
transform 1 0 20516 0 1 19040
box -38 -48 130 592
<< labels >>
rlabel metal3 s 21520 416 22000 536 6 address[0]
port 0 nsew default input
rlabel metal3 s 21520 1368 22000 1488 6 address[1]
port 1 nsew default input
rlabel metal3 s 0 824 480 944 6 address[2]
port 2 nsew default input
rlabel metal3 s 21520 2320 22000 2440 6 address[3]
port 3 nsew default input
rlabel metal3 s 21520 3272 22000 3392 6 address[4]
port 4 nsew default input
rlabel metal3 s 0 2592 480 2712 6 address[5]
port 5 nsew default input
rlabel metal3 s 21520 4224 22000 4344 6 address[6]
port 6 nsew default input
rlabel metal2 s 4894 0 4950 480 6 chany_bottom_in[0]
port 7 nsew default input
rlabel metal2 s 1214 21520 1270 22000 6 chany_bottom_in[1]
port 8 nsew default input
rlabel metal3 s 0 4496 480 4616 6 chany_bottom_in[2]
port 9 nsew default input
rlabel metal3 s 0 6264 480 6384 6 chany_bottom_in[3]
port 10 nsew default input
rlabel metal3 s 0 8168 480 8288 6 chany_bottom_in[4]
port 11 nsew default input
rlabel metal2 s 3606 21520 3662 22000 6 chany_bottom_in[5]
port 12 nsew default input
rlabel metal3 s 21520 5176 22000 5296 6 chany_bottom_in[6]
port 13 nsew default input
rlabel metal2 s 6090 21520 6146 22000 6 chany_bottom_in[7]
port 14 nsew default input
rlabel metal2 s 6918 0 6974 480 6 chany_bottom_in[8]
port 15 nsew default input
rlabel metal3 s 21520 6128 22000 6248 6 chany_bottom_out[0]
port 16 nsew default tristate
rlabel metal3 s 0 9936 480 10056 6 chany_bottom_out[1]
port 17 nsew default tristate
rlabel metal3 s 21520 7080 22000 7200 6 chany_bottom_out[2]
port 18 nsew default tristate
rlabel metal3 s 21520 8032 22000 8152 6 chany_bottom_out[3]
port 19 nsew default tristate
rlabel metal3 s 21520 8984 22000 9104 6 chany_bottom_out[4]
port 20 nsew default tristate
rlabel metal2 s 8482 21520 8538 22000 6 chany_bottom_out[5]
port 21 nsew default tristate
rlabel metal3 s 21520 9936 22000 10056 6 chany_bottom_out[6]
port 22 nsew default tristate
rlabel metal3 s 21520 10888 22000 11008 6 chany_bottom_out[7]
port 23 nsew default tristate
rlabel metal3 s 0 11840 480 11960 6 chany_bottom_out[8]
port 24 nsew default tristate
rlabel metal3 s 21520 11840 22000 11960 6 chany_top_in[0]
port 25 nsew default input
rlabel metal3 s 0 13608 480 13728 6 chany_top_in[1]
port 26 nsew default input
rlabel metal3 s 0 15512 480 15632 6 chany_top_in[2]
port 27 nsew default input
rlabel metal2 s 10966 21520 11022 22000 6 chany_top_in[3]
port 28 nsew default input
rlabel metal2 s 8850 0 8906 480 6 chany_top_in[4]
port 29 nsew default input
rlabel metal2 s 10874 0 10930 480 6 chany_top_in[5]
port 30 nsew default input
rlabel metal3 s 21520 12792 22000 12912 6 chany_top_in[6]
port 31 nsew default input
rlabel metal3 s 21520 13744 22000 13864 6 chany_top_in[7]
port 32 nsew default input
rlabel metal2 s 13358 21520 13414 22000 6 chany_top_in[8]
port 33 nsew default input
rlabel metal3 s 0 17280 480 17400 6 chany_top_out[0]
port 34 nsew default tristate
rlabel metal2 s 15842 21520 15898 22000 6 chany_top_out[1]
port 35 nsew default tristate
rlabel metal2 s 12898 0 12954 480 6 chany_top_out[2]
port 36 nsew default tristate
rlabel metal3 s 21520 14696 22000 14816 6 chany_top_out[3]
port 37 nsew default tristate
rlabel metal3 s 21520 15648 22000 15768 6 chany_top_out[4]
port 38 nsew default tristate
rlabel metal3 s 0 19184 480 19304 6 chany_top_out[5]
port 39 nsew default tristate
rlabel metal2 s 18234 21520 18290 22000 6 chany_top_out[6]
port 40 nsew default tristate
rlabel metal3 s 21520 16600 22000 16720 6 chany_top_out[7]
port 41 nsew default tristate
rlabel metal2 s 14922 0 14978 480 6 chany_top_out[8]
port 42 nsew default tristate
rlabel metal2 s 2870 0 2926 480 6 data_in
port 43 nsew default input
rlabel metal2 s 938 0 994 480 6 enable
port 44 nsew default input
rlabel metal2 s 16854 0 16910 480 6 left_grid_pin_0_
port 45 nsew default tristate
rlabel metal3 s 21520 19456 22000 19576 6 left_grid_pin_10_
port 46 nsew default tristate
rlabel metal3 s 21520 20408 22000 20528 6 left_grid_pin_12_
port 47 nsew default tristate
rlabel metal3 s 21520 21360 22000 21480 6 left_grid_pin_14_
port 48 nsew default tristate
rlabel metal3 s 21520 17552 22000 17672 6 left_grid_pin_2_
port 49 nsew default tristate
rlabel metal3 s 0 20952 480 21072 6 left_grid_pin_4_
port 50 nsew default tristate
rlabel metal3 s 21520 18504 22000 18624 6 left_grid_pin_6_
port 51 nsew default tristate
rlabel metal2 s 18878 0 18934 480 6 left_grid_pin_8_
port 52 nsew default tristate
rlabel metal2 s 20718 21520 20774 22000 6 right_grid_pin_3_
port 53 nsew default tristate
rlabel metal2 s 20902 0 20958 480 6 right_grid_pin_7_
port 54 nsew default tristate
rlabel metal4 s 4611 2128 4931 19632 6 vpwr
port 55 nsew default input
rlabel metal4 s 8277 2128 8597 19632 6 vgnd
port 56 nsew default input
<< end >>
