VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sb_3__1_
  CLASS BLOCK ;
  FOREIGN sb_3__1_ ;
  ORIGIN 0.000 0.000 ;
  SIZE 140.000 BY 140.000 ;
  PIN address[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2.850 137.600 3.130 140.000 ;
    END
  END address[0]
  PIN address[1]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 2.760 2.400 3.360 ;
    END
  END address[1]
  PIN address[2]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 3.440 140.000 4.040 ;
    END
  END address[2]
  PIN address[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 16.190 0.000 16.470 2.400 ;
    END
  END address[3]
  PIN address[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 8.830 137.600 9.110 140.000 ;
    END
  END address[4]
  PIN address[5]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 8.880 2.400 9.480 ;
    END
  END address[5]
  PIN address[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 15.270 137.600 15.550 140.000 ;
    END
  END address[6]
  PIN bottom_left_grid_pin_13_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 23.090 0.000 23.370 2.400 ;
    END
  END bottom_left_grid_pin_13_
  PIN bottom_right_grid_pin_11_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 21.800 2.400 22.400 ;
    END
  END bottom_right_grid_pin_11_
  PIN bottom_right_grid_pin_13_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 28.150 137.600 28.430 140.000 ;
    END
  END bottom_right_grid_pin_13_
  PIN bottom_right_grid_pin_15_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 34.590 137.600 34.870 140.000 ;
    END
  END bottom_right_grid_pin_15_
  PIN bottom_right_grid_pin_1_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 10.920 140.000 11.520 ;
    END
  END bottom_right_grid_pin_1_
  PIN bottom_right_grid_pin_3_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 18.400 140.000 19.000 ;
    END
  END bottom_right_grid_pin_3_
  PIN bottom_right_grid_pin_5_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 15.000 2.400 15.600 ;
    END
  END bottom_right_grid_pin_5_
  PIN bottom_right_grid_pin_7_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 21.710 137.600 21.990 140.000 ;
    END
  END bottom_right_grid_pin_7_
  PIN bottom_right_grid_pin_9_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 29.530 0.000 29.810 2.400 ;
    END
  END bottom_right_grid_pin_9_
  PIN chanx_left_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 27.920 2.400 28.520 ;
    END
  END chanx_left_in[0]
  PIN chanx_left_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 40.570 137.600 40.850 140.000 ;
    END
  END chanx_left_in[1]
  PIN chanx_left_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 26.560 140.000 27.160 ;
    END
  END chanx_left_in[2]
  PIN chanx_left_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 34.040 2.400 34.640 ;
    END
  END chanx_left_in[3]
  PIN chanx_left_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 36.430 0.000 36.710 2.400 ;
    END
  END chanx_left_in[4]
  PIN chanx_left_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 40.840 2.400 41.440 ;
    END
  END chanx_left_in[5]
  PIN chanx_left_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 46.960 2.400 47.560 ;
    END
  END chanx_left_in[6]
  PIN chanx_left_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 42.870 0.000 43.150 2.400 ;
    END
  END chanx_left_in[7]
  PIN chanx_left_in[8]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 34.040 140.000 34.640 ;
    END
  END chanx_left_in[8]
  PIN chanx_left_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 53.080 2.400 53.680 ;
    END
  END chanx_left_out[0]
  PIN chanx_left_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 47.010 137.600 47.290 140.000 ;
    END
  END chanx_left_out[1]
  PIN chanx_left_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 137.600 42.200 140.000 42.800 ;
    END
  END chanx_left_out[2]
  PIN chanx_left_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 137.600 49.680 140.000 50.280 ;
    END
  END chanx_left_out[3]
  PIN chanx_left_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 49.770 0.000 50.050 2.400 ;
    END
  END chanx_left_out[4]
  PIN chanx_left_out[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 59.880 2.400 60.480 ;
    END
  END chanx_left_out[5]
  PIN chanx_left_out[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 137.600 57.840 140.000 58.440 ;
    END
  END chanx_left_out[6]
  PIN chanx_left_out[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 53.450 137.600 53.730 140.000 ;
    END
  END chanx_left_out[7]
  PIN chanx_left_out[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 59.890 137.600 60.170 140.000 ;
    END
  END chanx_left_out[8]
  PIN chany_bottom_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 65.320 140.000 65.920 ;
    END
  END chany_bottom_in[0]
  PIN chany_bottom_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 66.000 2.400 66.600 ;
    END
  END chany_bottom_in[1]
  PIN chany_bottom_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 66.330 137.600 66.610 140.000 ;
    END
  END chany_bottom_in[2]
  PIN chany_bottom_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 56.210 0.000 56.490 2.400 ;
    END
  END chany_bottom_in[3]
  PIN chany_bottom_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 72.770 137.600 73.050 140.000 ;
    END
  END chany_bottom_in[4]
  PIN chany_bottom_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 63.110 0.000 63.390 2.400 ;
    END
  END chany_bottom_in[5]
  PIN chany_bottom_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 72.800 2.400 73.400 ;
    END
  END chany_bottom_in[6]
  PIN chany_bottom_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 78.920 2.400 79.520 ;
    END
  END chany_bottom_in[7]
  PIN chany_bottom_in[8]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 73.480 140.000 74.080 ;
    END
  END chany_bottom_in[8]
  PIN chany_bottom_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 69.550 0.000 69.830 2.400 ;
    END
  END chany_bottom_out[0]
  PIN chany_bottom_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 137.600 80.960 140.000 81.560 ;
    END
  END chany_bottom_out[1]
  PIN chany_bottom_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 85.040 2.400 85.640 ;
    END
  END chany_bottom_out[2]
  PIN chany_bottom_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 76.450 0.000 76.730 2.400 ;
    END
  END chany_bottom_out[3]
  PIN chany_bottom_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 82.890 0.000 83.170 2.400 ;
    END
  END chany_bottom_out[4]
  PIN chany_bottom_out[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 137.600 88.440 140.000 89.040 ;
    END
  END chany_bottom_out[5]
  PIN chany_bottom_out[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 91.840 2.400 92.440 ;
    END
  END chany_bottom_out[6]
  PIN chany_bottom_out[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 78.750 137.600 79.030 140.000 ;
    END
  END chany_bottom_out[7]
  PIN chany_bottom_out[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 89.790 0.000 90.070 2.400 ;
    END
  END chany_bottom_out[8]
  PIN chany_top_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 85.190 137.600 85.470 140.000 ;
    END
  END chany_top_in[0]
  PIN chany_top_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 96.230 0.000 96.510 2.400 ;
    END
  END chany_top_in[1]
  PIN chany_top_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 103.130 0.000 103.410 2.400 ;
    END
  END chany_top_in[2]
  PIN chany_top_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 96.600 140.000 97.200 ;
    END
  END chany_top_in[3]
  PIN chany_top_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 91.630 137.600 91.910 140.000 ;
    END
  END chany_top_in[4]
  PIN chany_top_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 98.070 137.600 98.350 140.000 ;
    END
  END chany_top_in[5]
  PIN chany_top_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 104.080 140.000 104.680 ;
    END
  END chany_top_in[6]
  PIN chany_top_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 112.240 140.000 112.840 ;
    END
  END chany_top_in[7]
  PIN chany_top_in[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 109.570 0.000 109.850 2.400 ;
    END
  END chany_top_in[8]
  PIN chany_top_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 137.600 119.720 140.000 120.320 ;
    END
  END chany_top_out[0]
  PIN chany_top_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 104.510 137.600 104.790 140.000 ;
    END
  END chany_top_out[1]
  PIN chany_top_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 110.490 137.600 110.770 140.000 ;
    END
  END chany_top_out[2]
  PIN chany_top_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 116.930 137.600 117.210 140.000 ;
    END
  END chany_top_out[3]
  PIN chany_top_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 97.960 2.400 98.560 ;
    END
  END chany_top_out[4]
  PIN chany_top_out[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 116.470 0.000 116.750 2.400 ;
    END
  END chany_top_out[5]
  PIN chany_top_out[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 104.080 2.400 104.680 ;
    END
  END chany_top_out[6]
  PIN chany_top_out[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 110.880 2.400 111.480 ;
    END
  END chany_top_out[7]
  PIN chany_top_out[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 122.910 0.000 123.190 2.400 ;
    END
  END chany_top_out[8]
  PIN data_in
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 9.750 0.000 10.030 2.400 ;
    END
  END data_in
  PIN enable
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 3.310 0.000 3.590 2.400 ;
    END
  END enable
  PIN left_bottom_grid_pin_12_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 123.370 137.600 123.650 140.000 ;
    END
  END left_bottom_grid_pin_12_
  PIN left_top_grid_pin_10_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 117.000 2.400 117.600 ;
    END
  END left_top_grid_pin_10_
  PIN top_left_grid_pin_13_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 129.810 137.600 130.090 140.000 ;
    END
  END top_left_grid_pin_13_
  PIN top_right_grid_pin_11_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 136.250 0.000 136.530 2.400 ;
    END
  END top_right_grid_pin_11_
  PIN top_right_grid_pin_13_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 135.360 140.000 135.960 ;
    END
  END top_right_grid_pin_13_
  PIN top_right_grid_pin_15_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 136.040 2.400 136.640 ;
    END
  END top_right_grid_pin_15_
  PIN top_right_grid_pin_1_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 129.810 0.000 130.090 2.400 ;
    END
  END top_right_grid_pin_1_
  PIN top_right_grid_pin_3_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 123.120 2.400 123.720 ;
    END
  END top_right_grid_pin_3_
  PIN top_right_grid_pin_5_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 129.920 2.400 130.520 ;
    END
  END top_right_grid_pin_5_
  PIN top_right_grid_pin_7_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 127.880 140.000 128.480 ;
    END
  END top_right_grid_pin_7_
  PIN top_right_grid_pin_9_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 136.250 137.600 136.530 140.000 ;
    END
  END top_right_grid_pin_9_
  PIN vpwr
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT 28.055 10.640 29.655 128.080 ;
    END
  END vpwr
  PIN vgnd
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT 51.385 10.640 52.985 128.080 ;
    END
  END vgnd
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 134.320 127.925 ;
      LAYER met1 ;
        RECT 0.070 0.380 138.390 137.660 ;
      LAYER met2 ;
        RECT 0.100 137.320 2.570 137.770 ;
        RECT 3.410 137.320 8.550 137.770 ;
        RECT 9.390 137.320 14.990 137.770 ;
        RECT 15.830 137.320 21.430 137.770 ;
        RECT 22.270 137.320 27.870 137.770 ;
        RECT 28.710 137.320 34.310 137.770 ;
        RECT 35.150 137.320 40.290 137.770 ;
        RECT 41.130 137.320 46.730 137.770 ;
        RECT 47.570 137.320 53.170 137.770 ;
        RECT 54.010 137.320 59.610 137.770 ;
        RECT 60.450 137.320 66.050 137.770 ;
        RECT 66.890 137.320 72.490 137.770 ;
        RECT 73.330 137.320 78.470 137.770 ;
        RECT 79.310 137.320 84.910 137.770 ;
        RECT 85.750 137.320 91.350 137.770 ;
        RECT 92.190 137.320 97.790 137.770 ;
        RECT 98.630 137.320 104.230 137.770 ;
        RECT 105.070 137.320 110.210 137.770 ;
        RECT 111.050 137.320 116.650 137.770 ;
        RECT 117.490 137.320 123.090 137.770 ;
        RECT 123.930 137.320 129.530 137.770 ;
        RECT 130.370 137.320 135.970 137.770 ;
        RECT 136.810 137.320 138.370 137.770 ;
        RECT 0.100 2.680 138.370 137.320 ;
        RECT 0.100 0.270 3.030 2.680 ;
        RECT 3.870 0.270 9.470 2.680 ;
        RECT 10.310 0.270 15.910 2.680 ;
        RECT 16.750 0.270 22.810 2.680 ;
        RECT 23.650 0.270 29.250 2.680 ;
        RECT 30.090 0.270 36.150 2.680 ;
        RECT 36.990 0.270 42.590 2.680 ;
        RECT 43.430 0.270 49.490 2.680 ;
        RECT 50.330 0.270 55.930 2.680 ;
        RECT 56.770 0.270 62.830 2.680 ;
        RECT 63.670 0.270 69.270 2.680 ;
        RECT 70.110 0.270 76.170 2.680 ;
        RECT 77.010 0.270 82.610 2.680 ;
        RECT 83.450 0.270 89.510 2.680 ;
        RECT 90.350 0.270 95.950 2.680 ;
        RECT 96.790 0.270 102.850 2.680 ;
        RECT 103.690 0.270 109.290 2.680 ;
        RECT 110.130 0.270 116.190 2.680 ;
        RECT 117.030 0.270 122.630 2.680 ;
        RECT 123.470 0.270 129.530 2.680 ;
        RECT 130.370 0.270 135.970 2.680 ;
        RECT 136.810 0.270 138.370 2.680 ;
      LAYER met3 ;
        RECT 2.800 135.640 137.200 136.040 ;
        RECT 0.270 134.960 137.200 135.640 ;
        RECT 0.270 130.920 138.650 134.960 ;
        RECT 2.800 129.520 138.650 130.920 ;
        RECT 0.270 128.880 138.650 129.520 ;
        RECT 0.270 127.480 137.200 128.880 ;
        RECT 0.270 124.120 138.650 127.480 ;
        RECT 2.800 122.720 138.650 124.120 ;
        RECT 0.270 120.720 138.650 122.720 ;
        RECT 0.270 119.320 137.200 120.720 ;
        RECT 0.270 118.000 138.650 119.320 ;
        RECT 2.800 116.600 138.650 118.000 ;
        RECT 0.270 113.240 138.650 116.600 ;
        RECT 0.270 111.880 137.200 113.240 ;
        RECT 2.800 111.840 137.200 111.880 ;
        RECT 2.800 110.480 138.650 111.840 ;
        RECT 0.270 105.080 138.650 110.480 ;
        RECT 2.800 103.680 137.200 105.080 ;
        RECT 0.270 98.960 138.650 103.680 ;
        RECT 2.800 97.600 138.650 98.960 ;
        RECT 2.800 97.560 137.200 97.600 ;
        RECT 0.270 96.200 137.200 97.560 ;
        RECT 0.270 92.840 138.650 96.200 ;
        RECT 2.800 91.440 138.650 92.840 ;
        RECT 0.270 89.440 138.650 91.440 ;
        RECT 0.270 88.040 137.200 89.440 ;
        RECT 0.270 86.040 138.650 88.040 ;
        RECT 2.800 84.640 138.650 86.040 ;
        RECT 0.270 81.960 138.650 84.640 ;
        RECT 0.270 80.560 137.200 81.960 ;
        RECT 0.270 79.920 138.650 80.560 ;
        RECT 2.800 78.520 138.650 79.920 ;
        RECT 0.270 74.480 138.650 78.520 ;
        RECT 0.270 73.800 137.200 74.480 ;
        RECT 2.800 73.080 137.200 73.800 ;
        RECT 2.800 72.400 138.650 73.080 ;
        RECT 0.270 67.000 138.650 72.400 ;
        RECT 2.800 66.320 138.650 67.000 ;
        RECT 2.800 65.600 137.200 66.320 ;
        RECT 0.270 64.920 137.200 65.600 ;
        RECT 0.270 60.880 138.650 64.920 ;
        RECT 2.800 59.480 138.650 60.880 ;
        RECT 0.270 58.840 138.650 59.480 ;
        RECT 0.270 57.440 137.200 58.840 ;
        RECT 0.270 54.080 138.650 57.440 ;
        RECT 2.800 52.680 138.650 54.080 ;
        RECT 0.270 50.680 138.650 52.680 ;
        RECT 0.270 49.280 137.200 50.680 ;
        RECT 0.270 47.960 138.650 49.280 ;
        RECT 2.800 46.560 138.650 47.960 ;
        RECT 0.270 43.200 138.650 46.560 ;
        RECT 0.270 41.840 137.200 43.200 ;
        RECT 2.800 41.800 137.200 41.840 ;
        RECT 2.800 40.440 138.650 41.800 ;
        RECT 0.270 35.040 138.650 40.440 ;
        RECT 2.800 33.640 137.200 35.040 ;
        RECT 0.270 28.920 138.650 33.640 ;
        RECT 2.800 27.560 138.650 28.920 ;
        RECT 2.800 27.520 137.200 27.560 ;
        RECT 0.270 26.160 137.200 27.520 ;
        RECT 0.270 22.800 138.650 26.160 ;
        RECT 2.800 21.400 138.650 22.800 ;
        RECT 0.270 19.400 138.650 21.400 ;
        RECT 0.270 18.000 137.200 19.400 ;
        RECT 0.270 16.000 138.650 18.000 ;
        RECT 2.800 14.600 138.650 16.000 ;
        RECT 0.270 11.920 138.650 14.600 ;
        RECT 0.270 10.520 137.200 11.920 ;
        RECT 0.270 9.880 138.650 10.520 ;
        RECT 2.800 8.480 138.650 9.880 ;
        RECT 0.270 4.440 138.650 8.480 ;
        RECT 0.270 3.760 137.200 4.440 ;
        RECT 2.800 3.360 137.200 3.760 ;
      LAYER met4 ;
        RECT 0.295 10.640 27.655 128.080 ;
        RECT 30.055 10.640 50.985 128.080 ;
        RECT 53.385 10.640 138.625 128.080 ;
      LAYER met5 ;
        RECT 7.020 51.900 21.500 53.500 ;
  END
END sb_3__1_
END LIBRARY

