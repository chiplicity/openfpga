* NGSPICE file created from grid_clb.ext - technology: EFS8A

* Black-box entry subcircuit for scs8hd_decap_8 abstract view
.subckt scs8hd_decap_8 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_fill_2 abstract view
.subckt scs8hd_fill_2 vpwr vgnd
.ends

* Black-box entry subcircuit for scs8hd_diode_2 abstract view
.subckt scs8hd_diode_2 DIODE vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_decap_4 abstract view
.subckt scs8hd_decap_4 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_ebufn_2 abstract view
.subckt scs8hd_ebufn_2 A TEB Z vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_decap_12 abstract view
.subckt scs8hd_decap_12 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_nor2_4 abstract view
.subckt scs8hd_nor2_4 A B Y vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_buf_1 abstract view
.subckt scs8hd_buf_1 A X vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_decap_6 abstract view
.subckt scs8hd_decap_6 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_fill_1 abstract view
.subckt scs8hd_fill_1 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_inv_1 abstract view
.subckt scs8hd_inv_1 A Y vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_decap_3 abstract view
.subckt scs8hd_decap_3 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_lpflow_inputisolatch_1 abstract view
.subckt scs8hd_lpflow_inputisolatch_1 D Q SLEEPB vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_or4_4 abstract view
.subckt scs8hd_or4_4 A B C D X vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_tapvpwrvgnd_1 abstract view
.subckt scs8hd_tapvpwrvgnd_1 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_conb_1 abstract view
.subckt scs8hd_conb_1 HI LO vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_or2_4 abstract view
.subckt scs8hd_or2_4 A B X vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_inv_8 abstract view
.subckt scs8hd_inv_8 A Y vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_or3_4 abstract view
.subckt scs8hd_or3_4 A B C X vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_dfbbp_1 abstract view
.subckt scs8hd_dfbbp_1 CLK D Q QN RESETB SETB vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_clkbuf_16 abstract view
.subckt scs8hd_clkbuf_16 A X vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_clkbuf_1 abstract view
.subckt scs8hd_clkbuf_1 A X vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_nand2_4 abstract view
.subckt scs8hd_nand2_4 A B Y vgnd vpwr
.ends

.subckt grid_clb address[0] address[1] address[2] address[3] address[4] address[5]
+ address[6] address[7] address[8] address[9] bottom_width_0_height_0__pin_10_ bottom_width_0_height_0__pin_14_
+ bottom_width_0_height_0__pin_2_ bottom_width_0_height_0__pin_6_ clk data_in enable
+ left_width_0_height_0__pin_11_ left_width_0_height_0__pin_3_ left_width_0_height_0__pin_7_
+ reset right_width_0_height_0__pin_13_ right_width_0_height_0__pin_1_ right_width_0_height_0__pin_5_
+ right_width_0_height_0__pin_9_ set top_width_0_height_0__pin_0_ top_width_0_height_0__pin_12_
+ top_width_0_height_0__pin_4_ top_width_0_height_0__pin_8_ vpwr vgnd
XFILLER_54_203 vgnd vpwr scs8hd_decap_8
XFILLER_27_406 vpwr vgnd scs8hd_fill_2
XFILLER_39_266 vpwr vgnd scs8hd_fill_2
XFILLER_39_277 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.buf4_2_.scs8hd_buf_1_A
+ ltile_clb_0.mux_fle_1_in_2.INVTX1_14_.scs8hd_inv_1/Y vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mem_fle_3_in_2.LATCH_7_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_42_409 vgnd vpwr scs8hd_decap_4
XFILLER_35_461 vpwr vgnd scs8hd_fill_2
XFILLER_50_420 vgnd vpwr scs8hd_decap_4
XFILLER_50_431 vgnd vpwr scs8hd_decap_8
Xltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_6_.TGATE_0_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_12_.scs8hd_inv_1/Y
+ _613_/Y ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_6_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_22_166 vgnd vpwr scs8hd_decap_8
XANTENNA_ltile_clb_0.mux_fle_2_in_3.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_2_in_3.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_77_15 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mem_fle_3_in_3.LATCH_5_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_77_59 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mem_fle_0_in_0.LATCH_7_.latch_SLEEPB _518_/Y vgnd vpwr scs8hd_diode_2
XFILLER_77_339 vpwr vgnd scs8hd_fill_2
XFILLER_73_501 vgnd vpwr scs8hd_decap_12
XFILLER_45_214 vpwr vgnd scs8hd_fill_2
XFILLER_45_236 vpwr vgnd scs8hd_fill_2
X_501_ _421_/A _495_/X _501_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_45_269 vpwr vgnd scs8hd_fill_2
X_432_ _432_/A _429_/X _432_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2_TEB
+ _621_/Y vgnd vpwr scs8hd_diode_2
X_363_ _374_/A _365_/B _363_/Y vgnd vpwr scs8hd_nor2_4
X_294_ _293_/X _569_/A vgnd vpwr scs8hd_buf_1
XFILLER_9_159 vgnd vpwr scs8hd_decap_12
XFILLER_5_398 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_3_.scs8hd_inv_1_A
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_68_328 vgnd vpwr scs8hd_decap_8
XFILLER_68_306 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_1_in_3.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_1_in_3.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_36_225 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_1_.TGATE_1_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_3_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_36_269 vgnd vpwr scs8hd_decap_6
XFILLER_17_472 vgnd vpwr scs8hd_decap_8
XFILLER_44_280 vgnd vpwr scs8hd_fill_1
Xltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_3_.scs8hd_inv_1
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_3_.latch/Q
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_32_486 vgnd vpwr scs8hd_fill_1
Xltile_clb_0.mux_fle_2_in_1.INVTX1_5_.scs8hd_inv_1 right_width_0_height_0__pin_5_
+ ltile_clb_0.mux_fle_2_in_1.INVTX1_5_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XANTENNA__304__A _304_/A vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_0_in_1.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_0_in_1.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2/Z
+ ltile_clb_0.mem_fle_0_in_1.LATCH_7_.latch/Q ltile_clb_0.mux_fle_0_in_1.INVTX1_14_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_67_372 vpwr vgnd scs8hd_fill_2
XANTENNA__396__D _346_/D vgnd vpwr scs8hd_diode_2
XFILLER_27_225 vpwr vgnd scs8hd_fill_2
XFILLER_82_342 vgnd vpwr scs8hd_decap_12
XFILLER_27_236 vpwr vgnd scs8hd_fill_2
XFILLER_27_258 vpwr vgnd scs8hd_fill_2
XFILLER_63_39 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_27_269 vpwr vgnd scs8hd_fill_2
XFILLER_82_397 vgnd vpwr scs8hd_decap_6
XANTENNA_ltile_clb_0.mux_fle_3_in_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_3_in_0.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_5_.scs8hd_inv_1/Y
+ _620_/Y ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_1_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_23_442 vgnd vpwr scs8hd_decap_3
XFILLER_50_272 vgnd vpwr scs8hd_fill_1
XFILLER_12_32 vgnd vpwr scs8hd_decap_12
XFILLER_6_129 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_14_.scs8hd_inv_1
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_14_.latch/Q
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_14_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_ltile_clb_0.mux_fle_0_in_2.INVTX1_7_.scs8hd_inv_1_A left_width_0_height_0__pin_7_
+ vgnd vpwr scs8hd_diode_2
XFILLER_2_335 vgnd vpwr scs8hd_fill_1
XFILLER_77_147 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_13_.scs8hd_inv_1_A
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_13_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_58_350 vgnd vpwr scs8hd_fill_1
Xltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_0_.latch
+ data_in ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_0_.latch/Q
+ _546_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_37_51 vgnd vpwr scs8hd_decap_8
XFILLER_46_512 vgnd vpwr scs8hd_decap_4
XFILLER_37_62 vgnd vpwr scs8hd_decap_12
XFILLER_73_397 vgnd vpwr scs8hd_fill_1
XFILLER_26_291 vgnd vpwr scs8hd_decap_3
X_415_ _328_/A _432_/A vgnd vpwr scs8hd_buf_1
X_346_ address[8] _369_/B _346_/C _346_/D _347_/A vgnd vpwr scs8hd_or4_4
Xltile_clb_0.mux_fle_2_in_2.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_2_in_2.INVTX1_9_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_2_in_2.LATCH_1_.latch/Q ltile_clb_0.mux_fle_2_in_2.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
Xltile_clb_0.mux_fle_0_in_2.mux_l1_in_3_.TGATE_2_.scs8hd_ebufn_2 _642_/HI ltile_clb_0.mem_fle_0_in_2.LATCH_2_.latch/Q
+ ltile_clb_0.mux_fle_0_in_2.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
X_277_ _267_/X _564_/A _277_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_4_.TGATE_0_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_8_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_3_in_2.INVTX1_0_.scs8hd_inv_1 top_width_0_height_0__pin_0_ ltile_clb_0.mux_fle_3_in_2.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_5_184 vgnd vpwr scs8hd_decap_12
XFILLER_78_80 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mux_fle_1_in_3.INVTX1_4_.scs8hd_inv_1_A top_width_0_height_0__pin_4_
+ vgnd vpwr scs8hd_diode_2
XFILLER_76_180 vgnd vpwr scs8hd_decap_12
XFILLER_52_515 vgnd vpwr scs8hd_fill_1
XFILLER_24_206 vgnd vpwr scs8hd_decap_4
XANTENNA_ltile_clb_0.mux_fle_2_in_0.INVTX1_0_.scs8hd_inv_1_A top_width_0_height_0__pin_0_
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_1_.latch_SLEEPB
+ _571_/Y vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_2_in_2.INVTX1_9_.scs8hd_inv_1 right_width_0_height_0__pin_9_
+ ltile_clb_0.mux_fle_2_in_2.INVTX1_9_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XFILLER_47_309 vpwr vgnd scs8hd_fill_2
XFILLER_74_117 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_8_.scs8hd_inv_1
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_8_.latch/Q
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_8_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_74_27 vgnd vpwr scs8hd_decap_4
XFILLER_43_515 vgnd vpwr scs8hd_fill_1
XPHY_702 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_55_397 vpwr vgnd scs8hd_fill_2
XFILLER_15_239 vgnd vpwr scs8hd_decap_3
XANTENNA_ltile_clb_0.mem_fle_0_in_3.LATCH_0_.latch_SLEEPB _492_/Y vgnd vpwr scs8hd_diode_2
XPHY_735 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_724 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_713 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_768 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_757 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_746 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_11_423 vpwr vgnd scs8hd_fill_2
XPHY_779 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_11_434 vpwr vgnd scs8hd_fill_2
XFILLER_23_86 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mux_fle_0_in_2.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_0_in_2.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mem_fle_0_in_1.LATCH_2_.latch data_in ltile_clb_0.mem_fle_0_in_1.LATCH_2_.latch/Q
+ _512_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_78_401 vgnd vpwr scs8hd_decap_6
XFILLER_2_154 vgnd vpwr scs8hd_decap_12
XANTENNA__598__B _580_/X vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_3_in_3.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_3_in_3.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_61_301 vpwr vgnd scs8hd_fill_2
XFILLER_73_194 vpwr vgnd scs8hd_fill_2
XFILLER_73_172 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.mem_fle_1_in_1.LATCH_1_.latch data_in ltile_clb_0.mem_fle_1_in_1.LATCH_1_.latch/Q
+ _469_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_64_93 vgnd vpwr scs8hd_decap_12
XFILLER_61_367 vgnd vpwr scs8hd_decap_8
XFILLER_61_356 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_5_.scs8hd_inv_1_A
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_5_.latch/Q
+ vgnd vpwr scs8hd_diode_2
X_329_ _374_/A _338_/B _329_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA_ltile_clb_0.mux_fle_3_in_3.INVTX1_10_.scs8hd_inv_1_A bottom_width_0_height_0__pin_10_
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_3_in_3.INVTX1_4_.scs8hd_inv_1 top_width_0_height_0__pin_4_ ltile_clb_0.mux_fle_3_in_3.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
Xltile_clb_0.mem_fle_2_in_1.LATCH_0_.latch data_in ltile_clb_0.mem_fle_2_in_1.LATCH_0_.latch/Q
+ _426_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_50_3 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_6_.TGATE_1_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_13_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__301__B _545_/A vgnd vpwr scs8hd_diode_2
XFILLER_29_309 vpwr vgnd scs8hd_fill_2
XFILLER_69_489 vgnd vpwr scs8hd_decap_12
XFILLER_56_117 vgnd vpwr scs8hd_decap_12
XFILLER_25_515 vgnd vpwr scs8hd_fill_1
XFILLER_37_353 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.mux_fle_0_in_0.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_0_in_0.INVTX1_8_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_0_in_0.LATCH_0_.latch/Q ltile_clb_0.mux_fle_0_in_0.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_52_312 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_0_in_3.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_0_in_3.INVTX1_8_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_69_27 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mux_fle_3_in_1.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_3_in_1.INVTX1_8_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mem_fle_1_in_2.LATCH_0_.latch_SLEEPB _459_/Y vgnd vpwr scs8hd_diode_2
Xltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_3_.TGATE_0_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_6_.TGATE_0_.scs8hd_ebufn_2/Z
+ _631_/Y ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_1_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_16_515 vgnd vpwr scs8hd_fill_1
XFILLER_43_301 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_1_.TGATE_1_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_1_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_28_386 vgnd vpwr scs8hd_decap_8
XFILLER_43_334 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_13_.latch_D
+ data_in vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mem_fle_0_in_3.LATCH_5_.latch data_in ltile_clb_0.mem_fle_0_in_3.LATCH_5_.latch/Q
+ _487_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XPHY_510 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_43_345 vgnd vpwr scs8hd_decap_4
Xltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.buf4_2_.scs8hd_buf_1
+ ltile_clb_0.mux_fle_1_in_2.INVTX1_14_.scs8hd_inv_1/Y _624_/A vgnd vpwr scs8hd_buf_1
XPHY_521 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_43_378 vgnd vpwr scs8hd_fill_1
XPHY_532 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_543 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xltile_clb_0.mux_fle_1_in_3.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_1_in_3.INVTX1_9_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_1_in_3.LATCH_1_.latch/Q ltile_clb_0.mux_fle_1_in_3.mux_l1_in_2_.TGATE_3_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
Xltile_clb_0.mux_fle_3_in_3.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_3_in_3.INVTX1_4_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_3_in_3.LATCH_0_.latch/Q ltile_clb_0.mux_fle_3_in_3.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_70_197 vgnd vpwr scs8hd_decap_6
XPHY_587 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_554 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_565 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_576 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_598 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_11_297 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
+ _617_/Y vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mem_fle_1_in_3.LATCH_4_.latch data_in ltile_clb_0.mem_fle_1_in_3.LATCH_4_.latch/Q
+ _444_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA__402__A _391_/A vgnd vpwr scs8hd_diode_2
XFILLER_38_117 vgnd vpwr scs8hd_decap_12
XFILLER_66_459 vgnd vpwr scs8hd_decap_6
XFILLER_19_342 vpwr vgnd scs8hd_fill_2
XFILLER_74_492 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.mem_fle_2_in_3.LATCH_3_.latch data_in ltile_clb_0.mem_fle_2_in_3.LATCH_3_.latch/Q
+ _392_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_46_172 vgnd vpwr scs8hd_fill_1
XFILLER_46_194 vgnd vpwr scs8hd_fill_1
XFILLER_34_367 vpwr vgnd scs8hd_fill_2
XFILLER_61_175 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.mem_fle_3_in_3.LATCH_2_.latch data_in ltile_clb_0.mem_fle_3_in_3.LATCH_2_.latch/Q
+ _338_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_6_290 vpwr vgnd scs8hd_fill_2
XANTENNA__312__A _603_/A vgnd vpwr scs8hd_diode_2
XFILLER_69_264 vpwr vgnd scs8hd_fill_2
XFILLER_57_404 vpwr vgnd scs8hd_fill_2
XFILLER_57_437 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.mux_fle_3_in_0.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_3_in_0.INVTX1_3_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_3_in_0.LATCH_3_.latch/Q ltile_clb_0.mux_fle_3_in_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_65_492 vpwr vgnd scs8hd_fill_2
XFILLER_25_301 vpwr vgnd scs8hd_fill_2
XFILLER_37_172 vgnd vpwr scs8hd_decap_4
XFILLER_80_440 vgnd vpwr scs8hd_fill_1
XFILLER_25_367 vgnd vpwr scs8hd_fill_1
XFILLER_80_495 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mem_fle_2_in_1.LATCH_0_.latch_SLEEPB _426_/Y vgnd vpwr scs8hd_diode_2
XFILLER_71_39 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_14_.scs8hd_inv_1
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_14_.latch/Q
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_14_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_ltile_clb_0.mux_fle_0_in_2.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_0_in_2.LATCH_7_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_20_32 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_4_.TGATE_0_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_8_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_75_212 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.mem_ble4_out_0.LATCH_0_.latch
+ data_in ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.mem_ble4_out_0.LATCH_0_.latch/Q
+ _577_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_75_245 vpwr vgnd scs8hd_fill_2
XFILLER_75_234 vpwr vgnd scs8hd_fill_2
XFILLER_29_74 vgnd vpwr scs8hd_decap_12
XFILLER_75_278 vpwr vgnd scs8hd_fill_2
XFILLER_75_267 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_6_.latch_SLEEPB
+ _285_/Y vgnd vpwr scs8hd_diode_2
XFILLER_16_312 vgnd vpwr scs8hd_fill_1
XFILLER_28_183 vpwr vgnd scs8hd_fill_2
XFILLER_71_440 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_2_in_2.INVTX1_14_.scs8hd_inv_1_A ltile_clb_0.mux_fle_2_in_2.INVTX1_14_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
X_594_ _542_/A _588_/X _594_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_45_51 vgnd vpwr scs8hd_decap_8
XFILLER_45_62 vgnd vpwr scs8hd_decap_12
XFILLER_71_473 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l4_in_0_.TGATE_0_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ _627_/Y ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_16_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_31_315 vgnd vpwr scs8hd_decap_4
XFILLER_43_164 vpwr vgnd scs8hd_fill_2
XFILLER_43_175 vpwr vgnd scs8hd_fill_2
XPHY_340 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_351 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_362 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_373 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_384 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_395 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_ltile_clb_0.mux_fle_3_in_0.INVTX1_6_.scs8hd_inv_1_A bottom_width_0_height_0__pin_6_
+ vgnd vpwr scs8hd_diode_2
XFILLER_6_56 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.mux_fle_1_in_0.INVTX1_13_.scs8hd_inv_1 right_width_0_height_0__pin_13_
+ ltile_clb_0.mux_fle_1_in_0.INVTX1_13_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XANTENNA_ltile_clb_0.mux_fle_3_in_2.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_3_in_2.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_13_3 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_7_.scs8hd_inv_1_A
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_7_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_66_267 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_7_.TGATE_1_.scs8hd_ebufn_2_TEB
+ _620_/Y vgnd vpwr scs8hd_diode_2
XFILLER_19_161 vpwr vgnd scs8hd_fill_2
XFILLER_47_470 vpwr vgnd scs8hd_fill_2
XFILLER_62_484 vgnd vpwr scs8hd_decap_8
Xltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.INVTX1_0_.scs8hd_inv_1/Y
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.mem_ble4_out_0.LATCH_0_.latch/Q
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_34_175 vgnd vpwr scs8hd_decap_8
XFILLER_62_495 vgnd vpwr scs8hd_decap_12
XFILLER_22_326 vgnd vpwr scs8hd_decap_8
XFILLER_22_337 vgnd vpwr scs8hd_decap_8
Xltile_clb_0.mux_fle_0_in_0.INVTX1_0_.scs8hd_inv_1 top_width_0_height_0__pin_0_ ltile_clb_0.mux_fle_0_in_0.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA__307__A address[4] vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_1_in_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_1_in_0.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_30_370 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_3_in_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_3_in_2.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_1_208 vgnd vpwr scs8hd_decap_4
XANTENNA_ltile_clb_0.mem_fle_3_in_0.LATCH_0_.latch_SLEEPB _379_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
+ _613_/Y vgnd vpwr scs8hd_diode_2
Xltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_1_.scs8hd_inv_1
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_1_.latch/Q
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_57_245 vpwr vgnd scs8hd_fill_2
XFILLER_57_234 vgnd vpwr scs8hd_fill_1
XFILLER_72_226 vpwr vgnd scs8hd_fill_2
XFILLER_82_27 vgnd vpwr scs8hd_decap_4
XFILLER_53_451 vpwr vgnd scs8hd_fill_2
XFILLER_13_315 vpwr vgnd scs8hd_fill_2
XFILLER_13_326 vpwr vgnd scs8hd_fill_2
XFILLER_13_337 vpwr vgnd scs8hd_fill_2
XFILLER_13_348 vpwr vgnd scs8hd_fill_2
XFILLER_15_98 vgnd vpwr scs8hd_decap_12
XFILLER_40_145 vgnd vpwr scs8hd_decap_8
XANTENNA_ltile_clb_0.mux_fle_3_in_1.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_3_in_1.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_31_86 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_6_.TGATE_1_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_13_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_0_274 vgnd vpwr scs8hd_decap_3
XFILLER_36_407 vgnd vpwr scs8hd_decap_12
XFILLER_63_204 vpwr vgnd scs8hd_fill_2
XFILLER_29_481 vgnd vpwr scs8hd_decap_4
XANTENNA_ltile_clb_0.mem_fle_0_in_1.LATCH_1_.latch_SLEEPB _513_/Y vgnd vpwr scs8hd_diode_2
X_646_ _646_/HI _646_/LO vgnd vpwr scs8hd_conb_1
X_577_ _603_/A _575_/B _577_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_31_123 vgnd vpwr scs8hd_decap_12
XFILLER_72_93 vgnd vpwr scs8hd_decap_12
XPHY_170 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_181 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_192 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ _607_/Y ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
Xltile_clb_0.mux_fle_2_in_1.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_2_in_1.INVTX1_3_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_2_in_1.LATCH_3_.latch/Q ltile_clb_0.mux_fle_2_in_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_39_256 vgnd vpwr scs8hd_fill_1
Xltile_clb_0.mux_fle_0_in_1.INVTX1_4_.scs8hd_inv_1 top_width_0_height_0__pin_4_ ltile_clb_0.mux_fle_0_in_1.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_35_484 vpwr vgnd scs8hd_fill_2
XFILLER_62_270 vpwr vgnd scs8hd_fill_2
XFILLER_50_454 vgnd vpwr scs8hd_decap_4
XFILLER_50_487 vgnd vpwr scs8hd_decap_8
XANTENNA_ltile_clb_0.mux_fle_1_in_0.mux_l1_in_2_.TGATE_3_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_1_in_0.INVTX1_11_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_77_27 vgnd vpwr scs8hd_decap_12
XFILLER_77_318 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_0_in_1.INVTX1_13_.scs8hd_inv_1_A right_width_0_height_0__pin_13_
+ vgnd vpwr scs8hd_diode_2
XFILLER_58_510 vgnd vpwr scs8hd_decap_6
XANTENNA__500__A _334_/A vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_0_in_0.INVTX1_4_.scs8hd_inv_1_A top_width_0_height_0__pin_4_
+ vgnd vpwr scs8hd_diode_2
XFILLER_73_513 vgnd vpwr scs8hd_decap_3
X_500_ _334_/A _495_/X _500_/Y vgnd vpwr scs8hd_nor2_4
X_431_ _431_/A _429_/X _431_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_26_462 vpwr vgnd scs8hd_fill_2
XFILLER_53_292 vpwr vgnd scs8hd_fill_2
XFILLER_53_281 vgnd vpwr scs8hd_decap_8
XFILLER_13_123 vgnd vpwr scs8hd_decap_12
XFILLER_41_421 vgnd vpwr scs8hd_decap_4
X_362_ _326_/A _365_/B _362_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_13_167 vgnd vpwr scs8hd_decap_3
XFILLER_13_189 vpwr vgnd scs8hd_fill_2
X_293_ _278_/X _333_/A _293_/X vgnd vpwr scs8hd_or2_4
XFILLER_41_498 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mux_fle_2_in_0.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_2_in_0.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_5_300 vgnd vpwr scs8hd_decap_3
XANTENNA_ltile_clb_0.mem_fle_1_in_0.LATCH_1_.latch_SLEEPB _480_/Y vgnd vpwr scs8hd_diode_2
XFILLER_5_344 vgnd vpwr scs8hd_fill_1
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
+ _631_/Y vgnd vpwr scs8hd_diode_2
XFILLER_68_318 vgnd vpwr scs8hd_fill_1
XANTENNA__410__A _409_/X vgnd vpwr scs8hd_diode_2
XFILLER_76_384 vpwr vgnd scs8hd_fill_2
XFILLER_76_373 vgnd vpwr scs8hd_decap_6
XFILLER_36_215 vgnd vpwr scs8hd_decap_6
XFILLER_36_248 vpwr vgnd scs8hd_fill_2
XFILLER_36_259 vgnd vpwr scs8hd_decap_4
X_629_ _629_/A _629_/Y vgnd vpwr scs8hd_inv_8
XFILLER_44_270 vgnd vpwr scs8hd_decap_4
XFILLER_32_454 vgnd vpwr scs8hd_fill_1
XANTENNA_ltile_clb_0.mux_fle_1_in_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_1_in_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_80_3 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mux_fle_1_in_1.INVTX1_1_.scs8hd_inv_1_A right_width_0_height_0__pin_1_
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_9_.scs8hd_inv_1_A
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_9_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__304__B _546_/A vgnd vpwr scs8hd_diode_2
XANTENNA__320__A address[8] vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_0_in_2.INVTX1_8_.scs8hd_inv_1 top_width_0_height_0__pin_8_ ltile_clb_0.mux_fle_0_in_2.INVTX1_8_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_55_502 vgnd vpwr scs8hd_decap_12
XFILLER_27_204 vgnd vpwr scs8hd_decap_4
XFILLER_82_354 vgnd vpwr scs8hd_decap_12
XFILLER_42_207 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_2_in_2.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_2_in_2.INVTX1_8_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_14_.scs8hd_inv_1
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_14_.latch/Q
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_14_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_42_229 vgnd vpwr scs8hd_decap_4
Xltile_clb_0.mux_fle_0_in_2.INVTX1_11_.scs8hd_inv_1 left_width_0_height_0__pin_11_
+ ltile_clb_0.mux_fle_0_in_2.INVTX1_11_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XFILLER_23_487 vgnd vpwr scs8hd_fill_1
XFILLER_23_498 vgnd vpwr scs8hd_decap_4
XFILLER_50_295 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.mux_fle_3_in_2.INVTX1_10_.scs8hd_inv_1 bottom_width_0_height_0__pin_10_
+ ltile_clb_0.mux_fle_3_in_2.INVTX1_10_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XFILLER_12_44 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_10_.latch_D
+ data_in vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_2_.scs8hd_inv_1_A
+ ltile_clb_0.mux_fle_1_in_2.INVTX1_14_.scs8hd_inv_1/Y vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_0_in_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_0_in_0.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__230__A _229_/Y vgnd vpwr scs8hd_diode_2
XFILLER_77_159 vgnd vpwr scs8hd_decap_12
XFILLER_73_310 vgnd vpwr scs8hd_fill_1
XFILLER_73_332 vpwr vgnd scs8hd_fill_2
XFILLER_37_74 vgnd vpwr scs8hd_decap_12
XFILLER_73_376 vpwr vgnd scs8hd_fill_2
XFILLER_33_218 vpwr vgnd scs8hd_fill_2
X_414_ _431_/A _412_/B _414_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_53_62 vgnd vpwr scs8hd_decap_12
XFILLER_53_51 vgnd vpwr scs8hd_decap_8
XFILLER_41_240 vpwr vgnd scs8hd_fill_2
X_345_ _345_/A _346_/D vgnd vpwr scs8hd_buf_1
X_276_ _276_/A _564_/A vgnd vpwr scs8hd_buf_1
XFILLER_41_295 vgnd vpwr scs8hd_decap_4
XANTENNA__405__A _394_/A vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_0_in_3.INVTX1_13_.scs8hd_inv_1 right_width_0_height_0__pin_13_
+ ltile_clb_0.mux_fle_0_in_3.INVTX1_13_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
Xltile_clb_0.mux_fle_1_in_2.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_1_in_2.INVTX1_3_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_1_in_2.LATCH_3_.latch/Q ltile_clb_0.mux_fle_1_in_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_5_196 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.mux_fle_3_in_3.INVTX1_12_.scs8hd_inv_1 top_width_0_height_0__pin_12_
+ ltile_clb_0.mux_fle_3_in_3.INVTX1_12_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
Xltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_0_.scs8hd_inv_1/Y
+ _629_/Y ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
Xltile_clb_0.mux_fle_1_in_3.INVTX1_3_.scs8hd_inv_1 left_width_0_height_0__pin_3_ ltile_clb_0.mux_fle_1_in_3.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
Xltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.mem_ble4_out_0.LATCH_0_.latch
+ data_in ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.mem_ble4_out_0.LATCH_0_.latch/Q
+ _312_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_49_362 vpwr vgnd scs8hd_fill_2
XFILLER_76_192 vgnd vpwr scs8hd_decap_3
XANTENNA_ltile_clb_0.mux_fle_2_in_3.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_2_in_3.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_64_321 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_3_in_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_3_in_0.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_64_398 vgnd vpwr scs8hd_fill_1
XFILLER_17_292 vpwr vgnd scs8hd_fill_2
XFILLER_20_413 vgnd vpwr scs8hd_decap_4
XFILLER_32_273 vpwr vgnd scs8hd_fill_2
XANTENNA__315__A address[9] vgnd vpwr scs8hd_diode_2
XFILLER_9_480 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.INVTX1_1_.scs8hd_inv_1
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.INVTX1_1_.scs8hd_inv_1/A
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.mem_ble4_out_0.LATCH_0_.latch_SLEEPB
+ _551_/Y vgnd vpwr scs8hd_diode_2
XFILLER_74_129 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_55_343 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_4_.TGATE_1_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_9_.scs8hd_inv_1/Y
+ _628_/Y ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_2_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_ltile_clb_0.mux_fle_1_in_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_1_in_1.LATCH_4_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_3_in_3.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_3_in_3.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_55_376 vpwr vgnd scs8hd_fill_2
XFILLER_70_357 vgnd vpwr scs8hd_decap_8
XFILLER_70_346 vgnd vpwr scs8hd_decap_8
XPHY_736 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_725 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_714 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_703 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_769 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_758 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_747 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_7_428 vgnd vpwr scs8hd_decap_3
XFILLER_23_98 vgnd vpwr scs8hd_decap_12
XFILLER_2_166 vgnd vpwr scs8hd_decap_12
XFILLER_78_468 vgnd vpwr scs8hd_decap_12
XFILLER_19_502 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mux_fle_0_in_0.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_0_in_0.INVTX1_13_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_46_332 vpwr vgnd scs8hd_fill_2
XFILLER_34_505 vgnd vpwr scs8hd_decap_8
XFILLER_46_365 vpwr vgnd scs8hd_fill_2
XFILLER_73_184 vgnd vpwr scs8hd_decap_3
XFILLER_61_313 vgnd vpwr scs8hd_decap_3
XFILLER_46_398 vgnd vpwr scs8hd_decap_4
XANTENNA_ltile_clb_0.mux_fle_2_in_0.INVTX1_11_.scs8hd_inv_1_A left_width_0_height_0__pin_11_
+ vgnd vpwr scs8hd_diode_2
XFILLER_14_284 vgnd vpwr scs8hd_decap_3
XFILLER_80_93 vgnd vpwr scs8hd_decap_12
X_328_ _328_/A _374_/A vgnd vpwr scs8hd_buf_1
XANTENNA_ltile_clb_0.mux_fle_2_in_3.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_2_in_3.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
X_259_ _258_/X _259_/B _286_/B _333_/A vgnd vpwr scs8hd_or3_4
XFILLER_6_472 vpwr vgnd scs8hd_fill_2
XFILLER_43_3 vgnd vpwr scs8hd_decap_12
XFILLER_56_129 vgnd vpwr scs8hd_decap_6
XANTENNA_ltile_clb_0.mux_fle_0_in_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_0_in_1.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_37_376 vpwr vgnd scs8hd_fill_2
XFILLER_37_387 vpwr vgnd scs8hd_fill_2
XFILLER_52_346 vgnd vpwr scs8hd_decap_3
Xltile_clb_0.mux_fle_3_in_0.INVTX1_0_.scs8hd_inv_1 top_width_0_height_0__pin_0_ ltile_clb_0.mux_fle_3_in_0.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_69_39 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_1_.scs8hd_inv_1
+ ltile_clb_0.mux_fle_2_in_1.INVTX1_14_.scs8hd_inv_1/Y _615_/A vgnd vpwr scs8hd_inv_1
XANTENNA_ltile_clb_0.mux_fle_3_in_3.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_3_in_3.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_15_.latch_SLEEPB
+ _244_/Y vgnd vpwr scs8hd_diode_2
XFILLER_18_32 vgnd vpwr scs8hd_decap_12
XFILLER_28_332 vpwr vgnd scs8hd_fill_2
XFILLER_55_140 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.mux_fle_2_in_0.INVTX1_9_.scs8hd_inv_1 right_width_0_height_0__pin_9_
+ ltile_clb_0.mux_fle_2_in_0.INVTX1_9_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XFILLER_28_376 vgnd vpwr scs8hd_decap_3
XFILLER_70_154 vpwr vgnd scs8hd_fill_2
XFILLER_55_195 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_2_.TGATE_1_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_2_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XPHY_500 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_511 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_522 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_533 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_544 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_11_221 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_1_.TGATE_1_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_3_.TGATE_1_.scs8hd_ebufn_2/Z
+ _624_/Y ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XPHY_555 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_566 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_577 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_599 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_588 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_7_236 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.mux_fle_0_in_3.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_0_in_3.INVTX1_3_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_0_in_3.LATCH_3_.latch/Q ltile_clb_0.mux_fle_0_in_3.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_ltile_clb_0.mux_fle_2_in_1.INVTX1_7_.scs8hd_inv_1_A left_width_0_height_0__pin_7_
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_1_in_0.mux_l1_in_3_.TGATE_2_.scs8hd_ebufn_2 _644_/HI ltile_clb_0.mem_fle_1_in_0.LATCH_2_.latch/Q
+ ltile_clb_0.mux_fle_1_in_0.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XFILLER_7_258 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_5_.TGATE_1_.scs8hd_ebufn_2_TEB
+ _612_/Y vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_3_in_0.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_3_in_0.INVTX1_9_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_3_in_0.LATCH_1_.latch/Q ltile_clb_0.mux_fle_3_in_0.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA__402__B _399_/B vgnd vpwr scs8hd_diode_2
XFILLER_78_276 vgnd vpwr scs8hd_decap_4
XFILLER_66_416 vpwr vgnd scs8hd_fill_2
XFILLER_38_129 vgnd vpwr scs8hd_decap_12
XFILLER_61_110 vgnd vpwr scs8hd_decap_12
XFILLER_19_376 vpwr vgnd scs8hd_fill_2
XFILLER_19_387 vpwr vgnd scs8hd_fill_2
XFILLER_19_398 vpwr vgnd scs8hd_fill_2
XFILLER_34_346 vgnd vpwr scs8hd_decap_3
XFILLER_34_357 vgnd vpwr scs8hd_fill_1
XFILLER_42_390 vgnd vpwr scs8hd_decap_6
XANTENNA__312__B _309_/X vgnd vpwr scs8hd_diode_2
XFILLER_57_449 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_3_in_2.INVTX1_4_.scs8hd_inv_1_A top_width_0_height_0__pin_4_
+ vgnd vpwr scs8hd_diode_2
XFILLER_37_151 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_14_.scs8hd_inv_1
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_14_.latch/Q
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_14_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_25_346 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.mux_fle_3_in_1.INVTX1_4_.scs8hd_inv_1 top_width_0_height_0__pin_4_ ltile_clb_0.mux_fle_3_in_1.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_52_165 vgnd vpwr scs8hd_decap_12
XFILLER_25_379 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_0_in_1.mux_l1_in_2_.TGATE_3_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_0_in_1.INVTX1_11_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_40_305 vpwr vgnd scs8hd_fill_2
XANTENNA__503__A _343_/A vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mem_fle_2_in_3.LATCH_7_.latch_SLEEPB _388_/Y vgnd vpwr scs8hd_diode_2
XFILLER_20_44 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mux_fle_2_in_2.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_2_in_2.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_29_86 vgnd vpwr scs8hd_decap_12
XFILLER_48_449 vpwr vgnd scs8hd_fill_2
XFILLER_56_493 vgnd vpwr scs8hd_decap_12
XFILLER_56_482 vgnd vpwr scs8hd_decap_8
X_593_ _541_/A _588_/X _593_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_28_195 vpwr vgnd scs8hd_fill_2
XFILLER_43_110 vgnd vpwr scs8hd_decap_12
XFILLER_45_74 vgnd vpwr scs8hd_decap_12
XFILLER_71_485 vgnd vpwr scs8hd_decap_3
Xltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_2_.scs8hd_inv_1
+ ltile_clb_0.mux_fle_0_in_2.INVTX1_14_.scs8hd_inv_1/Y _633_/A vgnd vpwr scs8hd_inv_1
XPHY_330 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_341 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_352 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_61_51 vgnd vpwr scs8hd_decap_8
XPHY_363 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_374 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_385 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_61_62 vgnd vpwr scs8hd_decap_12
XPHY_396 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_ltile_clb_0.mux_fle_2_in_1.mux_l1_in_2_.TGATE_3_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_2_in_1.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_3_.scs8hd_inv_1/Y
+ _604_/Y ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_6_68 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.mux_fle_0_in_0.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_0_in_0.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2/Z
+ ltile_clb_0.mem_fle_0_in_0.LATCH_7_.latch/Q ltile_clb_0.mux_fle_0_in_0.INVTX1_14_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA__413__A _325_/A vgnd vpwr scs8hd_diode_2
XFILLER_3_283 vgnd vpwr scs8hd_decap_8
XFILLER_66_202 vgnd vpwr scs8hd_fill_1
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.INVTX1_0_.scs8hd_inv_1_A
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.INVTX1_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_0_in_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_0_in_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_66_224 vgnd vpwr scs8hd_decap_12
XFILLER_39_449 vpwr vgnd scs8hd_fill_2
XFILLER_66_257 vgnd vpwr scs8hd_fill_1
XFILLER_19_173 vgnd vpwr scs8hd_decap_6
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_47_482 vgnd vpwr scs8hd_fill_1
XFILLER_19_184 vpwr vgnd scs8hd_fill_2
XFILLER_62_474 vgnd vpwr scs8hd_fill_1
XFILLER_34_154 vgnd vpwr scs8hd_decap_12
XFILLER_30_393 vgnd vpwr scs8hd_fill_1
XANTENNA__323__A _388_/A vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_1_in_3.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_1_in_3.INVTX1_8_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_57_213 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.mux_fle_3_in_2.INVTX1_8_.scs8hd_inv_1 top_width_0_height_0__pin_8_ ltile_clb_0.mux_fle_3_in_2.INVTX1_8_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_72_205 vgnd vpwr scs8hd_decap_8
XFILLER_38_471 vgnd vpwr scs8hd_fill_1
XFILLER_25_110 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mem_fle_3_in_2.LATCH_7_.latch_SLEEPB _349_/Y vgnd vpwr scs8hd_diode_2
XFILLER_53_496 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.mux_fle_0_in_1.mux_l1_in_3_.TGATE_2_.scs8hd_ebufn_2 _641_/HI ltile_clb_0.mem_fle_0_in_1.LATCH_2_.latch/Q
+ ltile_clb_0.mux_fle_0_in_1.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
Xltile_clb_0.mux_fle_2_in_1.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_2_in_1.INVTX1_9_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_2_in_1.LATCH_1_.latch/Q ltile_clb_0.mux_fle_2_in_1.mux_l1_in_2_.TGATE_3_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
Xltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_6_.latch
+ data_in ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_6_.latch/Q
+ _285_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_9_.latch_SLEEPB
+ _563_/Y vgnd vpwr scs8hd_diode_2
XANTENNA__233__A _232_/X vgnd vpwr scs8hd_diode_2
XFILLER_31_98 vgnd vpwr scs8hd_decap_12
XFILLER_48_202 vpwr vgnd scs8hd_fill_2
XFILLER_36_419 vgnd vpwr scs8hd_decap_6
XFILLER_48_279 vgnd vpwr scs8hd_decap_12
X_645_ _645_/HI _645_/LO vgnd vpwr scs8hd_conb_1
XFILLER_16_154 vgnd vpwr scs8hd_decap_12
X_576_ _270_/B _575_/B _576_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_44_474 vgnd vpwr scs8hd_decap_8
XANTENNA__408__A address[6] vgnd vpwr scs8hd_diode_2
XFILLER_16_187 vgnd vpwr scs8hd_decap_3
XPHY_160 vgnd vpwr scs8hd_decap_3
XFILLER_31_135 vgnd vpwr scs8hd_decap_12
XFILLER_12_371 vpwr vgnd scs8hd_fill_2
XPHY_171 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_182 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_193 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_31_179 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_0_in_2.INVTX1_2_.scs8hd_inv_1_A bottom_width_0_height_0__pin_2_
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_3_in_2.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_3_in_2.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_79_360 vgnd vpwr scs8hd_decap_4
XFILLER_79_393 vgnd vpwr scs8hd_decap_6
XFILLER_79_382 vpwr vgnd scs8hd_fill_2
XFILLER_27_419 vpwr vgnd scs8hd_fill_2
XFILLER_47_290 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_2_.TGATE_1_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_2_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_35_496 vpwr vgnd scs8hd_fill_2
XANTENNA__318__A enable vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_3_in_1.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_3_in_1.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.mem_ble4_out_0.LATCH_0_.latch_SLEEPB
+ _577_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__ff_0.DFFSRQ_0_.dff_SETB
+ set vgnd vpwr scs8hd_diode_2
XFILLER_77_39 vgnd vpwr scs8hd_decap_12
XANTENNA__500__B _495_/X vgnd vpwr scs8hd_diode_2
XFILLER_26_32 vgnd vpwr scs8hd_decap_12
XFILLER_38_290 vgnd vpwr scs8hd_decap_4
X_430_ _430_/A _429_/X _430_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_60_219 vgnd vpwr scs8hd_decap_8
XFILLER_41_400 vpwr vgnd scs8hd_fill_2
X_361_ _388_/A _365_/B _361_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA__228__A _227_/X vgnd vpwr scs8hd_diode_2
XFILLER_13_135 vgnd vpwr scs8hd_decap_12
XFILLER_41_444 vpwr vgnd scs8hd_fill_2
X_292_ _267_/X _542_/A _292_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_5_356 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_0_in_3.INVTX1_11_.scs8hd_inv_1_A left_width_0_height_0__pin_11_
+ vgnd vpwr scs8hd_diode_2
XFILLER_5_367 vgnd vpwr scs8hd_decap_3
XFILLER_76_341 vgnd vpwr scs8hd_decap_6
XFILLER_76_396 vgnd vpwr scs8hd_fill_1
X_628_ _628_/A _628_/Y vgnd vpwr scs8hd_inv_8
XFILLER_51_208 vpwr vgnd scs8hd_fill_2
X_559_ _559_/A _558_/B _559_/Y vgnd vpwr scs8hd_nor2_4
Xltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_2_.TGATE_0_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_4_.TGATE_1_.scs8hd_ebufn_2/Z
+ _615_/Y ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_1_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_73_3 vgnd vpwr scs8hd_decap_12
XANTENNA__601__A _575_/A vgnd vpwr scs8hd_diode_2
XANTENNA__320__B _369_/B vgnd vpwr scs8hd_diode_2
XFILLER_82_311 vgnd vpwr scs8hd_decap_12
XFILLER_55_514 vpwr vgnd scs8hd_fill_2
XFILLER_82_366 vgnd vpwr scs8hd_decap_6
XANTENNA_ltile_clb_0.mux_fle_2_in_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_2_in_0.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_6_.latch
+ data_in ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_6_.latch/Q
+ _592_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
Xltile_clb_0.mux_fle_1_in_2.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_1_in_2.INVTX1_9_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_1_in_2.LATCH_1_.latch/Q ltile_clb_0.mux_fle_1_in_2.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
Xltile_clb_0.mux_fle_3_in_2.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_3_in_2.INVTX1_4_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_3_in_2.LATCH_0_.latch/Q ltile_clb_0.mux_fle_3_in_2.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_23_455 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_0_.scs8hd_inv_1_A
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_10_105 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mux_fle_2_in_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_2_in_0.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_4_.scs8hd_inv_1
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_4_.latch/Q
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_12_56 vgnd vpwr scs8hd_decap_12
XFILLER_2_359 vgnd vpwr scs8hd_decap_6
XANTENNA__511__A _334_/A vgnd vpwr scs8hd_diode_2
XANTENNA__230__B address[5] vgnd vpwr scs8hd_diode_2
XFILLER_18_205 vgnd vpwr scs8hd_decap_8
XFILLER_58_396 vgnd vpwr scs8hd_fill_1
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_15_.scs8hd_inv_1_A
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_15_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_61_506 vgnd vpwr scs8hd_decap_8
XFILLER_37_86 vgnd vpwr scs8hd_decap_12
XFILLER_26_260 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_0_in_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_0_in_1.LATCH_5_.latch/Q
+ vgnd vpwr scs8hd_diode_2
X_413_ _325_/A _431_/A vgnd vpwr scs8hd_buf_1
XFILLER_14_433 vpwr vgnd scs8hd_fill_2
X_344_ _379_/A _341_/B _344_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_53_74 vgnd vpwr scs8hd_decap_12
XFILLER_41_274 vpwr vgnd scs8hd_fill_2
X_275_ _236_/X _342_/A _276_/A vgnd vpwr scs8hd_or2_4
XANTENNA__405__B _398_/A vgnd vpwr scs8hd_diode_2
XANTENNA__421__A _421_/A vgnd vpwr scs8hd_diode_2
XFILLER_78_93 vgnd vpwr scs8hd_decap_12
XFILLER_68_105 vgnd vpwr scs8hd_decap_12
XFILLER_49_341 vpwr vgnd scs8hd_fill_2
XFILLER_64_311 vpwr vgnd scs8hd_fill_2
XFILLER_17_271 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_14_.latch_SLEEPB
+ _583_/Y vgnd vpwr scs8hd_diode_2
XFILLER_32_285 vgnd vpwr scs8hd_decap_3
XANTENNA__331__A _331_/A vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_55_322 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2_TEB
+ _604_/Y vgnd vpwr scs8hd_diode_2
XFILLER_15_208 vpwr vgnd scs8hd_fill_2
XPHY_726 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_715 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_704 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_23_241 vgnd vpwr scs8hd_fill_1
XANTENNA_ltile_clb_0.mux_fle_2_in_0.mux_l1_in_2_.TGATE_3_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_2_in_0.INVTX1_11_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XPHY_759 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_748 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_737 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_11_447 vpwr vgnd scs8hd_fill_2
XFILLER_23_285 vpwr vgnd scs8hd_fill_2
XANTENNA__506__A _514_/B vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_0_in_0.INVTX1_8_.scs8hd_inv_1 top_width_0_height_0__pin_8_ ltile_clb_0.mux_fle_0_in_0.INVTX1_8_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_ltile_clb_0.mux_fle_1_in_2.INVTX1_8_.scs8hd_inv_1_A top_width_0_height_0__pin_8_
+ vgnd vpwr scs8hd_diode_2
XFILLER_3_3 vgnd vpwr scs8hd_decap_12
XANTENNA__241__A _286_/A vgnd vpwr scs8hd_diode_2
XFILLER_78_414 vgnd vpwr scs8hd_fill_1
XFILLER_2_178 vgnd vpwr scs8hd_decap_12
XFILLER_78_447 vgnd vpwr scs8hd_fill_1
XFILLER_19_514 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_2_in_3.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_2_in_3.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_0_15 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mux_fle_3_in_0.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_3_in_0.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.INVTX1_1_.scs8hd_inv_1/Y
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.mem_ble4_out_0.LATCH_1_.latch/Q
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
Xltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_9_.scs8hd_inv_1
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_9_.latch/Q
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_9_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_46_388 vgnd vpwr scs8hd_decap_8
XFILLER_14_263 vgnd vpwr scs8hd_decap_12
XANTENNA__416__A _432_/A vgnd vpwr scs8hd_diode_2
X_327_ _286_/X _328_/A vgnd vpwr scs8hd_buf_1
X_258_ address[2] _258_/X vgnd vpwr scs8hd_buf_1
XFILLER_10_491 vgnd vpwr scs8hd_fill_1
XFILLER_36_3 vgnd vpwr scs8hd_decap_12
XFILLER_69_447 vgnd vpwr scs8hd_decap_3
Xltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_6_.latch
+ data_in ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_6_.latch/Q
+ _566_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_ltile_clb_0.mux_fle_2_in_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_2_in_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_2_.latch_SLEEPB
+ _596_/Y vgnd vpwr scs8hd_diode_2
XFILLER_49_160 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.mux_fle_2_in_3.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_2_in_3.INVTX1_4_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_2_in_3.LATCH_0_.latch/Q ltile_clb_0.mux_fle_2_in_3.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_64_141 vgnd vpwr scs8hd_fill_1
XANTENNA_ltile_clb_0.mux_fle_3_in_2.INVTX1_14_.scs8hd_inv_1_A ltile_clb_0.mux_fle_3_in_2.INVTX1_14_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_0_in_3.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_0_in_3.INVTX1_9_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_0_in_3.LATCH_1_.latch/Q ltile_clb_0.mux_fle_0_in_3.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_ltile_clb_0.mux_fle_2_in_3.INVTX1_5_.scs8hd_inv_1_A right_width_0_height_0__pin_5_
+ vgnd vpwr scs8hd_diode_2
XFILLER_64_174 vgnd vpwr scs8hd_decap_6
XFILLER_40_509 vgnd vpwr scs8hd_decap_6
XANTENNA__326__A _326_/A vgnd vpwr scs8hd_diode_2
XFILLER_20_222 vgnd vpwr scs8hd_decap_3
XANTENNA_ltile_clb_0.mux_fle_3_in_0.INVTX1_1_.scs8hd_inv_1_A right_width_0_height_0__pin_1_
+ vgnd vpwr scs8hd_diode_2
XFILLER_20_255 vgnd vpwr scs8hd_decap_3
Xltile_clb_0.mux_fle_1_in_1.INVTX1_3_.scs8hd_inv_1 left_width_0_height_0__pin_3_ ltile_clb_0.mux_fle_1_in_1.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_ltile_clb_0.mux_fle_3_in_2.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_3_in_2.INVTX1_8_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_2_.scs8hd_inv_1_A
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_68_480 vgnd vpwr scs8hd_decap_12
XFILLER_18_44 vgnd vpwr scs8hd_decap_12
XFILLER_28_344 vgnd vpwr scs8hd_decap_6
XFILLER_55_163 vgnd vpwr scs8hd_decap_3
XPHY_501 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_43_358 vpwr vgnd scs8hd_fill_2
XFILLER_34_32 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mem_fle_0_in_0.LATCH_6_.latch_D data_in vgnd vpwr scs8hd_diode_2
XPHY_512 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_523 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_534 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__236__A _246_/A vgnd vpwr scs8hd_diode_2
XPHY_545 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_556 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_567 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_578 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_ltile_clb_0.mux_fle_1_in_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_1_in_0.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XPHY_589 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_3_421 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.mux_fle_2_in_0.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_2_in_0.INVTX1_3_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_2_in_0.LATCH_3_.latch/Q ltile_clb_0.mux_fle_2_in_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_59_62 vgnd vpwr scs8hd_decap_12
XFILLER_59_51 vgnd vpwr scs8hd_decap_8
XFILLER_3_487 vgnd vpwr scs8hd_fill_1
XANTENNA_ltile_clb_0.mem_fle_0_in_1.LATCH_4_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB
+ _622_/Y vgnd vpwr scs8hd_diode_2
XFILLER_46_141 vgnd vpwr scs8hd_fill_1
XANTENNA_ltile_clb_0.mux_fle_1_in_2.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_1_in_2.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_46_163 vgnd vpwr scs8hd_decap_3
XFILLER_61_144 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.mux_fle_3_in_0.INVTX1_14_.scs8hd_inv_1 ltile_clb_0.mux_fle_3_in_0.INVTX1_14_.scs8hd_inv_1/A
+ ltile_clb_0.mux_fle_3_in_0.INVTX1_14_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XFILLER_61_188 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mem_fle_0_in_2.LATCH_2_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_3_in_3.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_3_in_3.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_57_428 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.mem_ble4_out_0.LATCH_0_.latch_SLEEPB
+ _603_/Y vgnd vpwr scs8hd_diode_2
XFILLER_72_409 vgnd vpwr scs8hd_decap_4
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__ff_0.DFFSRQ_0_.dff_D
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.INVTX1_1_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_37_141 vgnd vpwr scs8hd_fill_1
XANTENNA_ltile_clb_0.mem_fle_0_in_3.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_25_358 vpwr vgnd scs8hd_fill_2
XFILLER_52_177 vgnd vpwr scs8hd_decap_3
XFILLER_40_317 vpwr vgnd scs8hd_fill_2
XFILLER_40_328 vgnd vpwr scs8hd_decap_3
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_6_.TGATE_0_.scs8hd_ebufn_2_TEB
+ _613_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_6_.latch_D
+ data_in vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_1_in_2.INVTX1_7_.scs8hd_inv_1 left_width_0_height_0__pin_7_ ltile_clb_0.mux_fle_1_in_2.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_4_229 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l4_in_0_.TGATE_0_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l4_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_20_56 vgnd vpwr scs8hd_decap_12
XANTENNA__503__B _502_/B vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mem_fle_1_in_0.LATCH_2_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_0_435 vgnd vpwr scs8hd_decap_4
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_13_.latch_D
+ data_in vgnd vpwr scs8hd_diode_2
XFILLER_28_141 vgnd vpwr scs8hd_decap_12
XFILLER_29_98 vgnd vpwr scs8hd_decap_12
XFILLER_56_472 vgnd vpwr scs8hd_fill_1
X_592_ _540_/A _588_/X _592_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_16_325 vgnd vpwr scs8hd_decap_6
XFILLER_16_358 vgnd vpwr scs8hd_decap_8
XFILLER_71_453 vpwr vgnd scs8hd_fill_2
XFILLER_45_86 vgnd vpwr scs8hd_decap_12
XPHY_320 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_331 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_342 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_31_339 vpwr vgnd scs8hd_fill_2
XFILLER_43_199 vgnd vpwr scs8hd_decap_4
Xltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_7_.TGATE_0_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_14_.scs8hd_inv_1/Y
+ _605_/Y ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_3_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XPHY_353 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_364 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_391 vgnd vpwr scs8hd_decap_4
XPHY_375 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_386 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_ltile_clb_0.mem_fle_1_in_1.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mem_fle_3_in_3.LATCH_1_.latch_SLEEPB _341_/Y vgnd vpwr scs8hd_diode_2
XFILLER_61_74 vgnd vpwr scs8hd_decap_12
XPHY_397 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_6_.latch
+ data_in ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_6_.latch/Q
+ _540_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_ltile_clb_0.mux_fle_1_in_0.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_1_in_0.INVTX1_13_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_3_262 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_1_in_1.INVTX1_13_.scs8hd_inv_1_A right_width_0_height_0__pin_13_
+ vgnd vpwr scs8hd_diode_2
XFILLER_39_406 vpwr vgnd scs8hd_fill_2
XFILLER_39_428 vpwr vgnd scs8hd_fill_2
XFILLER_62_442 vpwr vgnd scs8hd_fill_2
XFILLER_62_431 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_3_in_3.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_3_in_3.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_34_166 vgnd vpwr scs8hd_decap_6
XFILLER_15_391 vpwr vgnd scs8hd_fill_2
XFILLER_30_383 vpwr vgnd scs8hd_fill_2
XANTENNA__604__A _604_/A vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_2_in_3.INVTX1_2_.scs8hd_inv_1 bottom_width_0_height_0__pin_2_
+ ltile_clb_0.mux_fle_2_in_3.INVTX1_2_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XANTENNA__323__B _338_/B vgnd vpwr scs8hd_diode_2
Xltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_10_.latch
+ data_in ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_10_.latch/Q
+ _561_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_ltile_clb_0.mux_fle_1_in_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_1_in_1.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_2_in_2.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_2_in_2.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_57_269 vpwr vgnd scs8hd_fill_2
XFILLER_57_258 vpwr vgnd scs8hd_fill_2
XFILLER_53_475 vpwr vgnd scs8hd_fill_2
XFILLER_53_464 vpwr vgnd scs8hd_fill_2
XFILLER_80_272 vgnd vpwr scs8hd_decap_3
XFILLER_25_199 vpwr vgnd scs8hd_fill_2
XFILLER_21_350 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_2_in_1.mux_l1_in_3_.TGATE_2_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_2_in_1.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__514__A _343_/A vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_4_.scs8hd_inv_1_A
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_4_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_0_in_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_0_in_3.LATCH_4_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_1_in_1.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_1_in_1.INVTX1_3_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_1_in_1.LATCH_3_.latch/Q ltile_clb_0.mux_fle_1_in_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_2_.latch_D
+ data_in vgnd vpwr scs8hd_diode_2
X_644_ _644_/HI _644_/LO vgnd vpwr scs8hd_conb_1
XFILLER_29_472 vgnd vpwr scs8hd_decap_3
XFILLER_44_420 vgnd vpwr scs8hd_decap_8
XFILLER_44_431 vpwr vgnd scs8hd_fill_2
XFILLER_71_250 vpwr vgnd scs8hd_fill_2
XFILLER_16_166 vgnd vpwr scs8hd_decap_12
X_575_ _575_/A _575_/B _575_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_44_497 vgnd vpwr scs8hd_decap_4
XPHY_161 vgnd vpwr scs8hd_decap_3
XPHY_150 vgnd vpwr scs8hd_decap_3
Xltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_7_.scs8hd_inv_1/Y
+ _612_/Y ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_1_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_31_147 vgnd vpwr scs8hd_decap_12
XFILLER_12_361 vgnd vpwr scs8hd_fill_1
XFILLER_8_310 vpwr vgnd scs8hd_fill_2
XPHY_172 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_183 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_194 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__424__A _436_/A vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_2_in_1.INVTX1_10_.scs8hd_inv_1 bottom_width_0_height_0__pin_10_
+ ltile_clb_0.mux_fle_2_in_1.INVTX1_10_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XANTENNA_ltile_clb_0.mux_fle_3_in_3.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_3_in_3.LATCH_7_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_8_387 vgnd vpwr scs8hd_decap_8
Xltile_clb_0.mem_fle_1_in_1.LATCH_7_.latch data_in ltile_clb_0.mem_fle_1_in_1.LATCH_7_.latch/Q
+ _463_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_67_501 vgnd vpwr scs8hd_decap_12
XFILLER_39_214 vgnd vpwr scs8hd_decap_4
XFILLER_39_225 vpwr vgnd scs8hd_fill_2
XFILLER_39_236 vgnd vpwr scs8hd_decap_4
XFILLER_82_515 vgnd vpwr scs8hd_fill_1
XFILLER_54_228 vgnd vpwr scs8hd_decap_6
XFILLER_35_420 vgnd vpwr scs8hd_fill_1
Xltile_clb_0.mem_fle_2_in_1.LATCH_6_.latch data_in ltile_clb_0.mem_fle_2_in_1.LATCH_6_.latch/Q
+ _414_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_ltile_clb_0.mem_fle_1_in_3.LATCH_2_.latch_SLEEPB _446_/Y vgnd vpwr scs8hd_diode_2
XANTENNA__318__B address[5] vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__334__A _334_/A vgnd vpwr scs8hd_diode_2
XFILLER_2_508 vgnd vpwr scs8hd_decap_8
Xltile_clb_0.mux_fle_2_in_2.INVTX1_12_.scs8hd_inv_1 top_width_0_height_0__pin_12_
+ ltile_clb_0.mux_fle_2_in_2.INVTX1_12_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
Xltile_clb_0.mem_fle_3_in_1.LATCH_5_.latch data_in ltile_clb_0.mem_fle_3_in_1.LATCH_5_.latch/Q
+ _363_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_77_309 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_1_in_1.mux_l1_in_2_.TGATE_3_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_1_in_1.INVTX1_11_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_26_431 vpwr vgnd scs8hd_fill_2
XFILLER_53_250 vpwr vgnd scs8hd_fill_2
XFILLER_26_44 vgnd vpwr scs8hd_decap_12
XANTENNA__509__A _328_/A vgnd vpwr scs8hd_diode_2
X_360_ _368_/B _365_/B vgnd vpwr scs8hd_buf_1
XFILLER_13_147 vgnd vpwr scs8hd_decap_12
XFILLER_41_467 vpwr vgnd scs8hd_fill_2
X_291_ _290_/X _542_/A vgnd vpwr scs8hd_buf_1
XFILLER_42_32 vgnd vpwr scs8hd_decap_12
XANTENNA__244__A _248_/A vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_1_in_0.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_1_in_0.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_13_.latch_SLEEPB
+ _558_/Y vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_3_in_0.INVTX1_8_.scs8hd_inv_1 top_width_0_height_0__pin_8_ ltile_clb_0.mux_fle_3_in_0.INVTX1_8_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_3_15 vgnd vpwr scs8hd_decap_12
XFILLER_67_51 vgnd vpwr scs8hd_decap_8
XFILLER_3_59 vpwr vgnd scs8hd_fill_2
XFILLER_67_62 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.mux_fle_2_in_3.INVTX1_14_.scs8hd_inv_1 ltile_clb_0.mux_fle_2_in_3.INVTX1_14_.scs8hd_inv_1/A
+ ltile_clb_0.mux_fle_2_in_3.INVTX1_14_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XFILLER_64_515 vgnd vpwr scs8hd_fill_1
XFILLER_36_206 vpwr vgnd scs8hd_fill_2
XFILLER_29_280 vpwr vgnd scs8hd_fill_2
X_627_ _627_/A _627_/Y vgnd vpwr scs8hd_inv_8
XFILLER_17_442 vpwr vgnd scs8hd_fill_2
XANTENNA__419__A _334_/A vgnd vpwr scs8hd_diode_2
XFILLER_17_486 vpwr vgnd scs8hd_fill_2
X_558_ _250_/X _558_/B _558_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA_ltile_clb_0.mem_fle_1_in_3.LATCH_6_.latch_D data_in vgnd vpwr scs8hd_diode_2
X_489_ _334_/A _484_/X _489_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_12_180 vgnd vpwr scs8hd_decap_8
XFILLER_66_3 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mux_fle_1_in_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_1_in_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_0_.TGATE_1_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ _608_/Y ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l4_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l4_in_0_.TGATE_0_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l4_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mem_fle_2_in_2.LATCH_2_.latch_SLEEPB _404_/Y vgnd vpwr scs8hd_diode_2
XFILLER_59_309 vpwr vgnd scs8hd_fill_2
XANTENNA__601__B _600_/X vgnd vpwr scs8hd_diode_2
XANTENNA__320__C _346_/C vgnd vpwr scs8hd_diode_2
XFILLER_82_323 vgnd vpwr scs8hd_decap_12
XANTENNA__329__A _374_/A vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_3_in_0.INVTX1_11_.scs8hd_inv_1_A left_width_0_height_0__pin_11_
+ vgnd vpwr scs8hd_diode_2
XFILLER_23_423 vpwr vgnd scs8hd_fill_2
XFILLER_35_272 vgnd vpwr scs8hd_decap_4
XFILLER_10_117 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.mux_fle_0_in_2.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_0_in_2.INVTX1_3_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_0_in_2.LATCH_3_.latch/Q ltile_clb_0.mux_fle_0_in_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_ltile_clb_0.mem_fle_2_in_1.LATCH_6_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_2_in_3.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_2_in_3.INVTX1_8_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_12_68 vgnd vpwr scs8hd_decap_12
XFILLER_2_305 vpwr vgnd scs8hd_fill_2
XFILLER_2_327 vgnd vpwr scs8hd_decap_8
XANTENNA_ltile_clb_0.mux_fle_0_in_3.INVTX1_9_.scs8hd_inv_1_A right_width_0_height_0__pin_9_
+ vgnd vpwr scs8hd_diode_2
XANTENNA__511__B _511_/B vgnd vpwr scs8hd_diode_2
XFILLER_58_331 vpwr vgnd scs8hd_fill_2
XFILLER_73_301 vpwr vgnd scs8hd_fill_2
XFILLER_58_364 vgnd vpwr scs8hd_fill_1
XFILLER_58_353 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_1_in_0.INVTX1_5_.scs8hd_inv_1_A right_width_0_height_0__pin_5_
+ vgnd vpwr scs8hd_diode_2
XFILLER_18_228 vgnd vpwr scs8hd_fill_1
XANTENNA_ltile_clb_0.mux_fle_0_in_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_0_in_1.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_73_356 vpwr vgnd scs8hd_fill_2
XFILLER_73_345 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mem_fle_2_in_2.LATCH_4_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA__239__A _259_/B vgnd vpwr scs8hd_diode_2
XFILLER_37_98 vgnd vpwr scs8hd_decap_12
X_412_ _430_/A _412_/B _412_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_26_272 vgnd vpwr scs8hd_fill_1
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_41_220 vpwr vgnd scs8hd_fill_2
X_343_ _343_/A _379_/A vgnd vpwr scs8hd_buf_1
XFILLER_53_86 vgnd vpwr scs8hd_decap_12
X_274_ _258_/X _603_/A _342_/A vgnd vpwr scs8hd_or2_4
XFILLER_5_110 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mux_fle_2_in_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_2_in_1.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mem_fle_2_in_3.LATCH_2_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_68_117 vgnd vpwr scs8hd_decap_12
XFILLER_1_382 vgnd vpwr scs8hd_decap_3
XFILLER_49_375 vpwr vgnd scs8hd_fill_2
XFILLER_64_345 vpwr vgnd scs8hd_fill_2
XFILLER_64_389 vpwr vgnd scs8hd_fill_2
XFILLER_64_378 vgnd vpwr scs8hd_decap_8
XANTENNA_ltile_clb_0.mux_fle_1_in_3.mux_l1_in_2_.TGATE_3_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_1_in_3.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_2_in_0.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_2_in_0.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mem_fle_3_in_1.LATCH_2_.latch_SLEEPB _366_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mem_fle_3_in_0.LATCH_4_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_20_459 vgnd vpwr scs8hd_decap_3
XANTENNA_ltile_clb_0.mux_fle_2_in_1.INVTX1_2_.scs8hd_inv_1_A bottom_width_0_height_0__pin_2_
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.mem_ble4_out_0.LATCH_0_.latch_SLEEPB
+ _312_/Y vgnd vpwr scs8hd_diode_2
XANTENNA__612__A _612_/A vgnd vpwr scs8hd_diode_2
XFILLER_4_80 vgnd vpwr scs8hd_decap_12
XFILLER_28_515 vgnd vpwr scs8hd_fill_1
XANTENNA_ltile_clb_0.mem_fle_3_in_1.LATCH_2_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_67_161 vpwr vgnd scs8hd_fill_2
XFILLER_43_507 vpwr vgnd scs8hd_fill_2
XPHY_727 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_716 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_705 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_23_220 vpwr vgnd scs8hd_fill_2
XPHY_749 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_738 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_2_.scs8hd_inv_1_A
+ ltile_clb_0.mux_fle_0_in_2.INVTX1_14_.scs8hd_inv_1/Y vgnd vpwr scs8hd_diode_2
XFILLER_11_404 vpwr vgnd scs8hd_fill_2
XFILLER_23_297 vpwr vgnd scs8hd_fill_2
XFILLER_7_419 vgnd vpwr scs8hd_decap_6
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
+ _614_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mem_fle_3_in_2.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mem_fle_0_in_2.LATCH_3_.latch_SLEEPB _500_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_8_.latch_D
+ data_in vgnd vpwr scs8hd_diode_2
XANTENNA__522__A _334_/A vgnd vpwr scs8hd_diode_2
XANTENNA__241__B _282_/B vgnd vpwr scs8hd_diode_2
XFILLER_78_426 vpwr vgnd scs8hd_fill_2
XFILLER_73_153 vpwr vgnd scs8hd_fill_2
XFILLER_0_27 vgnd vpwr scs8hd_decap_4
XFILLER_61_337 vpwr vgnd scs8hd_fill_2
XFILLER_14_231 vpwr vgnd scs8hd_fill_2
XFILLER_14_242 vgnd vpwr scs8hd_decap_4
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_0_in_1.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_0_in_1.INVTX1_13_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
X_326_ _326_/A _338_/B _326_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA__416__B _412_/B vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
X_257_ _248_/A _559_/A _257_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_6_430 vpwr vgnd scs8hd_fill_2
XANTENNA__432__A _432_/A vgnd vpwr scs8hd_diode_2
XFILLER_6_485 vgnd vpwr scs8hd_decap_4
XFILLER_69_415 vpwr vgnd scs8hd_fill_2
XFILLER_29_3 vgnd vpwr scs8hd_decap_12
XFILLER_77_470 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ _630_/Y ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_4_.TGATE_0_.scs8hd_ebufn_2_TEB
+ _605_/Y vgnd vpwr scs8hd_diode_2
XFILLER_52_359 vgnd vpwr scs8hd_decap_4
XANTENNA__607__A _607_/A vgnd vpwr scs8hd_diode_2
XANTENNA__326__B _338_/B vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_2_in_0.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_2_in_0.INVTX1_9_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_2_in_0.LATCH_1_.latch/Q ltile_clb_0.mux_fle_2_in_0.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_20_201 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mux_fle_0_in_2.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_0_in_2.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_0_in_0.mux_l1_in_3_.TGATE_2_.scs8hd_ebufn_2 _640_/HI ltile_clb_0.mem_fle_0_in_0.LATCH_2_.latch/Q
+ ltile_clb_0.mux_fle_0_in_0.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XFILLER_20_267 vgnd vpwr scs8hd_decap_6
XANTENNA__342__A _342_/A vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_3_in_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_3_in_0.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_2_in_3.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_2_in_3.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mem_fle_0_in_0.LATCH_1_.latch data_in ltile_clb_0.mem_fle_0_in_0.LATCH_1_.latch/Q
+ _524_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_68_492 vgnd vpwr scs8hd_decap_12
XFILLER_28_312 vpwr vgnd scs8hd_fill_2
XFILLER_18_56 vgnd vpwr scs8hd_decap_12
XFILLER_28_356 vgnd vpwr scs8hd_fill_1
XFILLER_55_175 vpwr vgnd scs8hd_fill_2
XFILLER_43_315 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mem_fle_1_in_1.LATCH_3_.latch_SLEEPB _467_/Y vgnd vpwr scs8hd_diode_2
XFILLER_70_167 vpwr vgnd scs8hd_fill_2
XFILLER_34_44 vgnd vpwr scs8hd_decap_12
XPHY_502 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_513 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_524 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_535 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__517__A _516_/X vgnd vpwr scs8hd_diode_2
XFILLER_51_392 vpwr vgnd scs8hd_fill_2
XFILLER_51_370 vpwr vgnd scs8hd_fill_2
XPHY_546 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_557 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_568 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xltile_clb_0.mem_fle_1_in_0.LATCH_0_.latch data_in ltile_clb_0.mem_fle_1_in_0.LATCH_0_.latch/Q
+ _481_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_11_245 vgnd vpwr scs8hd_fill_1
XPHY_579 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_11_267 vgnd vpwr scs8hd_fill_1
XFILLER_50_32 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.mux_fle_3_in_3.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_3_in_3.INVTX1_10_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_3_in_3.LATCH_2_.latch/Q ltile_clb_0.mux_fle_3_in_3.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA__252__A _282_/C vgnd vpwr scs8hd_diode_2
XFILLER_3_455 vpwr vgnd scs8hd_fill_2
XFILLER_59_74 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_0_.scs8hd_inv_1
+ ltile_clb_0.mux_fle_1_in_0.INVTX1_14_.scs8hd_inv_1/Y _621_/A vgnd vpwr scs8hd_inv_1
XFILLER_78_267 vgnd vpwr scs8hd_decap_8
XFILLER_66_407 vgnd vpwr scs8hd_decap_3
XFILLER_59_492 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_4_.latch_D
+ data_in vgnd vpwr scs8hd_diode_2
XFILLER_19_301 vpwr vgnd scs8hd_fill_2
XFILLER_75_62 vgnd vpwr scs8hd_decap_12
XFILLER_75_51 vgnd vpwr scs8hd_decap_8
XFILLER_19_367 vpwr vgnd scs8hd_fill_2
XFILLER_34_304 vpwr vgnd scs8hd_fill_2
XFILLER_61_123 vgnd vpwr scs8hd_decap_6
XFILLER_46_186 vgnd vpwr scs8hd_decap_8
XFILLER_61_167 vpwr vgnd scs8hd_fill_2
XANTENNA__427__A _409_/A vgnd vpwr scs8hd_diode_2
XFILLER_42_381 vpwr vgnd scs8hd_fill_2
X_309_ _308_/X _309_/X vgnd vpwr scs8hd_buf_1
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_5_.latch_SLEEPB
+ _541_/Y vgnd vpwr scs8hd_diode_2
XFILLER_69_223 vpwr vgnd scs8hd_fill_2
XFILLER_69_256 vgnd vpwr scs8hd_fill_1
XFILLER_65_440 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.mux_fle_0_in_3.INVTX1_1_.scs8hd_inv_1 right_width_0_height_0__pin_1_
+ ltile_clb_0.mux_fle_0_in_3.INVTX1_1_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XFILLER_37_197 vgnd vpwr scs8hd_decap_4
XFILLER_52_145 vgnd vpwr scs8hd_decap_6
XANTENNA__337__A _421_/A vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mem_fle_0_in_2.LATCH_4_.latch data_in ltile_clb_0.mem_fle_0_in_2.LATCH_4_.latch/Q
+ _499_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_ltile_clb_0.mux_fle_0_in_2.mux_l1_in_2_.TGATE_3_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_0_in_2.INVTX1_11_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_20_68 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mem_fle_2_in_0.LATCH_3_.latch_SLEEPB _434_/Y vgnd vpwr scs8hd_diode_2
XFILLER_0_425 vgnd vpwr scs8hd_decap_3
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_3_.TGATE_0_.scs8hd_ebufn_2_TEB
+ _623_/Y vgnd vpwr scs8hd_diode_2
XFILLER_0_458 vgnd vpwr scs8hd_fill_1
XFILLER_0_469 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.mem_fle_1_in_2.LATCH_3_.latch data_in ltile_clb_0.mem_fle_1_in_2.LATCH_3_.latch/Q
+ _456_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_48_407 vpwr vgnd scs8hd_fill_2
XFILLER_75_204 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_1_in_2.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_1_in_2.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_3_in_0.mux_l1_in_2_.TGATE_3_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_3_in_0.INVTX1_11_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
X_591_ _539_/A _588_/X _591_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_16_315 vgnd vpwr scs8hd_fill_1
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_3_.scs8hd_inv_1_A
+ ltile_clb_0.mux_fle_3_in_3.INVTX1_14_.scs8hd_inv_1/Y vgnd vpwr scs8hd_diode_2
XFILLER_16_337 vgnd vpwr scs8hd_decap_4
XFILLER_43_123 vgnd vpwr scs8hd_decap_12
XPHY_310 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__247__A _246_/X vgnd vpwr scs8hd_diode_2
XFILLER_45_98 vgnd vpwr scs8hd_decap_12
XPHY_321 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_332 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_343 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_31_329 vgnd vpwr scs8hd_fill_1
Xltile_clb_0.mem_fle_2_in_2.LATCH_2_.latch data_in ltile_clb_0.mem_fle_2_in_2.LATCH_2_.latch/Q
+ _404_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XPHY_354 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_365 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_376 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_61_86 vgnd vpwr scs8hd_decap_12
XPHY_387 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_398 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_6_15 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_14_.latch
+ data_in ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_14_.latch/Q
+ _531_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_ltile_clb_0.mux_fle_3_in_1.INVTX1_8_.scs8hd_inv_1_A top_width_0_height_0__pin_8_
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mem_fle_3_in_2.LATCH_1_.latch data_in ltile_clb_0.mem_fle_3_in_2.LATCH_1_.latch/Q
+ _355_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_47_462 vgnd vpwr scs8hd_decap_4
XFILLER_62_465 vgnd vpwr scs8hd_decap_3
XANTENNA_ltile_clb_0.mux_fle_0_in_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_0_in_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_1_in_1.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_1_in_1.INVTX1_9_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_1_in_1.LATCH_1_.latch/Q ltile_clb_0.mux_fle_1_in_1.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
Xltile_clb_0.mux_fle_3_in_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_3_in_1.INVTX1_4_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_3_in_1.LATCH_0_.latch/Q ltile_clb_0.mux_fle_3_in_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_15_370 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_1_in_3.INVTX1_11_.scs8hd_inv_1_A left_width_0_height_0__pin_11_
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_3_in_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_3_in_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XANTENNA__620__A _620_/A vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_3_in_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_3_in_0.LATCH_6_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_12_.latch_SLEEPB
+ _533_/Y vgnd vpwr scs8hd_diode_2
XFILLER_57_237 vpwr vgnd scs8hd_fill_2
XFILLER_38_462 vgnd vpwr scs8hd_decap_6
XFILLER_25_123 vgnd vpwr scs8hd_decap_12
XFILLER_80_251 vgnd vpwr scs8hd_decap_8
XFILLER_53_443 vpwr vgnd scs8hd_fill_2
XFILLER_25_167 vpwr vgnd scs8hd_fill_2
XFILLER_53_487 vgnd vpwr scs8hd_fill_1
XFILLER_21_362 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
+ _628_/Y vgnd vpwr scs8hd_diode_2
XFILLER_21_384 vgnd vpwr scs8hd_decap_4
XANTENNA__514__B _514_/B vgnd vpwr scs8hd_diode_2
XANTENNA__530__A _556_/A vgnd vpwr scs8hd_diode_2
XFILLER_0_211 vgnd vpwr scs8hd_decap_4
XFILLER_0_255 vpwr vgnd scs8hd_fill_2
XFILLER_0_222 vgnd vpwr scs8hd_fill_1
X_643_ _643_/HI _643_/LO vgnd vpwr scs8hd_conb_1
XANTENNA_ltile_clb_0.mux_fle_2_in_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_2_in_0.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_71_240 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.mux_fle_1_in_0.INVTX1_7_.scs8hd_inv_1 left_width_0_height_0__pin_7_ ltile_clb_0.mux_fle_1_in_0.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
Xltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.buf4_2_.scs8hd_buf_1
+ ltile_clb_0.mux_fle_2_in_2.INVTX1_14_.scs8hd_inv_1/Y _616_/A vgnd vpwr scs8hd_buf_1
X_574_ _573_/X _575_/B vgnd vpwr scs8hd_buf_1
XFILLER_71_273 vgnd vpwr scs8hd_decap_3
XFILLER_16_178 vgnd vpwr scs8hd_decap_6
XPHY_151 vgnd vpwr scs8hd_decap_3
XPHY_140 vgnd vpwr scs8hd_decap_3
XFILLER_31_159 vgnd vpwr scs8hd_decap_4
XPHY_162 vgnd vpwr scs8hd_decap_3
XFILLER_12_351 vpwr vgnd scs8hd_fill_2
XPHY_173 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_184 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_195 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__424__B _410_/X vgnd vpwr scs8hd_diode_2
XFILLER_8_366 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mem_fle_0_in_0.LATCH_4_.latch_SLEEPB _521_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_2_in_2.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_2_in_2.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__440__A _447_/B vgnd vpwr scs8hd_diode_2
XFILLER_67_513 vgnd vpwr scs8hd_decap_3
XFILLER_11_3 vgnd vpwr scs8hd_decap_12
XFILLER_39_248 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_10_.scs8hd_inv_1_A
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_10_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_62_251 vgnd vpwr scs8hd_decap_4
XFILLER_35_443 vpwr vgnd scs8hd_fill_2
XFILLER_35_465 vgnd vpwr scs8hd_decap_4
XFILLER_50_402 vgnd vpwr scs8hd_decap_3
XANTENNA__615__A _615_/A vgnd vpwr scs8hd_diode_2
XFILLER_30_192 vgnd vpwr scs8hd_decap_8
XANTENNA__350__A _326_/A vgnd vpwr scs8hd_diode_2
Xltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_2_.scs8hd_inv_1/Y
+ _621_/Y ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
Xltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_0_.scs8hd_inv_1
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_0_.latch/Q
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_45_218 vgnd vpwr scs8hd_decap_4
XFILLER_26_410 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_0_in_1.INVTX1_6_.scs8hd_inv_1_A bottom_width_0_height_0__pin_6_
+ vgnd vpwr scs8hd_diode_2
XFILLER_53_240 vpwr vgnd scs8hd_fill_2
XFILLER_26_56 vgnd vpwr scs8hd_decap_12
XANTENNA__509__B _511_/B vgnd vpwr scs8hd_diode_2
XFILLER_26_443 vgnd vpwr scs8hd_decap_3
XFILLER_26_476 vpwr vgnd scs8hd_fill_2
XFILLER_41_413 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.mux_fle_2_in_1.INVTX1_2_.scs8hd_inv_1 bottom_width_0_height_0__pin_2_
+ ltile_clb_0.mux_fle_2_in_1.INVTX1_2_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
X_290_ _278_/X _330_/A _290_/X vgnd vpwr scs8hd_or2_4
XFILLER_13_159 vgnd vpwr scs8hd_decap_8
XFILLER_42_44 vgnd vpwr scs8hd_decap_12
XANTENNA__525__A _343_/A vgnd vpwr scs8hd_diode_2
XANTENNA__244__B _556_/A vgnd vpwr scs8hd_diode_2
XFILLER_5_336 vpwr vgnd scs8hd_fill_2
XANTENNA__260__A _236_/X vgnd vpwr scs8hd_diode_2
XFILLER_3_27 vgnd vpwr scs8hd_decap_12
XFILLER_49_513 vgnd vpwr scs8hd_decap_3
XFILLER_67_74 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.mux_fle_0_in_2.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_0_in_2.INVTX1_9_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_0_in_2.LATCH_1_.latch/Q ltile_clb_0.mux_fle_0_in_2.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_76_398 vgnd vpwr scs8hd_decap_8
Xltile_clb_0.mux_fle_2_in_2.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_2_in_2.INVTX1_4_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_2_in_2.LATCH_0_.latch/Q ltile_clb_0.mux_fle_2_in_2.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_36_229 vpwr vgnd scs8hd_fill_2
X_626_ _626_/A _626_/Y vgnd vpwr scs8hd_inv_8
Xltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_5_.TGATE_1_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_11_.scs8hd_inv_1/Y
+ _620_/Y ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_2_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
Xltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_11_.scs8hd_inv_1
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_11_.latch/Q
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_11_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
X_557_ _247_/X _558_/B _557_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_32_424 vgnd vpwr scs8hd_decap_4
XFILLER_32_457 vgnd vpwr scs8hd_fill_1
XFILLER_44_284 vgnd vpwr scs8hd_decap_4
XFILLER_44_295 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_2_in_0.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_2_in_0.INVTX1_13_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__435__A _435_/A vgnd vpwr scs8hd_diode_2
XFILLER_32_468 vgnd vpwr scs8hd_decap_8
XFILLER_32_479 vgnd vpwr scs8hd_decap_4
X_488_ _331_/A _484_/X _488_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_8_141 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mux_fle_1_in_2.INVTX1_3_.scs8hd_inv_1_A left_width_0_height_0__pin_3_
+ vgnd vpwr scs8hd_diode_2
XFILLER_59_3 vgnd vpwr scs8hd_decap_12
XANTENNA__320__D _358_/D vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_1_.TGATE_0_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_1_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_1_in_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_1_in_1.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_67_343 vpwr vgnd scs8hd_fill_2
XFILLER_82_335 vgnd vpwr scs8hd_decap_6
XFILLER_67_398 vpwr vgnd scs8hd_fill_2
XFILLER_67_387 vpwr vgnd scs8hd_fill_2
XFILLER_27_229 vgnd vpwr scs8hd_decap_4
XANTENNA__329__B _338_/B vgnd vpwr scs8hd_diode_2
XFILLER_23_402 vpwr vgnd scs8hd_fill_2
XFILLER_23_413 vgnd vpwr scs8hd_decap_4
XFILLER_35_284 vpwr vgnd scs8hd_fill_2
XFILLER_50_210 vpwr vgnd scs8hd_fill_2
XFILLER_50_232 vpwr vgnd scs8hd_fill_2
XANTENNA__345__A _345_/A vgnd vpwr scs8hd_diode_2
XFILLER_23_468 vpwr vgnd scs8hd_fill_2
XFILLER_50_243 vpwr vgnd scs8hd_fill_2
XFILLER_50_276 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_2_in_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_2_in_1.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_10_129 vgnd vpwr scs8hd_decap_12
XFILLER_50_287 vgnd vpwr scs8hd_decap_8
XANTENNA_ltile_clb_0.mux_fle_1_in_0.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_1_in_0.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_2_317 vgnd vpwr scs8hd_fill_1
XFILLER_73_313 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.mux_fle_2_in_2.INVTX1_6_.scs8hd_inv_1 bottom_width_0_height_0__pin_6_
+ ltile_clb_0.mux_fle_2_in_2.INVTX1_6_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XFILLER_58_398 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_2_in_3.INVTX1_0_.scs8hd_inv_1_A top_width_0_height_0__pin_0_
+ vgnd vpwr scs8hd_diode_2
XFILLER_26_240 vgnd vpwr scs8hd_decap_8
X_411_ _410_/X _412_/B vgnd vpwr scs8hd_buf_1
XFILLER_14_402 vgnd vpwr scs8hd_decap_4
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l4_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
+ _619_/Y vgnd vpwr scs8hd_diode_2
X_342_ _342_/A _343_/A vgnd vpwr scs8hd_buf_1
XFILLER_41_254 vgnd vpwr scs8hd_decap_3
XFILLER_53_98 vgnd vpwr scs8hd_decap_12
X_273_ _267_/X _272_/X _273_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA__255__A _236_/X vgnd vpwr scs8hd_diode_2
Xltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_5_.scs8hd_inv_1
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_5_.latch/Q
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_68_129 vgnd vpwr scs8hd_decap_12
X_609_ _609_/A _609_/Y vgnd vpwr scs8hd_inv_8
XFILLER_59_129 vgnd vpwr scs8hd_fill_1
XFILLER_67_140 vgnd vpwr scs8hd_decap_6
XFILLER_67_184 vpwr vgnd scs8hd_fill_2
XFILLER_82_187 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.mux_fle_3_in_3.INVTX1_1_.scs8hd_inv_1 right_width_0_height_0__pin_1_
+ ltile_clb_0.mux_fle_3_in_3.INVTX1_1_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XPHY_717 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_706 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_739 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_728 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_23_254 vpwr vgnd scs8hd_fill_2
XFILLER_23_265 vgnd vpwr scs8hd_decap_3
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.buf4_1_.scs8hd_buf_1_A
+ ltile_clb_0.mux_fle_2_in_1.INVTX1_14_.scs8hd_inv_1/Y vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_2_in_1.mux_l1_in_2_.TGATE_3_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_2_in_1.INVTX1_11_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__522__B _517_/X vgnd vpwr scs8hd_diode_2
XANTENNA__241__C _286_/B vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_1_in_3.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_1_in_3.INVTX1_4_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_1_in_3.LATCH_0_.latch/Q ltile_clb_0.mux_fle_1_in_3.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_48_32 vgnd vpwr scs8hd_decap_12
XFILLER_58_151 vpwr vgnd scs8hd_fill_2
XFILLER_73_110 vgnd vpwr scs8hd_decap_12
XFILLER_58_173 vgnd vpwr scs8hd_decap_6
XFILLER_73_143 vgnd vpwr scs8hd_decap_3
XFILLER_73_176 vgnd vpwr scs8hd_decap_6
XANTENNA_ltile_clb_0.mux_fle_1_in_3.mux_l1_in_3_.TGATE_2_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_1_in_3.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_2_in_0.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_2_in_0.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_14_221 vgnd vpwr scs8hd_fill_1
XFILLER_9_15 vgnd vpwr scs8hd_decap_12
XFILLER_9_59 vpwr vgnd scs8hd_fill_2
XFILLER_14_298 vgnd vpwr scs8hd_decap_8
X_325_ _325_/A _326_/A vgnd vpwr scs8hd_buf_1
Xltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_12_.latch
+ data_in ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_12_.latch/Q
+ _585_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_10_471 vpwr vgnd scs8hd_fill_2
X_256_ _255_/X _559_/A vgnd vpwr scs8hd_buf_1
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__ff_0.DFFSRQ_0_.dff_CLK
+ clkbuf_1_1_0_clk/X vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mem_fle_0_in_3.LATCH_0_.latch data_in ltile_clb_0.mem_fle_0_in_3.LATCH_0_.latch/Q
+ _492_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA__432__B _429_/X vgnd vpwr scs8hd_diode_2
XFILLER_37_335 vpwr vgnd scs8hd_fill_2
XFILLER_37_357 vpwr vgnd scs8hd_fill_2
XFILLER_49_195 vpwr vgnd scs8hd_fill_2
XFILLER_64_154 vpwr vgnd scs8hd_fill_2
XFILLER_52_316 vgnd vpwr scs8hd_decap_6
XANTENNA_ltile_clb_0.mux_fle_3_in_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_3_in_2.LATCH_5_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_2_in_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_2_in_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_20_213 vgnd vpwr scs8hd_fill_1
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
+ _615_/Y vgnd vpwr scs8hd_diode_2
XFILLER_60_393 vgnd vpwr scs8hd_decap_4
Xltile_clb_0.mux_fle_1_in_0.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_1_in_0.INVTX1_3_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_1_in_0.LATCH_3_.latch/Q ltile_clb_0.mux_fle_1_in_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA__623__A _623_/A vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_2_in_1.INVTX1_13_.scs8hd_inv_1_A right_width_0_height_0__pin_13_
+ vgnd vpwr scs8hd_diode_2
XFILLER_55_110 vgnd vpwr scs8hd_decap_12
XFILLER_18_68 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mux_fle_3_in_3.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_3_in_3.INVTX1_8_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.INVTX1_0_.scs8hd_inv_1_A
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.INVTX1_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XPHY_503 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_514 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_525 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_34_56 vgnd vpwr scs8hd_decap_12
XPHY_536 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_547 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_558 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_569 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_11_257 vpwr vgnd scs8hd_fill_2
XFILLER_11_279 vpwr vgnd scs8hd_fill_2
XFILLER_7_217 vpwr vgnd scs8hd_fill_2
XANTENNA__533__A _559_/A vgnd vpwr scs8hd_diode_2
XFILLER_50_44 vgnd vpwr scs8hd_decap_12
XANTENNA__252__B address[1] vgnd vpwr scs8hd_diode_2
XFILLER_3_434 vpwr vgnd scs8hd_fill_2
XFILLER_78_202 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mux_fle_2_in_2.INVTX1_9_.scs8hd_inv_1_A right_width_0_height_0__pin_9_
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_1_in_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_1_in_1.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_59_86 vgnd vpwr scs8hd_decap_12
XFILLER_3_489 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_1_.TGATE_0_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_1_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_11_.scs8hd_inv_1
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_11_.latch/Q
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_11_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_19_346 vpwr vgnd scs8hd_fill_2
XFILLER_19_357 vpwr vgnd scs8hd_fill_2
XFILLER_75_74 vgnd vpwr scs8hd_decap_12
XFILLER_34_327 vgnd vpwr scs8hd_decap_6
XANTENNA__427__B _427_/B vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_0_in_2.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_0_in_2.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_61_179 vpwr vgnd scs8hd_fill_2
X_308_ _599_/A _231_/X _308_/X vgnd vpwr scs8hd_or2_4
X_239_ _259_/B _282_/B vgnd vpwr scs8hd_buf_1
XANTENNA__443__A _432_/A vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_3_.latch_SLEEPB
+ _295_/Y vgnd vpwr scs8hd_diode_2
XFILLER_6_294 vgnd vpwr scs8hd_decap_4
XFILLER_6_272 vgnd vpwr scs8hd_decap_3
XFILLER_41_3 vgnd vpwr scs8hd_decap_12
XFILLER_69_268 vpwr vgnd scs8hd_fill_2
XFILLER_57_408 vpwr vgnd scs8hd_fill_2
XFILLER_69_279 vpwr vgnd scs8hd_fill_2
XFILLER_57_419 vpwr vgnd scs8hd_fill_2
XFILLER_37_110 vgnd vpwr scs8hd_decap_12
XFILLER_65_463 vpwr vgnd scs8hd_fill_2
XFILLER_25_316 vpwr vgnd scs8hd_fill_2
XFILLER_65_496 vgnd vpwr scs8hd_decap_12
XFILLER_25_327 vgnd vpwr scs8hd_decap_4
XANTENNA__618__A _618_/A vgnd vpwr scs8hd_diode_2
XFILLER_37_176 vgnd vpwr scs8hd_fill_1
XANTENNA_ltile_clb_0.mux_fle_3_in_3.INVTX1_6_.scs8hd_inv_1_A bottom_width_0_height_0__pin_6_
+ vgnd vpwr scs8hd_diode_2
XFILLER_33_360 vgnd vpwr scs8hd_decap_4
XFILLER_33_382 vpwr vgnd scs8hd_fill_2
XANTENNA__353__A _392_/A vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_1_in_0.INVTX1_10_.scs8hd_inv_1 bottom_width_0_height_0__pin_10_
+ ltile_clb_0.mux_fle_1_in_0.INVTX1_10_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XFILLER_0_404 vgnd vpwr scs8hd_decap_4
XFILLER_75_238 vpwr vgnd scs8hd_fill_2
XFILLER_68_290 vgnd vpwr scs8hd_decap_4
XFILLER_56_441 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mux_fle_2_in_0.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_2_in_0.LATCH_7_.latch/Q
+ vgnd vpwr scs8hd_diode_2
X_590_ _564_/A _588_/X _590_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_28_154 vgnd vpwr scs8hd_decap_12
XANTENNA__528__A _528_/A vgnd vpwr scs8hd_diode_2
XFILLER_28_187 vpwr vgnd scs8hd_fill_2
XPHY_300 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_43_135 vgnd vpwr scs8hd_decap_12
XFILLER_43_168 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
+ _633_/Y vgnd vpwr scs8hd_diode_2
XPHY_311 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_322 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_333 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_43_179 vpwr vgnd scs8hd_fill_2
XPHY_344 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_355 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_366 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_377 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_388 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_399 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_61_98 vgnd vpwr scs8hd_decap_12
XANTENNA__263__A _258_/X vgnd vpwr scs8hd_diode_2
XFILLER_6_27 vgnd vpwr scs8hd_decap_4
XFILLER_3_220 vgnd vpwr scs8hd_decap_4
Xltile_clb_0.mux_fle_1_in_1.INVTX1_12_.scs8hd_inv_1 top_width_0_height_0__pin_12_
+ ltile_clb_0.mux_fle_1_in_1.INVTX1_12_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XFILLER_10_80 vgnd vpwr scs8hd_decap_12
XFILLER_3_297 vpwr vgnd scs8hd_fill_2
XFILLER_39_419 vpwr vgnd scs8hd_fill_2
XFILLER_66_249 vgnd vpwr scs8hd_decap_8
XFILLER_19_110 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mux_fle_1_in_1.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_1_in_1.INVTX1_13_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_81_208 vgnd vpwr scs8hd_decap_12
XFILLER_19_165 vpwr vgnd scs8hd_fill_2
XFILLER_47_474 vgnd vpwr scs8hd_decap_8
XFILLER_62_422 vgnd vpwr scs8hd_decap_6
XANTENNA__438__A _380_/X vgnd vpwr scs8hd_diode_2
XFILLER_47_485 vgnd vpwr scs8hd_decap_3
XANTENNA_ltile_clb_0.mux_fle_1_in_3.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_1_in_3.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_0_in_0.INVTX1_12_.scs8hd_inv_1_A top_width_0_height_0__pin_12_
+ vgnd vpwr scs8hd_diode_2
XANTENNA_clkbuf_0_clk_A clk vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_0_in_1.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_0_in_1.INVTX1_3_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_0_in_1.LATCH_3_.latch/Q ltile_clb_0.mux_fle_0_in_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_30_396 vgnd vpwr scs8hd_fill_1
Xltile_clb_0.mux_fle_1_in_2.INVTX1_14_.scs8hd_inv_1 ltile_clb_0.mux_fle_1_in_2.INVTX1_14_.scs8hd_inv_1/A
+ ltile_clb_0.mux_fle_1_in_2.INVTX1_14_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XANTENNA_ltile_clb_0.mux_fle_1_in_2.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_1_in_2.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_38_441 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mux_fle_1_in_2.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_1_in_2.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_65_260 vgnd vpwr scs8hd_decap_4
XANTENNA__348__A _355_/B vgnd vpwr scs8hd_diode_2
XFILLER_53_422 vpwr vgnd scs8hd_fill_2
XFILLER_25_135 vgnd vpwr scs8hd_decap_12
XFILLER_13_319 vpwr vgnd scs8hd_fill_2
XFILLER_25_179 vpwr vgnd scs8hd_fill_2
XFILLER_40_105 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_3_.TGATE_0_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_3_.TGATE_0_.scs8hd_ebufn_2/A
+ _607_/Y ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_1_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_13_.latch_D
+ data_in vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_0_in_1.INVTX1_1_.scs8hd_inv_1 right_width_0_height_0__pin_1_
+ ltile_clb_0.mux_fle_0_in_1.INVTX1_1_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XANTENNA__530__B _529_/X vgnd vpwr scs8hd_diode_2
XFILLER_0_234 vpwr vgnd scs8hd_fill_2
XFILLER_56_32 vgnd vpwr scs8hd_decap_12
XFILLER_0_289 vpwr vgnd scs8hd_fill_2
XFILLER_48_227 vgnd vpwr scs8hd_decap_3
XFILLER_63_208 vpwr vgnd scs8hd_fill_2
X_642_ _642_/HI _642_/LO vgnd vpwr scs8hd_conb_1
XFILLER_29_485 vgnd vpwr scs8hd_fill_1
XANTENNA__258__A address[2] vgnd vpwr scs8hd_diode_2
X_573_ _599_/A _552_/X _573_/X vgnd vpwr scs8hd_or2_4
XPHY_152 vgnd vpwr scs8hd_decap_3
XPHY_141 vgnd vpwr scs8hd_decap_3
XPHY_130 vgnd vpwr scs8hd_decap_3
XPHY_163 vgnd vpwr scs8hd_decap_3
XFILLER_12_341 vgnd vpwr scs8hd_fill_1
XPHY_174 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_185 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_8_345 vgnd vpwr scs8hd_fill_1
XPHY_196 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_6_.TGATE_0_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_12_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_0_in_3.INVTX1_4_.scs8hd_inv_1_A top_width_0_height_0__pin_4_
+ vgnd vpwr scs8hd_diode_2
XFILLER_79_341 vgnd vpwr scs8hd_fill_1
XANTENNA_ltile_clb_0.mux_fle_1_in_0.INVTX1_0_.scs8hd_inv_1_A top_width_0_height_0__pin_0_
+ vgnd vpwr scs8hd_diode_2
XFILLER_47_282 vgnd vpwr scs8hd_decap_8
XFILLER_62_230 vgnd vpwr scs8hd_decap_8
XFILLER_62_274 vgnd vpwr scs8hd_fill_1
XFILLER_22_105 vgnd vpwr scs8hd_decap_12
XFILLER_62_285 vgnd vpwr scs8hd_decap_3
XANTENNA_ltile_clb_0.mux_fle_0_in_0.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_0_in_0.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
+ _629_/Y vgnd vpwr scs8hd_diode_2
XANTENNA__631__A _631_/A vgnd vpwr scs8hd_diode_2
XANTENNA__350__B _353_/B vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_0_in_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_0_in_1.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_38_260 vgnd vpwr scs8hd_fill_1
XFILLER_53_230 vgnd vpwr scs8hd_fill_1
XFILLER_53_263 vpwr vgnd scs8hd_fill_2
XFILLER_26_68 vgnd vpwr scs8hd_decap_12
XFILLER_26_466 vpwr vgnd scs8hd_fill_2
XFILLER_53_296 vgnd vpwr scs8hd_decap_3
XANTENNA_ltile_clb_0.mux_fle_1_in_2.mux_l1_in_2_.TGATE_3_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_1_in_2.INVTX1_11_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__525__B _516_/X vgnd vpwr scs8hd_diode_2
XFILLER_42_56 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_12_.scs8hd_inv_1_A
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_12_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_0_in_2.INVTX1_5_.scs8hd_inv_1 right_width_0_height_0__pin_5_
+ ltile_clb_0.mux_fle_0_in_2.INVTX1_5_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XFILLER_5_315 vpwr vgnd scs8hd_fill_2
XANTENNA__541__A _541_/A vgnd vpwr scs8hd_diode_2
XANTENNA__260__B _333_/A vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_0_in_0.mux_l1_in_2_.TGATE_3_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_0_in_0.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_3_39 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_11_.scs8hd_inv_1
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_11_.latch/Q
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_11_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_67_86 vgnd vpwr scs8hd_decap_12
XFILLER_76_388 vpwr vgnd scs8hd_fill_2
X_625_ _625_/A _625_/Y vgnd vpwr scs8hd_inv_8
XFILLER_17_455 vpwr vgnd scs8hd_fill_2
XFILLER_29_293 vpwr vgnd scs8hd_fill_2
X_556_ _556_/A _558_/B _556_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_44_274 vgnd vpwr scs8hd_fill_1
XFILLER_17_499 vgnd vpwr scs8hd_decap_12
XFILLER_32_436 vgnd vpwr scs8hd_fill_1
X_487_ _328_/A _484_/X _487_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA__435__B _429_/X vgnd vpwr scs8hd_diode_2
XFILLER_40_480 vpwr vgnd scs8hd_fill_2
XANTENNA__451__A _450_/X vgnd vpwr scs8hd_diode_2
XFILLER_79_171 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mux_fle_1_in_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_1_in_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_0_in_3.INVTX1_10_.scs8hd_inv_1 bottom_width_0_height_0__pin_10_
+ ltile_clb_0.mux_fle_0_in_3.INVTX1_10_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XANTENNA__626__A _626_/A vgnd vpwr scs8hd_diode_2
XFILLER_31_480 vpwr vgnd scs8hd_fill_2
XFILLER_12_15 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.mux_fle_3_in_2.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_3_in_2.INVTX1_10_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_3_in_2.LATCH_2_.latch/Q ltile_clb_0.mux_fle_3_in_2.mux_l1_in_2_.TGATE_3_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_9_.scs8hd_inv_1_A
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_9_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_1_in_3.INVTX1_0_.scs8hd_inv_1 top_width_0_height_0__pin_0_ ltile_clb_0.mux_fle_1_in_3.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA__361__A _388_/A vgnd vpwr scs8hd_diode_2
Xltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_6_.scs8hd_inv_1/Y
+ _629_/Y ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_1_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_58_388 vpwr vgnd scs8hd_fill_2
XFILLER_58_377 vpwr vgnd scs8hd_fill_2
X_410_ _409_/X _410_/X vgnd vpwr scs8hd_buf_1
X_341_ _394_/A _341_/B _341_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA__536__A _528_/X vgnd vpwr scs8hd_diode_2
XFILLER_26_296 vgnd vpwr scs8hd_decap_6
XFILLER_41_200 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_0_in_2.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_0_in_2.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_0_in_3.INVTX1_9_.scs8hd_inv_1 right_width_0_height_0__pin_9_
+ ltile_clb_0.mux_fle_0_in_3.INVTX1_9_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XANTENNA__255__B _330_/A vgnd vpwr scs8hd_diode_2
X_272_ _271_/X _272_/X vgnd vpwr scs8hd_buf_1
XFILLER_41_299 vgnd vpwr scs8hd_fill_1
XFILLER_22_491 vpwr vgnd scs8hd_fill_2
XFILLER_5_123 vgnd vpwr scs8hd_decap_12
XANTENNA__271__A _236_/X vgnd vpwr scs8hd_diode_2
XFILLER_1_362 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_1_in_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_1_in_1.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_3_in_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_3_in_0.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_7_.TGATE_1_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_15_.scs8hd_inv_1/Y
+ _628_/Y ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_7_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_76_141 vgnd vpwr scs8hd_decap_12
XFILLER_64_303 vpwr vgnd scs8hd_fill_2
XFILLER_49_388 vpwr vgnd scs8hd_fill_2
XFILLER_52_509 vgnd vpwr scs8hd_decap_6
X_608_ _608_/A _608_/Y vgnd vpwr scs8hd_inv_8
XANTENNA__446__A _435_/A vgnd vpwr scs8hd_diode_2
XFILLER_17_296 vgnd vpwr scs8hd_decap_3
X_539_ _539_/A _541_/B _539_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_20_439 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_1_in_0.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_1_in_0.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_71_3 vgnd vpwr scs8hd_decap_12
XFILLER_9_484 vpwr vgnd scs8hd_fill_2
XFILLER_4_93 vgnd vpwr scs8hd_decap_12
XFILLER_67_174 vgnd vpwr scs8hd_decap_3
XFILLER_55_358 vpwr vgnd scs8hd_fill_2
XFILLER_55_347 vpwr vgnd scs8hd_fill_2
XFILLER_70_306 vgnd vpwr scs8hd_decap_12
XFILLER_82_199 vgnd vpwr scs8hd_decap_12
XFILLER_70_328 vgnd vpwr scs8hd_decap_8
XPHY_718 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_707 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__356__A _379_/A vgnd vpwr scs8hd_diode_2
XFILLER_23_200 vpwr vgnd scs8hd_fill_2
XPHY_729 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_23_233 vpwr vgnd scs8hd_fill_2
XFILLER_11_428 vgnd vpwr scs8hd_decap_4
XANTENNA_ltile_clb_0.mux_fle_2_in_2.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_2_in_2.LATCH_6_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_6_.TGATE_0_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_12_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_0_.TGATE_0_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ _625_/Y ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_48_44 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mux_fle_2_in_0.INVTX1_6_.scs8hd_inv_1_A bottom_width_0_height_0__pin_6_
+ vgnd vpwr scs8hd_diode_2
XFILLER_64_32 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.mux_fle_1_in_0.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_1_in_0.INVTX1_9_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_1_in_0.LATCH_1_.latch/Q ltile_clb_0.mux_fle_1_in_0.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_46_369 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.mux_fle_3_in_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_3_in_0.INVTX1_4_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_3_in_0.LATCH_0_.latch/Q ltile_clb_0.mux_fle_3_in_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_54_391 vpwr vgnd scs8hd_fill_2
XFILLER_54_380 vpwr vgnd scs8hd_fill_2
XANTENNA__266__A _248_/A vgnd vpwr scs8hd_diode_2
XFILLER_9_27 vgnd vpwr scs8hd_decap_12
X_324_ _324_/A _325_/A vgnd vpwr scs8hd_buf_1
X_255_ _236_/X _330_/A _255_/X vgnd vpwr scs8hd_or2_4
XFILLER_10_450 vgnd vpwr scs8hd_decap_8
XANTENNA_ltile_clb_0.mux_fle_0_in_2.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_0_in_2.INVTX1_13_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_12_.latch_SLEEPB
+ _257_/Y vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_2_in_0.INVTX1_6_.scs8hd_inv_1 bottom_width_0_height_0__pin_6_
+ ltile_clb_0.mux_fle_2_in_0.INVTX1_6_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XFILLER_69_439 vpwr vgnd scs8hd_fill_2
XFILLER_49_141 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_3_in_0.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_3_in_0.INVTX1_13_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_52_328 vgnd vpwr scs8hd_decap_3
Xltile_clb_0.mux_fle_2_in_3.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_2_in_3.INVTX1_10_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_2_in_3.LATCH_2_.latch/Q ltile_clb_0.mux_fle_2_in_3.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_60_372 vpwr vgnd scs8hd_fill_2
XFILLER_9_292 vpwr vgnd scs8hd_fill_2
XFILLER_9_281 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_3_in_1.INVTX1_3_.scs8hd_inv_1_A left_width_0_height_0__pin_3_
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_0_in_3.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_0_in_3.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_68_450 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_55_155 vpwr vgnd scs8hd_fill_2
XFILLER_16_509 vgnd vpwr scs8hd_decap_6
XANTENNA_ltile_clb_0.mux_fle_3_in_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_3_in_1.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_55_199 vpwr vgnd scs8hd_fill_2
XPHY_504 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_515 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_526 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_34_68 vgnd vpwr scs8hd_decap_12
XPHY_537 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_548 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_559 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_11_236 vpwr vgnd scs8hd_fill_2
XFILLER_11_225 vgnd vpwr scs8hd_decap_6
XANTENNA_ltile_clb_0.mux_fle_2_in_3.INVTX1_11_.scs8hd_inv_1_A left_width_0_height_0__pin_11_
+ vgnd vpwr scs8hd_diode_2
XANTENNA__533__B _529_/X vgnd vpwr scs8hd_diode_2
XFILLER_50_56 vgnd vpwr scs8hd_decap_12
XFILLER_3_479 vpwr vgnd scs8hd_fill_2
XFILLER_3_468 vpwr vgnd scs8hd_fill_2
XFILLER_1_3 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_11_.scs8hd_inv_1
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_11_.latch/Q
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_11_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_59_98 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.mux_fle_3_in_1.INVTX1_1_.scs8hd_inv_1 right_width_0_height_0__pin_1_
+ ltile_clb_0.mux_fle_3_in_1.INVTX1_1_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XFILLER_59_483 vgnd vpwr scs8hd_decap_4
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_2_.TGATE_0_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_2_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_74_442 vgnd vpwr scs8hd_decap_4
XFILLER_19_336 vgnd vpwr scs8hd_fill_1
XFILLER_75_86 vgnd vpwr scs8hd_decap_12
XFILLER_27_380 vpwr vgnd scs8hd_fill_2
XANTENNA__427__C _384_/X vgnd vpwr scs8hd_diode_2
Xltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_8_.scs8hd_inv_1
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_8_.latch/Q
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_8_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
Xltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_0_.scs8hd_inv_1/Y
+ _605_/Y ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_ltile_clb_0.mem_fle_2_in_3.LATCH_4_.latch_SLEEPB _391_/Y vgnd vpwr scs8hd_diode_2
XFILLER_30_501 vgnd vpwr scs8hd_decap_12
X_307_ address[4] _599_/A vgnd vpwr scs8hd_inv_8
X_238_ address[1] _259_/B vgnd vpwr scs8hd_inv_8
XANTENNA__443__B _446_/B vgnd vpwr scs8hd_diode_2
XFILLER_69_214 vpwr vgnd scs8hd_fill_2
XFILLER_34_3 vgnd vpwr scs8hd_decap_12
XFILLER_69_236 vpwr vgnd scs8hd_fill_2
XFILLER_65_420 vgnd vpwr scs8hd_decap_4
XFILLER_25_306 vgnd vpwr scs8hd_fill_1
XFILLER_37_144 vgnd vpwr scs8hd_decap_4
XFILLER_37_155 vpwr vgnd scs8hd_fill_2
XFILLER_40_309 vgnd vpwr scs8hd_decap_4
XANTENNA__634__A _634_/A vgnd vpwr scs8hd_diode_2
Xltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_4_.TGATE_1_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_9_.scs8hd_inv_1/Y
+ _604_/Y ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_2_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA__353__B _353_/B vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_0_in_3.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_0_in_3.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_20_15 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mux_fle_0_in_3.mux_l1_in_2_.TGATE_3_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_0_in_3.INVTX1_11_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_75_217 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.mux_fle_2_in_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_2_in_1.INVTX1_4_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_2_in_1.LATCH_0_.latch/Q ltile_clb_0.mux_fle_2_in_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
Xltile_clb_0.mux_fle_0_in_1.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_0_in_1.INVTX1_9_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_0_in_1.LATCH_1_.latch/Q ltile_clb_0.mux_fle_0_in_1.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_56_453 vgnd vpwr scs8hd_decap_4
XFILLER_28_166 vgnd vpwr scs8hd_decap_6
XFILLER_71_423 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_0_in_2.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_0_in_2.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_5_.TGATE_1_.scs8hd_ebufn_2_TEB
+ _628_/Y vgnd vpwr scs8hd_diode_2
XPHY_301 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_71_489 vgnd vpwr scs8hd_decap_12
XPHY_312 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_323 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_334 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_ltile_clb_0.mux_fle_3_in_1.mux_l1_in_2_.TGATE_3_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_3_in_1.INVTX1_11_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XPHY_345 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_356 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_367 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_378 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__544__A _544_/A vgnd vpwr scs8hd_diode_2
XPHY_389 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__263__B _282_/B vgnd vpwr scs8hd_diode_2
XFILLER_79_501 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.mux_fle_3_in_2.INVTX1_5_.scs8hd_inv_1 right_width_0_height_0__pin_5_
+ ltile_clb_0.mux_fle_3_in_2.INVTX1_5_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
Xltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_1_.latch
+ data_in ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_1_.latch/Q
+ _301_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_66_206 vgnd vpwr scs8hd_decap_8
XANTENNA_ltile_clb_0.mem_fle_3_in_2.LATCH_4_.latch_SLEEPB _352_/Y vgnd vpwr scs8hd_diode_2
XFILLER_74_250 vgnd vpwr scs8hd_decap_6
XANTENNA_ltile_clb_0.mux_fle_0_in_1.INVTX1_1_.scs8hd_inv_1_A right_width_0_height_0__pin_1_
+ vgnd vpwr scs8hd_diode_2
XFILLER_62_401 vpwr vgnd scs8hd_fill_2
XANTENNA__438__B _226_/X vgnd vpwr scs8hd_diode_2
XFILLER_19_188 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_6_.latch_SLEEPB
+ _566_/Y vgnd vpwr scs8hd_diode_2
XFILLER_22_309 vpwr vgnd scs8hd_fill_2
XFILLER_30_331 vgnd vpwr scs8hd_decap_4
XANTENNA__454__A _432_/A vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_0_in_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_0_in_3.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_57_217 vpwr vgnd scs8hd_fill_2
XANTENNA__629__A _629_/A vgnd vpwr scs8hd_diode_2
XFILLER_38_453 vgnd vpwr scs8hd_decap_4
XANTENNA_ltile_clb_0.mux_fle_3_in_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_3_in_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_65_283 vgnd vpwr scs8hd_decap_3
XANTENNA_ltile_clb_0.mux_fle_0_in_2.INVTX1_10_.scs8hd_inv_1_A bottom_width_0_height_0__pin_10_
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mem_fle_0_in_3.LATCH_5_.latch_SLEEPB _487_/Y vgnd vpwr scs8hd_diode_2
XFILLER_38_475 vgnd vpwr scs8hd_decap_12
XFILLER_25_147 vgnd vpwr scs8hd_decap_12
XFILLER_80_264 vgnd vpwr scs8hd_decap_8
XFILLER_15_15 vgnd vpwr scs8hd_decap_12
XFILLER_40_117 vgnd vpwr scs8hd_decap_12
XFILLER_15_59 vpwr vgnd scs8hd_fill_2
XFILLER_21_331 vpwr vgnd scs8hd_fill_2
XANTENNA__364__A _391_/A vgnd vpwr scs8hd_diode_2
XFILLER_0_246 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_3_.scs8hd_inv_1_A
+ ltile_clb_0.mux_fle_2_in_3.INVTX1_14_.scs8hd_inv_1/Y vgnd vpwr scs8hd_diode_2
XFILLER_76_504 vgnd vpwr scs8hd_decap_12
XFILLER_48_206 vgnd vpwr scs8hd_decap_8
XFILLER_48_239 vgnd vpwr scs8hd_decap_12
XFILLER_56_44 vgnd vpwr scs8hd_decap_12
XANTENNA__539__A _539_/A vgnd vpwr scs8hd_diode_2
XFILLER_29_453 vpwr vgnd scs8hd_fill_2
X_641_ _641_/HI _641_/LO vgnd vpwr scs8hd_conb_1
X_572_ _546_/A _554_/X _572_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_72_32 vgnd vpwr scs8hd_decap_12
XFILLER_71_297 vpwr vgnd scs8hd_fill_2
XPHY_142 vgnd vpwr scs8hd_decap_3
XPHY_131 vgnd vpwr scs8hd_decap_3
XPHY_120 vgnd vpwr scs8hd_decap_3
XPHY_164 vgnd vpwr scs8hd_decap_3
XPHY_153 vgnd vpwr scs8hd_decap_3
XPHY_175 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_191 vgnd vpwr scs8hd_decap_8
XANTENNA__274__A _258_/X vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_3_in_3.INVTX1_9_.scs8hd_inv_1 right_width_0_height_0__pin_9_
+ ltile_clb_0.mux_fle_3_in_3.INVTX1_9_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XANTENNA_ltile_clb_0.mux_fle_2_in_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_2_in_1.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_12_375 vpwr vgnd scs8hd_fill_2
XPHY_186 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_197 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_ltile_clb_0.mux_fle_1_in_2.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_1_in_2.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_clkbuf_1_0_0_clk_A clkbuf_0_clk/X vgnd vpwr scs8hd_diode_2
XANTENNA__449__A _380_/X vgnd vpwr scs8hd_diode_2
XFILLER_35_423 vpwr vgnd scs8hd_fill_2
XFILLER_62_220 vgnd vpwr scs8hd_fill_1
XFILLER_35_456 vgnd vpwr scs8hd_decap_3
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_12_.scs8hd_inv_1_A
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_12_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XPHY_0 vgnd vpwr scs8hd_decap_3
XFILLER_22_117 vgnd vpwr scs8hd_decap_12
XFILLER_15_191 vgnd vpwr scs8hd_decap_4
XFILLER_30_172 vgnd vpwr scs8hd_decap_4
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_3_.TGATE_1_.scs8hd_ebufn_2_TEB
+ _606_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mem_fle_1_in_2.LATCH_5_.latch_SLEEPB _454_/Y vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_1_in_2.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_1_in_2.INVTX1_4_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_1_in_2.LATCH_0_.latch/Q ltile_clb_0.mux_fle_1_in_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.mem_ble4_out_0.LATCH_1_.latch_D
+ data_in vgnd vpwr scs8hd_diode_2
XANTENNA__359__A _358_/X vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_2_.TGATE_0_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_4_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_14_.latch
+ data_in ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_14_.latch/Q
+ _248_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
Xltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.INVTX1_0_.scs8hd_inv_1/Y
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.mem_ble4_out_0.LATCH_0_.latch/Q
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_41_459 vpwr vgnd scs8hd_fill_2
XFILLER_21_172 vpwr vgnd scs8hd_fill_2
XFILLER_42_68 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_1_.latch
+ data_in ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_1_.latch/Q
+ _597_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
Xltile_clb_0.mem_fle_0_in_0.LATCH_7_.latch data_in ltile_clb_0.mem_fle_0_in_0.LATCH_7_.latch/Q
+ _518_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA__541__B _541_/B vgnd vpwr scs8hd_diode_2
XFILLER_67_98 vgnd vpwr scs8hd_decap_12
XFILLER_64_507 vgnd vpwr scs8hd_decap_8
XANTENNA__269__A _269_/A vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mem_fle_1_in_0.LATCH_6_.latch data_in ltile_clb_0.mem_fle_1_in_0.LATCH_6_.latch/Q
+ _475_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_17_401 vpwr vgnd scs8hd_fill_2
X_624_ _624_/A _624_/Y vgnd vpwr scs8hd_inv_8
XFILLER_17_423 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_1_.scs8hd_inv_1
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_1_.latch/Q
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_17_489 vgnd vpwr scs8hd_decap_8
X_555_ _554_/X _558_/B vgnd vpwr scs8hd_buf_1
XFILLER_44_242 vgnd vpwr scs8hd_decap_12
XFILLER_16_80 vgnd vpwr scs8hd_decap_12
X_486_ _325_/A _484_/X _486_/Y vgnd vpwr scs8hd_nor2_4
Xltile_clb_0.mem_fle_2_in_0.LATCH_5_.latch data_in ltile_clb_0.mem_fle_2_in_0.LATCH_5_.latch/Q
+ _432_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_12_194 vgnd vpwr scs8hd_decap_8
XFILLER_8_154 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mux_fle_2_in_1.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_2_in_1.INVTX1_13_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_67_334 vgnd vpwr scs8hd_decap_3
XFILLER_67_301 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.mem_fle_3_in_0.LATCH_4_.latch data_in ltile_clb_0.mem_fle_3_in_0.LATCH_4_.latch/Q
+ _375_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_67_367 vgnd vpwr scs8hd_decap_3
XFILLER_67_356 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_0_in_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_0_in_1.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_82_304 vgnd vpwr scs8hd_decap_6
XFILLER_35_220 vpwr vgnd scs8hd_fill_2
XFILLER_35_231 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mem_fle_2_in_1.LATCH_5_.latch_SLEEPB _416_/Y vgnd vpwr scs8hd_diode_2
XFILLER_23_437 vgnd vpwr scs8hd_decap_3
XFILLER_23_448 vgnd vpwr scs8hd_decap_4
XFILLER_35_297 vpwr vgnd scs8hd_fill_2
XFILLER_12_27 vgnd vpwr scs8hd_decap_4
XANTENNA__361__B _365_/B vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_0_in_0.mux_l1_in_3_.TGATE_2_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_0_in_0.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_2_in_2.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_2_in_2.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_58_367 vgnd vpwr scs8hd_fill_1
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_11_.latch_SLEEPB
+ _586_/Y vgnd vpwr scs8hd_diode_2
XFILLER_73_326 vgnd vpwr scs8hd_decap_4
Xltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_1_.TGATE_1_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_1_.TGATE_1_.scs8hd_ebufn_2/A
+ _622_/Y ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_26_264 vgnd vpwr scs8hd_decap_8
XFILLER_81_370 vgnd vpwr scs8hd_decap_8
XFILLER_14_437 vgnd vpwr scs8hd_decap_4
XANTENNA_ltile_clb_0.mux_fle_1_in_1.INVTX1_7_.scs8hd_inv_1_A left_width_0_height_0__pin_7_
+ vgnd vpwr scs8hd_diode_2
X_340_ _423_/A _394_/A vgnd vpwr scs8hd_buf_1
XFILLER_14_459 vgnd vpwr scs8hd_decap_3
X_271_ _236_/X _339_/A _271_/X vgnd vpwr scs8hd_or2_4
XFILLER_41_278 vpwr vgnd scs8hd_fill_2
XANTENNA__552__A _380_/A vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_3_in_1.INVTX1_13_.scs8hd_inv_1_A right_width_0_height_0__pin_13_
+ vgnd vpwr scs8hd_diode_2
XFILLER_5_135 vgnd vpwr scs8hd_decap_12
XANTENNA__271__B _339_/A vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_1_in_2.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_1_in_2.LATCH_7_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_49_301 vpwr vgnd scs8hd_fill_2
XFILLER_49_323 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mem_fle_0_in_1.LATCH_7_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_49_345 vpwr vgnd scs8hd_fill_2
XFILLER_49_367 vgnd vpwr scs8hd_fill_1
XFILLER_64_337 vgnd vpwr scs8hd_fill_1
X_607_ _607_/A _607_/Y vgnd vpwr scs8hd_inv_8
XFILLER_72_392 vgnd vpwr scs8hd_fill_1
XANTENNA__446__B _446_/B vgnd vpwr scs8hd_diode_2
XFILLER_17_275 vpwr vgnd scs8hd_fill_2
XFILLER_32_201 vgnd vpwr scs8hd_decap_4
Xltile_clb_0.mux_fle_0_in_0.INVTX1_5_.scs8hd_inv_1 right_width_0_height_0__pin_5_
+ ltile_clb_0.mux_fle_0_in_0.INVTX1_5_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
X_538_ _564_/A _541_/B _538_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_32_234 vgnd vpwr scs8hd_decap_3
XFILLER_32_256 vpwr vgnd scs8hd_fill_2
XFILLER_32_267 vgnd vpwr scs8hd_decap_4
X_469_ _436_/A _461_/X _469_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_9_452 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.mem_fle_3_in_2.LATCH_7_.latch data_in ltile_clb_0.mem_fle_3_in_2.LATCH_7_.latch/Q
+ _349_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_9_463 vgnd vpwr scs8hd_fill_1
XANTENNA__462__A _461_/X vgnd vpwr scs8hd_diode_2
XFILLER_64_3 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mem_fle_0_in_2.LATCH_5_.latch_D data_in vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_0_in_3.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_0_in_3.INVTX1_4_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_0_in_3.LATCH_0_.latch/Q ltile_clb_0.mux_fle_0_in_3.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_ltile_clb_0.mux_fle_2_in_2.INVTX1_4_.scs8hd_inv_1_A top_width_0_height_0__pin_4_
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mem_fle_3_in_0.LATCH_5_.latch_SLEEPB _374_/Y vgnd vpwr scs8hd_diode_2
XFILLER_4_190 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_6_.scs8hd_inv_1
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_6_.latch/Q
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_ltile_clb_0.mux_fle_1_in_0.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_1_in_0.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_28_507 vgnd vpwr scs8hd_decap_8
XFILLER_67_197 vgnd vpwr scs8hd_decap_3
XFILLER_55_326 vpwr vgnd scs8hd_fill_2
XFILLER_82_156 vgnd vpwr scs8hd_decap_12
XFILLER_70_318 vgnd vpwr scs8hd_fill_1
XPHY_708 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_1_.latch
+ data_in ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_1_.latch/Q
+ _571_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_ltile_clb_0.mem_fle_0_in_3.LATCH_3_.latch_D data_in vgnd vpwr scs8hd_diode_2
XPHY_719 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__356__B _355_/B vgnd vpwr scs8hd_diode_2
XFILLER_23_15 vgnd vpwr scs8hd_decap_12
XFILLER_23_289 vgnd vpwr scs8hd_decap_3
XFILLER_23_59 vpwr vgnd scs8hd_fill_2
XANTENNA__372__A _388_/A vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_9_.latch_D
+ data_in vgnd vpwr scs8hd_diode_2
XFILLER_2_105 vgnd vpwr scs8hd_decap_12
XFILLER_78_407 vgnd vpwr scs8hd_fill_1
XANTENNA_ltile_clb_0.mem_fle_1_in_0.LATCH_5_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_48_56 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mux_fle_2_in_2.mux_l1_in_2_.TGATE_3_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_2_in_2.INVTX1_11_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_73_123 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mem_fle_0_in_1.LATCH_6_.latch_SLEEPB _508_/Y vgnd vpwr scs8hd_diode_2
XFILLER_46_348 vpwr vgnd scs8hd_fill_2
XFILLER_64_44 vgnd vpwr scs8hd_decap_12
XFILLER_61_318 vpwr vgnd scs8hd_fill_2
XANTENNA__547__A _599_/A vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_3_in_3.INVTX1_1_.scs8hd_inv_1_A right_width_0_height_0__pin_1_
+ vgnd vpwr scs8hd_diode_2
XANTENNA__266__B _535_/A vgnd vpwr scs8hd_diode_2
XFILLER_80_32 vgnd vpwr scs8hd_decap_12
X_323_ _388_/A _338_/B _323_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_9_39 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.mux_fle_1_in_1.INVTX1_0_.scs8hd_inv_1 top_width_0_height_0__pin_0_ ltile_clb_0.mux_fle_1_in_1.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
Xltile_clb_0.mux_fle_0_in_0.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_0_in_0.INVTX1_3_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_0_in_0.LATCH_3_.latch/Q ltile_clb_0.mux_fle_0_in_0.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
X_254_ _286_/A _603_/A _330_/A vgnd vpwr scs8hd_or2_4
XFILLER_10_440 vgnd vpwr scs8hd_fill_1
XFILLER_6_411 vpwr vgnd scs8hd_fill_2
XANTENNA__282__A _286_/A vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_0_in_0.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_0_in_0.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mem_fle_1_in_1.LATCH_3_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_10_495 vgnd vpwr scs8hd_decap_8
XFILLER_10_484 vgnd vpwr scs8hd_decap_4
XFILLER_1_171 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.mux_fle_0_in_1.INVTX1_9_.scs8hd_inv_1 right_width_0_height_0__pin_9_
+ ltile_clb_0.mux_fle_0_in_1.INVTX1_9_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XFILLER_37_315 vpwr vgnd scs8hd_fill_2
XFILLER_49_164 vgnd vpwr scs8hd_decap_8
XFILLER_49_175 vpwr vgnd scs8hd_fill_2
XFILLER_37_326 vpwr vgnd scs8hd_fill_2
XFILLER_64_145 vgnd vpwr scs8hd_decap_8
XANTENNA_ltile_clb_0.mem_fle_1_in_2.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA__457__A _435_/A vgnd vpwr scs8hd_diode_2
XFILLER_64_189 vpwr vgnd scs8hd_fill_2
XFILLER_33_510 vgnd vpwr scs8hd_decap_6
XFILLER_9_260 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_2_in_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_2_in_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2_TEB
+ _620_/Y vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_0_in_0.INVTX1_12_.scs8hd_inv_1 top_width_0_height_0__pin_12_
+ ltile_clb_0.mux_fle_0_in_0.INVTX1_12_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
Xltile_clb_0.mux_fle_3_in_0.INVTX1_11_.scs8hd_inv_1 left_width_0_height_0__pin_11_
+ ltile_clb_0.mux_fle_3_in_0.INVTX1_11_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XFILLER_18_15 vgnd vpwr scs8hd_decap_12
XFILLER_55_123 vgnd vpwr scs8hd_decap_4
XANTENNA__367__A _394_/A vgnd vpwr scs8hd_diode_2
XFILLER_28_359 vgnd vpwr scs8hd_decap_3
XANTENNA_ltile_clb_0.mux_fle_1_in_0.INVTX1_12_.scs8hd_inv_1_A top_width_0_height_0__pin_12_
+ vgnd vpwr scs8hd_diode_2
XPHY_505 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_516 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_ltile_clb_0.mem_fle_2_in_0.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_51_362 vgnd vpwr scs8hd_fill_1
XFILLER_11_204 vpwr vgnd scs8hd_fill_2
XPHY_527 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_538 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_549 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_3_403 vgnd vpwr scs8hd_decap_3
XANTENNA_ltile_clb_0.mem_fle_1_in_0.LATCH_6_.latch_SLEEPB _475_/Y vgnd vpwr scs8hd_diode_2
XFILLER_50_68 vgnd vpwr scs8hd_decap_12
XFILLER_3_425 vpwr vgnd scs8hd_fill_2
XFILLER_78_215 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_5_.latch_D
+ data_in vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_0_in_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_0_in_0.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_59_462 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.mux_fle_0_in_1.INVTX1_14_.scs8hd_inv_1 ltile_clb_0.mux_fle_0_in_1.INVTX1_14_.scs8hd_inv_1/A
+ ltile_clb_0.mux_fle_0_in_1.INVTX1_14_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XFILLER_74_432 vgnd vpwr scs8hd_fill_1
XFILLER_19_315 vpwr vgnd scs8hd_fill_2
XFILLER_19_326 vpwr vgnd scs8hd_fill_2
XFILLER_75_98 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.mux_fle_3_in_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_3_in_3.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ ltile_clb_0.mem_fle_3_in_3.LATCH_4_.latch/Q ltile_clb_0.mux_fle_3_in_3.INVTX1_14_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA__277__A _267_/X vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_1_in_2.INVTX1_4_.scs8hd_inv_1 top_width_0_height_0__pin_4_ ltile_clb_0.mux_fle_1_in_2.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_ltile_clb_0.mux_fle_1_in_2.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_1_in_2.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_46_145 vgnd vpwr scs8hd_decap_8
XFILLER_15_510 vgnd vpwr scs8hd_decap_6
XFILLER_61_159 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.mux_fle_3_in_1.INVTX1_13_.scs8hd_inv_1 right_width_0_height_0__pin_13_
+ ltile_clb_0.mux_fle_3_in_1.INVTX1_13_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XANTENNA__427__D _346_/D vgnd vpwr scs8hd_diode_2
XFILLER_30_513 vgnd vpwr scs8hd_decap_3
XFILLER_42_362 vpwr vgnd scs8hd_fill_2
X_306_ _305_/X _575_/A vgnd vpwr scs8hd_buf_1
XFILLER_24_80 vgnd vpwr scs8hd_decap_12
X_237_ address[2] _286_/A vgnd vpwr scs8hd_inv_8
XANTENNA_ltile_clb_0.mux_fle_3_in_0.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_3_in_0.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_69_248 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_1_.latch
+ data_in ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_1_.latch/Q
+ _545_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_27_3 vgnd vpwr scs8hd_decap_12
XFILLER_77_270 vpwr vgnd scs8hd_fill_2
XFILLER_65_410 vpwr vgnd scs8hd_fill_2
XFILLER_37_123 vgnd vpwr scs8hd_decap_12
XFILLER_1_62 vgnd vpwr scs8hd_decap_12
XFILLER_1_51 vgnd vpwr scs8hd_decap_8
XFILLER_80_424 vgnd vpwr scs8hd_decap_12
XFILLER_65_476 vpwr vgnd scs8hd_fill_2
XFILLER_33_340 vpwr vgnd scs8hd_fill_2
XFILLER_33_351 vgnd vpwr scs8hd_decap_3
XFILLER_33_395 vgnd vpwr scs8hd_decap_3
XFILLER_20_27 vgnd vpwr scs8hd_decap_4
XFILLER_56_465 vgnd vpwr scs8hd_decap_4
XFILLER_71_402 vpwr vgnd scs8hd_fill_2
XFILLER_71_457 vpwr vgnd scs8hd_fill_2
XPHY_302 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_313 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_324 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_351 vpwr vgnd scs8hd_fill_2
XPHY_335 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_346 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_357 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_368 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_51_170 vpwr vgnd scs8hd_fill_2
XPHY_379 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__544__B _528_/X vgnd vpwr scs8hd_diode_2
XANTENNA__263__C _282_/C vgnd vpwr scs8hd_diode_2
XANTENNA__560__A _261_/X vgnd vpwr scs8hd_diode_2
XFILLER_79_513 vgnd vpwr scs8hd_decap_3
XFILLER_3_266 vpwr vgnd scs8hd_fill_2
XFILLER_10_93 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.mux_fle_1_in_3.INVTX1_8_.scs8hd_inv_1 top_width_0_height_0__pin_8_ ltile_clb_0.mux_fle_1_in_3.INVTX1_8_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
Xltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_4_.scs8hd_inv_1/Y
+ _613_/Y ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_1_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_19_123 vgnd vpwr scs8hd_decap_12
XFILLER_47_432 vpwr vgnd scs8hd_fill_2
XFILLER_47_443 vpwr vgnd scs8hd_fill_2
XFILLER_47_454 vpwr vgnd scs8hd_fill_2
XANTENNA__438__C _384_/X vgnd vpwr scs8hd_diode_2
XFILLER_47_498 vpwr vgnd scs8hd_fill_2
XFILLER_62_446 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_1_.latch_D
+ data_in vgnd vpwr scs8hd_diode_2
XFILLER_15_362 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_1_in_2.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_1_in_2.INVTX1_13_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_15_395 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_0_in_3.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_0_in_3.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__454__B _451_/X vgnd vpwr scs8hd_diode_2
XFILLER_30_387 vgnd vpwr scs8hd_decap_6
Xltile_clb_0.mux_fle_3_in_1.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_3_in_1.INVTX1_10_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_3_in_1.LATCH_2_.latch/Q ltile_clb_0.mux_fle_3_in_1.mux_l1_in_2_.TGATE_3_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
Xltile_clb_0.mem_fle_0_in_1.LATCH_3_.latch data_in ltile_clb_0.mem_fle_0_in_1.LATCH_3_.latch/Q
+ _511_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA__470__A _437_/A vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.buf4_3_.scs8hd_buf_1_A
+ ltile_clb_0.mux_fle_1_in_3.INVTX1_14_.scs8hd_inv_1/Y vgnd vpwr scs8hd_diode_2
XFILLER_65_240 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_6_.TGATE_0_.scs8hd_ebufn_2_TEB
+ _629_/Y vgnd vpwr scs8hd_diode_2
XFILLER_38_487 vgnd vpwr scs8hd_fill_1
XANTENNA_ltile_clb_0.mux_fle_0_in_2.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_0_in_2.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mem_fle_1_in_1.LATCH_2_.latch data_in ltile_clb_0.mem_fle_1_in_1.LATCH_2_.latch/Q
+ _468_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
Xltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_6_.TGATE_1_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_13_.scs8hd_inv_1/Y
+ _612_/Y ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_6_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_80_276 vgnd vpwr scs8hd_decap_8
XFILLER_53_479 vpwr vgnd scs8hd_fill_2
XFILLER_53_468 vgnd vpwr scs8hd_decap_4
XFILLER_15_27 vgnd vpwr scs8hd_decap_12
XFILLER_25_159 vgnd vpwr scs8hd_decap_8
XFILLER_80_287 vgnd vpwr scs8hd_decap_8
XANTENNA_ltile_clb_0.mux_fle_3_in_3.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_3_in_3.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_40_129 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mux_fle_1_in_3.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_1_in_3.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__364__B _365_/B vgnd vpwr scs8hd_diode_2
XFILLER_21_376 vpwr vgnd scs8hd_fill_2
XFILLER_31_15 vgnd vpwr scs8hd_decap_12
XFILLER_31_59 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.mem_fle_2_in_1.LATCH_1_.latch data_in ltile_clb_0.mem_fle_2_in_1.LATCH_1_.latch/Q
+ _424_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA__380__A _380_/A vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_0_.TGATE_1_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_48_218 vpwr vgnd scs8hd_fill_2
XFILLER_56_56 vgnd vpwr scs8hd_decap_12
XANTENNA__539__B _541_/B vgnd vpwr scs8hd_diode_2
XFILLER_29_443 vgnd vpwr scs8hd_decap_6
X_640_ _640_/HI _640_/LO vgnd vpwr scs8hd_conb_1
XFILLER_56_251 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.mem_fle_3_in_1.LATCH_0_.latch data_in ltile_clb_0.mem_fle_3_in_1.LATCH_0_.latch/Q
+ _368_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
X_571_ _545_/A _554_/X _571_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_29_498 vpwr vgnd scs8hd_fill_2
XFILLER_71_221 vgnd vpwr scs8hd_decap_4
XFILLER_44_435 vgnd vpwr scs8hd_decap_4
XFILLER_72_44 vgnd vpwr scs8hd_decap_12
XFILLER_71_254 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mem_fle_2_in_2.LATCH_7_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_2_in_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_2_in_1.LATCH_4_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__555__A _554_/X vgnd vpwr scs8hd_diode_2
XFILLER_44_468 vgnd vpwr scs8hd_decap_4
XPHY_143 vgnd vpwr scs8hd_decap_3
XPHY_132 vgnd vpwr scs8hd_decap_3
XPHY_121 vgnd vpwr scs8hd_decap_3
XPHY_110 vgnd vpwr scs8hd_decap_3
XFILLER_52_490 vgnd vpwr scs8hd_decap_4
XPHY_165 vgnd vpwr scs8hd_decap_3
XPHY_154 vgnd vpwr scs8hd_decap_3
XPHY_176 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__274__B _603_/A vgnd vpwr scs8hd_diode_2
XFILLER_8_314 vgnd vpwr scs8hd_decap_4
XPHY_187 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_198 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_4_.scs8hd_inv_1_A
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_4_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__290__A _278_/X vgnd vpwr scs8hd_diode_2
XFILLER_79_321 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mem_fle_2_in_3.LATCH_5_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_79_376 vgnd vpwr scs8hd_decap_4
XANTENNA__449__B _226_/X vgnd vpwr scs8hd_diode_2
XFILLER_62_210 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.mem_fle_0_in_3.LATCH_6_.latch data_in ltile_clb_0.mem_fle_0_in_3.LATCH_6_.latch/Q
+ _486_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XPHY_1 vgnd vpwr scs8hd_decap_3
XFILLER_50_416 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_10_.latch_SLEEPB
+ _561_/Y vgnd vpwr scs8hd_diode_2
XFILLER_22_129 vgnd vpwr scs8hd_decap_12
XANTENNA__465__A _432_/A vgnd vpwr scs8hd_diode_2
XFILLER_50_427 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mem_fle_3_in_0.LATCH_7_.latch_D data_in vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_3_in_0.INVTX1_5_.scs8hd_inv_1 right_width_0_height_0__pin_5_
+ ltile_clb_0.mux_fle_3_in_0.INVTX1_5_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
Xltile_clb_0.mux_fle_2_in_3.INVTX1_11_.scs8hd_inv_1 left_width_0_height_0__pin_11_
+ ltile_clb_0.mux_fle_2_in_3.INVTX1_11_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XANTENNA_ltile_clb_0.mux_fle_0_in_1.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_0_in_1.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mem_fle_1_in_3.LATCH_5_.latch data_in ltile_clb_0.mem_fle_1_in_3.LATCH_5_.latch/Q
+ _443_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
Xltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__ff_0.DFFSRQ_0_.dff
+ clkbuf_1_1_0_clk/X ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.INVTX1_1_.scs8hd_inv_1/A
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.INVTX1_0_.scs8hd_inv_1/A
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__ff_0.DFFSRQ_0_.dff/QN
+ reset set vgnd vpwr scs8hd_dfbbp_1
XFILLER_26_15 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
+ _616_/Y vgnd vpwr scs8hd_diode_2
XFILLER_38_240 vpwr vgnd scs8hd_fill_2
XFILLER_38_251 vgnd vpwr scs8hd_decap_6
XANTENNA_ltile_clb_0.mem_fle_3_in_1.LATCH_5_.latch_D data_in vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mem_fle_2_in_3.LATCH_4_.latch data_in ltile_clb_0.mem_fle_2_in_3.LATCH_4_.latch/Q
+ _391_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_26_457 vgnd vpwr scs8hd_fill_1
XANTENNA__375__A _391_/A vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_0_in_2.INVTX1_8_.scs8hd_inv_1_A top_width_0_height_0__pin_8_
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_1_in_3.mux_l1_in_2_.TGATE_3_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_1_in_3.INVTX1_11_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mem_fle_3_in_3.LATCH_3_.latch data_in ltile_clb_0.mem_fle_3_in_3.LATCH_3_.latch/Q
+ _335_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_ltile_clb_0.mem_fle_3_in_2.LATCH_3_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_14_.scs8hd_inv_1_A
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_14_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_1_501 vgnd vpwr scs8hd_decap_12
XFILLER_49_505 vgnd vpwr scs8hd_decap_8
XFILLER_76_335 vgnd vpwr scs8hd_fill_1
X_623_ _623_/A _623_/Y vgnd vpwr scs8hd_inv_8
XFILLER_29_240 vgnd vpwr scs8hd_decap_4
X_554_ _553_/X _554_/X vgnd vpwr scs8hd_buf_1
XFILLER_44_254 vgnd vpwr scs8hd_decap_3
Xltile_clb_0.mux_fle_2_in_2.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_2_in_2.INVTX1_10_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_2_in_2.LATCH_2_.latch/Q ltile_clb_0.mux_fle_2_in_2.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA__285__A _267_/X vgnd vpwr scs8hd_diode_2
X_485_ _314_/A _484_/X _485_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_44_276 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mem_fle_3_in_3.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_8_166 vgnd vpwr scs8hd_decap_12
XFILLER_32_80 vgnd vpwr scs8hd_decap_12
XFILLER_8_199 vgnd vpwr scs8hd_decap_3
XFILLER_4_372 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_1_in_3.INVTX1_5_.scs8hd_inv_1_A right_width_0_height_0__pin_5_
+ vgnd vpwr scs8hd_diode_2
XFILLER_79_184 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.mem_ble4_out_0.LATCH_1_.latch
+ data_in ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.mem_ble4_out_0.LATCH_1_.latch/Q
+ _576_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_ltile_clb_0.mux_fle_2_in_0.INVTX1_1_.scs8hd_inv_1_A right_width_0_height_0__pin_1_
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_3_in_1.INVTX1_9_.scs8hd_inv_1 right_width_0_height_0__pin_9_
+ ltile_clb_0.mux_fle_3_in_1.INVTX1_9_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XANTENNA_ltile_clb_0.mux_fle_1_in_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_1_in_3.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_50_224 vgnd vpwr scs8hd_decap_8
XFILLER_31_471 vgnd vpwr scs8hd_decap_6
XFILLER_31_493 vgnd vpwr scs8hd_decap_12
XFILLER_2_309 vgnd vpwr scs8hd_decap_8
XFILLER_58_302 vgnd vpwr scs8hd_decap_6
XFILLER_58_346 vgnd vpwr scs8hd_decap_4
XFILLER_58_335 vgnd vpwr scs8hd_fill_1
XFILLER_73_349 vpwr vgnd scs8hd_fill_2
XFILLER_26_210 vgnd vpwr scs8hd_decap_4
XFILLER_81_382 vpwr vgnd scs8hd_fill_2
XFILLER_14_416 vgnd vpwr scs8hd_decap_8
XFILLER_26_276 vpwr vgnd scs8hd_fill_2
XFILLER_26_287 vpwr vgnd scs8hd_fill_2
XFILLER_41_213 vgnd vpwr scs8hd_decap_4
XFILLER_41_224 vgnd vpwr scs8hd_decap_3
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_5_.TGATE_1_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_11_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
X_270_ _258_/X _270_/B _339_/A vgnd vpwr scs8hd_or2_4
XANTENNA__552__B address[7] vgnd vpwr scs8hd_diode_2
XFILLER_5_147 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mux_fle_0_in_3.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_0_in_3.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_78_32 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mux_fle_0_in_1.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_0_in_1.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_76_154 vgnd vpwr scs8hd_decap_12
XFILLER_64_316 vgnd vpwr scs8hd_decap_3
XFILLER_37_508 vgnd vpwr scs8hd_decap_8
XFILLER_64_349 vgnd vpwr scs8hd_decap_3
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_7_.latch_D
+ data_in vgnd vpwr scs8hd_diode_2
Xltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.buf4_2_.scs8hd_buf_1
+ ltile_clb_0.mux_fle_3_in_2.INVTX1_14_.scs8hd_inv_1/Y _608_/A vgnd vpwr scs8hd_buf_1
XANTENNA_ltile_clb_0.mux_fle_3_in_2.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_3_in_2.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_3_in_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_3_in_1.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_6_.scs8hd_inv_1_A
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_6_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_17_232 vgnd vpwr scs8hd_decap_4
XFILLER_17_254 vpwr vgnd scs8hd_fill_2
X_606_ _606_/A _606_/Y vgnd vpwr scs8hd_inv_8
XFILLER_72_382 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.mem_ble4_out_0.LATCH_1_.latch_D
+ data_in vgnd vpwr scs8hd_diode_2
X_537_ _272_/X _541_/B _537_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
+ _612_/Y vgnd vpwr scs8hd_diode_2
XFILLER_32_213 vgnd vpwr scs8hd_fill_1
XANTENNA_ltile_clb_0.mem_fle_0_in_2.LATCH_0_.latch_SLEEPB _503_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_3_in_3.INVTX1_11_.scs8hd_inv_1_A left_width_0_height_0__pin_11_
+ vgnd vpwr scs8hd_diode_2
X_468_ _435_/A _462_/X _468_/Y vgnd vpwr scs8hd_nor2_4
X_399_ _388_/A _399_/B _399_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_9_431 vpwr vgnd scs8hd_fill_2
XFILLER_57_3 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_0_.TGATE_1_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.INVTX1_0_.scs8hd_inv_1_A
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.INVTX1_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_3_in_1.mux_l1_in_2_.TGATE_3_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_3_in_1.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_67_110 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.mux_fle_0_in_0.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_0_in_0.INVTX1_9_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_0_in_0.LATCH_1_.latch/Q ltile_clb_0.mux_fle_0_in_0.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
Xltile_clb_0.mux_fle_2_in_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_2_in_0.INVTX1_4_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_2_in_0.LATCH_0_.latch/Q ltile_clb_0.mux_fle_2_in_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_82_168 vgnd vpwr scs8hd_decap_12
XPHY_709 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_63_371 vpwr vgnd scs8hd_fill_2
XFILLER_11_419 vpwr vgnd scs8hd_fill_2
XFILLER_23_27 vgnd vpwr scs8hd_decap_12
XANTENNA__372__B _377_/B vgnd vpwr scs8hd_diode_2
XFILLER_2_117 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_3_.TGATE_1_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_7_.TGATE_0_.scs8hd_ebufn_2/Z
+ _630_/Y ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_1_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_58_154 vpwr vgnd scs8hd_fill_2
XFILLER_46_305 vpwr vgnd scs8hd_fill_2
XFILLER_48_68 vgnd vpwr scs8hd_decap_12
XFILLER_73_135 vgnd vpwr scs8hd_decap_8
XFILLER_58_198 vpwr vgnd scs8hd_fill_2
XFILLER_46_327 vgnd vpwr scs8hd_decap_3
XFILLER_73_168 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.mux_fle_1_in_3.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_1_in_3.INVTX1_10_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_1_in_3.LATCH_2_.latch/Q ltile_clb_0.mux_fle_1_in_3.mux_l1_in_2_.TGATE_3_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA__547__B _526_/X vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_3_in_3.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_3_in_3.INVTX1_5_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_3_in_3.LATCH_1_.latch/Q ltile_clb_0.mux_fle_3_in_3.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_64_56 vgnd vpwr scs8hd_decap_12
XFILLER_54_360 vgnd vpwr scs8hd_fill_1
XFILLER_42_511 vgnd vpwr scs8hd_decap_4
XFILLER_14_235 vgnd vpwr scs8hd_decap_4
X_322_ _341_/B _338_/B vgnd vpwr scs8hd_buf_1
XFILLER_14_279 vgnd vpwr scs8hd_decap_3
XFILLER_80_44 vgnd vpwr scs8hd_decap_12
XANTENNA__563__A _272_/X vgnd vpwr scs8hd_diode_2
X_253_ _252_/X _603_/A vgnd vpwr scs8hd_buf_1
XANTENNA__282__B _282_/B vgnd vpwr scs8hd_diode_2
XFILLER_10_463 vgnd vpwr scs8hd_fill_1
XFILLER_6_445 vgnd vpwr scs8hd_decap_12
XFILLER_69_419 vgnd vpwr scs8hd_decap_6
XANTENNA_ltile_clb_0.mem_fle_1_in_1.LATCH_0_.latch_SLEEPB _470_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_0_in_3.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_0_in_3.INVTX1_13_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_49_110 vgnd vpwr scs8hd_decap_12
XFILLER_77_474 vgnd vpwr scs8hd_decap_12
XFILLER_77_463 vpwr vgnd scs8hd_fill_2
XFILLER_37_349 vpwr vgnd scs8hd_fill_2
XANTENNA__457__B _451_/X vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_60_341 vgnd vpwr scs8hd_decap_4
XFILLER_45_382 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_3_in_1.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_3_in_1.INVTX1_13_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_20_227 vpwr vgnd scs8hd_fill_2
XANTENNA__473__A _481_/B vgnd vpwr scs8hd_diode_2
XFILLER_18_27 vgnd vpwr scs8hd_decap_4
XFILLER_28_316 vgnd vpwr scs8hd_decap_3
XANTENNA__367__B _368_/B vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
+ _630_/Y vgnd vpwr scs8hd_diode_2
XFILLER_70_105 vgnd vpwr scs8hd_decap_12
XFILLER_55_179 vpwr vgnd scs8hd_fill_2
XFILLER_55_168 vpwr vgnd scs8hd_fill_2
XFILLER_36_371 vgnd vpwr scs8hd_decap_4
XFILLER_43_319 vgnd vpwr scs8hd_decap_6
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_2_.latch_SLEEPB
+ _544_/Y vgnd vpwr scs8hd_diode_2
XFILLER_34_15 vgnd vpwr scs8hd_decap_12
XFILLER_36_393 vpwr vgnd scs8hd_fill_2
XPHY_506 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_517 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_51_374 vpwr vgnd scs8hd_fill_2
XPHY_528 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_539 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__383__A address[8] vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_3_in_2.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_3_in_2.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_78_227 vgnd vpwr scs8hd_decap_12
XFILLER_59_441 vpwr vgnd scs8hd_fill_2
XFILLER_59_496 vpwr vgnd scs8hd_fill_2
XANTENNA__558__A _250_/X vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_1_in_2.INVTX1_10_.scs8hd_inv_1_A bottom_width_0_height_0__pin_10_
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l4_in_0_.TGATE_1_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ _626_/Y ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_16_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA__277__B _564_/A vgnd vpwr scs8hd_diode_2
XFILLER_27_360 vpwr vgnd scs8hd_fill_2
XFILLER_34_308 vpwr vgnd scs8hd_fill_2
XFILLER_34_319 vgnd vpwr scs8hd_decap_6
XFILLER_46_168 vgnd vpwr scs8hd_decap_4
XFILLER_27_393 vgnd vpwr scs8hd_decap_4
XANTENNA_ltile_clb_0.mux_fle_3_in_0.INVTX1_7_.scs8hd_inv_1_A left_width_0_height_0__pin_7_
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.tap_buf4_0_.scs8hd_inv_1_A
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mem_fle_2_in_0.LATCH_0_.latch_SLEEPB _437_/Y vgnd vpwr scs8hd_diode_2
XANTENNA__293__A _278_/X vgnd vpwr scs8hd_diode_2
X_305_ _282_/C _282_/B _305_/X vgnd vpwr scs8hd_or2_4
XFILLER_42_396 vgnd vpwr scs8hd_fill_1
X_236_ _246_/A _236_/X vgnd vpwr scs8hd_buf_1
XFILLER_6_242 vgnd vpwr scs8hd_decap_3
XFILLER_6_264 vgnd vpwr scs8hd_decap_8
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_4_.TGATE_0_.scs8hd_ebufn_2_TEB
+ _621_/Y vgnd vpwr scs8hd_diode_2
XFILLER_40_80 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_8_.scs8hd_inv_1_A
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_8_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_1_in_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_1_in_1.INVTX1_4_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_1_in_1.LATCH_0_.latch/Q ltile_clb_0.mux_fle_1_in_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA__468__A _435_/A vgnd vpwr scs8hd_diode_2
XFILLER_65_444 vpwr vgnd scs8hd_fill_2
XFILLER_1_74 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.INVTX1_1_.scs8hd_inv_1/Y
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.mem_ble4_out_0.LATCH_1_.latch/Q
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_37_135 vgnd vpwr scs8hd_decap_6
XFILLER_80_403 vgnd vpwr scs8hd_decap_12
XFILLER_52_105 vgnd vpwr scs8hd_decap_12
XFILLER_18_371 vpwr vgnd scs8hd_fill_2
XFILLER_37_168 vpwr vgnd scs8hd_fill_2
XFILLER_37_179 vpwr vgnd scs8hd_fill_2
XFILLER_80_436 vpwr vgnd scs8hd_fill_2
XFILLER_18_382 vgnd vpwr scs8hd_decap_4
XFILLER_21_503 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_5_.TGATE_1_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_11_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_9_.scs8hd_inv_1
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_9_.latch/Q
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_9_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_ltile_clb_0.mux_fle_2_in_0.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_2_in_0.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_29_15 vgnd vpwr scs8hd_decap_12
XFILLER_75_208 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.mem_ble4_out_0.LATCH_1_.latch
+ data_in ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.mem_ble4_out_0.LATCH_1_.latch/Q
+ _311_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_29_59 vpwr vgnd scs8hd_fill_2
XFILLER_68_260 vpwr vgnd scs8hd_fill_2
XANTENNA__378__A _394_/A vgnd vpwr scs8hd_diode_2
XFILLER_56_411 vgnd vpwr scs8hd_decap_8
Xltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.INVTX1_0_.scs8hd_inv_1
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.INVTX1_0_.scs8hd_inv_1/A
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_16_308 vgnd vpwr scs8hd_decap_4
XFILLER_71_436 vpwr vgnd scs8hd_fill_2
XPHY_303 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_314 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_325 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_363 vpwr vgnd scs8hd_fill_2
XPHY_336 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_347 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_358 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_369 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_51_193 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_3_in_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_3_in_0.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__560__B _558_/B vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_3_in_2.mux_l1_in_2_.TGATE_3_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_3_in_2.INVTX1_11_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_3_245 vpwr vgnd scs8hd_fill_2
XFILLER_59_282 vpwr vgnd scs8hd_fill_2
XANTENNA__288__A _287_/X vgnd vpwr scs8hd_diode_2
XFILLER_47_400 vpwr vgnd scs8hd_fill_2
XFILLER_47_422 vgnd vpwr scs8hd_decap_4
XFILLER_19_135 vgnd vpwr scs8hd_decap_12
XANTENNA__438__D _358_/D vgnd vpwr scs8hd_diode_2
XFILLER_19_179 vgnd vpwr scs8hd_fill_1
XFILLER_34_105 vgnd vpwr scs8hd_decap_12
XFILLER_47_466 vgnd vpwr scs8hd_fill_1
XFILLER_74_296 vgnd vpwr scs8hd_decap_3
XANTENNA_ltile_clb_0.mux_fle_1_in_0.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_1_in_0.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_15_352 vpwr vgnd scs8hd_fill_2
XFILLER_15_374 vgnd vpwr scs8hd_decap_4
Xltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ _606_/Y ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_42_182 vgnd vpwr scs8hd_decap_4
XFILLER_30_344 vgnd vpwr scs8hd_decap_12
XFILLER_30_366 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_1_in_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_1_in_1.LATCH_5_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__470__B _461_/X vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_1_in_0.INVTX1_4_.scs8hd_inv_1 top_width_0_height_0__pin_4_ ltile_clb_0.mux_fle_1_in_0.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_53_414 vpwr vgnd scs8hd_fill_2
XFILLER_53_403 vpwr vgnd scs8hd_fill_2
XFILLER_53_447 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mem_fle_0_in_0.LATCH_1_.latch_SLEEPB _524_/Y vgnd vpwr scs8hd_diode_2
XFILLER_15_39 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mux_fle_3_in_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_3_in_2.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_31_27 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mux_fle_0_in_1.INVTX1_14_.scs8hd_inv_1_A ltile_clb_0.mux_fle_0_in_1.INVTX1_14_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_0_in_0.INVTX1_5_.scs8hd_inv_1_A right_width_0_height_0__pin_5_
+ vgnd vpwr scs8hd_diode_2
XFILLER_29_400 vgnd vpwr scs8hd_decap_4
XFILLER_71_200 vgnd vpwr scs8hd_fill_1
XFILLER_56_263 vgnd vpwr scs8hd_fill_1
XFILLER_56_68 vgnd vpwr scs8hd_decap_12
XFILLER_16_105 vgnd vpwr scs8hd_decap_12
X_570_ _544_/A _554_/X _570_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_29_477 vpwr vgnd scs8hd_fill_2
XFILLER_44_403 vpwr vgnd scs8hd_fill_2
XFILLER_56_285 vpwr vgnd scs8hd_fill_2
XPHY_100 vgnd vpwr scs8hd_decap_3
XFILLER_72_56 vgnd vpwr scs8hd_decap_12
XPHY_133 vgnd vpwr scs8hd_decap_3
XPHY_122 vgnd vpwr scs8hd_decap_3
XPHY_111 vgnd vpwr scs8hd_decap_3
XFILLER_12_311 vpwr vgnd scs8hd_fill_2
XPHY_155 vgnd vpwr scs8hd_decap_3
XPHY_144 vgnd vpwr scs8hd_decap_3
XFILLER_12_322 vgnd vpwr scs8hd_decap_12
XPHY_166 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_12_355 vgnd vpwr scs8hd_decap_6
XFILLER_8_337 vgnd vpwr scs8hd_decap_6
XPHY_177 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_188 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_199 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__571__A _545_/A vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_0_in_2.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_0_in_2.INVTX1_4_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_0_in_2.LATCH_0_.latch/Q ltile_clb_0.mux_fle_0_in_2.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA__290__B _330_/A vgnd vpwr scs8hd_diode_2
Xltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_4_.TGATE_0_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_8_.scs8hd_inv_1/Y
+ _621_/Y ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_2_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_ltile_clb_0.mux_fle_2_in_2.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_2_in_2.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_79_355 vgnd vpwr scs8hd_decap_3
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_7_.latch_SLEEPB
+ _591_/Y vgnd vpwr scs8hd_diode_2
XFILLER_82_509 vgnd vpwr scs8hd_decap_6
XANTENNA__449__C _384_/X vgnd vpwr scs8hd_diode_2
XFILLER_35_403 vpwr vgnd scs8hd_fill_2
XFILLER_47_263 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_3_in_3.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_3_in_3.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_62_266 vpwr vgnd scs8hd_fill_2
XPHY_2 vgnd vpwr scs8hd_decap_3
XANTENNA_ltile_clb_0.mux_fle_1_in_1.INVTX1_2_.scs8hd_inv_1_A bottom_width_0_height_0__pin_2_
+ vgnd vpwr scs8hd_diode_2
XFILLER_15_171 vgnd vpwr scs8hd_fill_1
XANTENNA__465__B _462_/X vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_0_in_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_0_in_0.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xclkbuf_0_clk clk clkbuf_0_clk/X vgnd vpwr scs8hd_clkbuf_16
XFILLER_30_141 vgnd vpwr scs8hd_decap_12
XANTENNA__481__A _437_/A vgnd vpwr scs8hd_diode_2
XFILLER_7_62 vgnd vpwr scs8hd_decap_12
XFILLER_7_51 vgnd vpwr scs8hd_decap_8
XFILLER_7_370 vgnd vpwr scs8hd_decap_4
Xltile_clb_0.mux_fle_1_in_1.INVTX1_8_.scs8hd_inv_1 top_width_0_height_0__pin_8_ ltile_clb_0.mux_fle_1_in_1.INVTX1_8_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_53_222 vpwr vgnd scs8hd_fill_2
XFILLER_26_27 vgnd vpwr scs8hd_decap_4
XFILLER_26_414 vgnd vpwr scs8hd_decap_4
XFILLER_38_274 vgnd vpwr scs8hd_fill_1
XFILLER_38_285 vgnd vpwr scs8hd_decap_3
XFILLER_38_296 vgnd vpwr scs8hd_fill_1
XANTENNA__375__B _377_/B vgnd vpwr scs8hd_diode_2
XFILLER_41_417 vpwr vgnd scs8hd_fill_2
XFILLER_41_428 vgnd vpwr scs8hd_decap_3
XFILLER_42_15 vgnd vpwr scs8hd_decap_12
XANTENNA__391__A _391_/A vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_3_.scs8hd_inv_1_A
+ ltile_clb_0.mux_fle_1_in_3.INVTX1_14_.scs8hd_inv_1/Y vgnd vpwr scs8hd_diode_2
XFILLER_1_513 vgnd vpwr scs8hd_decap_3
XFILLER_76_325 vpwr vgnd scs8hd_fill_2
XFILLER_76_358 vgnd vpwr scs8hd_decap_8
XFILLER_76_369 vpwr vgnd scs8hd_fill_2
X_622_ _622_/A _622_/Y vgnd vpwr scs8hd_inv_8
XFILLER_29_252 vpwr vgnd scs8hd_fill_2
XFILLER_29_263 vpwr vgnd scs8hd_fill_2
XANTENNA__566__A _540_/A vgnd vpwr scs8hd_diode_2
XFILLER_44_200 vgnd vpwr scs8hd_decap_3
XFILLER_44_222 vgnd vpwr scs8hd_decap_3
X_553_ address[4] _552_/X _553_/X vgnd vpwr scs8hd_or2_4
XANTENNA__285__B _540_/A vgnd vpwr scs8hd_diode_2
XFILLER_32_439 vpwr vgnd scs8hd_fill_2
XFILLER_44_266 vpwr vgnd scs8hd_fill_2
XFILLER_44_299 vgnd vpwr scs8hd_decap_4
X_484_ _492_/B _484_/X vgnd vpwr scs8hd_buf_1
XFILLER_16_93 vgnd vpwr scs8hd_decap_12
XFILLER_12_141 vgnd vpwr scs8hd_decap_12
XFILLER_8_178 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_1_.scs8hd_inv_1/Y
+ _628_/Y ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_4_340 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.mux_fle_2_in_2.INVTX1_3_.scs8hd_inv_1 left_width_0_height_0__pin_3_ ltile_clb_0.mux_fle_2_in_2.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_79_196 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mux_fle_2_in_2.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_2_in_2.INVTX1_13_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
+ _617_/Y vgnd vpwr scs8hd_diode_2
Xltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_1_.TGATE_0_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_1_.TGATE_0_.scs8hd_ebufn_2/A
+ _617_/Y ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l4_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_75_380 vgnd vpwr scs8hd_fill_1
XANTENNA__476__A _432_/A vgnd vpwr scs8hd_diode_2
XFILLER_35_255 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_2_in_2.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_2_in_2.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_2_.scs8hd_inv_1
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_2_.latch/Q
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_50_247 vpwr vgnd scs8hd_fill_2
XFILLER_31_450 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_0_in_0.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_0_in_0.INVTX1_9_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_37_15 vgnd vpwr scs8hd_decap_12
XFILLER_73_306 vgnd vpwr scs8hd_decap_4
Xltile_clb_0.mux_fle_3_in_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_3_in_2.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ ltile_clb_0.mem_fle_3_in_2.LATCH_4_.latch/Q ltile_clb_0.mux_fle_3_in_2.INVTX1_14_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_ltile_clb_0.mux_fle_2_in_3.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_2_in_3.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_37_59 vpwr vgnd scs8hd_fill_2
XANTENNA__386__A _385_/X vgnd vpwr scs8hd_diode_2
XFILLER_14_406 vgnd vpwr scs8hd_fill_1
Xltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.INVTX1_1_.scs8hd_inv_1
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.INVTX1_1_.scs8hd_inv_1/A
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_41_236 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mem_fle_3_in_3.LATCH_6_.latch_SLEEPB _326_/Y vgnd vpwr scs8hd_diode_2
XANTENNA__552__C _227_/X vgnd vpwr scs8hd_diode_2
XFILLER_5_159 vgnd vpwr scs8hd_decap_12
XFILLER_78_44 vgnd vpwr scs8hd_decap_12
XFILLER_1_387 vpwr vgnd scs8hd_fill_2
XFILLER_49_336 vgnd vpwr scs8hd_decap_3
XFILLER_49_358 vpwr vgnd scs8hd_fill_2
XFILLER_64_328 vgnd vpwr scs8hd_decap_8
XFILLER_57_380 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_2_in_0.INVTX1_12_.scs8hd_inv_1_A top_width_0_height_0__pin_12_
+ vgnd vpwr scs8hd_diode_2
XANTENNA__296__A _282_/C vgnd vpwr scs8hd_diode_2
X_605_ _605_/A _605_/Y vgnd vpwr scs8hd_inv_8
XFILLER_17_288 vpwr vgnd scs8hd_fill_2
X_536_ _528_/X _541_/B vgnd vpwr scs8hd_buf_1
XFILLER_20_409 vpwr vgnd scs8hd_fill_2
X_467_ _434_/A _462_/X _467_/Y vgnd vpwr scs8hd_nor2_4
X_398_ _398_/A _399_/B vgnd vpwr scs8hd_buf_1
Xltile_clb_0.mux_fle_2_in_3.INVTX1_7_.scs8hd_inv_1 left_width_0_height_0__pin_7_ ltile_clb_0.mux_fle_2_in_3.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
Xltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_7_.latch
+ data_in ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_7_.latch/Q
+ _281_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_9_498 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_1_.TGATE_1_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_1_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_82_125 vgnd vpwr scs8hd_decap_12
XFILLER_55_317 vgnd vpwr scs8hd_decap_3
Xltile_clb_0.mux_fle_2_in_0.INVTX1_13_.scs8hd_inv_1 right_width_0_height_0__pin_13_
+ ltile_clb_0.mux_fle_2_in_0.INVTX1_13_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XFILLER_23_258 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_1_in_1.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_1_in_1.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_23_39 vgnd vpwr scs8hd_decap_12
XFILLER_2_129 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l4_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
+ _635_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_3_in_2.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_3_in_2.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_46_317 vgnd vpwr scs8hd_fill_1
XFILLER_61_309 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB
+ _613_/Y vgnd vpwr scs8hd_diode_2
XFILLER_64_68 vgnd vpwr scs8hd_decap_12
XFILLER_54_372 vpwr vgnd scs8hd_fill_2
XFILLER_54_350 vgnd vpwr scs8hd_decap_4
XANTENNA_ltile_clb_0.mux_fle_2_in_3.mux_l1_in_2_.TGATE_3_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_2_in_3.INVTX1_11_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
X_321_ _320_/X _341_/B vgnd vpwr scs8hd_buf_1
XFILLER_80_56 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mux_fle_2_in_1.INVTX1_8_.scs8hd_inv_1_A top_width_0_height_0__pin_8_
+ vgnd vpwr scs8hd_diode_2
XANTENNA__563__B _564_/B vgnd vpwr scs8hd_diode_2
X_252_ _282_/C address[1] _252_/X vgnd vpwr scs8hd_or2_4
Xltile_clb_0.mux_fle_3_in_0.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_3_in_0.INVTX1_10_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_3_in_0.LATCH_2_.latch/Q ltile_clb_0.mux_fle_3_in_0.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA__282__C _282_/C vgnd vpwr scs8hd_diode_2
XFILLER_6_468 vpwr vgnd scs8hd_fill_2
XFILLER_6_457 vgnd vpwr scs8hd_fill_1
XFILLER_69_409 vgnd vpwr scs8hd_decap_4
XANTENNA_ltile_clb_0.mux_fle_0_in_1.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_0_in_1.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_3_in_1.mux_l1_in_3_.TGATE_2_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_3_in_1.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_77_431 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_1_in_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_1_in_3.LATCH_4_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_1_184 vgnd vpwr scs8hd_decap_12
XFILLER_77_442 vpwr vgnd scs8hd_fill_2
XFILLER_77_486 vpwr vgnd scs8hd_fill_2
XFILLER_37_339 vgnd vpwr scs8hd_fill_1
XFILLER_38_80 vgnd vpwr scs8hd_decap_12
XFILLER_49_199 vgnd vpwr scs8hd_decap_4
XFILLER_64_158 vgnd vpwr scs8hd_decap_3
XANTENNA_ltile_clb_0.mem_fle_1_in_3.LATCH_7_.latch_SLEEPB _441_/Y vgnd vpwr scs8hd_diode_2
X_519_ _325_/A _517_/X _519_/Y vgnd vpwr scs8hd_nor2_4
Xltile_clb_0.mux_fle_2_in_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_2_in_3.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ ltile_clb_0.mem_fle_2_in_3.LATCH_4_.latch/Q ltile_clb_0.mux_fle_2_in_3.INVTX1_14_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_68_420 vgnd vpwr scs8hd_decap_8
XANTENNA_ltile_clb_0.mux_fle_3_in_2.INVTX1_5_.scs8hd_inv_1_A right_width_0_height_0__pin_5_
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_2_in_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_2_in_3.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_28_328 vpwr vgnd scs8hd_fill_2
XFILLER_55_136 vpwr vgnd scs8hd_fill_2
XFILLER_70_117 vgnd vpwr scs8hd_decap_12
XFILLER_34_27 vgnd vpwr scs8hd_decap_4
XPHY_507 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_0_.latch_SLEEPB
+ _304_/Y vgnd vpwr scs8hd_diode_2
XPHY_518 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_529 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__383__B _369_/B vgnd vpwr scs8hd_diode_2
XFILLER_50_15 vgnd vpwr scs8hd_decap_12
XFILLER_3_438 vpwr vgnd scs8hd_fill_2
XFILLER_78_239 vgnd vpwr scs8hd_decap_8
XFILLER_74_401 vgnd vpwr scs8hd_decap_4
XFILLER_59_475 vpwr vgnd scs8hd_fill_2
XANTENNA__558__B _558_/B vgnd vpwr scs8hd_diode_2
Xltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_7_.latch
+ data_in ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_7_.latch/Q
+ _591_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_54_191 vgnd vpwr scs8hd_decap_8
XANTENNA__574__A _573_/X vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_1_in_3.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_1_in_3.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
X_304_ _304_/A _546_/A _304_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA__293__B _333_/A vgnd vpwr scs8hd_diode_2
XFILLER_42_375 vgnd vpwr scs8hd_decap_4
XFILLER_42_386 vpwr vgnd scs8hd_fill_2
X_235_ address[3] _246_/A vgnd vpwr scs8hd_inv_8
XFILLER_24_93 vgnd vpwr scs8hd_decap_12
XFILLER_10_272 vgnd vpwr scs8hd_decap_3
XFILLER_6_276 vgnd vpwr scs8hd_decap_3
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.INVTX1_1_.scs8hd_inv_1_A
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.INVTX1_1_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_69_206 vgnd vpwr scs8hd_decap_8
XANTENNA_ltile_clb_0.mem_fle_2_in_2.LATCH_7_.latch_SLEEPB _399_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_2_in_0.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_2_in_0.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_77_283 vpwr vgnd scs8hd_fill_2
XANTENNA__468__B _462_/X vgnd vpwr scs8hd_diode_2
XFILLER_77_294 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
+ _631_/Y vgnd vpwr scs8hd_diode_2
XFILLER_80_415 vgnd vpwr scs8hd_decap_6
XFILLER_1_86 vgnd vpwr scs8hd_decap_12
XFILLER_80_459 vgnd vpwr scs8hd_decap_12
XFILLER_52_128 vgnd vpwr scs8hd_decap_8
XFILLER_52_117 vgnd vpwr scs8hd_decap_8
XANTENNA__484__A _492_/B vgnd vpwr scs8hd_diode_2
XFILLER_60_150 vgnd vpwr scs8hd_decap_3
XFILLER_21_515 vgnd vpwr scs8hd_fill_1
XANTENNA_ltile_clb_0.mux_fle_0_in_1.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_0_in_1.LATCH_6_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_29_27 vgnd vpwr scs8hd_decap_12
XANTENNA__378__B _379_/B vgnd vpwr scs8hd_diode_2
XFILLER_68_294 vgnd vpwr scs8hd_fill_1
XFILLER_45_15 vgnd vpwr scs8hd_decap_12
XFILLER_45_59 vpwr vgnd scs8hd_fill_2
XANTENNA__394__A _394_/A vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_2_in_1.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_2_in_1.INVTX1_10_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_2_in_1.LATCH_2_.latch/Q ltile_clb_0.mux_fle_2_in_1.mux_l1_in_2_.TGATE_3_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XPHY_304 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_315 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_12_504 vgnd vpwr scs8hd_decap_12
XPHY_326 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_337 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_348 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_359 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_8_508 vgnd vpwr scs8hd_decap_8
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.mem_ble4_out_0.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_1_in_2.INVTX1_11_.scs8hd_inv_1 left_width_0_height_0__pin_11_
+ ltile_clb_0.mux_fle_1_in_2.INVTX1_11_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XFILLER_3_235 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.buf4_0_.scs8hd_buf_1_A
+ ltile_clb_0.mux_fle_3_in_0.INVTX1_14_.scs8hd_inv_1/Y vgnd vpwr scs8hd_diode_2
XFILLER_3_279 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_1_.TGATE_1_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_1_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XANTENNA__569__A _569_/A vgnd vpwr scs8hd_diode_2
XFILLER_19_147 vgnd vpwr scs8hd_decap_12
XFILLER_19_169 vpwr vgnd scs8hd_fill_2
XFILLER_34_117 vgnd vpwr scs8hd_decap_12
XFILLER_62_459 vgnd vpwr scs8hd_decap_3
XFILLER_30_312 vgnd vpwr scs8hd_decap_8
XANTENNA_ltile_clb_0.mux_fle_0_in_2.INVTX1_3_.scs8hd_inv_1_A left_width_0_height_0__pin_3_
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mem_fle_3_in_1.LATCH_7_.latch_SLEEPB _361_/Y vgnd vpwr scs8hd_diode_2
XFILLER_30_356 vgnd vpwr scs8hd_fill_1
XANTENNA_ltile_clb_0.mux_fle_1_in_3.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_1_in_3.INVTX1_13_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_32_3 vgnd vpwr scs8hd_decap_12
XANTENNA__479__A _435_/A vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_3_in_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_3_in_1.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_1_in_3.INVTX1_13_.scs8hd_inv_1 right_width_0_height_0__pin_13_
+ ltile_clb_0.mux_fle_1_in_3.INVTX1_13_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XFILLER_38_401 vgnd vpwr scs8hd_decap_8
XFILLER_38_412 vgnd vpwr scs8hd_decap_3
XFILLER_65_275 vpwr vgnd scs8hd_fill_2
XFILLER_65_297 vpwr vgnd scs8hd_fill_2
XFILLER_53_426 vgnd vpwr scs8hd_fill_1
XFILLER_61_481 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_2_in_3.mux_l1_in_2_.TGATE_3_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_2_in_3.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_31_39 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mux_fle_3_in_0.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_3_in_0.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_1_in_3.INVTX1_0_.scs8hd_inv_1_A top_width_0_height_0__pin_0_
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_7_.latch
+ data_in ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_7_.latch/Q
+ _565_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA__389__A _326_/A vgnd vpwr scs8hd_diode_2
XFILLER_0_249 vgnd vpwr scs8hd_decap_4
XFILLER_0_238 vgnd vpwr scs8hd_decap_8
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__ff_0.DFFSRQ_0_.dff_CLK
+ clkbuf_1_1_0_clk/X vgnd vpwr scs8hd_diode_2
XFILLER_29_423 vpwr vgnd scs8hd_fill_2
XFILLER_71_212 vgnd vpwr scs8hd_decap_3
XFILLER_16_117 vgnd vpwr scs8hd_decap_12
XFILLER_71_245 vpwr vgnd scs8hd_fill_2
XFILLER_72_68 vgnd vpwr scs8hd_decap_12
XFILLER_71_278 vgnd vpwr scs8hd_decap_6
XPHY_134 vgnd vpwr scs8hd_decap_3
XPHY_123 vgnd vpwr scs8hd_decap_3
XPHY_112 vgnd vpwr scs8hd_decap_3
XFILLER_12_301 vgnd vpwr scs8hd_fill_1
XPHY_101 vgnd vpwr scs8hd_decap_3
XPHY_156 vgnd vpwr scs8hd_decap_3
XPHY_145 vgnd vpwr scs8hd_decap_3
XFILLER_12_334 vpwr vgnd scs8hd_fill_2
XPHY_167 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_178 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_189 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_ltile_clb_0.mux_fle_0_in_3.INVTX1_12_.scs8hd_inv_1_A top_width_0_height_0__pin_12_
+ vgnd vpwr scs8hd_diode_2
XFILLER_12_389 vgnd vpwr scs8hd_decap_8
XFILLER_8_349 vgnd vpwr scs8hd_decap_8
XANTENNA__571__B _554_/X vgnd vpwr scs8hd_diode_2
XFILLER_79_301 vpwr vgnd scs8hd_fill_2
XANTENNA__299__A _286_/B vgnd vpwr scs8hd_diode_2
XANTENNA__449__D _346_/D vgnd vpwr scs8hd_diode_2
Xltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_2_.TGATE_1_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_2_.TGATE_1_.scs8hd_ebufn_2/A
+ _614_/Y ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_1_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
Xltile_clb_0.mux_fle_0_in_2.INVTX1_2_.scs8hd_inv_1 bottom_width_0_height_0__pin_2_
+ ltile_clb_0.mux_fle_0_in_2.INVTX1_2_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XFILLER_47_297 vpwr vgnd scs8hd_fill_2
XPHY_3 vgnd vpwr scs8hd_decap_3
XFILLER_46_80 vgnd vpwr scs8hd_decap_12
XFILLER_43_492 vpwr vgnd scs8hd_fill_2
XPHY_690 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__481__B _481_/B vgnd vpwr scs8hd_diode_2
XFILLER_7_74 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mux_fle_0_in_2.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_0_in_2.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_1_in_2.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_1_in_2.INVTX1_10_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_1_in_2.LATCH_2_.latch/Q ltile_clb_0.mux_fle_1_in_2.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_38_264 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.mux_fle_3_in_2.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_3_in_2.INVTX1_5_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_3_in_2.LATCH_1_.latch/Q ltile_clb_0.mux_fle_3_in_2.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_1_.scs8hd_inv_1_A
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_53_245 vgnd vpwr scs8hd_decap_3
XFILLER_53_267 vgnd vpwr scs8hd_decap_3
XFILLER_42_27 vgnd vpwr scs8hd_decap_4
XANTENNA_ltile_clb_0.mux_fle_3_in_0.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_3_in_0.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XANTENNA__391__B _388_/B vgnd vpwr scs8hd_diode_2
XFILLER_5_319 vgnd vpwr scs8hd_decap_4
XFILLER_76_304 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_16_.scs8hd_inv_1_A
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_16_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_76_337 vpwr vgnd scs8hd_fill_2
XFILLER_29_220 vpwr vgnd scs8hd_fill_2
X_621_ _621_/A _621_/Y vgnd vpwr scs8hd_inv_8
XFILLER_29_231 vgnd vpwr scs8hd_decap_3
XFILLER_17_437 vgnd vpwr scs8hd_decap_3
XFILLER_29_297 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_3_in_3.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_3_in_3.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
X_552_ _380_/A address[7] _227_/X _345_/A _552_/X vgnd vpwr scs8hd_or4_4
XANTENNA__566__B _564_/B vgnd vpwr scs8hd_diode_2
XFILLER_17_459 vpwr vgnd scs8hd_fill_2
XFILLER_32_407 vgnd vpwr scs8hd_decap_6
X_483_ _482_/X _492_/B vgnd vpwr scs8hd_buf_1
XFILLER_25_481 vgnd vpwr scs8hd_fill_1
XANTENNA__582__A _556_/A vgnd vpwr scs8hd_diode_2
XFILLER_40_451 vgnd vpwr scs8hd_decap_6
Xltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_6_.TGATE_0_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_12_.scs8hd_inv_1/Y
+ _629_/Y ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_6_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_40_484 vgnd vpwr scs8hd_decap_4
XFILLER_32_93 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mux_fle_2_in_0.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_2_in_0.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_67_315 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_6_.TGATE_1_.scs8hd_ebufn_2_TEB
+ _612_/Y vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_0_in_3.INVTX1_6_.scs8hd_inv_1 bottom_width_0_height_0__pin_6_
+ ltile_clb_0.mux_fle_0_in_3.INVTX1_6_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XANTENNA__476__B _479_/B vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_12_.latch_D
+ data_in vgnd vpwr scs8hd_diode_2
XFILLER_35_245 vgnd vpwr scs8hd_fill_1
XFILLER_35_278 vgnd vpwr scs8hd_decap_4
XFILLER_16_481 vgnd vpwr scs8hd_fill_1
XANTENNA__492__A _343_/A vgnd vpwr scs8hd_diode_2
XFILLER_31_484 vgnd vpwr scs8hd_decap_4
Xltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_7_.latch
+ data_in ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_7_.latch/Q
+ _539_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
+ _605_/Y vgnd vpwr scs8hd_diode_2
XFILLER_37_27 vgnd vpwr scs8hd_decap_12
XFILLER_66_381 vgnd vpwr scs8hd_decap_4
XFILLER_53_15 vgnd vpwr scs8hd_decap_12
XFILLER_53_59 vpwr vgnd scs8hd_fill_2
XFILLER_41_259 vpwr vgnd scs8hd_fill_2
XANTENNA__552__D _345_/A vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_1_in_2.INVTX1_9_.scs8hd_inv_1_A right_width_0_height_0__pin_9_
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_11_.latch
+ data_in ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_11_.latch/Q
+ _560_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_78_56 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.mux_fle_1_in_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_1_in_0.INVTX1_4_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_1_in_0.LATCH_0_.latch/Q ltile_clb_0.mux_fle_1_in_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_1_333 vgnd vpwr scs8hd_decap_4
XFILLER_49_315 vgnd vpwr scs8hd_decap_6
Xltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
+ _639_/HI ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.mem_ble4_out_0.LATCH_2_.latch/Q
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_64_307 vpwr vgnd scs8hd_fill_2
XANTENNA__577__A _603_/A vgnd vpwr scs8hd_diode_2
XFILLER_17_201 vpwr vgnd scs8hd_fill_2
XFILLER_17_212 vgnd vpwr scs8hd_decap_4
XANTENNA__296__B _282_/B vgnd vpwr scs8hd_diode_2
X_604_ _604_/A _604_/Y vgnd vpwr scs8hd_inv_8
X_535_ _535_/A _529_/X _535_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_72_395 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_2_in_2.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_2_in_2.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_32_226 vgnd vpwr scs8hd_decap_8
XFILLER_32_248 vgnd vpwr scs8hd_decap_8
X_466_ _433_/A _462_/X _466_/Y vgnd vpwr scs8hd_nor2_4
X_397_ _397_/A _398_/A vgnd vpwr scs8hd_buf_1
XFILLER_9_422 vpwr vgnd scs8hd_fill_2
XFILLER_9_411 vpwr vgnd scs8hd_fill_2
XFILLER_13_462 vpwr vgnd scs8hd_fill_2
XFILLER_13_484 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_3_in_2.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_3_in_2.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_9_466 vgnd vpwr scs8hd_decap_3
Xltile_clb_0.mux_fle_2_in_3.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_2_in_3.INVTX1_5_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_2_in_3.LATCH_1_.latch/Q ltile_clb_0.mux_fle_2_in_3.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_67_123 vgnd vpwr scs8hd_decap_6
Xltile_clb_0.mux_fle_0_in_3.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_0_in_3.INVTX1_10_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_0_in_3.LATCH_2_.latch/Q ltile_clb_0.mux_fle_0_in_3.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_ltile_clb_0.mux_fle_2_in_3.INVTX1_6_.scs8hd_inv_1_A bottom_width_0_height_0__pin_6_
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_2_in_2.INVTX1_10_.scs8hd_inv_1_A bottom_width_0_height_0__pin_10_
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_1_in_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_1_in_0.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__487__A _328_/A vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_0_in_3.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_0_in_3.LATCH_5_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_48_370 vpwr vgnd scs8hd_fill_2
XFILLER_82_137 vgnd vpwr scs8hd_decap_12
XFILLER_48_381 vgnd vpwr scs8hd_decap_3
XFILLER_51_502 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_3_in_0.INVTX1_2_.scs8hd_inv_1_A bottom_width_0_height_0__pin_2_
+ vgnd vpwr scs8hd_diode_2
XFILLER_63_384 vpwr vgnd scs8hd_fill_2
XFILLER_23_215 vgnd vpwr scs8hd_decap_3
XFILLER_23_237 vgnd vpwr scs8hd_decap_4
Xltile_clb_0.mux_fle_2_in_0.INVTX1_3_.scs8hd_inv_1 left_width_0_height_0__pin_3_ ltile_clb_0.mux_fle_2_in_0.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_31_281 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_3_.scs8hd_inv_1_A
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_48_15 vgnd vpwr scs8hd_decap_12
XANTENNA__397__A _397_/A vgnd vpwr scs8hd_diode_2
XFILLER_58_134 vgnd vpwr scs8hd_decap_12
XFILLER_14_204 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.mem_fle_2_in_1.LATCH_7_.latch data_in ltile_clb_0.mem_fle_2_in_1.LATCH_7_.latch/Q
+ _412_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
X_320_ address[8] _369_/B _346_/C _358_/D _320_/X vgnd vpwr scs8hd_or4_4
XFILLER_54_395 vpwr vgnd scs8hd_fill_2
XFILLER_14_215 vgnd vpwr scs8hd_decap_6
XFILLER_14_259 vpwr vgnd scs8hd_fill_2
XFILLER_14_248 vpwr vgnd scs8hd_fill_2
X_251_ _248_/A _250_/X _251_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_80_68 vgnd vpwr scs8hd_decap_12
XFILLER_13_51 vgnd vpwr scs8hd_decap_8
XFILLER_13_62 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.mem_fle_3_in_1.LATCH_6_.latch data_in ltile_clb_0.mem_fle_3_in_1.LATCH_6_.latch/Q
+ _362_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_49_123 vgnd vpwr scs8hd_decap_6
XFILLER_1_196 vgnd vpwr scs8hd_decap_12
XFILLER_49_145 vpwr vgnd scs8hd_fill_2
XFILLER_45_362 vpwr vgnd scs8hd_fill_2
XFILLER_45_395 vpwr vgnd scs8hd_fill_2
XFILLER_54_80 vgnd vpwr scs8hd_decap_12
X_518_ _314_/A _517_/X _518_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_60_398 vgnd vpwr scs8hd_decap_3
XFILLER_60_376 vgnd vpwr scs8hd_decap_4
X_449_ _380_/X _226_/X _384_/X _346_/D _449_/X vgnd vpwr scs8hd_or4_4
XFILLER_20_218 vpwr vgnd scs8hd_fill_2
XFILLER_13_281 vgnd vpwr scs8hd_fill_1
XFILLER_9_285 vgnd vpwr scs8hd_decap_4
XFILLER_62_3 vgnd vpwr scs8hd_decap_12
XFILLER_9_296 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_3_in_2.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_3_in_2.INVTX1_13_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_68_454 vgnd vpwr scs8hd_decap_4
XFILLER_68_443 vgnd vpwr scs8hd_decap_4
Xltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_5_.scs8hd_inv_1
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_5_.latch/Q
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_ltile_clb_0.mem_fle_2_in_3.LATCH_1_.latch_SLEEPB _394_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_3_in_2.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_3_in_2.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_6_.scs8hd_inv_1/Y
+ _605_/Y ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_1_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_55_159 vpwr vgnd scs8hd_fill_2
XFILLER_70_129 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.mux_fle_2_in_1.INVTX1_7_.scs8hd_inv_1 left_width_0_height_0__pin_7_ ltile_clb_0.mux_fle_2_in_1.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_ltile_clb_0.mux_fle_1_in_0.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_1_in_0.INVTX1_9_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_24_513 vgnd vpwr scs8hd_decap_3
XFILLER_36_384 vpwr vgnd scs8hd_fill_2
XPHY_508 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_51_365 vgnd vpwr scs8hd_fill_1
XFILLER_51_343 vgnd vpwr scs8hd_decap_4
XPHY_519 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_50_27 vgnd vpwr scs8hd_decap_4
Xltile_clb_0.mux_fle_0_in_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_0_in_1.INVTX1_4_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_0_in_1.LATCH_0_.latch/Q ltile_clb_0.mux_fle_0_in_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_3_417 vpwr vgnd scs8hd_fill_2
XFILLER_3_428 vgnd vpwr scs8hd_decap_3
XANTENNA_ltile_clb_0.mux_fle_3_in_3.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_3_in_3.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_59_487 vgnd vpwr scs8hd_fill_1
XFILLER_74_457 vgnd vpwr scs8hd_fill_1
XFILLER_74_446 vgnd vpwr scs8hd_fill_1
XFILLER_74_468 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_16_.scs8hd_inv_1
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_16_.scs8hd_inv_1/A
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.INVTX1_1_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_inv_1
XFILLER_82_490 vgnd vpwr scs8hd_decap_6
Xltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_7_.TGATE_1_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_15_.scs8hd_inv_1/Y
+ _604_/Y ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_3_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_42_354 vgnd vpwr scs8hd_fill_1
X_303_ _302_/X _546_/A vgnd vpwr scs8hd_buf_1
X_234_ _304_/A _248_/A vgnd vpwr scs8hd_buf_1
XANTENNA__590__A _564_/A vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_1_in_1.INVTX1_14_.scs8hd_inv_1_A ltile_clb_0.mux_fle_1_in_1.INVTX1_14_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_0_in_0.INVTX1_0_.scs8hd_inv_1_A top_width_0_height_0__pin_0_
+ vgnd vpwr scs8hd_diode_2
XFILLER_40_93 vgnd vpwr scs8hd_decap_12
XFILLER_2_450 vgnd vpwr scs8hd_decap_8
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.mem_ble4_out_0.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_2_472 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mem_fle_0_in_0.LATCH_2_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_65_424 vgnd vpwr scs8hd_fill_1
XFILLER_65_457 vgnd vpwr scs8hd_decap_4
XFILLER_1_98 vgnd vpwr scs8hd_decap_12
XFILLER_33_321 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.mux_fle_3_in_2.INVTX1_2_.scs8hd_inv_1 bottom_width_0_height_0__pin_2_
+ ltile_clb_0.mux_fle_3_in_2.INVTX1_2_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XFILLER_60_184 vgnd vpwr scs8hd_decap_4
XANTENNA_ltile_clb_0.mem_fle_0_in_1.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mem_fle_3_in_2.LATCH_1_.latch_SLEEPB _355_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_3_.latch_SLEEPB
+ _569_/Y vgnd vpwr scs8hd_diode_2
XFILLER_29_39 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mux_fle_2_in_1.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_2_in_1.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_56_457 vgnd vpwr scs8hd_fill_1
XFILLER_56_424 vgnd vpwr scs8hd_decap_8
XANTENNA_ltile_clb_0.mux_fle_2_in_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_2_in_1.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_45_27 vgnd vpwr scs8hd_decap_12
XFILLER_24_310 vpwr vgnd scs8hd_fill_2
XANTENNA__394__B _387_/A vgnd vpwr scs8hd_diode_2
XPHY_305 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_316 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_332 vpwr vgnd scs8hd_fill_2
XFILLER_61_15 vgnd vpwr scs8hd_decap_12
XPHY_327 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_338 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_349 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_376 vgnd vpwr scs8hd_decap_8
XFILLER_24_387 vpwr vgnd scs8hd_fill_2
XFILLER_61_59 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_5_.scs8hd_inv_1_A
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_5_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_2_in_0.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_2_in_0.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mem_fle_0_in_3.LATCH_2_.latch_SLEEPB _490_/Y vgnd vpwr scs8hd_diode_2
XFILLER_59_240 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__569__B _554_/X vgnd vpwr scs8hd_diode_2
XFILLER_59_262 vgnd vpwr scs8hd_fill_1
XANTENNA_ltile_clb_0.mux_fle_3_in_3.mux_l1_in_2_.TGATE_3_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_3_in_3.INVTX1_11_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_59_295 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_2_.latch_D
+ data_in vgnd vpwr scs8hd_diode_2
XFILLER_62_405 vpwr vgnd scs8hd_fill_2
XFILLER_74_276 vgnd vpwr scs8hd_decap_3
XANTENNA__585__A _559_/A vgnd vpwr scs8hd_diode_2
XFILLER_15_310 vpwr vgnd scs8hd_fill_2
XFILLER_34_129 vgnd vpwr scs8hd_decap_12
XFILLER_42_151 vpwr vgnd scs8hd_fill_2
XFILLER_30_335 vgnd vpwr scs8hd_fill_1
XANTENNA_ltile_clb_0.mux_fle_1_in_1.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_1_in_1.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__479__B _479_/B vgnd vpwr scs8hd_diode_2
XFILLER_25_3 vgnd vpwr scs8hd_decap_12
XFILLER_65_221 vgnd vpwr scs8hd_decap_4
XFILLER_38_424 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.mux_fle_3_in_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_3_in_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ ltile_clb_0.mem_fle_3_in_1.LATCH_4_.latch/Q ltile_clb_0.mux_fle_3_in_1.INVTX1_14_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_38_457 vgnd vpwr scs8hd_fill_1
XFILLER_38_468 vgnd vpwr scs8hd_fill_1
XFILLER_80_202 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.mux_fle_3_in_3.INVTX1_6_.scs8hd_inv_1 bottom_width_0_height_0__pin_6_
+ ltile_clb_0.mux_fle_3_in_3.INVTX1_6_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XANTENNA__495__A _502_/B vgnd vpwr scs8hd_diode_2
XFILLER_61_460 vpwr vgnd scs8hd_fill_2
XFILLER_21_302 vgnd vpwr scs8hd_decap_3
XFILLER_21_313 vgnd vpwr scs8hd_fill_1
XFILLER_21_335 vpwr vgnd scs8hd_fill_2
XFILLER_21_346 vpwr vgnd scs8hd_fill_2
XFILLER_33_195 vpwr vgnd scs8hd_fill_2
XFILLER_21_357 vgnd vpwr scs8hd_decap_3
XANTENNA_ltile_clb_0.mux_fle_3_in_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_3_in_3.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XANTENNA__389__B _388_/B vgnd vpwr scs8hd_diode_2
XFILLER_56_210 vgnd vpwr scs8hd_decap_4
XFILLER_56_15 vgnd vpwr scs8hd_decap_12
XFILLER_29_457 vpwr vgnd scs8hd_fill_2
XFILLER_16_129 vgnd vpwr scs8hd_decap_12
XPHY_124 vgnd vpwr scs8hd_decap_3
XPHY_113 vgnd vpwr scs8hd_decap_3
XPHY_102 vgnd vpwr scs8hd_decap_3
XPHY_157 vgnd vpwr scs8hd_decap_3
XPHY_146 vgnd vpwr scs8hd_decap_3
XPHY_135 vgnd vpwr scs8hd_decap_3
XANTENNA_ltile_clb_0.mem_fle_1_in_2.LATCH_2_.latch_SLEEPB _457_/Y vgnd vpwr scs8hd_diode_2
XFILLER_12_379 vgnd vpwr scs8hd_fill_1
XFILLER_8_328 vgnd vpwr scs8hd_decap_8
XPHY_168 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_179 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_4_.TGATE_1_.scs8hd_ebufn_2_TEB
+ _604_/Y vgnd vpwr scs8hd_diode_2
XFILLER_21_51 vgnd vpwr scs8hd_decap_8
XFILLER_21_62 vgnd vpwr scs8hd_decap_12
XANTENNA__299__B address[1] vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mem_fle_0_in_0.LATCH_2_.latch data_in ltile_clb_0.mem_fle_0_in_0.LATCH_2_.latch/Q
+ _523_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_ltile_clb_0.mux_fle_2_in_3.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_2_in_3.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_62_202 vgnd vpwr scs8hd_decap_8
XFILLER_35_416 vgnd vpwr scs8hd_decap_4
XPHY_4 vgnd vpwr scs8hd_decap_3
XANTENNA_ltile_clb_0.mux_fle_2_in_3.mux_l1_in_3_.TGATE_2_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_2_in_3.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mem_fle_1_in_0.LATCH_1_.latch data_in ltile_clb_0.mem_fle_1_in_0.LATCH_1_.latch/Q
+ _480_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_15_184 vpwr vgnd scs8hd_fill_2
XPHY_680 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_62_80 vgnd vpwr scs8hd_decap_12
XFILLER_30_154 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mux_fle_3_in_0.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_3_in_0.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XPHY_691 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_30_176 vgnd vpwr scs8hd_fill_1
XANTENNA_ltile_clb_0.mux_fle_0_in_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_0_in_1.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_7_86 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mem_fle_2_in_0.LATCH_0_.latch data_in ltile_clb_0.mem_fle_2_in_0.LATCH_0_.latch/Q
+ _437_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_ltile_clb_0.mux_fle_3_in_0.INVTX1_12_.scs8hd_inv_1_A top_width_0_height_0__pin_12_
+ vgnd vpwr scs8hd_diode_2
XFILLER_53_202 vgnd vpwr scs8hd_decap_4
XFILLER_26_427 vpwr vgnd scs8hd_fill_2
XFILLER_26_438 vgnd vpwr scs8hd_decap_3
XFILLER_26_449 vgnd vpwr scs8hd_decap_8
XFILLER_21_110 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mem_fle_0_in_3.LATCH_6_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_34_493 vgnd vpwr scs8hd_decap_12
XFILLER_21_165 vgnd vpwr scs8hd_fill_1
XFILLER_21_176 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ _623_/Y ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_ltile_clb_0.mux_fle_1_in_0.INVTX1_6_.scs8hd_inv_1_A bottom_width_0_height_0__pin_6_
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mem_fle_2_in_1.LATCH_2_.latch_SLEEPB _422_/Y vgnd vpwr scs8hd_diode_2
Xltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_16_.scs8hd_inv_1
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_16_.scs8hd_inv_1/A
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.INVTX1_1_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_inv_1
X_620_ _620_/A _620_/Y vgnd vpwr scs8hd_inv_8
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.INVTX1_0_.scs8hd_inv_1_A
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.INVTX1_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_17_405 vgnd vpwr scs8hd_decap_3
X_551_ _603_/A _548_/X _551_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_29_276 vpwr vgnd scs8hd_fill_2
XFILLER_44_213 vgnd vpwr scs8hd_fill_1
X_482_ _380_/X _427_/B _228_/X _526_/D _482_/X vgnd vpwr scs8hd_or4_4
XFILLER_25_471 vpwr vgnd scs8hd_fill_2
XFILLER_12_154 vgnd vpwr scs8hd_decap_12
XANTENNA__582__B _585_/B vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mem_fle_0_in_2.LATCH_5_.latch data_in ltile_clb_0.mem_fle_0_in_2.LATCH_5_.latch/Q
+ _498_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_8_.latch_SLEEPB
+ _277_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mem_fle_1_in_1.LATCH_6_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_4_364 vgnd vpwr scs8hd_decap_6
XFILLER_79_110 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.mux_fle_2_in_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_2_in_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ ltile_clb_0.mem_fle_2_in_2.LATCH_4_.latch/Q ltile_clb_0.mux_fle_2_in_2.INVTX1_14_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
Xltile_clb_0.mem_fle_1_in_2.LATCH_4_.latch data_in ltile_clb_0.mem_fle_1_in_2.LATCH_4_.latch/Q
+ _455_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_75_393 vpwr vgnd scs8hd_fill_2
XFILLER_35_224 vpwr vgnd scs8hd_fill_2
XFILLER_35_235 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mem_fle_1_in_2.LATCH_4_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_23_419 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_2_in_3.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_2_in_3.INVTX1_13_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_3_.TGATE_1_.scs8hd_ebufn_2_TEB
+ _622_/Y vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mem_fle_2_in_2.LATCH_3_.latch data_in ltile_clb_0.mem_fle_2_in_2.LATCH_3_.latch/Q
+ _403_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_ltile_clb_0.mux_fle_2_in_1.INVTX1_3_.scs8hd_inv_1_A left_width_0_height_0__pin_3_
+ vgnd vpwr scs8hd_diode_2
XANTENNA__492__B _492_/B vgnd vpwr scs8hd_diode_2
XFILLER_31_463 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_1_in_2.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_1_in_2.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_15_.latch
+ data_in ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_15_.latch/Q
+ _530_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
Xltile_clb_0.mem_fle_3_in_2.LATCH_2_.latch data_in ltile_clb_0.mem_fle_3_in_2.LATCH_2_.latch/Q
+ _354_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_ltile_clb_0.mem_fle_1_in_3.LATCH_2_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_0_in_1.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_0_in_1.INVTX1_9_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_0_in_0.INVTX1_2_.scs8hd_inv_1 bottom_width_0_height_0__pin_2_
+ ltile_clb_0.mux_fle_0_in_0.INVTX1_2_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XFILLER_58_327 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_37_39 vgnd vpwr scs8hd_decap_12
XFILLER_66_360 vgnd vpwr scs8hd_decap_8
XFILLER_81_330 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_3_.scs8hd_inv_1_A
+ ltile_clb_0.mux_fle_0_in_3.INVTX1_14_.scs8hd_inv_1/Y vgnd vpwr scs8hd_diode_2
XFILLER_53_27 vgnd vpwr scs8hd_decap_12
XFILLER_34_290 vgnd vpwr scs8hd_fill_1
XANTENNA_ltile_clb_0.mem_fle_3_in_0.LATCH_2_.latch_SLEEPB _377_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mem_fle_2_in_0.LATCH_4_.latch_D data_in vgnd vpwr scs8hd_diode_2
Xltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_3_.scs8hd_inv_1
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_3_.latch/Q
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_ltile_clb_0.mux_fle_0_in_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_0_in_0.LATCH_4_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_1_301 vpwr vgnd scs8hd_fill_2
XFILLER_78_68 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mux_fle_3_in_2.INVTX1_0_.scs8hd_inv_1_A top_width_0_height_0__pin_0_
+ vgnd vpwr scs8hd_diode_2
XFILLER_1_345 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_7_.TGATE_0_.scs8hd_ebufn_2_TEB
+ _613_/Y vgnd vpwr scs8hd_diode_2
XFILLER_1_378 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_8_.latch_D
+ data_in vgnd vpwr scs8hd_diode_2
XANTENNA__577__B _575_/B vgnd vpwr scs8hd_diode_2
XFILLER_76_168 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mem_fle_2_in_1.LATCH_2_.latch_D data_in vgnd vpwr scs8hd_diode_2
X_603_ _603_/A _600_/X _603_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_57_393 vpwr vgnd scs8hd_fill_2
XANTENNA__296__C address[3] vgnd vpwr scs8hd_diode_2
X_534_ _261_/X _529_/X _534_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA__593__A _541_/A vgnd vpwr scs8hd_diode_2
X_465_ _432_/A _462_/X _465_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA_ltile_clb_0.mux_fle_3_in_0.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_3_in_0.LATCH_7_.latch/Q
+ vgnd vpwr scs8hd_diode_2
X_396_ _380_/X _427_/B _384_/X _346_/D _397_/A vgnd vpwr scs8hd_or4_4
XFILLER_40_271 vgnd vpwr scs8hd_decap_4
XFILLER_40_293 vgnd vpwr scs8hd_fill_1
XANTENNA_ltile_clb_0.mem_fle_2_in_2.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mem_fle_0_in_1.LATCH_3_.latch_SLEEPB _511_/Y vgnd vpwr scs8hd_diode_2
XFILLER_4_32 vgnd vpwr scs8hd_decap_12
XFILLER_67_157 vpwr vgnd scs8hd_fill_2
XANTENNA__487__B _484_/X vgnd vpwr scs8hd_diode_2
XFILLER_67_179 vpwr vgnd scs8hd_fill_2
XFILLER_36_511 vgnd vpwr scs8hd_decap_4
XFILLER_82_149 vgnd vpwr scs8hd_decap_6
Xltile_clb_0.mux_fle_2_in_0.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_2_in_0.INVTX1_10_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_2_in_0.LATCH_2_.latch/Q ltile_clb_0.mux_fle_2_in_0.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_51_514 vpwr vgnd scs8hd_fill_2
XFILLER_31_260 vgnd vpwr scs8hd_decap_6
XANTENNA_ltile_clb_0.mux_fle_2_in_3.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_2_in_3.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_0_in_1.INVTX1_6_.scs8hd_inv_1 bottom_width_0_height_0__pin_6_
+ ltile_clb_0.mux_fle_0_in_1.INVTX1_6_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XANTENNA_ltile_clb_0.mux_fle_1_in_2.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_1_in_2.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_48_27 vgnd vpwr scs8hd_decap_4
XANTENNA_ltile_clb_0.mem_fle_3_in_0.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_58_146 vgnd vpwr scs8hd_decap_3
XFILLER_73_149 vpwr vgnd scs8hd_fill_2
XFILLER_64_15 vgnd vpwr scs8hd_decap_12
XFILLER_39_382 vgnd vpwr scs8hd_decap_4
XANTENNA_ltile_clb_0.mux_fle_2_in_2.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_2_in_2.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_81_171 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.mux_fle_3_in_3.mux_l1_in_2_.TGATE_3_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_3_in_3.INVTX1_11_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_3_in_3.LATCH_3_.latch/Q ltile_clb_0.mux_fle_3_in_3.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_10_411 vgnd vpwr scs8hd_decap_4
X_250_ _250_/A _250_/X vgnd vpwr scs8hd_buf_1
XFILLER_22_293 vgnd vpwr scs8hd_fill_1
XFILLER_13_74 vgnd vpwr scs8hd_decap_12
XFILLER_6_426 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.mux_fle_1_in_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_1_in_3.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ ltile_clb_0.mem_fle_1_in_3.LATCH_4_.latch/Q ltile_clb_0.mux_fle_1_in_3.INVTX1_14_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_10_488 vgnd vpwr scs8hd_fill_1
XFILLER_77_400 vgnd vpwr scs8hd_decap_6
XANTENNA__588__A _580_/X vgnd vpwr scs8hd_diode_2
XFILLER_64_105 vgnd vpwr scs8hd_decap_12
XFILLER_37_319 vpwr vgnd scs8hd_fill_2
XFILLER_49_179 vpwr vgnd scs8hd_fill_2
XFILLER_38_93 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mux_fle_0_in_2.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_0_in_2.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_4_.latch_D
+ data_in vgnd vpwr scs8hd_diode_2
X_517_ _516_/X _517_/X vgnd vpwr scs8hd_buf_1
XANTENNA_ltile_clb_0.mem_fle_1_in_0.LATCH_3_.latch_SLEEPB _478_/Y vgnd vpwr scs8hd_diode_2
X_448_ _437_/A _447_/B _448_/Y vgnd vpwr scs8hd_nor2_4
X_379_ _379_/A _379_/B _379_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_9_242 vpwr vgnd scs8hd_fill_2
XFILLER_70_80 vgnd vpwr scs8hd_decap_12
XFILLER_9_264 vgnd vpwr scs8hd_decap_6
XANTENNA_ltile_clb_0.mux_fle_3_in_0.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_3_in_0.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_55_3 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.buf4_1_.scs8hd_buf_1
+ ltile_clb_0.mux_fle_0_in_1.INVTX1_14_.scs8hd_inv_1/Y _630_/A vgnd vpwr scs8hd_buf_1
Xltile_clb_0.mux_fle_0_in_1.INVTX1_11_.scs8hd_inv_1 left_width_0_height_0__pin_11_
+ ltile_clb_0.mux_fle_0_in_1.INVTX1_11_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
Xltile_clb_0.mux_fle_1_in_2.INVTX1_1_.scs8hd_inv_1 right_width_0_height_0__pin_1_
+ ltile_clb_0.mux_fle_1_in_2.INVTX1_1_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
Xltile_clb_0.mux_fle_3_in_1.INVTX1_10_.scs8hd_inv_1 bottom_width_0_height_0__pin_10_
+ ltile_clb_0.mux_fle_3_in_1.INVTX1_10_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XANTENNA__498__A _328_/A vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.mem_ble4_out_0.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_51_322 vpwr vgnd scs8hd_fill_2
XPHY_509 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_51_388 vpwr vgnd scs8hd_fill_2
XFILLER_11_208 vpwr vgnd scs8hd_fill_2
XFILLER_51_399 vpwr vgnd scs8hd_fill_2
XFILLER_59_15 vgnd vpwr scs8hd_decap_12
XFILLER_59_59 vpwr vgnd scs8hd_fill_2
XFILLER_59_400 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_16_.scs8hd_inv_1
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_16_.scs8hd_inv_1/A
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.INVTX1_1_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_inv_1
Xltile_clb_0.mux_fle_0_in_2.INVTX1_13_.scs8hd_inv_1 right_width_0_height_0__pin_13_
+ ltile_clb_0.mux_fle_0_in_2.INVTX1_13_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XFILLER_19_319 vpwr vgnd scs8hd_fill_2
XFILLER_46_105 vgnd vpwr scs8hd_decap_12
XFILLER_74_425 vgnd vpwr scs8hd_decap_4
Xltile_clb_0.mux_fle_3_in_2.INVTX1_12_.scs8hd_inv_1 top_width_0_height_0__pin_12_
+ ltile_clb_0.mux_fle_3_in_2.INVTX1_12_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XANTENNA_ltile_clb_0.mux_fle_1_in_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_1_in_1.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
X_302_ _278_/X _342_/A _302_/X vgnd vpwr scs8hd_or2_4
X_233_ _232_/X _304_/A vgnd vpwr scs8hd_buf_1
XANTENNA__590__B _588_/X vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_3_in_1.INVTX1_9_.scs8hd_inv_1_A right_width_0_height_0__pin_9_
+ vgnd vpwr scs8hd_diode_2
XFILLER_10_285 vpwr vgnd scs8hd_fill_2
XFILLER_6_223 vgnd vpwr scs8hd_decap_4
XFILLER_69_219 vpwr vgnd scs8hd_fill_2
XFILLER_2_484 vgnd vpwr scs8hd_decap_12
XFILLER_77_274 vgnd vpwr scs8hd_decap_3
XFILLER_65_414 vgnd vpwr scs8hd_decap_4
XANTENNA_ltile_clb_0.mux_fle_1_in_0.mux_l1_in_2_.TGATE_3_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_1_in_0.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_1_in_1.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_1_in_1.INVTX1_10_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_1_in_1.LATCH_2_.latch/Q ltile_clb_0.mux_fle_1_in_1.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
Xltile_clb_0.mux_fle_3_in_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_3_in_1.INVTX1_5_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_3_in_1.LATCH_1_.latch/Q ltile_clb_0.mux_fle_3_in_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_18_352 vpwr vgnd scs8hd_fill_2
XFILLER_18_363 vpwr vgnd scs8hd_fill_2
XFILLER_60_174 vgnd vpwr scs8hd_decap_8
Xltile_clb_0.mux_fle_3_in_3.INVTX1_14_.scs8hd_inv_1 ltile_clb_0.mux_fle_3_in_3.INVTX1_14_.scs8hd_inv_1/A
+ ltile_clb_0.mux_fle_3_in_3.INVTX1_14_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XANTENNA_ltile_clb_0.mux_fle_1_in_3.INVTX1_12_.scs8hd_inv_1_A top_width_0_height_0__pin_12_
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_1_in_3.INVTX1_5_.scs8hd_inv_1 right_width_0_height_0__pin_5_
+ ltile_clb_0.mux_fle_1_in_3.INVTX1_5_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_0_.latch_D
+ data_in vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_2_in_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_2_in_0.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l4_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
+ _618_/Y vgnd vpwr scs8hd_diode_2
Xltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_5_.TGATE_0_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_10_.scs8hd_inv_1/Y
+ _613_/Y ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_2_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_28_105 vgnd vpwr scs8hd_decap_12
XFILLER_71_406 vpwr vgnd scs8hd_fill_2
XFILLER_56_469 vgnd vpwr scs8hd_fill_1
XFILLER_71_428 vgnd vpwr scs8hd_decap_3
XFILLER_45_39 vgnd vpwr scs8hd_decap_12
XPHY_306 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_322 vgnd vpwr scs8hd_decap_3
XPHY_317 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_328 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_339 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_355 vgnd vpwr scs8hd_fill_1
XFILLER_61_27 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.mem_ble4_out_0.LATCH_2_.latch_SLEEPB
+ _549_/Y vgnd vpwr scs8hd_diode_2
XFILLER_51_174 vgnd vpwr scs8hd_decap_3
XANTENNA_ltile_clb_0.mem_fle_3_in_2.LATCH_6_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_59_252 vpwr vgnd scs8hd_fill_2
XFILLER_47_414 vpwr vgnd scs8hd_fill_2
XFILLER_59_274 vgnd vpwr scs8hd_decap_8
XFILLER_19_51 vgnd vpwr scs8hd_decap_8
XFILLER_19_62 vgnd vpwr scs8hd_decap_12
XFILLER_47_447 vpwr vgnd scs8hd_fill_2
XFILLER_47_458 vpwr vgnd scs8hd_fill_2
XFILLER_74_288 vgnd vpwr scs8hd_decap_8
XFILLER_62_428 vgnd vpwr scs8hd_fill_1
XANTENNA__585__B _585_/B vgnd vpwr scs8hd_diode_2
XFILLER_15_333 vpwr vgnd scs8hd_fill_2
XFILLER_27_193 vgnd vpwr scs8hd_decap_4
XFILLER_70_450 vgnd vpwr scs8hd_decap_8
XFILLER_42_141 vgnd vpwr scs8hd_decap_8
XPHY_840 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_ltile_clb_0.mem_fle_3_in_3.LATCH_4_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_11_.scs8hd_inv_1_A
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_11_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_2_in_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_2_in_1.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_18_3 vgnd vpwr scs8hd_decap_12
XFILLER_53_428 vgnd vpwr scs8hd_decap_4
XFILLER_61_494 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_13_.latch
+ data_in ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_13_.latch/Q
+ _584_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
Xltile_clb_0.mem_fle_0_in_3.LATCH_1_.latch data_in ltile_clb_0.mem_fle_0_in_3.LATCH_1_.latch/Q
+ _491_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_ltile_clb_0.mux_fle_2_in_0.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_2_in_0.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_3_.scs8hd_inv_1/Y
+ _620_/Y ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_0_218 vgnd vpwr scs8hd_decap_4
XANTENNA_ltile_clb_0.mux_fle_2_in_0.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_2_in_0.INVTX1_9_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_0_in_1.INVTX1_7_.scs8hd_inv_1_A left_width_0_height_0__pin_7_
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mem_fle_1_in_3.LATCH_0_.latch data_in ltile_clb_0.mem_fle_1_in_3.LATCH_0_.latch/Q
+ _448_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_56_27 vgnd vpwr scs8hd_decap_4
Xltile_clb_0.mux_fle_3_in_0.INVTX1_2_.scs8hd_inv_1 bottom_width_0_height_0__pin_2_
+ ltile_clb_0.mux_fle_3_in_0.INVTX1_2_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XFILLER_72_15 vgnd vpwr scs8hd_decap_12
XFILLER_71_236 vpwr vgnd scs8hd_fill_2
XFILLER_71_269 vpwr vgnd scs8hd_fill_2
XPHY_125 vgnd vpwr scs8hd_decap_3
XPHY_114 vgnd vpwr scs8hd_decap_3
XFILLER_52_450 vgnd vpwr scs8hd_decap_4
XPHY_103 vgnd vpwr scs8hd_decap_3
XFILLER_24_141 vgnd vpwr scs8hd_decap_12
XPHY_158 vgnd vpwr scs8hd_decap_3
XPHY_147 vgnd vpwr scs8hd_decap_3
XPHY_136 vgnd vpwr scs8hd_decap_3
XFILLER_52_494 vgnd vpwr scs8hd_fill_1
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_0_.TGATE_0_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_3_.scs8hd_inv_1
+ ltile_clb_0.mux_fle_2_in_3.INVTX1_14_.scs8hd_inv_1/Y _619_/A vgnd vpwr scs8hd_inv_1
XFILLER_8_318 vgnd vpwr scs8hd_fill_1
XPHY_169 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_21_74 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mux_fle_3_in_2.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_3_in_2.LATCH_6_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_79_325 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
+ _614_/Y vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_0_in_2.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_0_in_2.INVTX1_10_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_0_in_2.LATCH_2_.latch/Q ltile_clb_0.mux_fle_0_in_2.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
Xltile_clb_0.mux_fle_2_in_2.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_2_in_2.INVTX1_5_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_2_in_2.LATCH_1_.latch/Q ltile_clb_0.mux_fle_2_in_2.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA__299__C address[3] vgnd vpwr scs8hd_diode_2
XANTENNA__596__A _544_/A vgnd vpwr scs8hd_diode_2
XFILLER_47_255 vpwr vgnd scs8hd_fill_2
XFILLER_62_247 vpwr vgnd scs8hd_fill_2
XFILLER_28_491 vpwr vgnd scs8hd_fill_2
XFILLER_35_439 vpwr vgnd scs8hd_fill_2
XFILLER_46_93 vgnd vpwr scs8hd_decap_12
XFILLER_62_258 vgnd vpwr scs8hd_decap_8
XPHY_5 vgnd vpwr scs8hd_decap_3
XFILLER_15_163 vgnd vpwr scs8hd_fill_1
XFILLER_43_472 vpwr vgnd scs8hd_fill_2
XFILLER_43_483 vpwr vgnd scs8hd_fill_2
XPHY_670 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_ltile_clb_0.mux_fle_1_in_2.INVTX1_4_.scs8hd_inv_1_A top_width_0_height_0__pin_4_
+ vgnd vpwr scs8hd_diode_2
XPHY_692 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_681 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_30_188 vpwr vgnd scs8hd_fill_2
XFILLER_7_362 vpwr vgnd scs8hd_fill_2
XFILLER_7_98 vgnd vpwr scs8hd_decap_12
XFILLER_38_244 vpwr vgnd scs8hd_fill_2
XFILLER_81_501 vgnd vpwr scs8hd_decap_12
XFILLER_53_236 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_0_in_3.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_0_in_3.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.buf4_0_.scs8hd_buf_1_A
+ ltile_clb_0.mux_fle_0_in_0.INVTX1_14_.scs8hd_inv_1/Y vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_5_.TGATE_0_.scs8hd_ebufn_2_TEB
+ _605_/Y vgnd vpwr scs8hd_diode_2
Xltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_16_.scs8hd_inv_1
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_16_.scs8hd_inv_1/A
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.INVTX1_1_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_inv_1
XANTENNA_ltile_clb_0.mux_fle_3_in_1.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_3_in_1.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_67_15 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mux_fle_3_in_2.INVTX1_10_.scs8hd_inv_1_A bottom_width_0_height_0__pin_10_
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_3_in_1.INVTX1_6_.scs8hd_inv_1 bottom_width_0_height_0__pin_6_
+ ltile_clb_0.mux_fle_3_in_1.INVTX1_6_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XANTENNA_ltile_clb_0.mux_fle_2_in_3.INVTX1_1_.scs8hd_inv_1_A right_width_0_height_0__pin_1_
+ vgnd vpwr scs8hd_diode_2
XFILLER_67_59 vpwr vgnd scs8hd_fill_2
X_550_ _270_/B _548_/X _550_/Y vgnd vpwr scs8hd_nor2_4
X_481_ _437_/A _481_/B _481_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_25_461 vgnd vpwr scs8hd_fill_1
XFILLER_12_166 vgnd vpwr scs8hd_decap_12
XFILLER_12_188 vgnd vpwr scs8hd_decap_3
XFILLER_40_497 vgnd vpwr scs8hd_decap_12
XFILLER_4_321 vpwr vgnd scs8hd_fill_2
XFILLER_4_376 vgnd vpwr scs8hd_decap_4
XFILLER_4_398 vgnd vpwr scs8hd_decap_3
XFILLER_67_339 vpwr vgnd scs8hd_fill_2
XFILLER_75_383 vgnd vpwr scs8hd_fill_1
XANTENNA_ltile_clb_0.mux_fle_2_in_1.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_2_in_1.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_23_409 vpwr vgnd scs8hd_fill_2
XFILLER_50_206 vpwr vgnd scs8hd_fill_2
XFILLER_43_291 vgnd vpwr scs8hd_fill_1
Xltile_clb_0.mux_fle_0_in_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_0_in_0.INVTX1_4_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_0_in_0.LATCH_0_.latch/Q ltile_clb_0.mux_fle_0_in_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
+ _632_/Y vgnd vpwr scs8hd_diode_2
XFILLER_81_342 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.buf4_2_.scs8hd_buf_1_A
+ ltile_clb_0.mux_fle_2_in_2.INVTX1_14_.scs8hd_inv_1/Y vgnd vpwr scs8hd_diode_2
XFILLER_81_386 vgnd vpwr scs8hd_decap_12
XFILLER_53_39 vgnd vpwr scs8hd_decap_12
XFILLER_41_217 vgnd vpwr scs8hd_fill_1
XFILLER_22_431 vgnd vpwr scs8hd_decap_4
XFILLER_22_442 vgnd vpwr scs8hd_decap_4
XFILLER_22_453 vgnd vpwr scs8hd_decap_3
Xltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_2_.TGATE_0_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_2_.TGATE_0_.scs8hd_ebufn_2/A
+ _631_/Y ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_1_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_ltile_clb_0.mux_fle_1_in_3.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_1_in_3.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_1_in_3.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_1_in_3.INVTX1_5_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_1_in_3.LATCH_1_.latch/Q ltile_clb_0.mux_fle_1_in_3.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
Xltile_clb_0.mux_fle_3_in_3.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_3_in_3.INVTX1_0_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_3_in_3.LATCH_0_.latch/Q ltile_clb_0.mux_fle_3_in_3.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
X_602_ _270_/B _600_/X _602_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_72_320 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.INVTX1_0_.scs8hd_inv_1/Y
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.mem_ble4_out_0.LATCH_0_.latch/Q
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_17_236 vgnd vpwr scs8hd_fill_1
XANTENNA__296__D _258_/X vgnd vpwr scs8hd_diode_2
XFILLER_27_51 vgnd vpwr scs8hd_decap_8
XFILLER_27_62 vgnd vpwr scs8hd_decap_12
X_533_ _559_/A _529_/X _533_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_17_258 vpwr vgnd scs8hd_fill_2
XFILLER_72_386 vgnd vpwr scs8hd_decap_6
XANTENNA__593__B _588_/X vgnd vpwr scs8hd_diode_2
X_464_ _431_/A _462_/X _464_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_13_431 vpwr vgnd scs8hd_fill_2
XFILLER_25_291 vgnd vpwr scs8hd_decap_4
X_395_ _379_/A _387_/A _395_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_9_435 vpwr vgnd scs8hd_fill_2
XFILLER_13_475 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_1_in_2.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_1_in_2.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_40_250 vgnd vpwr scs8hd_decap_6
XANTENNA_ltile_clb_0.mux_fle_3_in_3.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_3_in_3.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_4_44 vgnd vpwr scs8hd_decap_12
XFILLER_68_80 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_12_.latch_D
+ data_in vgnd vpwr scs8hd_diode_2
XFILLER_82_106 vgnd vpwr scs8hd_decap_12
XFILLER_63_331 vpwr vgnd scs8hd_fill_2
XFILLER_75_191 vpwr vgnd scs8hd_fill_2
XFILLER_63_375 vpwr vgnd scs8hd_fill_2
XFILLER_16_291 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_1_in_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_1_in_1.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_0_.TGATE_0_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_2_in_1.INVTX1_14_.scs8hd_inv_1_A ltile_clb_0.mux_fle_2_in_1.INVTX1_14_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.mem_ble4_out_0.LATCH_2_.latch_SLEEPB
+ _575_/Y vgnd vpwr scs8hd_diode_2
XFILLER_58_158 vgnd vpwr scs8hd_decap_4
XFILLER_46_309 vgnd vpwr scs8hd_decap_8
XFILLER_64_27 vgnd vpwr scs8hd_decap_4
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.INVTX1_1_.scs8hd_inv_1_A
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.INVTX1_1_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_42_515 vgnd vpwr scs8hd_fill_1
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.mem_ble4_out_0.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_80_15 vgnd vpwr scs8hd_decap_12
XFILLER_10_467 vpwr vgnd scs8hd_fill_2
XFILLER_13_86 vgnd vpwr scs8hd_decap_12
XFILLER_1_110 vgnd vpwr scs8hd_decap_12
XFILLER_77_423 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
+ _628_/Y vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_3_in_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_3_in_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ ltile_clb_0.mem_fle_3_in_0.LATCH_4_.latch/Q ltile_clb_0.mux_fle_3_in_0.INVTX1_14_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_77_489 vgnd vpwr scs8hd_decap_12
XFILLER_64_117 vgnd vpwr scs8hd_decap_12
X_516_ _516_/A _516_/X vgnd vpwr scs8hd_buf_1
XFILLER_60_345 vgnd vpwr scs8hd_fill_1
XFILLER_54_93 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_0_.scs8hd_inv_1_A
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_60_389 vpwr vgnd scs8hd_fill_2
X_447_ _436_/A _447_/B _447_/Y vgnd vpwr scs8hd_nor2_4
X_378_ _394_/A _379_/B _378_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_9_232 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_0_in_1.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_0_in_1.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_48_3 vgnd vpwr scs8hd_decap_12
XFILLER_68_401 vgnd vpwr scs8hd_decap_8
XANTENNA__498__B _495_/X vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_3_in_3.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_3_in_3.INVTX1_13_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_3_in_3.INVTX1_7_.scs8hd_inv_1_A left_width_0_height_0__pin_7_
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_2_in_2.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_2_in_2.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_51_378 vgnd vpwr scs8hd_fill_1
XANTENNA_ltile_clb_0.mux_fle_1_in_1.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_1_in_1.INVTX1_9_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_59_27 vgnd vpwr scs8hd_decap_12
XFILLER_59_445 vpwr vgnd scs8hd_fill_2
XFILLER_59_423 vpwr vgnd scs8hd_fill_2
XFILLER_75_15 vgnd vpwr scs8hd_decap_12
XFILLER_75_59 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_6_.scs8hd_inv_1
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_6_.latch/Q
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_46_117 vgnd vpwr scs8hd_decap_12
XFILLER_27_331 vpwr vgnd scs8hd_fill_2
XFILLER_27_364 vpwr vgnd scs8hd_fill_2
XFILLER_27_397 vgnd vpwr scs8hd_fill_1
X_301_ _304_/A _545_/A _301_/Y vgnd vpwr scs8hd_nor2_4
X_232_ address[4] _231_/X _232_/X vgnd vpwr scs8hd_or2_4
XFILLER_10_253 vgnd vpwr scs8hd_decap_4
XFILLER_6_202 vgnd vpwr scs8hd_decap_12
XANTENNA__599__A _599_/A vgnd vpwr scs8hd_diode_2
XFILLER_77_231 vgnd vpwr scs8hd_decap_12
XFILLER_2_496 vgnd vpwr scs8hd_decap_12
XFILLER_77_253 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_0_in_0.INVTX1_13_.scs8hd_inv_1_A right_width_0_height_0__pin_13_
+ vgnd vpwr scs8hd_diode_2
XFILLER_33_301 vpwr vgnd scs8hd_fill_2
XFILLER_33_356 vpwr vgnd scs8hd_fill_2
XFILLER_33_378 vpwr vgnd scs8hd_fill_2
XANTENNA__302__A _278_/X vgnd vpwr scs8hd_diode_2
XFILLER_68_286 vpwr vgnd scs8hd_fill_2
XFILLER_28_117 vgnd vpwr scs8hd_decap_12
XFILLER_56_459 vgnd vpwr scs8hd_decap_3
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_5_.TGATE_0_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_10_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_3_.TGATE_1_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_3_.TGATE_1_.scs8hd_ebufn_2/A
+ _606_/Y ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_1_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_36_161 vpwr vgnd scs8hd_fill_2
XPHY_307 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_ltile_clb_0.mux_fle_1_in_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_1_in_1.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XPHY_318 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_329 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_51_131 vpwr vgnd scs8hd_fill_2
XFILLER_51_142 vpwr vgnd scs8hd_fill_2
XFILLER_51_153 vgnd vpwr scs8hd_fill_1
XANTENNA_ltile_clb_0.mux_fle_2_in_2.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_2_in_2.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_61_39 vgnd vpwr scs8hd_decap_12
XFILLER_51_197 vgnd vpwr scs8hd_decap_4
Xltile_clb_0.mux_fle_1_in_0.INVTX1_1_.scs8hd_inv_1 right_width_0_height_0__pin_1_
+ ltile_clb_0.mux_fle_1_in_0.INVTX1_1_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XFILLER_10_32 vgnd vpwr scs8hd_decap_12
XFILLER_3_249 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.mux_fle_2_in_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_2_in_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ ltile_clb_0.mem_fle_2_in_1.LATCH_4_.latch/Q ltile_clb_0.mux_fle_2_in_1.INVTX1_14_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_59_231 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_1_in_0.mux_l1_in_3_.TGATE_2_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_1_in_0.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_47_404 vgnd vpwr scs8hd_fill_1
XFILLER_74_212 vpwr vgnd scs8hd_fill_2
XFILLER_59_286 vgnd vpwr scs8hd_decap_4
XFILLER_19_74 vgnd vpwr scs8hd_decap_12
XFILLER_47_426 vgnd vpwr scs8hd_fill_1
XFILLER_74_267 vgnd vpwr scs8hd_decap_8
XFILLER_15_301 vpwr vgnd scs8hd_fill_2
XFILLER_35_51 vgnd vpwr scs8hd_decap_8
XFILLER_70_462 vgnd vpwr scs8hd_decap_12
XFILLER_15_356 vgnd vpwr scs8hd_decap_4
XFILLER_35_62 vgnd vpwr scs8hd_decap_12
XPHY_841 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_830 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_42_186 vgnd vpwr scs8hd_fill_1
XANTENNA_ltile_clb_0.mux_fle_0_in_3.INVTX1_5_.scs8hd_inv_1_A right_width_0_height_0__pin_5_
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_1_in_0.INVTX1_1_.scs8hd_inv_1_A right_width_0_height_0__pin_1_
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_1_in_2.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_1_in_2.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_2_in_2.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_2_in_2.LATCH_7_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_76_80 vgnd vpwr scs8hd_decap_12
XFILLER_65_256 vpwr vgnd scs8hd_fill_2
XFILLER_80_215 vgnd vpwr scs8hd_decap_12
XFILLER_53_418 vpwr vgnd scs8hd_fill_2
XFILLER_46_470 vpwr vgnd scs8hd_fill_2
XFILLER_80_259 vgnd vpwr scs8hd_decap_3
XFILLER_33_175 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_7_.TGATE_0_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_14_.scs8hd_inv_1/Y
+ _621_/Y ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_7_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_4_.latch_SLEEPB
+ _594_/Y vgnd vpwr scs8hd_diode_2
XFILLER_56_289 vgnd vpwr scs8hd_decap_8
XFILLER_56_267 vgnd vpwr scs8hd_decap_6
XFILLER_44_407 vgnd vpwr scs8hd_decap_4
XFILLER_37_492 vpwr vgnd scs8hd_fill_2
XFILLER_72_27 vgnd vpwr scs8hd_decap_4
XPHY_115 vgnd vpwr scs8hd_decap_3
XFILLER_52_462 vgnd vpwr scs8hd_decap_8
XPHY_104 vgnd vpwr scs8hd_decap_3
Xltile_clb_0.mux_fle_1_in_1.INVTX1_5_.scs8hd_inv_1 right_width_0_height_0__pin_5_
+ ltile_clb_0.mux_fle_1_in_1.INVTX1_5_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XPHY_148 vgnd vpwr scs8hd_decap_3
XPHY_137 vgnd vpwr scs8hd_decap_3
XPHY_126 vgnd vpwr scs8hd_decap_3
XFILLER_12_315 vgnd vpwr scs8hd_decap_4
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_7_.TGATE_1_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_15_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_13_.scs8hd_inv_1_A
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_13_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XPHY_159 vgnd vpwr scs8hd_decap_3
XFILLER_12_337 vgnd vpwr scs8hd_decap_4
XFILLER_20_392 vgnd vpwr scs8hd_decap_4
XFILLER_4_514 vpwr vgnd scs8hd_fill_2
XFILLER_21_86 vgnd vpwr scs8hd_decap_12
XFILLER_79_337 vgnd vpwr scs8hd_decap_4
XANTENNA__299__D _258_/X vgnd vpwr scs8hd_diode_2
XANTENNA__596__B _580_/X vgnd vpwr scs8hd_diode_2
XFILLER_47_234 vpwr vgnd scs8hd_fill_2
XFILLER_47_245 vgnd vpwr scs8hd_fill_1
XFILLER_62_215 vgnd vpwr scs8hd_decap_3
XFILLER_47_278 vpwr vgnd scs8hd_fill_2
XPHY_6 vgnd vpwr scs8hd_decap_3
XFILLER_43_451 vpwr vgnd scs8hd_fill_2
XFILLER_15_175 vpwr vgnd scs8hd_fill_2
XFILLER_70_292 vgnd vpwr scs8hd_decap_3
XPHY_671 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_660 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_15_197 vpwr vgnd scs8hd_fill_2
XPHY_693 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_682 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_62_93 vgnd vpwr scs8hd_decap_12
XFILLER_30_3 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mux_fle_0_in_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_0_in_2.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_78_370 vpwr vgnd scs8hd_fill_2
XFILLER_66_510 vgnd vpwr scs8hd_decap_6
XFILLER_38_223 vpwr vgnd scs8hd_fill_2
XFILLER_81_513 vgnd vpwr scs8hd_decap_3
XFILLER_53_226 vgnd vpwr scs8hd_decap_4
XFILLER_19_481 vgnd vpwr scs8hd_decap_4
XANTENNA_ltile_clb_0.mux_fle_3_in_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_3_in_0.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_3_in_2.mux_l1_in_2_.TGATE_3_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_3_in_2.INVTX1_11_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_3_in_2.LATCH_3_.latch/Q ltile_clb_0.mux_fle_3_in_2.mux_l1_in_2_.TGATE_3_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_61_281 vgnd vpwr scs8hd_decap_4
Xltile_clb_0.mux_fle_2_in_2.INVTX1_0_.scs8hd_inv_1 top_width_0_height_0__pin_0_ ltile_clb_0.mux_fle_2_in_2.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_21_123 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_7_.scs8hd_inv_1/Y
+ _628_/Y ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_1_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.mem_ble4_out_0.LATCH_2_.latch_SLEEPB
+ _601_/Y vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_1_in_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_1_in_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ ltile_clb_0.mem_fle_1_in_2.LATCH_4_.latch/Q ltile_clb_0.mux_fle_1_in_2.INVTX1_14_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB
+ _615_/Y vgnd vpwr scs8hd_diode_2
XFILLER_67_27 vgnd vpwr scs8hd_decap_12
XFILLER_76_329 vgnd vpwr scs8hd_decap_6
XFILLER_69_392 vgnd vpwr scs8hd_decap_6
Xltile_clb_0.mux_fle_1_in_2.INVTX1_9_.scs8hd_inv_1 right_width_0_height_0__pin_9_
+ ltile_clb_0.mux_fle_1_in_2.INVTX1_9_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
X_480_ _436_/A _481_/B _480_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_52_270 vpwr vgnd scs8hd_fill_2
XFILLER_25_484 vpwr vgnd scs8hd_fill_2
XFILLER_8_105 vgnd vpwr scs8hd_decap_12
XFILLER_4_311 vgnd vpwr scs8hd_decap_6
XFILLER_4_344 vgnd vpwr scs8hd_decap_3
XFILLER_79_123 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mux_fle_0_in_3.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_0_in_3.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__400__A _326_/A vgnd vpwr scs8hd_diode_2
XFILLER_75_362 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mem_fle_3_in_3.LATCH_3_.latch_SLEEPB _335_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_1_in_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_1_in_0.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_35_204 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_5_.TGATE_0_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_10_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_35_259 vpwr vgnd scs8hd_fill_2
XFILLER_16_473 vgnd vpwr scs8hd_decap_8
XFILLER_78_3 vgnd vpwr scs8hd_decap_12
XPHY_490 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_7_171 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mux_fle_0_in_2.mux_l1_in_2_.TGATE_3_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_0_in_2.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_2_.latch
+ data_in ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_2_.latch/Q
+ _298_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA__310__A _575_/A vgnd vpwr scs8hd_diode_2
XFILLER_26_215 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_0_in_2.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_0_in_2.INVTX1_9_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_81_354 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.mux_fle_2_in_3.INVTX1_4_.scs8hd_inv_1 top_width_0_height_0__pin_4_ ltile_clb_0.mux_fle_2_in_3.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_26_248 vgnd vpwr scs8hd_decap_3
XFILLER_81_398 vgnd vpwr scs8hd_decap_12
XFILLER_22_410 vgnd vpwr scs8hd_decap_8
XFILLER_22_487 vpwr vgnd scs8hd_fill_2
XFILLER_22_498 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mux_fle_3_in_0.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_3_in_0.INVTX1_9_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_78_15 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_0_.TGATE_1_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ _624_/Y ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_1_314 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.mux_fle_2_in_0.INVTX1_10_.scs8hd_inv_1 bottom_width_0_height_0__pin_10_
+ ltile_clb_0.mux_fle_2_in_0.INVTX1_10_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XFILLER_1_358 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_2_in_0.INVTX1_7_.scs8hd_inv_1_A left_width_0_height_0__pin_7_
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_1_in_0.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_1_in_0.INVTX1_10_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_1_in_0.LATCH_2_.latch/Q ltile_clb_0.mux_fle_1_in_0.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
Xltile_clb_0.mux_fle_3_in_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_3_in_0.INVTX1_5_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_3_in_0.LATCH_1_.latch/Q ltile_clb_0.mux_fle_3_in_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_57_362 vpwr vgnd scs8hd_fill_2
X_601_ _575_/A _600_/X _601_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_45_502 vpwr vgnd scs8hd_fill_2
XFILLER_72_365 vpwr vgnd scs8hd_fill_2
X_532_ _250_/X _529_/X _532_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_27_74 vgnd vpwr scs8hd_decap_12
XFILLER_72_398 vpwr vgnd scs8hd_fill_2
XFILLER_13_410 vpwr vgnd scs8hd_fill_2
XFILLER_32_207 vgnd vpwr scs8hd_decap_6
X_463_ _430_/A _462_/X _463_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_13_443 vgnd vpwr scs8hd_decap_4
X_394_ _394_/A _387_/A _394_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_43_51 vgnd vpwr scs8hd_decap_8
XFILLER_43_62 vgnd vpwr scs8hd_decap_12
XFILLER_13_498 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
+ _633_/Y vgnd vpwr scs8hd_diode_2
XFILLER_4_141 vgnd vpwr scs8hd_decap_12
XFILLER_4_56 vgnd vpwr scs8hd_decap_12
XFILLER_48_351 vpwr vgnd scs8hd_fill_2
XFILLER_82_118 vgnd vpwr scs8hd_decap_6
Xltile_clb_0.mux_fle_2_in_1.INVTX1_12_.scs8hd_inv_1 top_width_0_height_0__pin_12_
+ ltile_clb_0.mux_fle_2_in_1.INVTX1_12_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XFILLER_48_395 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.mux_fle_2_in_3.mux_l1_in_2_.TGATE_3_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_2_in_3.INVTX1_11_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_2_in_3.LATCH_3_.latch/Q ltile_clb_0.mux_fle_2_in_3.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_63_354 vpwr vgnd scs8hd_fill_2
XFILLER_16_281 vgnd vpwr scs8hd_fill_1
XFILLER_31_240 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.mux_fle_0_in_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_0_in_3.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ ltile_clb_0.mem_fle_0_in_3.LATCH_4_.latch/Q ltile_clb_0.mux_fle_0_in_3.INVTX1_14_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_ltile_clb_0.mux_fle_3_in_1.INVTX1_4_.scs8hd_inv_1_A top_width_0_height_0__pin_4_
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_7_.TGATE_1_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_15_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_1_.TGATE_0_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_1_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_8_491 vpwr vgnd scs8hd_fill_2
XANTENNA__305__A _282_/C vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_1_in_3.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_1_in_3.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mem_fle_1_in_3.LATCH_4_.latch_SLEEPB _444_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_1_in_3.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_1_in_3.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_39_351 vpwr vgnd scs8hd_fill_2
XFILLER_54_332 vpwr vgnd scs8hd_fill_2
XFILLER_54_387 vpwr vgnd scs8hd_fill_2
XFILLER_54_376 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_2_in_3.INVTX1_12_.scs8hd_inv_1_A top_width_0_height_0__pin_12_
+ vgnd vpwr scs8hd_diode_2
XFILLER_81_184 vgnd vpwr scs8hd_decap_12
XFILLER_54_398 vgnd vpwr scs8hd_decap_3
XANTENNA_ltile_clb_0.mux_fle_1_in_2.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_1_in_2.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_80_27 vgnd vpwr scs8hd_decap_4
Xltile_clb_0.mux_fle_2_in_2.INVTX1_14_.scs8hd_inv_1 ltile_clb_0.mux_fle_2_in_2.INVTX1_14_.scs8hd_inv_1/A
+ ltile_clb_0.mux_fle_2_in_2.INVTX1_14_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XFILLER_10_435 vgnd vpwr scs8hd_decap_3
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__ff_0.DFFSRQ_0_.dff_SETB
+ set vgnd vpwr scs8hd_diode_2
XFILLER_13_98 vgnd vpwr scs8hd_decap_12
XFILLER_8_3 vgnd vpwr scs8hd_decap_12
XFILLER_77_446 vpwr vgnd scs8hd_fill_2
XFILLER_77_435 vpwr vgnd scs8hd_fill_2
XFILLER_64_129 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_1_.scs8hd_inv_1/Y
+ _604_/Y ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
Xltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_15_.latch
+ data_in ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_15_.latch/Q
+ _244_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_45_332 vgnd vpwr scs8hd_decap_4
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_15_.latch_SLEEPB
+ _556_/Y vgnd vpwr scs8hd_diode_2
X_515_ _409_/A _381_/Y _228_/X _345_/A _516_/A vgnd vpwr scs8hd_or4_4
XFILLER_60_357 vgnd vpwr scs8hd_decap_8
X_446_ _435_/A _446_/B _446_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_13_240 vpwr vgnd scs8hd_fill_2
X_377_ _338_/A _377_/B _377_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_13_284 vpwr vgnd scs8hd_fill_2
XFILLER_9_211 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_0_in_3.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_0_in_3.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_2_.latch
+ data_in ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_2_.latch/Q
+ _596_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_9_255 vgnd vpwr scs8hd_decap_3
XANTENNA_ltile_clb_0.mux_fle_3_in_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_3_in_1.LATCH_4_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_70_93 vgnd vpwr scs8hd_decap_12
XFILLER_5_472 vgnd vpwr scs8hd_decap_4
XFILLER_5_461 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_3_in_1.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_3_in_1.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_68_468 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.mem_fle_1_in_0.LATCH_7_.latch data_in ltile_clb_0.mem_fle_1_in_0.LATCH_7_.latch/Q
+ _474_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_55_129 vpwr vgnd scs8hd_fill_2
XFILLER_36_310 vpwr vgnd scs8hd_fill_2
XFILLER_24_505 vgnd vpwr scs8hd_decap_8
XFILLER_63_184 vgnd vpwr scs8hd_decap_3
Xltile_clb_0.mem_fle_2_in_0.LATCH_6_.latch data_in ltile_clb_0.mem_fle_2_in_0.LATCH_6_.latch/Q
+ _431_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_ltile_clb_0.mem_fle_2_in_2.LATCH_4_.latch_SLEEPB _402_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_3_.TGATE_1_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_7_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_59_39 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.mux_fle_2_in_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_2_in_1.INVTX1_5_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_2_in_1.LATCH_1_.latch/Q ltile_clb_0.mux_fle_2_in_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB
+ _629_/Y vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_0_in_1.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_0_in_1.INVTX1_10_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_0_in_1.LATCH_2_.latch/Q ltile_clb_0.mux_fle_0_in_1.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
Xltile_clb_0.mem_fle_3_in_0.LATCH_5_.latch data_in ltile_clb_0.mem_fle_3_in_0.LATCH_5_.latch/Q
+ _374_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_75_27 vgnd vpwr scs8hd_decap_12
XFILLER_74_405 vgnd vpwr scs8hd_fill_1
XFILLER_59_479 vpwr vgnd scs8hd_fill_2
XFILLER_74_449 vgnd vpwr scs8hd_decap_8
XFILLER_46_129 vgnd vpwr scs8hd_decap_12
XFILLER_27_376 vpwr vgnd scs8hd_fill_2
X_300_ _300_/A _545_/A vgnd vpwr scs8hd_buf_1
XFILLER_42_313 vgnd vpwr scs8hd_decap_6
XFILLER_42_346 vgnd vpwr scs8hd_decap_8
XFILLER_10_210 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_0_in_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_0_in_1.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
X_231_ address[6] _226_/X _228_/X _345_/A _231_/X vgnd vpwr scs8hd_or4_4
XFILLER_6_247 vgnd vpwr scs8hd_decap_3
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.mem_ble4_out_0.LATCH_2_.latch_D
+ data_in vgnd vpwr scs8hd_diode_2
XANTENNA__599__B _578_/X vgnd vpwr scs8hd_diode_2
XFILLER_77_210 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mux_fle_0_in_1.INVTX1_2_.scs8hd_inv_1_A bottom_width_0_height_0__pin_2_
+ vgnd vpwr scs8hd_diode_2
XFILLER_77_243 vgnd vpwr scs8hd_fill_1
XFILLER_77_298 vpwr vgnd scs8hd_fill_2
XFILLER_18_398 vgnd vpwr scs8hd_fill_1
XFILLER_33_313 vpwr vgnd scs8hd_fill_2
XFILLER_45_195 vpwr vgnd scs8hd_fill_2
X_429_ _428_/X _429_/X vgnd vpwr scs8hd_buf_1
XFILLER_60_3 vgnd vpwr scs8hd_decap_12
XANTENNA__302__B _342_/A vgnd vpwr scs8hd_diode_2
XFILLER_68_265 vpwr vgnd scs8hd_fill_2
XFILLER_68_254 vgnd vpwr scs8hd_decap_4
XFILLER_68_243 vgnd vpwr scs8hd_decap_8
XFILLER_68_232 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mem_fle_3_in_1.LATCH_4_.latch_SLEEPB _364_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_0_in_2.INVTX1_11_.scs8hd_inv_1_A left_width_0_height_0__pin_11_
+ vgnd vpwr scs8hd_diode_2
XFILLER_68_276 vgnd vpwr scs8hd_fill_1
XANTENNA_ltile_clb_0.mux_fle_2_in_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_2_in_1.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_28_129 vgnd vpwr scs8hd_decap_12
XFILLER_71_419 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.mem_ble4_out_0.LATCH_2_.latch_SLEEPB
+ _310_/Y vgnd vpwr scs8hd_diode_2
XFILLER_51_110 vgnd vpwr scs8hd_decap_12
XPHY_308 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_319 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_346 vgnd vpwr scs8hd_decap_3
Xltile_clb_0.mux_fle_1_in_3.INVTX1_10_.scs8hd_inv_1 bottom_width_0_height_0__pin_10_
+ ltile_clb_0.mux_fle_1_in_3.INVTX1_10_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XFILLER_10_44 vgnd vpwr scs8hd_decap_12
XFILLER_3_239 vgnd vpwr scs8hd_decap_3
Xltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_1_.scs8hd_inv_1
+ ltile_clb_0.mux_fle_3_in_1.INVTX1_14_.scs8hd_inv_1/Y _607_/A vgnd vpwr scs8hd_inv_1
XFILLER_74_235 vgnd vpwr scs8hd_decap_12
XFILLER_19_86 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_2_.latch
+ data_in ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_2_.latch/Q
+ _570_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_70_430 vgnd vpwr scs8hd_decap_8
XANTENNA_ltile_clb_0.mem_fle_0_in_2.LATCH_5_.latch_SLEEPB _498_/Y vgnd vpwr scs8hd_diode_2
XPHY_820 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_35_74 vgnd vpwr scs8hd_decap_12
XPHY_842 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_831 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_70_474 vgnd vpwr scs8hd_decap_12
XFILLER_30_327 vpwr vgnd scs8hd_fill_2
XFILLER_42_165 vpwr vgnd scs8hd_fill_2
XFILLER_51_51 vgnd vpwr scs8hd_decap_8
XFILLER_51_62 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_1_.TGATE_0_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_1_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XANTENNA__403__A _392_/A vgnd vpwr scs8hd_diode_2
Xltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_1_.TGATE_0_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_1_.TGATE_0_.scs8hd_ebufn_2/A
+ _615_/Y ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_2_250 vgnd vpwr scs8hd_decap_3
XFILLER_2_272 vgnd vpwr scs8hd_decap_3
XFILLER_65_213 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_13_.scs8hd_inv_1_A
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_13_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_65_279 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_1_in_1.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_1_in_1.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_80_227 vgnd vpwr scs8hd_decap_12
XFILLER_33_110 vgnd vpwr scs8hd_decap_12
XFILLER_73_290 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_15_.latch_D
+ data_in vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
+ _607_/Y vgnd vpwr scs8hd_diode_2
XFILLER_61_485 vgnd vpwr scs8hd_decap_3
XFILLER_21_316 vpwr vgnd scs8hd_fill_2
XFILLER_33_165 vgnd vpwr scs8hd_fill_1
Xltile_clb_0.mux_fle_3_in_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_3_in_2.INVTX1_0_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_3_in_2.LATCH_0_.latch/Q ltile_clb_0.mux_fle_3_in_2.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA__313__A _313_/A vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_1_in_2.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_1_in_2.INVTX1_5_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_1_in_2.LATCH_1_.latch/Q ltile_clb_0.mux_fle_1_in_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
Xltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.INVTX1_1_.scs8hd_inv_1/Y
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.mem_ble4_out_0.LATCH_1_.latch/Q
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_56_224 vgnd vpwr scs8hd_decap_12
XFILLER_29_449 vgnd vpwr scs8hd_fill_1
XANTENNA_ltile_clb_0.mux_fle_2_in_1.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_2_in_1.INVTX1_9_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_64_290 vgnd vpwr scs8hd_decap_4
XPHY_116 vgnd vpwr scs8hd_decap_3
XPHY_105 vgnd vpwr scs8hd_decap_3
XFILLER_52_430 vgnd vpwr scs8hd_decap_4
XPHY_149 vgnd vpwr scs8hd_decap_3
XPHY_138 vgnd vpwr scs8hd_decap_3
XPHY_127 vgnd vpwr scs8hd_decap_3
XFILLER_24_154 vgnd vpwr scs8hd_decap_12
XFILLER_20_371 vpwr vgnd scs8hd_fill_2
XFILLER_21_98 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mem_fle_1_in_1.LATCH_5_.latch_SLEEPB _465_/Y vgnd vpwr scs8hd_diode_2
XFILLER_47_213 vpwr vgnd scs8hd_fill_2
XFILLER_15_110 vgnd vpwr scs8hd_decap_12
XPHY_7 vgnd vpwr scs8hd_decap_3
XFILLER_43_496 vgnd vpwr scs8hd_decap_4
XPHY_661 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_650 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_694 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_683 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_672 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_2_.scs8hd_inv_1
+ ltile_clb_0.mux_fle_1_in_2.INVTX1_14_.scs8hd_inv_1/Y _625_/A vgnd vpwr scs8hd_inv_1
XFILLER_30_168 vpwr vgnd scs8hd_fill_2
XFILLER_11_382 vgnd vpwr scs8hd_decap_3
XFILLER_7_331 vpwr vgnd scs8hd_fill_2
XFILLER_7_397 vgnd vpwr scs8hd_fill_1
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_3_.TGATE_1_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_3_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_23_3 vgnd vpwr scs8hd_decap_12
XFILLER_38_257 vgnd vpwr scs8hd_fill_1
XFILLER_38_268 vgnd vpwr scs8hd_decap_6
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_7_.latch_SLEEPB
+ _539_/Y vgnd vpwr scs8hd_diode_2
XFILLER_19_471 vpwr vgnd scs8hd_fill_2
XFILLER_34_430 vgnd vpwr scs8hd_decap_4
XANTENNA_ltile_clb_0.mux_fle_0_in_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_0_in_0.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_61_260 vpwr vgnd scs8hd_fill_2
XFILLER_21_135 vgnd vpwr scs8hd_decap_12
XANTENNA__308__A _599_/A vgnd vpwr scs8hd_diode_2
XFILLER_21_168 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.mux_fle_0_in_3.INVTX1_3_.scs8hd_inv_1 left_width_0_height_0__pin_3_ ltile_clb_0.mux_fle_0_in_3.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_67_39 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_2_.latch
+ data_in ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_2_.latch/Q
+ _544_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_76_308 vgnd vpwr scs8hd_decap_6
XFILLER_69_371 vgnd vpwr scs8hd_fill_1
XFILLER_72_514 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_3_in_2.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_3_in_2.mux_l1_in_3_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_17_419 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_1_in_1.INVTX1_8_.scs8hd_inv_1_A top_width_0_height_0__pin_8_
+ vgnd vpwr scs8hd_diode_2
XFILLER_44_205 vgnd vpwr scs8hd_decap_8
XFILLER_44_227 vpwr vgnd scs8hd_fill_2
XFILLER_16_32 vgnd vpwr scs8hd_decap_12
XFILLER_25_441 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mem_fle_2_in_0.LATCH_5_.latch_SLEEPB _432_/Y vgnd vpwr scs8hd_diode_2
XFILLER_40_433 vgnd vpwr scs8hd_decap_3
XFILLER_8_117 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mux_fle_3_in_1.INVTX1_14_.scs8hd_inv_1_A ltile_clb_0.mux_fle_3_in_1.INVTX1_14_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_4_389 vgnd vpwr scs8hd_decap_6
XFILLER_79_135 vgnd vpwr scs8hd_decap_12
XFILLER_67_319 vpwr vgnd scs8hd_fill_2
XANTENNA__400__B _399_/B vgnd vpwr scs8hd_diode_2
XFILLER_75_352 vpwr vgnd scs8hd_fill_2
XFILLER_35_216 vgnd vpwr scs8hd_fill_1
XFILLER_16_441 vgnd vpwr scs8hd_decap_4
XFILLER_16_463 vgnd vpwr scs8hd_fill_1
XFILLER_16_485 vgnd vpwr scs8hd_decap_12
XPHY_480 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_ltile_clb_0.mux_fle_2_in_2.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_2_in_2.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XPHY_491 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xltile_clb_0.mux_fle_0_in_3.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_0_in_3.INVTX1_5_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_0_in_3.LATCH_1_.latch/Q ltile_clb_0.mux_fle_0_in_3.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
Xltile_clb_0.mux_fle_2_in_3.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_2_in_3.INVTX1_0_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_2_in_3.LATCH_0_.latch/Q ltile_clb_0.mux_fle_2_in_3.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_ltile_clb_0.mux_fle_2_in_2.INVTX1_5_.scs8hd_inv_1_A right_width_0_height_0__pin_5_
+ vgnd vpwr scs8hd_diode_2
XFILLER_58_319 vgnd vpwr scs8hd_decap_6
XANTENNA__310__B _309_/X vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_0_in_0.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_0_in_0.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_78_190 vgnd vpwr scs8hd_decap_12
XFILLER_66_385 vgnd vpwr scs8hd_fill_1
XFILLER_22_477 vgnd vpwr scs8hd_fill_1
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_14_.latch_SLEEPB
+ _531_/Y vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mem_fle_0_in_1.LATCH_4_.latch data_in ltile_clb_0.mem_fle_0_in_1.LATCH_4_.latch/Q
+ _510_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_78_27 vgnd vpwr scs8hd_decap_4
XANTENNA__501__A _421_/A vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_0_in_3.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_0_in_3.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_76_105 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mux_fle_3_in_3.INVTX1_2_.scs8hd_inv_1_A bottom_width_0_height_0__pin_2_
+ vgnd vpwr scs8hd_diode_2
X_600_ _599_/X _600_/X vgnd vpwr scs8hd_buf_1
Xltile_clb_0.mux_fle_2_in_0.INVTX1_0_.scs8hd_inv_1 top_width_0_height_0__pin_0_ ltile_clb_0.mux_fle_2_in_0.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
X_531_ _247_/X _529_/X _531_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_17_205 vpwr vgnd scs8hd_fill_2
XFILLER_17_216 vgnd vpwr scs8hd_fill_1
Xltile_clb_0.mem_fle_1_in_1.LATCH_3_.latch data_in ltile_clb_0.mem_fle_1_in_1.LATCH_3_.latch/Q
+ _467_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_45_514 vpwr vgnd scs8hd_fill_2
XFILLER_27_86 vgnd vpwr scs8hd_decap_12
X_462_ _461_/X _462_/X vgnd vpwr scs8hd_buf_1
X_393_ _338_/A _388_/B _393_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_25_271 vgnd vpwr scs8hd_fill_1
XFILLER_9_426 vgnd vpwr scs8hd_fill_1
XFILLER_43_74 vgnd vpwr scs8hd_decap_12
XFILLER_9_459 vgnd vpwr scs8hd_decap_4
XFILLER_9_448 vpwr vgnd scs8hd_fill_2
XFILLER_40_285 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.mem_fle_2_in_1.LATCH_2_.latch data_in ltile_clb_0.mem_fle_2_in_1.LATCH_2_.latch/Q
+ _422_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_ltile_clb_0.mux_fle_0_in_2.mux_l1_in_3_.TGATE_2_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_0_in_2.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_6_.TGATE_1_.scs8hd_ebufn_2_TEB
+ _628_/Y vgnd vpwr scs8hd_diode_2
XANTENNA__411__A _410_/X vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_1_in_0.INVTX1_9_.scs8hd_inv_1 right_width_0_height_0__pin_9_
+ ltile_clb_0.mux_fle_1_in_0.INVTX1_9_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XFILLER_4_68 vgnd vpwr scs8hd_decap_12
XFILLER_68_93 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mem_fle_0_in_0.LATCH_5_.latch_D data_in vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mem_fle_3_in_1.LATCH_1_.latch data_in ltile_clb_0.mem_fle_3_in_1.LATCH_1_.latch/Q
+ _367_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_ltile_clb_0.mem_fle_0_in_0.LATCH_6_.latch_SLEEPB _519_/Y vgnd vpwr scs8hd_diode_2
XFILLER_48_374 vgnd vpwr scs8hd_decap_4
XFILLER_51_506 vgnd vpwr scs8hd_decap_8
XFILLER_63_399 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
+ _621_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__ff_0.DFFSRQ_0_.dff_CLK
+ clkbuf_1_0_0_clk/X vgnd vpwr scs8hd_diode_2
XFILLER_31_285 vgnd vpwr scs8hd_decap_3
XANTENNA_ltile_clb_0.mem_fle_0_in_1.LATCH_3_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA__305__B _282_/B vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_1_in_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_1_in_2.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_2_in_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_2_in_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ ltile_clb_0.mem_fle_2_in_0.LATCH_4_.latch/Q ltile_clb_0.mux_fle_2_in_0.INVTX1_14_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_ltile_clb_0.mux_fle_2_in_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_2_in_1.LATCH_5_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__321__A _320_/X vgnd vpwr scs8hd_diode_2
XFILLER_58_105 vgnd vpwr scs8hd_decap_12
XFILLER_39_330 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_1_in_0.INVTX1_13_.scs8hd_inv_1_A right_width_0_height_0__pin_13_
+ vgnd vpwr scs8hd_diode_2
XFILLER_39_363 vgnd vpwr scs8hd_decap_3
Xltile_clb_0.mem_fle_0_in_3.LATCH_7_.latch data_in ltile_clb_0.mem_fle_0_in_3.LATCH_7_.latch/Q
+ _485_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_ltile_clb_0.mem_fle_0_in_2.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_14_208 vgnd vpwr scs8hd_decap_6
XFILLER_81_196 vgnd vpwr scs8hd_decap_12
XFILLER_22_274 vgnd vpwr scs8hd_fill_1
XFILLER_6_407 vpwr vgnd scs8hd_fill_2
XFILLER_22_296 vgnd vpwr scs8hd_decap_4
Xltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_2_.scs8hd_inv_1
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_2_.latch/Q
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
Xltile_clb_0.mem_fle_1_in_3.LATCH_6_.latch data_in ltile_clb_0.mem_fle_1_in_3.LATCH_6_.latch/Q
+ _442_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_1_123 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_6_.TGATE_0_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_12_.scs8hd_inv_1/Y
+ _605_/Y ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_3_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA__231__A address[6] vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_3_in_3.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_3_in_3.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ ltile_clb_0.mem_fle_3_in_3.LATCH_5_.latch/Q ltile_clb_0.mux_fle_3_in_3.INVTX1_14_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
Xltile_clb_0.mux_fle_2_in_1.INVTX1_4_.scs8hd_inv_1 top_width_0_height_0__pin_4_ ltile_clb_0.mux_fle_2_in_1.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
Xltile_clb_0.mem_fle_2_in_3.LATCH_5_.latch data_in ltile_clb_0.mem_fle_2_in_3.LATCH_5_.latch/Q
+ _390_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_57_171 vgnd vpwr scs8hd_fill_1
XFILLER_18_514 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_5_.latch_D
+ data_in vgnd vpwr scs8hd_diode_2
XFILLER_72_163 vgnd vpwr scs8hd_decap_4
XFILLER_72_141 vgnd vpwr scs8hd_decap_12
X_514_ _343_/A _514_/B _514_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_45_399 vpwr vgnd scs8hd_fill_2
X_445_ _434_/A _446_/B _445_/Y vgnd vpwr scs8hd_nor2_4
X_376_ _392_/A _377_/B _376_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA_ltile_clb_0.mem_fle_1_in_0.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_9_201 vgnd vpwr scs8hd_fill_1
XANTENNA__406__A _379_/A vgnd vpwr scs8hd_diode_2
XFILLER_9_245 vgnd vpwr scs8hd_decap_4
Xltile_clb_0.mem_fle_3_in_3.LATCH_4_.latch data_in ltile_clb_0.mem_fle_3_in_3.LATCH_4_.latch/Q
+ _332_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_12_.latch_D
+ data_in vgnd vpwr scs8hd_diode_2
Xltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_13_.scs8hd_inv_1
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_13_.latch/Q
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_13_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_ltile_clb_0.mux_fle_0_in_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_0_in_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_76_480 vgnd vpwr scs8hd_decap_12
XFILLER_36_333 vgnd vpwr scs8hd_decap_3
XFILLER_63_163 vpwr vgnd scs8hd_fill_2
XFILLER_63_196 vpwr vgnd scs8hd_fill_2
XFILLER_63_174 vgnd vpwr scs8hd_decap_3
XFILLER_36_388 vgnd vpwr scs8hd_decap_3
XFILLER_51_358 vgnd vpwr scs8hd_decap_4
XANTENNA__316__A address[6] vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_0_in_3.INVTX1_0_.scs8hd_inv_1_A top_width_0_height_0__pin_0_
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.mem_ble4_out_0.LATCH_2_.latch
+ data_in ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.mem_ble4_out_0.LATCH_2_.latch/Q
+ _575_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_ltile_clb_0.mux_fle_1_in_2.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_1_in_2.INVTX1_9_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_59_458 vpwr vgnd scs8hd_fill_2
XFILLER_75_39 vgnd vpwr scs8hd_decap_12
XFILLER_27_344 vpwr vgnd scs8hd_fill_2
XFILLER_39_193 vgnd vpwr scs8hd_decap_3
XFILLER_82_450 vgnd vpwr scs8hd_decap_12
XFILLER_54_163 vpwr vgnd scs8hd_fill_2
XFILLER_27_355 vgnd vpwr scs8hd_decap_3
XFILLER_54_174 vgnd vpwr scs8hd_decap_8
XFILLER_24_32 vgnd vpwr scs8hd_decap_12
XFILLER_42_358 vpwr vgnd scs8hd_fill_2
X_230_ _229_/Y address[5] _345_/A vgnd vpwr scs8hd_or2_4
XANTENNA__226__A address[7] vgnd vpwr scs8hd_diode_2
XFILLER_6_215 vgnd vpwr scs8hd_decap_4
XFILLER_6_259 vgnd vpwr scs8hd_decap_3
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_0_.latch_SLEEPB
+ _572_/Y vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_2_in_2.INVTX1_8_.scs8hd_inv_1 top_width_0_height_0__pin_8_ ltile_clb_0.mux_fle_2_in_2.INVTX1_8_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_2_432 vgnd vpwr scs8hd_decap_6
Xltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_5_.scs8hd_inv_1/Y
+ _612_/Y ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_1_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_77_222 vpwr vgnd scs8hd_fill_2
XFILLER_49_51 vgnd vpwr scs8hd_decap_8
XFILLER_49_62 vgnd vpwr scs8hd_decap_12
XFILLER_65_428 vgnd vpwr scs8hd_decap_3
XFILLER_18_322 vgnd vpwr scs8hd_decap_12
XFILLER_73_461 vgnd vpwr scs8hd_decap_3
XFILLER_45_152 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_7_.scs8hd_inv_1
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_7_.latch/Q
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_33_336 vpwr vgnd scs8hd_fill_2
XFILLER_60_133 vgnd vpwr scs8hd_decap_3
Xltile_clb_0.mux_fle_3_in_1.mux_l1_in_2_.TGATE_3_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_3_in_1.INVTX1_11_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_3_in_1.LATCH_3_.latch/Q ltile_clb_0.mux_fle_3_in_1.mux_l1_in_2_.TGATE_3_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_33_347 vpwr vgnd scs8hd_fill_2
X_428_ _428_/A _428_/X vgnd vpwr scs8hd_buf_1
XFILLER_60_188 vgnd vpwr scs8hd_fill_1
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_1_.latch_D
+ data_in vgnd vpwr scs8hd_diode_2
XFILLER_41_380 vgnd vpwr scs8hd_decap_3
X_359_ _358_/X _368_/B vgnd vpwr scs8hd_buf_1
Xltile_clb_0.mux_fle_1_in_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_1_in_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ ltile_clb_0.mem_fle_1_in_1.LATCH_4_.latch/Q ltile_clb_0.mux_fle_1_in_1.INVTX1_14_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_53_3 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mux_fle_0_in_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_0_in_2.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_5_292 vpwr vgnd scs8hd_fill_2
XFILLER_68_211 vgnd vpwr scs8hd_decap_3
XFILLER_49_480 vpwr vgnd scs8hd_fill_2
XFILLER_64_450 vgnd vpwr scs8hd_decap_8
XFILLER_36_141 vgnd vpwr scs8hd_decap_12
XFILLER_24_314 vgnd vpwr scs8hd_decap_8
XFILLER_36_174 vgnd vpwr scs8hd_decap_8
XFILLER_36_185 vpwr vgnd scs8hd_fill_2
XPHY_309 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_ltile_clb_0.mux_fle_0_in_1.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_0_in_1.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_51_166 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_3_in_2.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_3_in_2.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_2_in_3.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_2_in_3.mux_l1_in_3_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_3_in_3.INVTX1_3_.scs8hd_inv_1 left_width_0_height_0__pin_3_ ltile_clb_0.mux_fle_3_in_3.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_10_56 vgnd vpwr scs8hd_decap_12
XFILLER_59_222 vgnd vpwr scs8hd_decap_3
XFILLER_47_428 vpwr vgnd scs8hd_fill_2
XFILLER_59_299 vpwr vgnd scs8hd_fill_2
XFILLER_19_98 vgnd vpwr scs8hd_decap_12
XFILLER_62_409 vpwr vgnd scs8hd_fill_2
XFILLER_82_280 vgnd vpwr scs8hd_decap_12
XFILLER_55_483 vgnd vpwr scs8hd_decap_3
XFILLER_15_314 vpwr vgnd scs8hd_fill_2
XPHY_810 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_843 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_832 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_821 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_70_486 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_5_.scs8hd_inv_1_A
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_5_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_35_86 vgnd vpwr scs8hd_decap_12
XFILLER_23_380 vpwr vgnd scs8hd_fill_2
XFILLER_42_199 vgnd vpwr scs8hd_decap_6
XFILLER_7_502 vgnd vpwr scs8hd_decap_12
XFILLER_51_74 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__403__B _399_/B vgnd vpwr scs8hd_diode_2
XFILLER_2_240 vgnd vpwr scs8hd_decap_8
XFILLER_2_262 vpwr vgnd scs8hd_fill_2
XFILLER_38_428 vpwr vgnd scs8hd_fill_2
XFILLER_76_93 vgnd vpwr scs8hd_decap_12
XFILLER_65_236 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_1_in_3.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_1_in_3.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_18_141 vgnd vpwr scs8hd_decap_12
XFILLER_46_450 vgnd vpwr scs8hd_decap_8
XFILLER_80_239 vgnd vpwr scs8hd_decap_12
XFILLER_46_483 vgnd vpwr scs8hd_decap_6
XFILLER_61_431 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mem_fle_1_in_2.LATCH_7_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_61_464 vpwr vgnd scs8hd_fill_2
XFILLER_33_199 vgnd vpwr scs8hd_decap_4
Xltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.buf4_1_.scs8hd_buf_1
+ ltile_clb_0.mux_fle_1_in_1.INVTX1_14_.scs8hd_inv_1/Y _622_/A vgnd vpwr scs8hd_buf_1
XANTENNA_ltile_clb_0.mem_fle_1_in_3.LATCH_5_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_29_406 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.mem_ble4_out_0.LATCH_2_.latch_D
+ data_in vgnd vpwr scs8hd_diode_2
XFILLER_56_236 vgnd vpwr scs8hd_decap_4
XFILLER_29_439 vpwr vgnd scs8hd_fill_2
XFILLER_71_217 vpwr vgnd scs8hd_fill_2
XFILLER_52_420 vgnd vpwr scs8hd_decap_8
XFILLER_37_483 vgnd vpwr scs8hd_decap_4
XANTENNA_ltile_clb_0.mux_fle_0_in_2.INVTX1_9_.scs8hd_inv_1_A right_width_0_height_0__pin_9_
+ vgnd vpwr scs8hd_diode_2
XPHY_106 vgnd vpwr scs8hd_decap_3
XPHY_139 vgnd vpwr scs8hd_decap_3
XPHY_128 vgnd vpwr scs8hd_decap_3
XPHY_117 vgnd vpwr scs8hd_decap_3
XFILLER_24_166 vgnd vpwr scs8hd_decap_12
XFILLER_52_497 vgnd vpwr scs8hd_decap_12
XFILLER_24_199 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mem_fle_2_in_0.LATCH_7_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_15_.scs8hd_inv_1_A
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_15_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_20_361 vgnd vpwr scs8hd_fill_1
XANTENNA__504__A _409_/A vgnd vpwr scs8hd_diode_2
XFILLER_79_317 vpwr vgnd scs8hd_fill_2
XFILLER_75_501 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.mux_fle_2_in_2.mux_l1_in_2_.TGATE_3_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_2_in_2.INVTX1_11_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_2_in_2.LATCH_3_.latch/Q ltile_clb_0.mux_fle_2_in_2.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_ltile_clb_0.mem_fle_2_in_1.LATCH_5_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_28_483 vgnd vpwr scs8hd_decap_6
XPHY_8 vgnd vpwr scs8hd_decap_3
XFILLER_43_420 vgnd vpwr scs8hd_decap_6
XFILLER_43_442 vpwr vgnd scs8hd_fill_2
XPHY_662 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_651 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_640 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xltile_clb_0.mux_fle_0_in_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_0_in_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ ltile_clb_0.mem_fle_0_in_2.LATCH_4_.latch/Q ltile_clb_0.mux_fle_0_in_2.INVTX1_14_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XPHY_695 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_684 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_673 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_3_.TGATE_0_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_3_.TGATE_0_.scs8hd_ebufn_2/A
+ _623_/Y ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_3_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA__414__A _431_/A vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_1_in_3.INVTX1_6_.scs8hd_inv_1_A bottom_width_0_height_0__pin_6_
+ vgnd vpwr scs8hd_diode_2
XFILLER_7_376 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_13_.scs8hd_inv_1
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_13_.latch/Q
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_13_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
Xltile_clb_0.mem_fle_0_in_2.LATCH_0_.latch data_in ltile_clb_0.mem_fle_0_in_2.LATCH_0_.latch/Q
+ _503_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_ltile_clb_0.mem_fle_2_in_2.LATCH_3_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_4_.TGATE_1_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_9_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_2_in_0.INVTX1_2_.scs8hd_inv_1_A bottom_width_0_height_0__pin_2_
+ vgnd vpwr scs8hd_diode_2
XFILLER_16_3 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mux_fle_2_in_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_2_in_3.LATCH_4_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_53_206 vgnd vpwr scs8hd_fill_1
XANTENNA_ltile_clb_0.mux_fle_0_in_3.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_0_in_3.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_5_.latch_SLEEPB
+ _289_/Y vgnd vpwr scs8hd_diode_2
XANTENNA__308__B _231_/X vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mem_fle_2_in_3.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_21_147 vgnd vpwr scs8hd_decap_12
XANTENNA__324__A _324_/A vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_3_in_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_3_in_1.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_10_.latch
+ data_in ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_10_.latch/Q
+ _535_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_57_501 vgnd vpwr scs8hd_decap_12
XFILLER_29_203 vpwr vgnd scs8hd_fill_2
XFILLER_29_236 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mem_fle_3_in_0.LATCH_3_.latch_D data_in vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_1_in_0.INVTX1_12_.scs8hd_inv_1 top_width_0_height_0__pin_12_
+ ltile_clb_0.mux_fle_1_in_0.INVTX1_12_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_4_.TGATE_1_.scs8hd_ebufn_2_TEB
+ _620_/Y vgnd vpwr scs8hd_diode_2
XFILLER_16_44 vgnd vpwr scs8hd_decap_12
XFILLER_25_420 vgnd vpwr scs8hd_decap_4
XFILLER_25_475 vgnd vpwr scs8hd_decap_6
XFILLER_40_467 vpwr vgnd scs8hd_fill_2
XFILLER_8_129 vgnd vpwr scs8hd_decap_12
XFILLER_32_32 vgnd vpwr scs8hd_decap_12
XANTENNA__234__A _304_/A vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mem_fle_3_in_1.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_4_335 vgnd vpwr scs8hd_fill_1
XFILLER_79_147 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.mem_ble4_out_0.LATCH_2_.latch
+ data_in ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.mem_ble4_out_0.LATCH_2_.latch/Q
+ _310_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_48_501 vgnd vpwr scs8hd_decap_12
XFILLER_57_62 vgnd vpwr scs8hd_decap_12
XFILLER_57_51 vgnd vpwr scs8hd_decap_8
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_7_.scs8hd_inv_1_A
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_7_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_75_397 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_0_.scs8hd_inv_1
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_0_.latch/Q
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_ltile_clb_0.mux_fle_3_in_3.INVTX1_12_.scs8hd_inv_1_A top_width_0_height_0__pin_12_
+ vgnd vpwr scs8hd_diode_2
XANTENNA__409__A _409_/A vgnd vpwr scs8hd_diode_2
XFILLER_35_239 vgnd vpwr scs8hd_decap_3
XANTENNA_ltile_clb_0.mux_fle_0_in_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_0_in_0.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_7_.latch_D
+ data_in vgnd vpwr scs8hd_diode_2
XFILLER_16_497 vgnd vpwr scs8hd_decap_12
XFILLER_31_412 vpwr vgnd scs8hd_fill_2
XFILLER_31_423 vgnd vpwr scs8hd_decap_4
XFILLER_31_434 vgnd vpwr scs8hd_fill_1
Xltile_clb_0.mux_fle_1_in_1.INVTX1_14_.scs8hd_inv_1 ltile_clb_0.mux_fle_1_in_1.INVTX1_14_.scs8hd_inv_1/A
+ ltile_clb_0.mux_fle_1_in_1.INVTX1_14_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XFILLER_43_283 vgnd vpwr scs8hd_decap_8
XFILLER_31_467 vpwr vgnd scs8hd_fill_2
XPHY_470 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.INVTX1_1_.scs8hd_inv_1_A
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.INVTX1_1_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_31_489 vpwr vgnd scs8hd_fill_2
XPHY_481 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_492 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_11_191 vpwr vgnd scs8hd_fill_2
XFILLER_7_184 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l4_in_0_.TGATE_0_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l4_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ _619_/Y ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_16_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
Xltile_clb_0.mux_fle_0_in_0.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_0_in_0.INVTX1_10_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_0_in_0.LATCH_2_.latch/Q ltile_clb_0.mux_fle_0_in_0.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
Xltile_clb_0.mux_fle_2_in_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_2_in_0.INVTX1_5_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_2_in_0.LATCH_1_.latch/Q ltile_clb_0.mux_fle_2_in_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_3_390 vgnd vpwr scs8hd_decap_6
XANTENNA_ltile_clb_0.mux_fle_3_in_0.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_3_in_0.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_26_206 vpwr vgnd scs8hd_fill_2
XANTENNA__319__A _526_/D vgnd vpwr scs8hd_diode_2
XFILLER_81_378 vgnd vpwr scs8hd_fill_1
XANTENNA_ltile_clb_0.mem_fle_0_in_1.LATCH_0_.latch_SLEEPB _514_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_0_in_3.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_0_in_3.INVTX1_9_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__501__B _495_/X vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_1_in_1.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_1_in_1.LATCH_6_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_76_117 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.mux_fle_1_in_3.mux_l1_in_2_.TGATE_3_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_1_in_3.INVTX1_11_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_1_in_3.LATCH_3_.latch/Q ltile_clb_0.mux_fle_1_in_3.mux_l1_in_2_.TGATE_3_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_ltile_clb_0.mux_fle_3_in_1.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_3_in_1.INVTX1_9_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_3_in_3.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_3_in_3.INVTX1_6_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_3_in_3.LATCH_2_.latch/Q ltile_clb_0.mux_fle_3_in_3.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_69_191 vpwr vgnd scs8hd_fill_2
XFILLER_57_342 vpwr vgnd scs8hd_fill_2
X_530_ _556_/A _529_/X _530_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_57_397 vpwr vgnd scs8hd_fill_2
XFILLER_17_239 vgnd vpwr scs8hd_decap_3
XFILLER_27_98 vgnd vpwr scs8hd_decap_12
X_461_ _460_/X _461_/X vgnd vpwr scs8hd_buf_1
XANTENNA__229__A enable vgnd vpwr scs8hd_diode_2
X_392_ _392_/A _388_/B _392_/Y vgnd vpwr scs8hd_nor2_4
Xltile_clb_0.mux_fle_0_in_1.INVTX1_3_.scs8hd_inv_1 left_width_0_height_0__pin_3_ ltile_clb_0.mux_fle_0_in_1.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_43_86 vgnd vpwr scs8hd_decap_12
XFILLER_4_154 vgnd vpwr scs8hd_decap_12
XFILLER_36_515 vgnd vpwr scs8hd_fill_1
XFILLER_63_323 vpwr vgnd scs8hd_fill_2
XFILLER_63_367 vgnd vpwr scs8hd_fill_1
XFILLER_31_297 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_3_.latch_D
+ data_in vgnd vpwr scs8hd_diode_2
XANTENNA__602__A _270_/B vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_0_in_3.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_0_in_3.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mem_fle_1_in_0.LATCH_0_.latch_SLEEPB _481_/Y vgnd vpwr scs8hd_diode_2
XFILLER_58_117 vgnd vpwr scs8hd_decap_12
XFILLER_66_172 vpwr vgnd scs8hd_fill_2
XFILLER_66_150 vgnd vpwr scs8hd_decap_3
XFILLER_54_301 vpwr vgnd scs8hd_fill_2
XFILLER_66_194 vgnd vpwr scs8hd_decap_6
XFILLER_39_397 vgnd vpwr scs8hd_decap_3
XFILLER_54_356 vgnd vpwr scs8hd_decap_4
XFILLER_10_415 vgnd vpwr scs8hd_fill_1
XFILLER_10_459 vgnd vpwr scs8hd_decap_4
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_7_.TGATE_0_.scs8hd_ebufn_2_TEB
+ _629_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_3_in_3.mux_l1_in_2_.TGATE_3_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_3_in_3.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__512__A _421_/A vgnd vpwr scs8hd_diode_2
XFILLER_1_135 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mux_fle_1_in_2.INVTX1_11_.scs8hd_inv_1_A left_width_0_height_0__pin_11_
+ vgnd vpwr scs8hd_diode_2
XANTENNA__231__B _226_/X vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_4_.TGATE_1_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_9_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_77_459 vpwr vgnd scs8hd_fill_2
XFILLER_57_150 vpwr vgnd scs8hd_fill_2
XFILLER_45_301 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_3_in_0.INVTX1_8_.scs8hd_inv_1_A top_width_0_height_0__pin_8_
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_0_in_2.INVTX1_7_.scs8hd_inv_1 left_width_0_height_0__pin_7_ ltile_clb_0.mux_fle_0_in_2.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_45_345 vpwr vgnd scs8hd_fill_2
XFILLER_60_304 vgnd vpwr scs8hd_decap_12
X_513_ _423_/A _514_/B _513_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_45_378 vpwr vgnd scs8hd_fill_2
XFILLER_60_337 vpwr vgnd scs8hd_fill_2
X_444_ _433_/A _446_/B _444_/Y vgnd vpwr scs8hd_nor2_4
X_375_ _391_/A _377_/B _375_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA__406__B _398_/A vgnd vpwr scs8hd_diode_2
XFILLER_13_297 vgnd vpwr scs8hd_decap_6
Xltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_13_.scs8hd_inv_1
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_13_.latch/Q
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_13_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_ltile_clb_0.mem_fle_3_in_3.LATCH_7_.latch_D data_in vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_0_in_2.INVTX1_10_.scs8hd_inv_1 bottom_width_0_height_0__pin_10_
+ ltile_clb_0.mux_fle_0_in_2.INVTX1_10_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_9_.scs8hd_inv_1_A
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_9_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_1_in_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_1_in_1.INVTX1_5_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_1_in_1.LATCH_1_.latch/Q ltile_clb_0.mux_fle_1_in_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA__422__A _435_/A vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_3_in_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_3_in_1.INVTX1_0_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_3_in_1.LATCH_0_.latch/Q ltile_clb_0.mux_fle_3_in_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_5_452 vgnd vpwr scs8hd_decap_3
XFILLER_5_441 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
+ _638_/HI ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.mem_ble4_out_0.LATCH_2_.latch/Q
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_76_492 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mux_fle_3_in_2.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_3_in_2.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_63_142 vpwr vgnd scs8hd_fill_2
XFILLER_36_367 vpwr vgnd scs8hd_fill_2
XFILLER_51_326 vpwr vgnd scs8hd_fill_2
XANTENNA__332__A _391_/A vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_1_in_0.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_1_in_0.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_59_404 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.mux_fle_0_in_3.INVTX1_12_.scs8hd_inv_1 top_width_0_height_0__pin_12_
+ ltile_clb_0.mux_fle_0_in_3.INVTX1_12_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XFILLER_74_429 vgnd vpwr scs8hd_fill_1
Xltile_clb_0.mux_fle_3_in_3.INVTX1_11_.scs8hd_inv_1 left_width_0_height_0__pin_11_
+ ltile_clb_0.mux_fle_3_in_3.INVTX1_11_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XFILLER_27_301 vpwr vgnd scs8hd_fill_2
XFILLER_27_323 vgnd vpwr scs8hd_fill_1
XFILLER_82_462 vgnd vpwr scs8hd_decap_3
Xltile_clb_0.mux_fle_1_in_3.INVTX1_2_.scs8hd_inv_1 bottom_width_0_height_0__pin_2_
+ ltile_clb_0.mux_fle_1_in_3.INVTX1_2_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XFILLER_24_44 vgnd vpwr scs8hd_decap_12
XANTENNA__507__A _314_/A vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
+ _616_/Y vgnd vpwr scs8hd_diode_2
XFILLER_10_267 vgnd vpwr scs8hd_decap_3
XFILLER_10_289 vgnd vpwr scs8hd_decap_4
XFILLER_40_32 vgnd vpwr scs8hd_decap_12
XANTENNA__242__A _236_/X vgnd vpwr scs8hd_diode_2
Xltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.INVTX1_0_.scs8hd_inv_1
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.INVTX1_0_.scs8hd_inv_1/A
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_77_245 vpwr vgnd scs8hd_fill_2
XFILLER_49_74 vgnd vpwr scs8hd_decap_12
XFILLER_1_15 vgnd vpwr scs8hd_decap_12
XFILLER_65_51 vgnd vpwr scs8hd_decap_8
XFILLER_1_59 vpwr vgnd scs8hd_fill_2
XFILLER_18_312 vgnd vpwr scs8hd_fill_1
XFILLER_18_334 vpwr vgnd scs8hd_fill_2
XFILLER_65_62 vgnd vpwr scs8hd_decap_12
XFILLER_18_367 vpwr vgnd scs8hd_fill_2
XFILLER_73_473 vpwr vgnd scs8hd_fill_2
XFILLER_18_378 vpwr vgnd scs8hd_fill_2
XFILLER_18_389 vgnd vpwr scs8hd_decap_6
XFILLER_45_175 vpwr vgnd scs8hd_fill_2
X_427_ _409_/A _427_/B _384_/X _346_/D _428_/A vgnd vpwr scs8hd_or4_4
XANTENNA__417__A _331_/A vgnd vpwr scs8hd_diode_2
X_358_ address[8] _369_/B _369_/C _358_/D _358_/X vgnd vpwr scs8hd_or4_4
X_289_ _267_/X _541_/A _289_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_5_271 vpwr vgnd scs8hd_fill_2
XFILLER_46_3 vgnd vpwr scs8hd_decap_12
XFILLER_56_407 vpwr vgnd scs8hd_fill_2
XFILLER_64_440 vpwr vgnd scs8hd_fill_2
XFILLER_64_495 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mux_fle_2_in_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_2_in_2.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_24_359 vpwr vgnd scs8hd_fill_2
XFILLER_51_123 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_0_.scs8hd_inv_1/Y
+ _621_/Y ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA__327__A _286_/X vgnd vpwr scs8hd_diode_2
XFILLER_51_156 vgnd vpwr scs8hd_fill_1
Xltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_8_.latch
+ data_in ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_8_.latch/Q
+ _277_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_ltile_clb_0.mux_fle_0_in_0.INVTX1_6_.scs8hd_inv_1_A bottom_width_0_height_0__pin_6_
+ vgnd vpwr scs8hd_diode_2
XFILLER_3_208 vgnd vpwr scs8hd_decap_12
XFILLER_10_68 vgnd vpwr scs8hd_decap_12
XFILLER_74_204 vgnd vpwr scs8hd_decap_8
XFILLER_59_256 vgnd vpwr scs8hd_decap_6
XFILLER_47_418 vpwr vgnd scs8hd_fill_2
XFILLER_55_462 vpwr vgnd scs8hd_fill_2
XFILLER_27_175 vpwr vgnd scs8hd_fill_2
XFILLER_82_292 vgnd vpwr scs8hd_decap_12
XPHY_811 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_800 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_15_348 vpwr vgnd scs8hd_fill_2
XPHY_844 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_833 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_822 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__237__A address[2] vgnd vpwr scs8hd_diode_2
XFILLER_35_98 vgnd vpwr scs8hd_decap_12
XFILLER_70_498 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.mux_fle_0_in_2.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_0_in_2.INVTX1_5_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_0_in_2.LATCH_1_.latch/Q ltile_clb_0.mux_fle_0_in_2.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_42_189 vgnd vpwr scs8hd_fill_1
Xltile_clb_0.mux_fle_2_in_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_2_in_2.INVTX1_0_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_2_in_2.LATCH_0_.latch/Q ltile_clb_0.mux_fle_2_in_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_7_514 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_4_.TGATE_1_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_9_.scs8hd_inv_1/Y
+ _620_/Y ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_2_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_51_86 vgnd vpwr scs8hd_decap_12
XFILLER_2_285 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_0_.scs8hd_inv_1
+ ltile_clb_0.mux_fle_2_in_0.INVTX1_14_.scs8hd_inv_1/Y _613_/A vgnd vpwr scs8hd_inv_1
XANTENNA_ltile_clb_0.mux_fle_1_in_1.INVTX1_3_.scs8hd_inv_1_A left_width_0_height_0__pin_3_
+ vgnd vpwr scs8hd_diode_2
XFILLER_46_440 vgnd vpwr scs8hd_fill_1
XFILLER_46_462 vgnd vpwr scs8hd_decap_8
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_14_.latch_SLEEPB
+ _248_/Y vgnd vpwr scs8hd_diode_2
XFILLER_33_123 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mux_fle_0_in_1.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_0_in_1.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l4_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
+ _634_/Y vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_2_in_0.INVTX1_8_.scs8hd_inv_1 top_width_0_height_0__pin_8_ ltile_clb_0.mux_fle_2_in_0.INVTX1_8_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_ltile_clb_0.mux_fle_3_in_2.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_3_in_2.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB
+ _612_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_1_in_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_1_in_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XANTENNA__610__A _610_/A vgnd vpwr scs8hd_diode_2
XFILLER_2_80 vgnd vpwr scs8hd_decap_12
XFILLER_37_440 vpwr vgnd scs8hd_fill_2
XFILLER_64_270 vgnd vpwr scs8hd_decap_4
XPHY_107 vgnd vpwr scs8hd_decap_3
XPHY_129 vgnd vpwr scs8hd_decap_3
XPHY_118 vgnd vpwr scs8hd_decap_3
XFILLER_52_454 vgnd vpwr scs8hd_fill_1
XFILLER_24_178 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_1_in_3.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_1_in_3.LATCH_5_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_2_in_2.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_2_in_2.INVTX1_9_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_2_in_2.INVTX1_0_.scs8hd_inv_1_A top_width_0_height_0__pin_0_
+ vgnd vpwr scs8hd_diode_2
XANTENNA__504__B _381_/Y vgnd vpwr scs8hd_diode_2
XFILLER_4_506 vgnd vpwr scs8hd_decap_8
XANTENNA__520__A _328_/A vgnd vpwr scs8hd_diode_2
XFILLER_75_513 vgnd vpwr scs8hd_decap_3
XANTENNA_ltile_clb_0.mux_fle_0_in_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_0_in_0.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_28_440 vgnd vpwr scs8hd_decap_12
XFILLER_47_259 vpwr vgnd scs8hd_fill_2
XFILLER_28_462 vpwr vgnd scs8hd_fill_2
XFILLER_55_281 vpwr vgnd scs8hd_fill_2
XPHY_9 vgnd vpwr scs8hd_decap_3
XFILLER_15_123 vgnd vpwr scs8hd_decap_12
XFILLER_28_495 vgnd vpwr scs8hd_decap_12
XFILLER_43_432 vgnd vpwr scs8hd_fill_1
XFILLER_15_167 vpwr vgnd scs8hd_fill_2
XFILLER_43_487 vgnd vpwr scs8hd_fill_1
XPHY_652 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_641 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_630 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_13_.scs8hd_inv_1
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_13_.latch/Q
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_13_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XPHY_696 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_685 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_674 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_663 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xltile_clb_0.mux_fle_3_in_1.INVTX1_3_.scs8hd_inv_1 left_width_0_height_0__pin_3_ ltile_clb_0.mux_fle_3_in_1.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA__414__B _412_/B vgnd vpwr scs8hd_diode_2
XFILLER_7_344 vpwr vgnd scs8hd_fill_2
XANTENNA__430__A _430_/A vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_1_.TGATE_1_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_1_.TGATE_1_.scs8hd_ebufn_2/A
+ _616_/Y ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l4_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_ltile_clb_0.mem_fle_2_in_3.LATCH_6_.latch_SLEEPB _389_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_15_.latch_D
+ data_in vgnd vpwr scs8hd_diode_2
XFILLER_38_204 vpwr vgnd scs8hd_fill_2
XFILLER_38_215 vgnd vpwr scs8hd_decap_4
Xltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_8_.latch
+ data_in ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_8_.latch/Q
+ _590_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_53_218 vpwr vgnd scs8hd_fill_2
XFILLER_61_240 vpwr vgnd scs8hd_fill_2
XFILLER_34_476 vgnd vpwr scs8hd_decap_8
XFILLER_21_159 vgnd vpwr scs8hd_decap_6
Xltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_1_.scs8hd_inv_1
+ ltile_clb_0.mux_fle_0_in_1.INVTX1_14_.scs8hd_inv_1/Y _631_/A vgnd vpwr scs8hd_inv_1
XANTENNA__605__A _605_/A vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_3_in_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_3_in_2.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2/Z
+ ltile_clb_0.mem_fle_3_in_2.LATCH_5_.latch/Q ltile_clb_0.mux_fle_3_in_2.INVTX1_14_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA__340__A _423_/A vgnd vpwr scs8hd_diode_2
XFILLER_69_362 vpwr vgnd scs8hd_fill_2
XFILLER_57_513 vgnd vpwr scs8hd_decap_3
XFILLER_29_248 vpwr vgnd scs8hd_fill_2
XFILLER_29_259 vpwr vgnd scs8hd_fill_2
XFILLER_44_218 vpwr vgnd scs8hd_fill_2
XFILLER_52_262 vgnd vpwr scs8hd_decap_8
XFILLER_52_251 vgnd vpwr scs8hd_decap_3
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_16_56 vgnd vpwr scs8hd_decap_12
XFILLER_25_454 vgnd vpwr scs8hd_decap_4
Xltile_clb_0.mux_fle_1_in_3.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_1_in_3.INVTX1_0_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_1_in_3.LATCH_0_.latch/Q ltile_clb_0.mux_fle_1_in_3.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_25_498 vgnd vpwr scs8hd_decap_3
XANTENNA_ltile_clb_0.mux_fle_3_in_3.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_3_in_3.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_40_457 vgnd vpwr scs8hd_fill_1
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
+ _630_/Y vgnd vpwr scs8hd_diode_2
XFILLER_32_44 vgnd vpwr scs8hd_decap_12
XANTENNA__515__A _409_/A vgnd vpwr scs8hd_diode_2
XFILLER_4_325 vpwr vgnd scs8hd_fill_2
XANTENNA__250__A _250_/A vgnd vpwr scs8hd_diode_2
XFILLER_79_159 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.INVTX1_1_.scs8hd_inv_1
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.INVTX1_1_.scs8hd_inv_1/A
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_ltile_clb_0.mux_fle_2_in_0.INVTX1_13_.scs8hd_inv_1_A right_width_0_height_0__pin_13_
+ vgnd vpwr scs8hd_diode_2
XFILLER_48_513 vgnd vpwr scs8hd_decap_3
XFILLER_57_74 vgnd vpwr scs8hd_decap_12
XFILLER_75_376 vgnd vpwr scs8hd_decap_4
XANTENNA_ltile_clb_0.mux_fle_0_in_1.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_0_in_1.LATCH_7_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_73_62 vgnd vpwr scs8hd_decap_12
XFILLER_73_51 vgnd vpwr scs8hd_decap_8
Xltile_clb_0.mux_fle_3_in_2.INVTX1_7_.scs8hd_inv_1 left_width_0_height_0__pin_7_ ltile_clb_0.mux_fle_3_in_2.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA__409__B _427_/B vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_0_in_0.mux_l1_in_3_.TGATE_2_.scs8hd_ebufn_2_A _640_/HI
+ vgnd vpwr scs8hd_diode_2
XFILLER_31_446 vpwr vgnd scs8hd_fill_2
XPHY_460 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_471 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_ltile_clb_0.mem_fle_3_in_2.LATCH_6_.latch_SLEEPB _350_/Y vgnd vpwr scs8hd_diode_2
XPHY_482 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_493 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__425__A _343_/A vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_3_in_3.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_3_in_3.INVTX1_12_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_3_in_3.LATCH_0_.latch/Q ltile_clb_0.mux_fle_3_in_3.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_ltile_clb_0.mux_fle_2_in_3.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_2_in_3.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_8_.latch_SLEEPB
+ _564_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.mem_ble4_out_0.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_66_332 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_5_.TGATE_0_.scs8hd_ebufn_2_TEB
+ _621_/Y vgnd vpwr scs8hd_diode_2
XFILLER_26_229 vgnd vpwr scs8hd_decap_8
XANTENNA_ltile_clb_0.mux_fle_0_in_1.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_0_in_1.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__335__A _392_/A vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mem_fle_0_in_3.LATCH_7_.latch_SLEEPB _485_/Y vgnd vpwr scs8hd_diode_2
XFILLER_1_339 vgnd vpwr scs8hd_decap_4
XFILLER_76_129 vgnd vpwr scs8hd_decap_12
XFILLER_57_376 vpwr vgnd scs8hd_fill_2
XFILLER_72_335 vgnd vpwr scs8hd_fill_1
XANTENNA_ltile_clb_0.mux_fle_2_in_1.INVTX1_9_.scs8hd_inv_1_A right_width_0_height_0__pin_9_
+ vgnd vpwr scs8hd_diode_2
XFILLER_60_508 vgnd vpwr scs8hd_decap_8
X_460_ _409_/A _226_/X _384_/A _358_/D _460_/X vgnd vpwr scs8hd_or4_4
Xltile_clb_0.mux_fle_3_in_0.mux_l1_in_2_.TGATE_3_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_3_in_0.INVTX1_11_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_3_in_0.LATCH_3_.latch/Q ltile_clb_0.mux_fle_3_in_0.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
X_391_ _391_/A _388_/B _391_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA_ltile_clb_0.mux_fle_3_in_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_3_in_1.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_13_435 vpwr vgnd scs8hd_fill_2
XFILLER_13_479 vgnd vpwr scs8hd_decap_3
XANTENNA__245__A address[0] vgnd vpwr scs8hd_diode_2
XFILLER_43_98 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.mux_fle_1_in_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_1_in_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ ltile_clb_0.mem_fle_1_in_0.LATCH_4_.latch/Q ltile_clb_0.mux_fle_1_in_0.INVTX1_14_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_4_166 vgnd vpwr scs8hd_decap_12
XFILLER_4_15 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_8_.latch
+ data_in ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_8_.latch/Q
+ _564_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_ltile_clb_0.mux_fle_3_in_0.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_3_in_0.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_48_321 vgnd vpwr scs8hd_decap_4
XFILLER_48_332 vgnd vpwr scs8hd_decap_4
XFILLER_63_302 vgnd vpwr scs8hd_decap_3
XFILLER_48_387 vgnd vpwr scs8hd_decap_8
XFILLER_63_335 vpwr vgnd scs8hd_fill_2
XFILLER_63_379 vgnd vpwr scs8hd_decap_3
X_589_ _272_/X _588_/X _589_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_16_295 vgnd vpwr scs8hd_decap_4
XFILLER_31_221 vpwr vgnd scs8hd_fill_2
XFILLER_76_3 vgnd vpwr scs8hd_decap_12
XPHY_290 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xltile_clb_0.mux_fle_2_in_3.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_2_in_3.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ ltile_clb_0.mem_fle_2_in_3.LATCH_5_.latch/Q ltile_clb_0.mux_fle_2_in_3.INVTX1_14_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_ltile_clb_0.mux_fle_3_in_2.INVTX1_6_.scs8hd_inv_1_A bottom_width_0_height_0__pin_6_
+ vgnd vpwr scs8hd_diode_2
XANTENNA__602__B _600_/X vgnd vpwr scs8hd_diode_2
XFILLER_58_129 vgnd vpwr scs8hd_decap_3
XANTENNA_ltile_clb_0.mux_fle_1_in_3.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_1_in_3.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_39_343 vgnd vpwr scs8hd_fill_1
XFILLER_39_376 vgnd vpwr scs8hd_decap_4
XFILLER_81_110 vgnd vpwr scs8hd_decap_12
XFILLER_54_346 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mem_fle_1_in_2.LATCH_7_.latch_SLEEPB _452_/Y vgnd vpwr scs8hd_diode_2
XFILLER_22_276 vpwr vgnd scs8hd_fill_2
XFILLER_10_427 vgnd vpwr scs8hd_decap_8
XANTENNA__512__B _511_/B vgnd vpwr scs8hd_diode_2
XFILLER_1_147 vgnd vpwr scs8hd_decap_12
XANTENNA__231__C _228_/X vgnd vpwr scs8hd_diode_2
XFILLER_49_129 vgnd vpwr scs8hd_fill_1
XFILLER_38_32 vgnd vpwr scs8hd_decap_12
XFILLER_57_184 vgnd vpwr scs8hd_decap_3
XFILLER_72_154 vpwr vgnd scs8hd_fill_2
X_512_ _421_/A _511_/B _512_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_72_176 vgnd vpwr scs8hd_decap_12
X_443_ _432_/A _446_/B _443_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_13_221 vgnd vpwr scs8hd_fill_1
X_374_ _374_/A _377_/B _374_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_13_265 vgnd vpwr scs8hd_fill_1
XFILLER_9_236 vgnd vpwr scs8hd_decap_4
XANTENNA__422__B _412_/B vgnd vpwr scs8hd_diode_2
XFILLER_5_486 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_3_.scs8hd_inv_1
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_3_.latch/Q
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_0_180 vgnd vpwr scs8hd_decap_6
XFILLER_48_151 vpwr vgnd scs8hd_fill_2
XFILLER_63_110 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mux_fle_0_in_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_0_in_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_0_.scs8hd_inv_1_A
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_3_in_3.mux_l1_in_3_.TGATE_2_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_3_in_3.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_8_280 vpwr vgnd scs8hd_fill_2
XANTENNA__613__A _613_/A vgnd vpwr scs8hd_diode_2
XANTENNA__332__B _338_/B vgnd vpwr scs8hd_diode_2
Xltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_2_.TGATE_0_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_2_.TGATE_0_.scs8hd_ebufn_2/A
+ _607_/Y ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_1_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_ltile_clb_0.mem_fle_2_in_1.LATCH_7_.latch_SLEEPB _412_/Y vgnd vpwr scs8hd_diode_2
XFILLER_74_408 vgnd vpwr scs8hd_decap_6
XFILLER_67_471 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.mux_fle_2_in_1.mux_l1_in_2_.TGATE_3_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_2_in_1.INVTX1_11_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_2_in_1.LATCH_3_.latch/Q ltile_clb_0.mux_fle_2_in_1.mux_l1_in_2_.TGATE_3_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_39_162 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_1_in_3.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_1_in_3.INVTX1_9_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_0_in_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_0_in_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ ltile_clb_0.mem_fle_0_in_1.LATCH_4_.latch/Q ltile_clb_0.mux_fle_0_in_1.INVTX1_14_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_24_56 vgnd vpwr scs8hd_decap_12
XANTENNA__507__B _511_/B vgnd vpwr scs8hd_diode_2
XFILLER_50_360 vpwr vgnd scs8hd_fill_2
XFILLER_10_224 vgnd vpwr scs8hd_decap_12
XFILLER_10_202 vgnd vpwr scs8hd_decap_8
Xltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_8_.latch
+ data_in ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_8_.latch/Q
+ _538_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_50_382 vpwr vgnd scs8hd_fill_2
XFILLER_50_393 vpwr vgnd scs8hd_fill_2
XFILLER_10_257 vgnd vpwr scs8hd_fill_1
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_13_.latch_SLEEPB
+ _584_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__ff_0.DFFSRQ_0_.dff_D
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.INVTX1_1_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.buf4_1_.scs8hd_buf_1_A
+ ltile_clb_0.mux_fle_3_in_1.INVTX1_14_.scs8hd_inv_1/Y vgnd vpwr scs8hd_diode_2
XANTENNA__523__A _421_/A vgnd vpwr scs8hd_diode_2
XFILLER_40_44 vgnd vpwr scs8hd_decap_12
XANTENNA__242__B _313_/A vgnd vpwr scs8hd_diode_2
XFILLER_6_3 vgnd vpwr scs8hd_decap_12
XFILLER_49_86 vgnd vpwr scs8hd_decap_12
XFILLER_77_279 vpwr vgnd scs8hd_fill_2
XFILLER_77_257 vpwr vgnd scs8hd_fill_2
XFILLER_1_27 vgnd vpwr scs8hd_decap_12
XFILLER_58_471 vpwr vgnd scs8hd_fill_2
XFILLER_18_302 vgnd vpwr scs8hd_decap_4
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
+ _604_/Y vgnd vpwr scs8hd_diode_2
XFILLER_45_110 vgnd vpwr scs8hd_decap_12
XFILLER_65_74 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mux_fle_0_in_2.INVTX1_4_.scs8hd_inv_1_A top_width_0_height_0__pin_4_
+ vgnd vpwr scs8hd_diode_2
XFILLER_73_485 vgnd vpwr scs8hd_decap_3
XFILLER_60_146 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_12_.latch_D
+ data_in vgnd vpwr scs8hd_diode_2
XFILLER_26_390 vpwr vgnd scs8hd_fill_2
XFILLER_81_62 vgnd vpwr scs8hd_decap_12
XFILLER_81_51 vgnd vpwr scs8hd_decap_8
X_426_ _437_/A _410_/X _426_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_60_157 vgnd vpwr scs8hd_decap_6
X_357_ address[6] address[7] _369_/C vgnd vpwr scs8hd_or2_4
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_10_.scs8hd_inv_1_A
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_10_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__433__A _433_/A vgnd vpwr scs8hd_diode_2
X_288_ _287_/X _541_/A vgnd vpwr scs8hd_buf_1
Xltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_12_.latch
+ data_in ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_12_.latch/Q
+ _559_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_39_3 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.mux_fle_0_in_0.INVTX1_7_.scs8hd_inv_1 left_width_0_height_0__pin_7_ ltile_clb_0.mux_fle_0_in_0.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_56_419 vpwr vgnd scs8hd_fill_2
XFILLER_49_493 vgnd vpwr scs8hd_fill_1
XANTENNA__608__A _608_/A vgnd vpwr scs8hd_diode_2
XFILLER_36_165 vgnd vpwr scs8hd_decap_6
XANTENNA_ltile_clb_0.mem_fle_3_in_0.LATCH_7_.latch_SLEEPB _372_/Y vgnd vpwr scs8hd_diode_2
XFILLER_51_179 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_8_.scs8hd_inv_1
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_8_.latch/Q
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_8_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_32_382 vpwr vgnd scs8hd_fill_2
XANTENNA__343__A _343_/A vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_1_in_3.INVTX1_1_.scs8hd_inv_1_A right_width_0_height_0__pin_1_
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_2_in_2.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_2_in_2.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_27_110 vgnd vpwr scs8hd_decap_12
XPHY_801 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_70_422 vgnd vpwr scs8hd_decap_6
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_1_.latch_SLEEPB
+ _597_/Y vgnd vpwr scs8hd_diode_2
XANTENNA__518__A _314_/A vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_0_in_3.INVTX1_13_.scs8hd_inv_1_A right_width_0_height_0__pin_13_
+ vgnd vpwr scs8hd_diode_2
XPHY_845 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_834 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_823 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_812 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__253__A _252_/X vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_0_in_3.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_0_in_3.LATCH_6_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_1_in_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_1_in_0.LATCH_4_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_51_98 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.mux_fle_1_in_1.INVTX1_2_.scs8hd_inv_1 bottom_width_0_height_0__pin_2_
+ ltile_clb_0.mux_fle_1_in_1.INVTX1_2_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XFILLER_46_430 vgnd vpwr scs8hd_decap_4
XFILLER_18_154 vgnd vpwr scs8hd_decap_12
XANTENNA__428__A _428_/A vgnd vpwr scs8hd_diode_2
XFILLER_33_135 vgnd vpwr scs8hd_decap_12
XFILLER_61_477 vpwr vgnd scs8hd_fill_2
XFILLER_33_168 vpwr vgnd scs8hd_fill_2
XFILLER_33_179 vpwr vgnd scs8hd_fill_2
X_409_ _409_/A _427_/B _384_/X _358_/D _409_/X vgnd vpwr scs8hd_or4_4
XFILLER_14_382 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.mem_fle_3_in_1.LATCH_7_.latch data_in ltile_clb_0.mem_fle_3_in_1.LATCH_7_.latch/Q
+ _361_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
Xltile_clb_0.mux_fle_1_in_2.mux_l1_in_2_.TGATE_3_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_1_in_2.INVTX1_11_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_1_in_2.LATCH_3_.latch/Q ltile_clb_0.mux_fle_1_in_2.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
Xltile_clb_0.mux_fle_3_in_2.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_3_in_2.INVTX1_6_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_3_in_2.LATCH_2_.latch/Q ltile_clb_0.mux_fle_3_in_2.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_2_.scs8hd_inv_1_A
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_29_419 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_4_.scs8hd_inv_1/Y
+ _629_/Y ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_1_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_37_452 vgnd vpwr scs8hd_fill_1
XFILLER_64_260 vgnd vpwr scs8hd_decap_3
XANTENNA__338__A _338_/A vgnd vpwr scs8hd_diode_2
XFILLER_37_496 vgnd vpwr scs8hd_decap_12
XPHY_119 vgnd vpwr scs8hd_decap_3
XPHY_108 vgnd vpwr scs8hd_decap_3
Xltile_clb_0.mux_fle_0_in_0.INVTX1_14_.scs8hd_inv_1 ltile_clb_0.mux_fle_0_in_0.INVTX1_14_.scs8hd_inv_1/A
+ ltile_clb_0.mux_fle_0_in_0.INVTX1_14_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XANTENNA_ltile_clb_0.mux_fle_2_in_0.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_2_in_0.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_20_341 vgnd vpwr scs8hd_fill_1
XFILLER_32_190 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.mux_fle_3_in_0.INVTX1_13_.scs8hd_inv_1 right_width_0_height_0__pin_13_
+ ltile_clb_0.mux_fle_3_in_0.INVTX1_13_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XFILLER_20_396 vgnd vpwr scs8hd_fill_1
XANTENNA__504__C _228_/X vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_3_in_3.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_3_in_3.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__520__B _517_/X vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_7_.TGATE_0_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_14_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_46_32 vgnd vpwr scs8hd_decap_12
XFILLER_47_238 vgnd vpwr scs8hd_decap_4
XFILLER_28_452 vgnd vpwr scs8hd_decap_6
XANTENNA__248__A _248_/A vgnd vpwr scs8hd_diode_2
XFILLER_15_135 vgnd vpwr scs8hd_decap_12
XPHY_620 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_6_.TGATE_1_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_13_.scs8hd_inv_1/Y
+ _628_/Y ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_6_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_43_455 vpwr vgnd scs8hd_fill_2
XPHY_653 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_642 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_631 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_15_179 vpwr vgnd scs8hd_fill_2
XFILLER_30_105 vgnd vpwr scs8hd_decap_12
XPHY_686 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_675 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_ltile_clb_0.mux_fle_3_in_2.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_3_in_2.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XPHY_664 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_11_341 vgnd vpwr scs8hd_fill_1
XPHY_697 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_7_15 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2_TEB
+ _613_/Y vgnd vpwr scs8hd_diode_2
XFILLER_11_396 vpwr vgnd scs8hd_fill_2
XFILLER_7_59 vpwr vgnd scs8hd_fill_2
XFILLER_7_389 vgnd vpwr scs8hd_decap_8
Xltile_clb_0.mux_fle_1_in_2.INVTX1_6_.scs8hd_inv_1 bottom_width_0_height_0__pin_6_
+ ltile_clb_0.mux_fle_1_in_2.INVTX1_6_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XANTENNA__430__B _429_/X vgnd vpwr scs8hd_diode_2
XFILLER_78_374 vgnd vpwr scs8hd_decap_6
Xltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.tap_buf4_0_.scs8hd_inv_1
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.tap_buf4_0_.scs8hd_inv_1/A
+ right_width_0_height_0__pin_13_ vgnd vpwr scs8hd_inv_1
XFILLER_38_227 vgnd vpwr scs8hd_decap_4
XFILLER_19_441 vpwr vgnd scs8hd_fill_2
XFILLER_19_485 vgnd vpwr scs8hd_fill_1
XFILLER_46_271 vgnd vpwr scs8hd_decap_4
XFILLER_46_293 vgnd vpwr scs8hd_fill_1
XFILLER_61_252 vgnd vpwr scs8hd_decap_3
XFILLER_61_285 vgnd vpwr scs8hd_fill_1
XANTENNA_ltile_clb_0.mem_fle_3_in_3.LATCH_0_.latch_SLEEPB _344_/Y vgnd vpwr scs8hd_diode_2
XANTENNA__621__A _621_/A vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_3_in_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_3_in_2.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_29_216 vpwr vgnd scs8hd_fill_2
XFILLER_29_227 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__ff_0.DFFSRQ_0_.dff
+ clkbuf_1_0_0_clk/X ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.INVTX1_1_.scs8hd_inv_1/A
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.INVTX1_0_.scs8hd_inv_1/A
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__ff_0.DFFSRQ_0_.dff/QN
+ reset set vgnd vpwr scs8hd_dfbbp_1
XFILLER_72_506 vgnd vpwr scs8hd_decap_8
XFILLER_25_411 vgnd vpwr scs8hd_decap_3
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_16_68 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.mem_ble4_out_0.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_52_285 vgnd vpwr scs8hd_decap_12
XFILLER_52_274 vgnd vpwr scs8hd_fill_1
XFILLER_12_105 vgnd vpwr scs8hd_decap_12
XFILLER_40_447 vpwr vgnd scs8hd_fill_2
XFILLER_32_56 vgnd vpwr scs8hd_decap_12
XANTENNA__515__B _381_/Y vgnd vpwr scs8hd_diode_2
XFILLER_20_193 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.mux_fle_3_in_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_3_in_0.INVTX1_0_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_3_in_0.LATCH_0_.latch/Q ltile_clb_0.mux_fle_3_in_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
Xltile_clb_0.mux_fle_1_in_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_1_in_0.INVTX1_5_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_1_in_0.LATCH_1_.latch/Q ltile_clb_0.mux_fle_1_in_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA__531__A _247_/X vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_2_in_3.INVTX1_1_.scs8hd_inv_1 right_width_0_height_0__pin_1_
+ ltile_clb_0.mux_fle_2_in_3.INVTX1_1_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XFILLER_57_86 vgnd vpwr scs8hd_decap_12
XFILLER_35_208 vgnd vpwr scs8hd_decap_8
XFILLER_28_271 vpwr vgnd scs8hd_fill_2
XFILLER_28_293 vgnd vpwr scs8hd_fill_1
XFILLER_73_74 vgnd vpwr scs8hd_decap_12
XANTENNA__409__C _384_/X vgnd vpwr scs8hd_diode_2
XFILLER_43_252 vgnd vpwr scs8hd_decap_4
XFILLER_31_403 vpwr vgnd scs8hd_fill_2
XFILLER_43_263 vgnd vpwr scs8hd_fill_1
XPHY_450 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_461 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_472 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_483 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_494 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_ltile_clb_0.mux_fle_2_in_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_2_in_1.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_11_171 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.mux_fle_2_in_3.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_2_in_3.INVTX1_6_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_2_in_3.LATCH_2_.latch/Q ltile_clb_0.mux_fle_2_in_3.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
Xltile_clb_0.mux_fle_0_in_3.mux_l1_in_2_.TGATE_3_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_0_in_3.INVTX1_11_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_0_in_3.LATCH_3_.latch/Q ltile_clb_0.mux_fle_0_in_3.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA__441__A _430_/A vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_2_in_3.INVTX1_7_.scs8hd_inv_1_A left_width_0_height_0__pin_7_
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_2_in_2.INVTX1_11_.scs8hd_inv_1_A left_width_0_height_0__pin_11_
+ vgnd vpwr scs8hd_diode_2
XFILLER_21_3 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mux_fle_3_in_0.INVTX1_3_.scs8hd_inv_1_A left_width_0_height_0__pin_3_
+ vgnd vpwr scs8hd_diode_2
XFILLER_66_377 vpwr vgnd scs8hd_fill_2
XFILLER_26_219 vgnd vpwr scs8hd_fill_1
XANTENNA_ltile_clb_0.mux_fle_2_in_0.mux_l1_in_2_.TGATE_3_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_2_in_0.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_34_252 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mux_fle_2_in_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_2_in_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB
+ _631_/Y vgnd vpwr scs8hd_diode_2
XANTENNA__616__A _616_/A vgnd vpwr scs8hd_diode_2
XANTENNA__335__B _338_/B vgnd vpwr scs8hd_diode_2
XFILLER_22_469 vgnd vpwr scs8hd_decap_8
XFILLER_8_80 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_4_.scs8hd_inv_1_A
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_4_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__351__A _374_/A vgnd vpwr scs8hd_diode_2
XFILLER_1_318 vpwr vgnd scs8hd_fill_2
XFILLER_69_182 vgnd vpwr scs8hd_fill_1
XFILLER_57_322 vgnd vpwr scs8hd_decap_4
XFILLER_72_303 vgnd vpwr scs8hd_decap_4
XFILLER_17_219 vpwr vgnd scs8hd_fill_2
XFILLER_45_506 vgnd vpwr scs8hd_decap_8
XFILLER_72_369 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_3_in_2.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_3_in_2.INVTX1_9_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
X_390_ _374_/A _388_/B _390_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_13_403 vpwr vgnd scs8hd_fill_2
XFILLER_13_414 vpwr vgnd scs8hd_fill_2
XFILLER_25_252 vpwr vgnd scs8hd_fill_2
XFILLER_25_274 vpwr vgnd scs8hd_fill_2
XFILLER_80_391 vgnd vpwr scs8hd_decap_6
XFILLER_9_407 vpwr vgnd scs8hd_fill_2
XFILLER_13_458 vpwr vgnd scs8hd_fill_2
XFILLER_40_233 vpwr vgnd scs8hd_fill_2
XANTENNA__526__A _380_/A vgnd vpwr scs8hd_diode_2
XFILLER_9_418 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mem_fle_1_in_3.LATCH_1_.latch_SLEEPB _447_/Y vgnd vpwr scs8hd_diode_2
XFILLER_21_480 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_1_in_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_1_in_0.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__261__A _260_/X vgnd vpwr scs8hd_diode_2
XFILLER_4_178 vgnd vpwr scs8hd_decap_12
XFILLER_4_27 vgnd vpwr scs8hd_decap_4
XFILLER_0_351 vpwr vgnd scs8hd_fill_2
XFILLER_0_362 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.mux_fle_2_in_2.INVTX1_11_.scs8hd_inv_1 left_width_0_height_0__pin_11_
+ ltile_clb_0.mux_fle_2_in_2.INVTX1_11_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XFILLER_0_384 vpwr vgnd scs8hd_fill_2
XFILLER_0_395 vpwr vgnd scs8hd_fill_2
XFILLER_75_163 vgnd vpwr scs8hd_fill_1
XFILLER_48_355 vgnd vpwr scs8hd_decap_4
XFILLER_63_358 vgnd vpwr scs8hd_decap_6
X_588_ _580_/X _588_/X vgnd vpwr scs8hd_buf_1
XFILLER_16_274 vgnd vpwr scs8hd_fill_1
XFILLER_31_200 vgnd vpwr scs8hd_decap_8
XANTENNA__436__A _436_/A vgnd vpwr scs8hd_diode_2
XPHY_280 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_10_.latch
+ data_in ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_10_.latch/Q
+ _266_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XPHY_291 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_8_473 vgnd vpwr scs8hd_decap_3
XFILLER_69_3 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_12_.latch_SLEEPB
+ _559_/Y vgnd vpwr scs8hd_diode_2
Xltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_7_.scs8hd_inv_1/Y
+ _604_/Y ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_1_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
Xltile_clb_0.mem_fle_0_in_0.LATCH_3_.latch data_in ltile_clb_0.mem_fle_0_in_0.LATCH_3_.latch/Q
+ _522_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
Xltile_clb_0.mux_fle_3_in_0.INVTX1_7_.scs8hd_inv_1 left_width_0_height_0__pin_7_ ltile_clb_0.mux_fle_3_in_0.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_54_325 vgnd vpwr scs8hd_decap_4
XFILLER_54_314 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_7_.TGATE_0_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_14_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_2_in_3.INVTX1_13_.scs8hd_inv_1 right_width_0_height_0__pin_13_
+ ltile_clb_0.mux_fle_2_in_3.INVTX1_13_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
Xltile_clb_0.mem_fle_1_in_0.LATCH_2_.latch data_in ltile_clb_0.mem_fle_1_in_0.LATCH_2_.latch/Q
+ _479_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_ltile_clb_0.mux_fle_3_in_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_3_in_1.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__346__A address[8] vgnd vpwr scs8hd_diode_2
XFILLER_22_266 vgnd vpwr scs8hd_decap_8
Xltile_clb_0.mux_fle_0_in_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_0_in_1.INVTX1_5_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_0_in_1.LATCH_1_.latch/Q ltile_clb_0.mux_fle_0_in_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
Xltile_clb_0.mux_fle_2_in_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_2_in_1.INVTX1_0_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_2_in_1.LATCH_0_.latch/Q ltile_clb_0.mux_fle_2_in_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
Xltile_clb_0.mem_fle_2_in_0.LATCH_1_.latch data_in ltile_clb_0.mem_fle_2_in_0.LATCH_1_.latch/Q
+ _436_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA__231__D _345_/A vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_3_in_0.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_3_in_0.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_1_159 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l4_in_0_.TGATE_1_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l4_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_38_44 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mem_fle_2_in_2.LATCH_1_.latch_SLEEPB _405_/Y vgnd vpwr scs8hd_diode_2
XFILLER_18_506 vgnd vpwr scs8hd_decap_8
XFILLER_57_196 vpwr vgnd scs8hd_fill_2
XFILLER_57_163 vpwr vgnd scs8hd_fill_2
XFILLER_45_336 vgnd vpwr scs8hd_fill_1
XFILLER_54_32 vgnd vpwr scs8hd_decap_12
X_511_ _334_/A _511_/B _511_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_45_358 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.mem_fle_3_in_0.LATCH_0_.latch data_in ltile_clb_0.mem_fle_3_in_0.LATCH_0_.latch/Q
+ _379_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_72_188 vpwr vgnd scs8hd_fill_2
XFILLER_60_328 vgnd vpwr scs8hd_decap_8
XFILLER_13_200 vpwr vgnd scs8hd_fill_2
X_442_ _431_/A _446_/B _442_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA__256__A _255_/X vgnd vpwr scs8hd_diode_2
X_373_ _326_/A _377_/B _373_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_13_255 vpwr vgnd scs8hd_fill_2
XFILLER_9_215 vpwr vgnd scs8hd_fill_2
XFILLER_13_277 vgnd vpwr scs8hd_decap_4
XANTENNA_ltile_clb_0.mux_fle_0_in_1.INVTX1_10_.scs8hd_inv_1_A bottom_width_0_height_0__pin_10_
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_0_in_0.INVTX1_1_.scs8hd_inv_1_A right_width_0_height_0__pin_1_
+ vgnd vpwr scs8hd_diode_2
XFILLER_79_62 vgnd vpwr scs8hd_decap_12
XFILLER_79_51 vgnd vpwr scs8hd_decap_8
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
+ _609_/Y vgnd vpwr scs8hd_diode_2
XFILLER_68_439 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_1_in_0.mux_l1_in_3_.TGATE_2_.scs8hd_ebufn_2_A _644_/HI
+ vgnd vpwr scs8hd_diode_2
XFILLER_76_450 vpwr vgnd scs8hd_fill_2
XFILLER_36_314 vgnd vpwr scs8hd_decap_4
XFILLER_48_185 vpwr vgnd scs8hd_fill_2
XFILLER_51_317 vgnd vpwr scs8hd_decap_3
XFILLER_51_339 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.mem_fle_0_in_2.LATCH_6_.latch data_in ltile_clb_0.mem_fle_0_in_2.LATCH_6_.latch/Q
+ _497_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_3_in_3.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_3_in_3.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mem_fle_1_in_2.LATCH_5_.latch data_in ltile_clb_0.mem_fle_1_in_2.LATCH_5_.latch/Q
+ _454_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_59_428 vpwr vgnd scs8hd_fill_2
XFILLER_67_461 vgnd vpwr scs8hd_decap_3
XANTENNA_ltile_clb_0.mux_fle_1_in_1.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_1_in_1.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_67_483 vgnd vpwr scs8hd_decap_4
XFILLER_82_497 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_6_.scs8hd_inv_1_A
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_6_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_42_328 vgnd vpwr scs8hd_decap_6
Xltile_clb_0.mem_fle_2_in_2.LATCH_4_.latch data_in ltile_clb_0.mem_fle_2_in_2.LATCH_4_.latch/Q
+ _402_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_54_199 vgnd vpwr scs8hd_fill_1
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__ff_0.DFFSRQ_0_.dff_RESETB
+ reset vgnd vpwr scs8hd_diode_2
XFILLER_24_68 vgnd vpwr scs8hd_decap_12
XFILLER_10_236 vgnd vpwr scs8hd_decap_4
XFILLER_6_229 vpwr vgnd scs8hd_fill_2
XANTENNA__523__B _517_/X vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mem_fle_3_in_1.LATCH_1_.latch_SLEEPB _367_/Y vgnd vpwr scs8hd_diode_2
XFILLER_40_56 vgnd vpwr scs8hd_decap_12
XFILLER_2_413 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.mem_fle_3_in_2.LATCH_3_.latch data_in ltile_clb_0.mem_fle_3_in_2.LATCH_3_.latch/Q
+ _353_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_2_468 vpwr vgnd scs8hd_fill_2
XFILLER_49_98 vgnd vpwr scs8hd_decap_12
XFILLER_1_39 vgnd vpwr scs8hd_decap_12
XFILLER_65_86 vgnd vpwr scs8hd_decap_12
XFILLER_33_317 vpwr vgnd scs8hd_fill_2
XFILLER_45_199 vpwr vgnd scs8hd_fill_2
X_425_ _343_/A _437_/A vgnd vpwr scs8hd_buf_1
XFILLER_81_74 vgnd vpwr scs8hd_decap_12
X_356_ _379_/A _355_/B _356_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_41_361 vgnd vpwr scs8hd_decap_3
XANTENNA__433__B _429_/X vgnd vpwr scs8hd_diode_2
X_287_ _278_/X _286_/X _287_/X vgnd vpwr scs8hd_or2_4
XFILLER_5_240 vpwr vgnd scs8hd_fill_2
XFILLER_68_203 vgnd vpwr scs8hd_decap_8
XANTENNA_ltile_clb_0.mem_fle_0_in_2.LATCH_2_.latch_SLEEPB _501_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_0_in_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_0_in_0.LATCH_5_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_3_in_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_3_in_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ ltile_clb_0.mem_fle_3_in_1.LATCH_5_.latch/Q ltile_clb_0.mux_fle_3_in_1.INVTX1_14_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_68_236 vgnd vpwr scs8hd_decap_4
XFILLER_68_269 vgnd vpwr scs8hd_decap_6
XFILLER_49_461 vpwr vgnd scs8hd_fill_2
XFILLER_76_291 vgnd vpwr scs8hd_decap_4
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_7_.TGATE_1_.scs8hd_ebufn_2_TEB
+ _612_/Y vgnd vpwr scs8hd_diode_2
XFILLER_24_328 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.mux_fle_1_in_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_1_in_2.INVTX1_0_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_1_in_2.LATCH_0_.latch/Q ltile_clb_0.mux_fle_1_in_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA__624__A _624_/A vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_2_in_3.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_2_in_3.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_10_15 vgnd vpwr scs8hd_decap_12
XFILLER_59_236 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
+ _605_/Y vgnd vpwr scs8hd_diode_2
XFILLER_55_420 vgnd vpwr scs8hd_fill_1
XFILLER_82_261 vgnd vpwr scs8hd_decap_12
XFILLER_70_412 vgnd vpwr scs8hd_fill_1
XFILLER_15_306 vgnd vpwr scs8hd_fill_1
XPHY_802 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_27_199 vpwr vgnd scs8hd_fill_2
XANTENNA__518__B _517_/X vgnd vpwr scs8hd_diode_2
XPHY_835 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_824 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_813 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_42_169 vpwr vgnd scs8hd_fill_2
XANTENNA__534__A _261_/X vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_3_in_2.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_3_in_2.INVTX1_12_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_3_in_2.LATCH_0_.latch/Q ltile_clb_0.mux_fle_3_in_2.mux_l1_in_3_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.mem_ble4_out_0.LATCH_0_.latch_D
+ data_in vgnd vpwr scs8hd_diode_2
XFILLER_2_221 vgnd vpwr scs8hd_decap_4
XANTENNA_ltile_clb_0.mux_fle_2_in_3.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_2_in_3.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_38_409 vgnd vpwr scs8hd_fill_1
XFILLER_65_217 vpwr vgnd scs8hd_fill_2
XFILLER_18_166 vgnd vpwr scs8hd_decap_8
XFILLER_61_423 vpwr vgnd scs8hd_fill_2
XFILLER_21_309 vgnd vpwr scs8hd_decap_4
XFILLER_33_147 vgnd vpwr scs8hd_decap_12
XFILLER_61_489 vgnd vpwr scs8hd_decap_3
X_408_ address[6] _409_/A vgnd vpwr scs8hd_buf_1
XANTENNA_ltile_clb_0.mem_fle_1_in_1.LATCH_2_.latch_SLEEPB _468_/Y vgnd vpwr scs8hd_diode_2
XANTENNA__444__A _433_/A vgnd vpwr scs8hd_diode_2
X_339_ _339_/A _423_/A vgnd vpwr scs8hd_buf_1
XANTENNA_ltile_clb_0.mux_fle_2_in_2.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_2_in_2.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_51_3 vgnd vpwr scs8hd_decap_12
XFILLER_69_501 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mux_fle_3_in_0.INVTX1_13_.scs8hd_inv_1_A right_width_0_height_0__pin_13_
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_1_in_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_1_in_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_56_206 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l4_in_0_.TGATE_1_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l4_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_2_93 vgnd vpwr scs8hd_decap_12
XANTENNA__619__A _619_/A vgnd vpwr scs8hd_diode_2
XFILLER_49_291 vgnd vpwr scs8hd_fill_1
XFILLER_52_401 vgnd vpwr scs8hd_decap_4
XFILLER_37_464 vpwr vgnd scs8hd_fill_2
XFILLER_37_475 vpwr vgnd scs8hd_fill_2
XANTENNA__338__B _338_/B vgnd vpwr scs8hd_diode_2
XPHY_109 vgnd vpwr scs8hd_decap_3
XANTENNA__354__A _338_/A vgnd vpwr scs8hd_diode_2
Xltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ _622_/Y ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_20_353 vpwr vgnd scs8hd_fill_2
XFILLER_20_375 vgnd vpwr scs8hd_decap_4
XANTENNA__504__D _526_/D vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_1_in_0.INVTX1_7_.scs8hd_inv_1_A left_width_0_height_0__pin_7_
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_2_in_3.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_2_in_3.INVTX1_9_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_4_.latch_SLEEPB
+ _542_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.INVTX1_1_.scs8hd_inv_1_A
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.INVTX1_1_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_47_217 vgnd vpwr scs8hd_decap_6
XANTENNA__529__A _528_/X vgnd vpwr scs8hd_diode_2
XFILLER_28_420 vpwr vgnd scs8hd_fill_2
XFILLER_46_44 vgnd vpwr scs8hd_decap_12
XFILLER_55_294 vgnd vpwr scs8hd_decap_3
XANTENNA__248__B _247_/X vgnd vpwr scs8hd_diode_2
XFILLER_43_412 vpwr vgnd scs8hd_fill_2
XPHY_610 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_15_147 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.mux_fle_0_in_3.INVTX1_0_.scs8hd_inv_1 top_width_0_height_0__pin_0_ ltile_clb_0.mux_fle_0_in_3.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_62_32 vgnd vpwr scs8hd_decap_12
XPHY_643 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_632 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_621 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_30_117 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mux_fle_0_in_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_0_in_1.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XPHY_687 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_676 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_665 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_654 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_11_320 vpwr vgnd scs8hd_fill_2
XANTENNA__264__A _236_/X vgnd vpwr scs8hd_diode_2
XPHY_698 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_11_364 vpwr vgnd scs8hd_fill_2
XFILLER_7_313 vgnd vpwr scs8hd_fill_1
XFILLER_7_27 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.mem_ble4_out_0.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_7_335 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.mux_fle_2_in_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_2_in_2.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2/Z
+ ltile_clb_0.mem_fle_2_in_2.LATCH_5_.latch/Q ltile_clb_0.mux_fle_2_in_2.INVTX1_14_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_78_331 vgnd vpwr scs8hd_decap_4
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
+ _623_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mem_fle_2_in_0.LATCH_2_.latch_SLEEPB _435_/Y vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_0_in_3.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_0_in_3.INVTX1_0_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_0_in_3.LATCH_0_.latch/Q ltile_clb_0.mux_fle_0_in_3.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_19_475 vgnd vpwr scs8hd_decap_4
XANTENNA__439__A _438_/X vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_2_in_1.INVTX1_4_.scs8hd_inv_1_A top_width_0_height_0__pin_4_
+ vgnd vpwr scs8hd_diode_2
XFILLER_34_412 vgnd vpwr scs8hd_decap_3
XFILLER_61_231 vgnd vpwr scs8hd_decap_6
XFILLER_34_445 vpwr vgnd scs8hd_fill_2
XFILLER_61_264 vpwr vgnd scs8hd_fill_2
XFILLER_61_297 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_3_.TGATE_0_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_3_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mem_fle_0_in_1.LATCH_6_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_1_in_1.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_1_in_1.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_69_375 vpwr vgnd scs8hd_fill_2
XANTENNA__349__A _388_/A vgnd vpwr scs8hd_diode_2
XFILLER_37_272 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mem_fle_0_in_2.LATCH_4_.latch_D data_in vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_2_in_3.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_2_in_3.INVTX1_12_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_2_in_3.LATCH_0_.latch/Q ltile_clb_0.mux_fle_2_in_3.mux_l1_in_3_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_ltile_clb_0.mux_fle_3_in_2.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_3_in_2.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_12_117 vgnd vpwr scs8hd_decap_12
XFILLER_52_297 vgnd vpwr scs8hd_decap_4
XFILLER_40_459 vgnd vpwr scs8hd_decap_8
XANTENNA__515__C _228_/X vgnd vpwr scs8hd_diode_2
XFILLER_32_68 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mux_fle_3_in_2.INVTX1_1_.scs8hd_inv_1_A right_width_0_height_0__pin_1_
+ vgnd vpwr scs8hd_diode_2
XFILLER_4_349 vgnd vpwr scs8hd_decap_4
XANTENNA__531__B _529_/X vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mem_fle_0_in_3.LATCH_2_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_75_301 vpwr vgnd scs8hd_fill_2
XFILLER_75_323 vgnd vpwr scs8hd_decap_12
XFILLER_75_356 vgnd vpwr scs8hd_decap_4
XFILLER_57_98 vgnd vpwr scs8hd_decap_12
XANTENNA__259__A _258_/X vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_11_.latch_SLEEPB
+ _534_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_8_.latch_D
+ data_in vgnd vpwr scs8hd_diode_2
XANTENNA__409__D _358_/D vgnd vpwr scs8hd_diode_2
XFILLER_16_445 vgnd vpwr scs8hd_fill_1
XFILLER_16_456 vpwr vgnd scs8hd_fill_2
XFILLER_43_231 vpwr vgnd scs8hd_fill_2
XFILLER_73_86 vgnd vpwr scs8hd_decap_12
XPHY_440 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_451 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_462 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_43_297 vpwr vgnd scs8hd_fill_2
XPHY_473 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_484 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_495 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_ltile_clb_0.mem_fle_1_in_0.LATCH_4_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_7_110 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mux_fle_0_in_1.mux_l1_in_3_.TGATE_2_.scs8hd_ebufn_2_A _641_/HI
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_15_.latch_D
+ data_in vgnd vpwr scs8hd_diode_2
XFILLER_7_198 vpwr vgnd scs8hd_fill_2
XANTENNA__441__B _446_/B vgnd vpwr scs8hd_diode_2
XFILLER_3_360 vgnd vpwr scs8hd_decap_4
XFILLER_14_3 vgnd vpwr scs8hd_decap_12
XFILLER_81_304 vgnd vpwr scs8hd_fill_1
Xltile_clb_0.mux_fle_2_in_0.mux_l1_in_2_.TGATE_3_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_2_in_0.INVTX1_11_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_2_in_0.LATCH_3_.latch/Q ltile_clb_0.mux_fle_2_in_0.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_66_356 vgnd vpwr scs8hd_fill_1
XFILLER_66_389 vgnd vpwr scs8hd_decap_8
XFILLER_19_283 vgnd vpwr scs8hd_decap_3
XANTENNA_ltile_clb_0.mem_fle_1_in_1.LATCH_2_.latch_D data_in vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_0_in_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_0_in_0.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2/Z
+ ltile_clb_0.mem_fle_0_in_0.LATCH_4_.latch/Q ltile_clb_0.mux_fle_0_in_0.INVTX1_14_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_22_459 vgnd vpwr scs8hd_fill_1
Xltile_clb_0.mux_fle_1_in_0.INVTX1_6_.scs8hd_inv_1 bottom_width_0_height_0__pin_6_
+ ltile_clb_0.mux_fle_1_in_0.INVTX1_6_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
Xltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.buf4_1_.scs8hd_buf_1
+ ltile_clb_0.mux_fle_2_in_1.INVTX1_14_.scs8hd_inv_1/Y _614_/A vgnd vpwr scs8hd_buf_1
XANTENNA__632__A _632_/A vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_0_in_2.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_0_in_2.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__351__B _353_/B vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mem_fle_1_in_2.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mem_fle_0_in_0.LATCH_3_.latch_SLEEPB _522_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_3_in_0.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_3_in_0.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_72_337 vgnd vpwr scs8hd_decap_6
Xltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_1_.TGATE_0_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_1_.TGATE_0_.scs8hd_ebufn_2/A
+ _633_/Y ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l4_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_72_348 vgnd vpwr scs8hd_decap_8
Xltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_14_.latch
+ data_in ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_14_.latch/Q
+ _583_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_13_426 vgnd vpwr scs8hd_fill_1
XFILLER_25_297 vpwr vgnd scs8hd_fill_2
XFILLER_40_223 vgnd vpwr scs8hd_fill_1
XANTENNA__526__B address[7] vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_2_in_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_2_in_1.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_40_267 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.mem_fle_0_in_3.LATCH_2_.latch data_in ltile_clb_0.mem_fle_0_in_3.LATCH_2_.latch/Q
+ _490_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
Xltile_clb_0.mux_fle_1_in_3.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_1_in_3.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ ltile_clb_0.mem_fle_1_in_3.LATCH_5_.latch/Q ltile_clb_0.mux_fle_1_in_3.INVTX1_14_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_40_289 vgnd vpwr scs8hd_decap_4
XANTENNA__542__A _542_/A vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mem_fle_1_in_3.LATCH_1_.latch data_in ltile_clb_0.mem_fle_1_in_3.LATCH_1_.latch/Q
+ _447_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_ltile_clb_0.mem_fle_2_in_0.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_48_312 vpwr vgnd scs8hd_fill_2
XFILLER_48_378 vgnd vpwr scs8hd_fill_1
XFILLER_75_175 vgnd vpwr scs8hd_decap_8
XANTENNA_ltile_clb_0.mux_fle_2_in_0.mux_l1_in_3_.TGATE_2_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_2_in_0.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_63_348 vgnd vpwr scs8hd_decap_4
X_587_ _535_/A _585_/B _587_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA_ltile_clb_0.mux_fle_0_in_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_0_in_2.LATCH_4_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__436__B _428_/X vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mem_fle_2_in_3.LATCH_0_.latch data_in ltile_clb_0.mem_fle_2_in_3.LATCH_0_.latch/Q
+ _395_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XPHY_270 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_31_256 vpwr vgnd scs8hd_fill_2
XPHY_281 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_292 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xltile_clb_0.mux_fle_2_in_1.INVTX1_1_.scs8hd_inv_1 right_width_0_height_0__pin_1_
+ ltile_clb_0.mux_fle_2_in_1.INVTX1_1_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XFILLER_8_441 vgnd vpwr scs8hd_decap_4
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_9_.latch_SLEEPB
+ _589_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_4_.latch_D
+ data_in vgnd vpwr scs8hd_diode_2
XFILLER_8_496 vgnd vpwr scs8hd_decap_12
XFILLER_8_485 vgnd vpwr scs8hd_decap_4
XANTENNA__452__A _430_/A vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__ff_0.DFFSRQ_0_.dff_RESETB
+ reset vgnd vpwr scs8hd_diode_2
XFILLER_39_301 vpwr vgnd scs8hd_fill_2
XFILLER_39_334 vgnd vpwr scs8hd_decap_3
XFILLER_66_164 vpwr vgnd scs8hd_fill_2
XFILLER_81_123 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mux_fle_3_in_2.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_3_in_2.LATCH_7_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__627__A _627_/A vgnd vpwr scs8hd_diode_2
XANTENNA__346__B _369_/B vgnd vpwr scs8hd_diode_2
XFILLER_13_15 vgnd vpwr scs8hd_decap_12
XFILLER_10_407 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_10_.scs8hd_inv_1
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_10_.latch/Q
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_10_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_22_289 vgnd vpwr scs8hd_decap_4
XFILLER_13_59 vpwr vgnd scs8hd_fill_2
XANTENNA__362__A _326_/A vgnd vpwr scs8hd_diode_2
XFILLER_38_56 vgnd vpwr scs8hd_decap_12
XFILLER_57_175 vpwr vgnd scs8hd_fill_2
X_510_ _331_/A _511_/B _510_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_45_315 vpwr vgnd scs8hd_fill_2
XFILLER_60_318 vgnd vpwr scs8hd_fill_1
XFILLER_54_44 vgnd vpwr scs8hd_decap_12
XANTENNA__537__A _272_/X vgnd vpwr scs8hd_diode_2
X_441_ _430_/A _446_/B _441_/Y vgnd vpwr scs8hd_nor2_4
X_372_ _388_/A _377_/B _372_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_53_370 vpwr vgnd scs8hd_fill_2
XFILLER_41_510 vgnd vpwr scs8hd_decap_6
XFILLER_13_245 vgnd vpwr scs8hd_fill_1
Xltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_2_.scs8hd_inv_1/Y
+ _613_/Y ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_70_32 vgnd vpwr scs8hd_decap_12
XFILLER_9_249 vgnd vpwr scs8hd_fill_1
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_3_.TGATE_0_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_3_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XANTENNA__272__A _271_/X vgnd vpwr scs8hd_diode_2
XFILLER_79_74 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_5_.TGATE_1_.scs8hd_ebufn_2_TEB
+ _604_/Y vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_1_in_1.mux_l1_in_2_.TGATE_3_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_1_in_1.INVTX1_11_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_1_in_1.LATCH_3_.latch/Q ltile_clb_0.mux_fle_1_in_1.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
Xltile_clb_0.mux_fle_3_in_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_3_in_1.INVTX1_6_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_3_in_1.LATCH_2_.latch/Q ltile_clb_0.mux_fle_3_in_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_63_123 vgnd vpwr scs8hd_decap_12
XFILLER_36_348 vgnd vpwr scs8hd_decap_8
XANTENNA__447__A _436_/A vgnd vpwr scs8hd_diode_2
X_639_ _639_/HI _639_/LO vgnd vpwr scs8hd_conb_1
XANTENNA_ltile_clb_0.mux_fle_1_in_3.INVTX1_13_.scs8hd_inv_1_A right_width_0_height_0__pin_13_
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_2_in_2.INVTX1_5_.scs8hd_inv_1 right_width_0_height_0__pin_5_
+ ltile_clb_0.mux_fle_2_in_2.INVTX1_5_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XFILLER_81_3 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mux_fle_0_in_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_0_in_2.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_5_.TGATE_1_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_11_.scs8hd_inv_1/Y
+ _612_/Y ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_2_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_8_293 vgnd vpwr scs8hd_decap_6
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_0_.latch_D
+ data_in vgnd vpwr scs8hd_diode_2
Xltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_4_.scs8hd_inv_1
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_4_.latch/Q
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_ltile_clb_0.mux_fle_3_in_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_3_in_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_27_315 vpwr vgnd scs8hd_fill_2
XFILLER_39_175 vpwr vgnd scs8hd_fill_2
XFILLER_54_145 vpwr vgnd scs8hd_fill_2
XFILLER_27_348 vpwr vgnd scs8hd_fill_2
XANTENNA__357__A address[6] vgnd vpwr scs8hd_diode_2
XFILLER_54_167 vgnd vpwr scs8hd_decap_4
XFILLER_35_381 vgnd vpwr scs8hd_decap_3
XFILLER_50_373 vgnd vpwr scs8hd_decap_3
XFILLER_6_219 vgnd vpwr scs8hd_fill_1
XFILLER_40_68 vgnd vpwr scs8hd_decap_12
XFILLER_58_451 vgnd vpwr scs8hd_decap_4
XFILLER_73_443 vpwr vgnd scs8hd_fill_2
XFILLER_18_337 vgnd vpwr scs8hd_decap_4
XFILLER_18_348 vpwr vgnd scs8hd_fill_2
XFILLER_45_123 vgnd vpwr scs8hd_decap_12
XFILLER_65_98 vgnd vpwr scs8hd_decap_12
XANTENNA__267__A _304_/A vgnd vpwr scs8hd_diode_2
XFILLER_45_156 vpwr vgnd scs8hd_fill_2
X_424_ _436_/A _410_/X _424_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_41_340 vpwr vgnd scs8hd_fill_2
XFILLER_81_86 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.mux_fle_3_in_3.INVTX1_0_.scs8hd_inv_1 top_width_0_height_0__pin_0_ ltile_clb_0.mux_fle_3_in_3.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_ltile_clb_0.mux_fle_2_in_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_2_in_0.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
X_355_ _394_/A _355_/B _355_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_14_80 vgnd vpwr scs8hd_decap_12
X_286_ _286_/A _286_/B address[1] _286_/X vgnd vpwr scs8hd_or3_4
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_12_.scs8hd_inv_1_A
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_12_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_5_296 vpwr vgnd scs8hd_fill_2
XFILLER_68_215 vgnd vpwr scs8hd_decap_6
XANTENNA_ltile_clb_0.mem_fle_2_in_2.LATCH_6_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_49_484 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.mux_fle_2_in_3.INVTX1_9_.scs8hd_inv_1 right_width_0_height_0__pin_9_
+ ltile_clb_0.mux_fle_2_in_3.INVTX1_9_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XFILLER_64_421 vgnd vpwr scs8hd_decap_8
XANTENNA_ltile_clb_0.mux_fle_1_in_3.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_1_in_3.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_2_in_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_2_in_0.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_17_381 vgnd vpwr scs8hd_decap_4
XFILLER_36_189 vgnd vpwr scs8hd_decap_8
XFILLER_32_340 vgnd vpwr scs8hd_decap_8
XFILLER_32_351 vgnd vpwr scs8hd_decap_8
XFILLER_20_513 vgnd vpwr scs8hd_decap_3
XFILLER_32_373 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mem_fle_2_in_3.LATCH_4_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_10_27 vgnd vpwr scs8hd_decap_4
XANTENNA_ltile_clb_0.mux_fle_0_in_1.INVTX1_8_.scs8hd_inv_1_A top_width_0_height_0__pin_8_
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_1_in_2.mux_l1_in_2_.TGATE_3_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_1_in_2.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_59_248 vpwr vgnd scs8hd_fill_2
XFILLER_74_218 vgnd vpwr scs8hd_decap_6
XANTENNA_ltile_clb_0.mem_fle_3_in_0.LATCH_6_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_55_443 vpwr vgnd scs8hd_fill_2
XFILLER_27_123 vgnd vpwr scs8hd_decap_12
XFILLER_70_402 vgnd vpwr scs8hd_decap_8
XFILLER_27_167 vgnd vpwr scs8hd_decap_3
XFILLER_82_273 vgnd vpwr scs8hd_decap_6
XFILLER_55_498 vpwr vgnd scs8hd_fill_2
XFILLER_15_329 vpwr vgnd scs8hd_fill_2
XPHY_836 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_825 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_814 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_803 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_23_362 vpwr vgnd scs8hd_fill_2
XFILLER_23_384 vpwr vgnd scs8hd_fill_2
XANTENNA__534__B _529_/X vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_0_in_2.mux_l1_in_2_.TGATE_3_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_0_in_2.INVTX1_11_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_0_in_2.LATCH_3_.latch/Q ltile_clb_0.mux_fle_0_in_2.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
Xltile_clb_0.mux_fle_2_in_2.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_2_in_2.INVTX1_6_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_2_in_2.LATCH_2_.latch/Q ltile_clb_0.mux_fle_2_in_2.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_ltile_clb_0.mem_fle_3_in_1.LATCH_4_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA__550__A _270_/B vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__ff_0.DFFSRQ_0_.dff_CLK
+ clkbuf_1_0_0_clk/X vgnd vpwr scs8hd_diode_2
XFILLER_2_266 vgnd vpwr scs8hd_decap_4
XFILLER_46_410 vgnd vpwr scs8hd_decap_4
XFILLER_73_273 vpwr vgnd scs8hd_fill_2
XFILLER_61_435 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_1_in_2.INVTX1_5_.scs8hd_inv_1_A right_width_0_height_0__pin_5_
+ vgnd vpwr scs8hd_diode_2
XFILLER_33_159 vgnd vpwr scs8hd_decap_6
XANTENNA_ltile_clb_0.mem_fle_3_in_2.LATCH_2_.latch_D data_in vgnd vpwr scs8hd_diode_2
XPHY_90 vgnd vpwr scs8hd_decap_3
X_407_ _314_/A _430_/A vgnd vpwr scs8hd_buf_1
X_338_ _338_/A _338_/B _338_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_14_395 vpwr vgnd scs8hd_fill_2
XANTENNA__444__B _446_/B vgnd vpwr scs8hd_diode_2
X_269_ _269_/A _270_/B vgnd vpwr scs8hd_buf_1
XANTENNA_ltile_clb_0.mux_fle_2_in_0.mux_l1_in_3_.TGATE_2_.scs8hd_ebufn_2_A _648_/HI
+ vgnd vpwr scs8hd_diode_2
XANTENNA__460__A _409_/A vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.mem_ble4_out_0.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_44_3 vgnd vpwr scs8hd_decap_12
XFILLER_69_513 vgnd vpwr scs8hd_decap_3
XANTENNA_ltile_clb_0.mem_fle_3_in_3.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_49_281 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_1_.TGATE_1_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_1_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.buf4_1_.scs8hd_buf_1_A
+ ltile_clb_0.mux_fle_0_in_1.INVTX1_14_.scs8hd_inv_1/Y vgnd vpwr scs8hd_diode_2
XFILLER_37_487 vgnd vpwr scs8hd_fill_1
XFILLER_52_457 vgnd vpwr scs8hd_fill_1
XFILLER_52_446 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_10_.scs8hd_inv_1
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_10_.latch/Q
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_10_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_52_479 vgnd vpwr scs8hd_decap_8
XANTENNA__635__A _635_/A vgnd vpwr scs8hd_diode_2
XANTENNA__354__B _353_/B vgnd vpwr scs8hd_diode_2
XFILLER_20_398 vpwr vgnd scs8hd_fill_2
XFILLER_21_15 vgnd vpwr scs8hd_decap_12
XFILLER_21_59 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_3_in_2.INVTX1_11_.scs8hd_inv_1_A left_width_0_height_0__pin_11_
+ vgnd vpwr scs8hd_diode_2
XANTENNA__370__A _370_/A vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_2_in_1.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_2_in_1.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_2_in_3.INVTX1_2_.scs8hd_inv_1_A bottom_width_0_height_0__pin_2_
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_2_in_3.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_2_in_3.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_2_.latch_SLEEPB
+ _298_/Y vgnd vpwr scs8hd_diode_2
XFILLER_46_56 vgnd vpwr scs8hd_decap_12
XFILLER_55_262 vpwr vgnd scs8hd_fill_2
XFILLER_43_402 vgnd vpwr scs8hd_fill_1
XFILLER_70_254 vpwr vgnd scs8hd_fill_2
XFILLER_70_221 vpwr vgnd scs8hd_fill_2
XPHY_611 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_600 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_15_159 vgnd vpwr scs8hd_decap_4
XFILLER_43_446 vgnd vpwr scs8hd_decap_3
XFILLER_43_468 vpwr vgnd scs8hd_fill_2
XFILLER_70_287 vgnd vpwr scs8hd_decap_3
XFILLER_70_276 vpwr vgnd scs8hd_fill_2
XFILLER_62_44 vgnd vpwr scs8hd_decap_12
XPHY_644 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_633 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_622 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__545__A _545_/A vgnd vpwr scs8hd_diode_2
XFILLER_43_479 vpwr vgnd scs8hd_fill_2
XPHY_677 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_666 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_655 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_23_181 vpwr vgnd scs8hd_fill_2
XFILLER_23_192 vgnd vpwr scs8hd_fill_1
XFILLER_30_129 vgnd vpwr scs8hd_decap_12
XPHY_699 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_688 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_7_303 vpwr vgnd scs8hd_fill_2
XANTENNA__264__B _263_/X vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_2_in_2.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_2_in_2.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_11_376 vgnd vpwr scs8hd_decap_4
XFILLER_7_39 vgnd vpwr scs8hd_decap_12
XFILLER_7_358 vpwr vgnd scs8hd_fill_2
XANTENNA__280__A _279_/X vgnd vpwr scs8hd_diode_2
XFILLER_78_354 vgnd vpwr scs8hd_decap_3
XFILLER_19_454 vpwr vgnd scs8hd_fill_2
XFILLER_19_498 vpwr vgnd scs8hd_fill_2
XFILLER_34_424 vgnd vpwr scs8hd_decap_4
XFILLER_34_457 vgnd vpwr scs8hd_fill_1
XANTENNA__455__A _433_/A vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_0_in_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_0_in_0.INVTX1_5_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_0_in_0.LATCH_1_.latch/Q ltile_clb_0.mux_fle_0_in_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
Xltile_clb_0.mux_fle_2_in_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_2_in_0.INVTX1_0_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_2_in_0.LATCH_0_.latch/Q ltile_clb_0.mux_fle_2_in_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_6_391 vgnd vpwr scs8hd_decap_6
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_6_.latch_D
+ data_in vgnd vpwr scs8hd_diode_2
XFILLER_69_343 vgnd vpwr scs8hd_decap_4
XFILLER_69_332 vgnd vpwr scs8hd_decap_4
XFILLER_69_321 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.mem_ble4_out_0.LATCH_0_.latch_D
+ data_in vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_1_in_1.INVTX1_11_.scs8hd_inv_1 left_width_0_height_0__pin_11_
+ ltile_clb_0.mux_fle_1_in_1.INVTX1_11_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.buf4_3_.scs8hd_buf_1_A
+ ltile_clb_0.mux_fle_2_in_3.INVTX1_14_.scs8hd_inv_1/Y vgnd vpwr scs8hd_diode_2
XANTENNA__349__B _353_/B vgnd vpwr scs8hd_diode_2
XFILLER_37_240 vpwr vgnd scs8hd_fill_2
XFILLER_16_15 vgnd vpwr scs8hd_decap_12
XFILLER_25_424 vgnd vpwr scs8hd_fill_1
Xltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_2_.TGATE_1_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_5_.TGATE_0_.scs8hd_ebufn_2/Z
+ _630_/Y ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_1_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_ltile_clb_0.mux_fle_3_in_3.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_3_in_3.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__365__A _392_/A vgnd vpwr scs8hd_diode_2
XFILLER_12_129 vgnd vpwr scs8hd_decap_12
XANTENNA__515__D _345_/A vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_1_in_3.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_1_in_3.INVTX1_6_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_1_in_3.LATCH_2_.latch/Q ltile_clb_0.mux_fle_1_in_3.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_20_162 vgnd vpwr scs8hd_fill_1
Xltile_clb_0.mux_fle_3_in_3.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_3_in_3.INVTX1_1_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_3_in_3.LATCH_1_.latch/Q ltile_clb_0.mux_fle_3_in_3.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_4_317 vgnd vpwr scs8hd_fill_1
Xltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.INVTX1_1_.scs8hd_inv_1/Y
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.mem_ble4_out_0.LATCH_1_.latch/Q
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_75_335 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__ff_0.DFFSRQ_0_.dff_RESETB
+ reset vgnd vpwr scs8hd_diode_2
XFILLER_63_508 vgnd vpwr scs8hd_decap_8
XANTENNA__259__B _259_/B vgnd vpwr scs8hd_diode_2
XFILLER_16_402 vgnd vpwr scs8hd_decap_4
XFILLER_43_243 vgnd vpwr scs8hd_fill_1
Xltile_clb_0.mux_fle_1_in_2.INVTX1_13_.scs8hd_inv_1 right_width_0_height_0__pin_13_
+ ltile_clb_0.mux_fle_1_in_2.INVTX1_13_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XFILLER_73_98 vgnd vpwr scs8hd_decap_12
XANTENNA__275__A _236_/X vgnd vpwr scs8hd_diode_2
XPHY_430 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_441 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_452 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_463 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_474 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_485 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_496 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_11_184 vgnd vpwr scs8hd_decap_4
XFILLER_22_80 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mux_fle_1_in_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_1_in_1.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_0_in_1.INVTX1_0_.scs8hd_inv_1 top_width_0_height_0__pin_0_ ltile_clb_0.mux_fle_0_in_1.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_54_508 vgnd vpwr scs8hd_decap_8
XFILLER_34_243 vgnd vpwr scs8hd_fill_1
XFILLER_22_427 vpwr vgnd scs8hd_fill_2
XFILLER_22_438 vpwr vgnd scs8hd_fill_2
XFILLER_22_449 vpwr vgnd scs8hd_fill_2
XFILLER_34_287 vgnd vpwr scs8hd_fill_1
XANTENNA_ltile_clb_0.mux_fle_1_in_1.INVTX1_10_.scs8hd_inv_1_A bottom_width_0_height_0__pin_10_
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_2_in_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_2_in_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_8_93 vgnd vpwr scs8hd_decap_12
XFILLER_1_309 vgnd vpwr scs8hd_decap_3
XFILLER_69_151 vgnd vpwr scs8hd_fill_1
XFILLER_69_184 vgnd vpwr scs8hd_decap_4
XFILLER_57_346 vgnd vpwr scs8hd_decap_3
XFILLER_72_327 vgnd vpwr scs8hd_decap_8
XFILLER_72_316 vpwr vgnd scs8hd_fill_2
XFILLER_65_390 vgnd vpwr scs8hd_decap_4
XFILLER_25_221 vpwr vgnd scs8hd_fill_2
XFILLER_25_243 vgnd vpwr scs8hd_fill_1
XFILLER_25_287 vpwr vgnd scs8hd_fill_2
XFILLER_40_213 vgnd vpwr scs8hd_fill_1
XANTENNA__526__C _228_/X vgnd vpwr scs8hd_diode_2
XFILLER_21_471 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_3_in_3.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_3_in_3.INVTX1_9_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__542__B _541_/B vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_3_in_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_3_in_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2/Z
+ ltile_clb_0.mem_fle_3_in_0.LATCH_5_.latch/Q ltile_clb_0.mux_fle_3_in_0.INVTX1_14_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_68_32 vgnd vpwr scs8hd_decap_12
XFILLER_0_320 vpwr vgnd scs8hd_fill_2
XFILLER_0_331 vgnd vpwr scs8hd_decap_4
XFILLER_75_110 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mux_fle_1_in_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_1_in_1.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_48_346 vgnd vpwr scs8hd_decap_3
XFILLER_75_187 vpwr vgnd scs8hd_fill_2
XFILLER_63_327 vgnd vpwr scs8hd_fill_1
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_1_.scs8hd_inv_1_A
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
X_655_ _655_/HI _655_/LO vgnd vpwr scs8hd_conb_1
XFILLER_56_390 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_1_.TGATE_1_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_1_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
X_586_ _261_/X _585_/B _586_/Y vgnd vpwr scs8hd_nor2_4
Xltile_clb_0.mux_fle_1_in_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_1_in_1.INVTX1_0_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_1_in_1.LATCH_0_.latch/Q ltile_clb_0.mux_fle_1_in_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_71_371 vpwr vgnd scs8hd_fill_2
XFILLER_16_276 vgnd vpwr scs8hd_decap_3
XPHY_260 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_31_268 vpwr vgnd scs8hd_fill_2
XPHY_271 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_8_420 vgnd vpwr scs8hd_decap_8
XPHY_282 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_293 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_12_493 vgnd vpwr scs8hd_decap_8
XANTENNA__452__B _451_/X vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_0_in_2.INVTX1_4_.scs8hd_inv_1 top_width_0_height_0__pin_4_ ltile_clb_0.mux_fle_0_in_2.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_ltile_clb_0.mux_fle_3_in_3.INVTX1_8_.scs8hd_inv_1_A top_width_0_height_0__pin_8_
+ vgnd vpwr scs8hd_diode_2
XFILLER_66_154 vgnd vpwr scs8hd_fill_1
XFILLER_27_508 vgnd vpwr scs8hd_decap_8
XFILLER_81_135 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_10_.scs8hd_inv_1
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_10_.latch/Q
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_10_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_62_393 vgnd vpwr scs8hd_decap_4
XANTENNA__346__C _346_/C vgnd vpwr scs8hd_diode_2
XFILLER_22_224 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_2_in_1.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_2_in_1.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_13_27 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.mux_fle_3_in_1.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_3_in_1.INVTX1_12_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_3_in_1.LATCH_0_.latch/Q ltile_clb_0.mux_fle_3_in_1.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA__362__B _365_/B vgnd vpwr scs8hd_diode_2
XFILLER_77_419 vpwr vgnd scs8hd_fill_2
XFILLER_57_110 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.mem_ble4_out_0.LATCH_0_.latch
+ data_in ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.mem_ble4_out_0.LATCH_0_.latch/Q
+ _551_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_38_68 vgnd vpwr scs8hd_decap_12
X_440_ _447_/B _446_/B vgnd vpwr scs8hd_buf_1
XFILLER_54_56 vgnd vpwr scs8hd_decap_12
XANTENNA__537__B _541_/B vgnd vpwr scs8hd_diode_2
X_371_ _379_/B _377_/B vgnd vpwr scs8hd_buf_1
XFILLER_13_224 vpwr vgnd scs8hd_fill_2
XFILLER_80_190 vgnd vpwr scs8hd_decap_12
XFILLER_70_44 vgnd vpwr scs8hd_decap_12
XFILLER_9_228 vpwr vgnd scs8hd_fill_2
XANTENNA__553__A address[4] vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_4_.TGATE_0_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_8_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_5_445 vpwr vgnd scs8hd_fill_2
XFILLER_5_423 vpwr vgnd scs8hd_fill_2
XFILLER_5_489 vgnd vpwr scs8hd_decap_12
XFILLER_5_478 vgnd vpwr scs8hd_decap_8
XFILLER_79_86 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mux_fle_0_in_0.INVTX1_14_.scs8hd_inv_1_A ltile_clb_0.mux_fle_0_in_0.INVTX1_14_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_36_327 vgnd vpwr scs8hd_decap_4
XFILLER_48_154 vpwr vgnd scs8hd_fill_2
XFILLER_63_135 vgnd vpwr scs8hd_decap_4
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB
+ _614_/Y vgnd vpwr scs8hd_diode_2
XFILLER_63_179 vpwr vgnd scs8hd_fill_2
XFILLER_63_157 vgnd vpwr scs8hd_decap_4
XANTENNA__447__B _447_/B vgnd vpwr scs8hd_diode_2
X_638_ _638_/HI _638_/LO vgnd vpwr scs8hd_conb_1
XANTENNA_ltile_clb_0.mux_fle_1_in_1.mux_l1_in_3_.TGATE_2_.scs8hd_ebufn_2_A _645_/HI
+ vgnd vpwr scs8hd_diode_2
XFILLER_44_371 vgnd vpwr scs8hd_decap_4
X_569_ _569_/A _554_/X _569_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA__463__A _430_/A vgnd vpwr scs8hd_diode_2
XFILLER_74_3 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.mux_fle_0_in_3.INVTX1_8_.scs8hd_inv_1 top_width_0_height_0__pin_8_ ltile_clb_0.mux_fle_0_in_3.INVTX1_8_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_59_419 vpwr vgnd scs8hd_fill_2
XFILLER_39_110 vgnd vpwr scs8hd_decap_12
XFILLER_39_143 vpwr vgnd scs8hd_fill_2
XFILLER_54_135 vgnd vpwr scs8hd_fill_1
XFILLER_27_327 vpwr vgnd scs8hd_fill_2
XFILLER_39_198 vgnd vpwr scs8hd_decap_3
XFILLER_82_466 vgnd vpwr scs8hd_decap_12
XANTENNA__357__B address[7] vgnd vpwr scs8hd_diode_2
XFILLER_24_15 vgnd vpwr scs8hd_decap_12
XFILLER_35_371 vgnd vpwr scs8hd_decap_4
XANTENNA_ltile_clb_0.mux_fle_1_in_2.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_1_in_2.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_0_in_3.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_0_in_3.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_50_341 vgnd vpwr scs8hd_decap_4
XANTENNA__373__A _326_/A vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_1_in_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_1_in_0.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_10_249 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.mux_fle_2_in_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_2_in_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ ltile_clb_0.mem_fle_2_in_1.LATCH_5_.latch/Q ltile_clb_0.mux_fle_2_in_1.INVTX1_14_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_6_.TGATE_0_.scs8hd_ebufn_2_TEB
+ _605_/Y vgnd vpwr scs8hd_diode_2
Xltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_3_.latch
+ data_in ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_3_.latch/Q
+ _295_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_77_227 vpwr vgnd scs8hd_fill_2
XFILLER_77_249 vgnd vpwr scs8hd_fill_1
XFILLER_73_400 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.mux_fle_0_in_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_0_in_2.INVTX1_0_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_0_in_2.LATCH_0_.latch/Q ltile_clb_0.mux_fle_0_in_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
Xltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_6_.scs8hd_inv_1/Y
+ _621_/Y ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_1_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA__548__A _547_/X vgnd vpwr scs8hd_diode_2
XFILLER_45_135 vpwr vgnd scs8hd_fill_2
XFILLER_73_477 vgnd vpwr scs8hd_decap_8
XFILLER_60_105 vgnd vpwr scs8hd_decap_12
XFILLER_45_179 vpwr vgnd scs8hd_fill_2
X_423_ _423_/A _436_/A vgnd vpwr scs8hd_buf_1
XFILLER_60_138 vgnd vpwr scs8hd_decap_8
XANTENNA_ltile_clb_0.mux_fle_0_in_3.INVTX1_6_.scs8hd_inv_1_A bottom_width_0_height_0__pin_6_
+ vgnd vpwr scs8hd_diode_2
X_354_ _338_/A _353_/B _354_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_41_385 vpwr vgnd scs8hd_fill_2
XFILLER_81_98 vgnd vpwr scs8hd_decap_12
X_285_ _267_/X _540_/A _285_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA__283__A _278_/X vgnd vpwr scs8hd_diode_2
XFILLER_41_396 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_1_in_0.INVTX1_2_.scs8hd_inv_1_A bottom_width_0_height_0__pin_2_
+ vgnd vpwr scs8hd_diode_2
XFILLER_5_275 vpwr vgnd scs8hd_fill_2
XFILLER_30_80 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_6_.TGATE_1_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_13_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_64_444 vgnd vpwr scs8hd_decap_4
XANTENNA__458__A _436_/A vgnd vpwr scs8hd_diode_2
XFILLER_36_157 vpwr vgnd scs8hd_fill_2
XFILLER_51_127 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.mux_fle_2_in_2.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_2_in_2.INVTX1_12_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_2_in_2.LATCH_0_.latch/Q ltile_clb_0.mux_fle_2_in_2.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_51_138 vpwr vgnd scs8hd_fill_2
XFILLER_51_149 vgnd vpwr scs8hd_decap_4
Xltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_7_.TGATE_1_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_15_.scs8hd_inv_1/Y
+ _620_/Y ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_7_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_59_227 vpwr vgnd scs8hd_fill_2
XFILLER_59_205 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_11_.latch_SLEEPB
+ _262_/Y vgnd vpwr scs8hd_diode_2
XFILLER_19_15 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.mux_fle_2_in_0.INVTX1_5_.scs8hd_inv_1 right_width_0_height_0__pin_5_
+ ltile_clb_0.mux_fle_2_in_0.INVTX1_5_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XFILLER_19_59 vpwr vgnd scs8hd_fill_2
XANTENNA__368__A _379_/A vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
+ _632_/Y vgnd vpwr scs8hd_diode_2
XFILLER_27_135 vgnd vpwr scs8hd_decap_12
XFILLER_82_230 vgnd vpwr scs8hd_decap_12
XFILLER_55_466 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_14_.scs8hd_inv_1_A
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_14_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_27_179 vpwr vgnd scs8hd_fill_2
XFILLER_42_105 vgnd vpwr scs8hd_decap_12
XPHY_826 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_815 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_804 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_23_341 vpwr vgnd scs8hd_fill_2
XPHY_837 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_11_503 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.tap_buf4_0_.scs8hd_inv_1
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.tap_buf4_0_.scs8hd_inv_1/A
+ top_width_0_height_0__pin_12_ vgnd vpwr scs8hd_inv_1
XANTENNA__550__B _548_/X vgnd vpwr scs8hd_diode_2
XFILLER_4_3 vgnd vpwr scs8hd_decap_12
XFILLER_2_289 vgnd vpwr scs8hd_decap_3
XFILLER_76_32 vgnd vpwr scs8hd_decap_12
XANTENNA__278__A address[3] vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_1_in_3.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_1_in_3.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_73_252 vpwr vgnd scs8hd_fill_2
XFILLER_61_403 vgnd vpwr scs8hd_fill_1
X_406_ _379_/A _398_/A _406_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_14_341 vgnd vpwr scs8hd_decap_4
XFILLER_14_352 vgnd vpwr scs8hd_decap_12
XPHY_80 vgnd vpwr scs8hd_decap_3
XPHY_91 vgnd vpwr scs8hd_decap_3
Xltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_0_.TGATE_0_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ _617_/Y ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l4_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_41_171 vpwr vgnd scs8hd_fill_2
X_337_ _421_/A _338_/A vgnd vpwr scs8hd_buf_1
X_268_ _286_/B address[1] _269_/A vgnd vpwr scs8hd_or2_4
XANTENNA__460__B _226_/X vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_1_in_2.mux_l1_in_3_.TGATE_2_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_1_in_2.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_37_3 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_10_.scs8hd_inv_1
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_10_.latch/Q
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_10_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
Xclkbuf_1_1_0_clk clkbuf_0_clk/X clkbuf_1_1_0_clk/X vgnd vpwr scs8hd_clkbuf_1
XFILLER_37_400 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.mux_fle_3_in_1.INVTX1_0_.scs8hd_inv_1 top_width_0_height_0__pin_0_ ltile_clb_0.mux_fle_3_in_1.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_37_444 vgnd vpwr scs8hd_decap_8
XFILLER_64_274 vgnd vpwr scs8hd_fill_1
XFILLER_24_105 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mux_fle_1_in_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_1_in_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_52_436 vgnd vpwr scs8hd_fill_1
Xltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_3_.latch
+ data_in ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_3_.latch/Q
+ _595_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_20_311 vgnd vpwr scs8hd_decap_4
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__ff_0.DFFSRQ_0_.dff_RESETB
+ reset vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_1_in_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_1_in_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ ltile_clb_0.mem_fle_1_in_2.LATCH_5_.latch/Q ltile_clb_0.mux_fle_1_in_2.INVTX1_14_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_20_388 vpwr vgnd scs8hd_fill_2
XFILLER_21_27 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_7_.scs8hd_inv_1
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_7_.latch/Q
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_ltile_clb_0.mem_fle_2_in_3.LATCH_3_.latch_SLEEPB _392_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_4_.TGATE_0_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_8_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_2_in_1.INVTX1_9_.scs8hd_inv_1 right_width_0_height_0__pin_9_
+ ltile_clb_0.mux_fle_2_in_1.INVTX1_9_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XANTENNA_ltile_clb_0.mux_fle_3_in_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_3_in_1.LATCH_5_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_28_466 vgnd vpwr scs8hd_decap_8
XFILLER_46_68 vgnd vpwr scs8hd_decap_12
XPHY_601 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_634 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_623 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_612 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__545__B _528_/X vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mem_fle_2_in_0.LATCH_7_.latch data_in ltile_clb_0.mem_fle_2_in_0.LATCH_7_.latch/Q
+ _430_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XPHY_678 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_62_56 vgnd vpwr scs8hd_decap_12
XPHY_667 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_656 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_645 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_51_480 vpwr vgnd scs8hd_fill_2
XFILLER_23_171 vgnd vpwr scs8hd_decap_8
XPHY_689 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_11_344 vgnd vpwr scs8hd_decap_3
XFILLER_7_348 vgnd vpwr scs8hd_fill_1
XANTENNA__561__A _535_/A vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_0_in_2.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_0_in_2.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mem_fle_3_in_0.LATCH_6_.latch data_in ltile_clb_0.mem_fle_3_in_0.LATCH_6_.latch/Q
+ _373_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_78_366 vpwr vgnd scs8hd_fill_2
XFILLER_38_208 vgnd vpwr scs8hd_decap_6
XFILLER_38_219 vgnd vpwr scs8hd_fill_1
Xltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.mem_ble4_out_0.LATCH_0_.latch
+ data_in ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.mem_ble4_out_0.LATCH_0_.latch/Q
+ _603_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_ltile_clb_0.mux_fle_3_in_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_3_in_0.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_1_in_3.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_1_in_3.INVTX1_12_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_1_in_3.LATCH_0_.latch/Q ltile_clb_0.mux_fle_1_in_3.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_46_285 vgnd vpwr scs8hd_decap_8
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB
+ _628_/Y vgnd vpwr scs8hd_diode_2
XFILLER_61_277 vpwr vgnd scs8hd_fill_2
XANTENNA__455__B _451_/X vgnd vpwr scs8hd_diode_2
XANTENNA__471__A _409_/A vgnd vpwr scs8hd_diode_2
XFILLER_69_300 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_0_in_1.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_0_in_1.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_3_in_2.INVTX1_4_.scs8hd_inv_1 top_width_0_height_0__pin_4_ ltile_clb_0.mux_fle_3_in_2.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_ltile_clb_0.mem_fle_3_in_2.LATCH_3_.latch_SLEEPB _353_/Y vgnd vpwr scs8hd_diode_2
XFILLER_52_211 vgnd vpwr scs8hd_decap_3
XFILLER_16_27 vgnd vpwr scs8hd_decap_4
XFILLER_25_458 vgnd vpwr scs8hd_fill_1
XANTENNA__365__B _365_/B vgnd vpwr scs8hd_diode_2
XFILLER_33_480 vpwr vgnd scs8hd_fill_2
XFILLER_40_428 vgnd vpwr scs8hd_decap_3
XFILLER_20_141 vgnd vpwr scs8hd_decap_12
XFILLER_32_15 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_5_.latch_SLEEPB
+ _567_/Y vgnd vpwr scs8hd_diode_2
XANTENNA__381__A _226_/X vgnd vpwr scs8hd_diode_2
XFILLER_4_307 vpwr vgnd scs8hd_fill_2
XFILLER_4_329 vgnd vpwr scs8hd_decap_6
XANTENNA_ltile_clb_0.mux_fle_2_in_0.INVTX1_8_.scs8hd_inv_1_A top_width_0_height_0__pin_8_
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_1_in_0.mux_l1_in_2_.TGATE_3_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_1_in_0.INVTX1_11_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_1_in_0.LATCH_3_.latch/Q ltile_clb_0.mux_fle_1_in_0.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
Xltile_clb_0.mux_fle_3_in_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_3_in_0.INVTX1_6_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_3_in_0.LATCH_2_.latch/Q ltile_clb_0.mux_fle_3_in_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_6_.TGATE_1_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_13_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XANTENNA__259__C _286_/B vgnd vpwr scs8hd_diode_2
XANTENNA__556__A _556_/A vgnd vpwr scs8hd_diode_2
XFILLER_28_285 vpwr vgnd scs8hd_fill_2
XANTENNA__275__B _342_/A vgnd vpwr scs8hd_diode_2
XFILLER_43_277 vgnd vpwr scs8hd_decap_4
XFILLER_24_480 vgnd vpwr scs8hd_decap_4
XPHY_420 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_31_428 vgnd vpwr scs8hd_decap_6
XPHY_431 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_442 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_453 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_ltile_clb_0.mem_fle_0_in_3.LATCH_4_.latch_SLEEPB _488_/Y vgnd vpwr scs8hd_diode_2
XPHY_464 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_475 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_486 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_7_123 vgnd vpwr scs8hd_decap_12
XPHY_497 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__291__A _290_/X vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_0_.scs8hd_inv_1_A
+ ltile_clb_0.mux_fle_3_in_0.INVTX1_14_.scs8hd_inv_1/Y vgnd vpwr scs8hd_diode_2
XFILLER_3_373 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_0_in_2.mux_l1_in_3_.TGATE_2_.scs8hd_ebufn_2_A _642_/HI
+ vgnd vpwr scs8hd_diode_2
XFILLER_78_141 vgnd vpwr scs8hd_decap_12
XFILLER_81_306 vgnd vpwr scs8hd_decap_12
XFILLER_19_252 vpwr vgnd scs8hd_fill_2
XFILLER_19_263 vgnd vpwr scs8hd_decap_4
Xltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_3_.latch
+ data_in ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_3_.latch/Q
+ _569_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_34_222 vgnd vpwr scs8hd_decap_8
XFILLER_34_233 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.mux_fle_0_in_3.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_0_in_3.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ ltile_clb_0.mem_fle_0_in_3.LATCH_5_.latch/Q ltile_clb_0.mux_fle_0_in_3.INVTX1_14_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA__466__A _433_/A vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_3_in_1.INVTX1_5_.scs8hd_inv_1_A right_width_0_height_0__pin_5_
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_3_in_0.mux_l1_in_3_.TGATE_2_.scs8hd_ebufn_2_A _652_/HI
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_3_in_3.INVTX1_8_.scs8hd_inv_1 top_width_0_height_0__pin_8_ ltile_clb_0.mux_fle_3_in_3.INVTX1_8_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_ltile_clb_0.mux_fle_1_in_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_1_in_2.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_0_in_3.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_0_in_3.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_69_174 vpwr vgnd scs8hd_fill_2
XFILLER_57_358 vpwr vgnd scs8hd_fill_2
XFILLER_27_15 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mux_fle_2_in_3.INVTX1_13_.scs8hd_inv_1_A right_width_0_height_0__pin_13_
+ vgnd vpwr scs8hd_diode_2
XFILLER_27_59 vpwr vgnd scs8hd_fill_2
XANTENNA__376__A _392_/A vgnd vpwr scs8hd_diode_2
XFILLER_80_383 vpwr vgnd scs8hd_fill_2
XFILLER_13_439 vpwr vgnd scs8hd_fill_2
XANTENNA__526__D _526_/D vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_3_in_1.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_3_in_1.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_1_in_1.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_1_in_1.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
+ _606_/Y vgnd vpwr scs8hd_diode_2
XFILLER_68_44 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mem_fle_1_in_2.LATCH_4_.latch_SLEEPB _455_/Y vgnd vpwr scs8hd_diode_2
XFILLER_48_303 vgnd vpwr scs8hd_decap_3
X_654_ _654_/HI _654_/LO vgnd vpwr scs8hd_conb_1
XFILLER_63_306 vpwr vgnd scs8hd_fill_2
XFILLER_56_380 vgnd vpwr scs8hd_decap_4
XFILLER_16_211 vgnd vpwr scs8hd_decap_3
XANTENNA__286__A _286_/A vgnd vpwr scs8hd_diode_2
X_585_ _559_/A _585_/B _585_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_2_.TGATE_1_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_5_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_16_266 vgnd vpwr scs8hd_decap_8
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_15_.latch_D
+ data_in vgnd vpwr scs8hd_diode_2
XFILLER_31_225 vpwr vgnd scs8hd_fill_2
XPHY_261 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_250 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_31_236 vpwr vgnd scs8hd_fill_2
XFILLER_12_472 vgnd vpwr scs8hd_decap_12
XFILLER_12_450 vpwr vgnd scs8hd_fill_2
XPHY_272 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_283 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_294 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_79_461 vgnd vpwr scs8hd_decap_4
XFILLER_79_472 vgnd vpwr scs8hd_decap_12
XFILLER_66_133 vgnd vpwr scs8hd_decap_12
XFILLER_39_347 vpwr vgnd scs8hd_fill_2
XFILLER_39_358 vgnd vpwr scs8hd_decap_3
XFILLER_66_177 vgnd vpwr scs8hd_decap_6
XFILLER_81_147 vgnd vpwr scs8hd_decap_12
XANTENNA__346__D _346_/D vgnd vpwr scs8hd_diode_2
Xltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_0_.scs8hd_inv_1
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_0_.latch/Q
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_13_39 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.mux_fle_2_in_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_2_in_1.INVTX1_6_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_2_in_1.LATCH_2_.latch/Q ltile_clb_0.mux_fle_2_in_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
Xltile_clb_0.mux_fle_0_in_1.mux_l1_in_2_.TGATE_3_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_0_in_1.INVTX1_11_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_0_in_1.LATCH_3_.latch/Q ltile_clb_0.mux_fle_0_in_1.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_45_339 vgnd vpwr scs8hd_decap_4
X_370_ _370_/A _379_/B vgnd vpwr scs8hd_buf_1
XFILLER_54_68 vgnd vpwr scs8hd_decap_12
XFILLER_13_236 vpwr vgnd scs8hd_fill_2
XFILLER_70_56 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mem_fle_2_in_1.LATCH_4_.latch_SLEEPB _418_/Y vgnd vpwr scs8hd_diode_2
XANTENNA__553__B _552_/X vgnd vpwr scs8hd_diode_2
XFILLER_5_402 vpwr vgnd scs8hd_fill_2
XFILLER_5_457 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_0_in_1.INVTX1_3_.scs8hd_inv_1_A left_width_0_height_0__pin_3_
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_0_in_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_0_in_0.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_3_.latch
+ data_in ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_3_.latch/Q
+ _543_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_79_98 vgnd vpwr scs8hd_decap_12
XFILLER_28_80 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_10_.latch_SLEEPB
+ _587_/Y vgnd vpwr scs8hd_diode_2
X_637_ _637_/HI _637_/LO vgnd vpwr scs8hd_conb_1
X_568_ _542_/A _564_/B _568_/Y vgnd vpwr scs8hd_nor2_4
X_499_ _331_/A _495_/X _499_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA__463__B _462_/X vgnd vpwr scs8hd_diode_2
XFILLER_12_291 vpwr vgnd scs8hd_fill_2
XFILLER_67_3 vgnd vpwr scs8hd_decap_12
XFILLER_5_62 vgnd vpwr scs8hd_decap_12
XFILLER_5_51 vgnd vpwr scs8hd_decap_8
XANTENNA_ltile_clb_0.mux_fle_0_in_3.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_0_in_3.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_0_in_2.INVTX1_12_.scs8hd_inv_1_A top_width_0_height_0__pin_12_
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_82_478 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mux_fle_1_in_2.INVTX1_0_.scs8hd_inv_1_A top_width_0_height_0__pin_0_
+ vgnd vpwr scs8hd_diode_2
XFILLER_42_309 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_3_in_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_3_in_3.LATCH_4_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_62_191 vgnd vpwr scs8hd_decap_4
XFILLER_24_27 vgnd vpwr scs8hd_decap_4
XANTENNA_ltile_clb_0.mux_fle_3_in_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_3_in_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XANTENNA__373__B _377_/B vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_0_in_0.INVTX1_4_.scs8hd_inv_1 top_width_0_height_0__pin_4_ ltile_clb_0.mux_fle_0_in_0.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_40_15 vgnd vpwr scs8hd_decap_12
XFILLER_2_438 vgnd vpwr scs8hd_fill_1
XFILLER_58_442 vgnd vpwr scs8hd_decap_6
XFILLER_58_431 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mem_fle_3_in_0.LATCH_4_.latch_SLEEPB _375_/Y vgnd vpwr scs8hd_diode_2
XFILLER_58_475 vgnd vpwr scs8hd_decap_8
Xltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_5_.scs8hd_inv_1
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_5_.latch/Q
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_73_423 vpwr vgnd scs8hd_fill_2
XFILLER_58_486 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_3_.TGATE_0_.scs8hd_ebufn_2_TEB
+ _615_/Y vgnd vpwr scs8hd_diode_2
XFILLER_73_456 vgnd vpwr scs8hd_decap_3
XFILLER_45_169 vgnd vpwr scs8hd_decap_4
XFILLER_73_489 vgnd vpwr scs8hd_decap_12
X_422_ _435_/A _412_/B _422_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_60_117 vgnd vpwr scs8hd_decap_12
XFILLER_26_383 vgnd vpwr scs8hd_fill_1
XANTENNA__564__A _564_/A vgnd vpwr scs8hd_diode_2
XFILLER_26_394 vgnd vpwr scs8hd_decap_3
X_353_ _392_/A _353_/B _353_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA__283__B _324_/A vgnd vpwr scs8hd_diode_2
X_284_ _284_/A _540_/A vgnd vpwr scs8hd_buf_1
XFILLER_14_93 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_1_.TGATE_1_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_1_.TGATE_1_.scs8hd_ebufn_2/A
+ _614_/Y ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
Xltile_clb_0.mem_fle_0_in_1.LATCH_5_.latch data_in ltile_clb_0.mem_fle_0_in_1.LATCH_5_.latch/Q
+ _509_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_5_254 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_2_in_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_2_in_1.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_14_.scs8hd_inv_1_A
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_14_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_1_460 vpwr vgnd scs8hd_fill_2
XFILLER_76_261 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.mem_fle_1_in_1.LATCH_4_.latch data_in ltile_clb_0.mem_fle_1_in_1.LATCH_4_.latch/Q
+ _466_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_76_283 vpwr vgnd scs8hd_fill_2
XANTENNA__458__B _450_/X vgnd vpwr scs8hd_diode_2
XFILLER_64_478 vgnd vpwr scs8hd_decap_8
XFILLER_64_467 vpwr vgnd scs8hd_fill_2
XFILLER_17_361 vgnd vpwr scs8hd_decap_3
XANTENNA__474__A _430_/A vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mem_fle_0_in_1.LATCH_5_.latch_SLEEPB _509_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_0_in_3.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_0_in_3.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_1_in_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_1_in_0.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mem_fle_2_in_1.LATCH_3_.latch data_in ltile_clb_0.mem_fle_2_in_1.LATCH_3_.latch/Q
+ _420_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
Xltile_clb_0.mux_fle_1_in_2.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_1_in_2.INVTX1_6_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_1_in_2.LATCH_2_.latch/Q ltile_clb_0.mux_fle_1_in_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
Xltile_clb_0.mux_fle_3_in_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_3_in_2.INVTX1_1_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_3_in_2.LATCH_1_.latch/Q ltile_clb_0.mux_fle_3_in_2.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
Xltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
+ _637_/HI ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.mem_ble4_out_0.LATCH_2_.latch/Q
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_19_27 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.mem_fle_3_in_1.LATCH_2_.latch data_in ltile_clb_0.mem_fle_3_in_1.LATCH_2_.latch/Q
+ _366_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_67_283 vgnd vpwr scs8hd_decap_3
XFILLER_55_423 vpwr vgnd scs8hd_fill_2
XFILLER_55_412 vpwr vgnd scs8hd_fill_2
XANTENNA__368__B _368_/B vgnd vpwr scs8hd_diode_2
XFILLER_82_242 vgnd vpwr scs8hd_decap_6
XFILLER_27_147 vgnd vpwr scs8hd_decap_12
XFILLER_35_15 vgnd vpwr scs8hd_decap_12
XFILLER_42_117 vgnd vpwr scs8hd_decap_12
XPHY_827 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_816 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_805 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__384__A _384_/A vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_2_.TGATE_1_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_2_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_35_59 vpwr vgnd scs8hd_fill_2
XFILLER_35_191 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.mux_fle_0_in_1.INVTX1_8_.scs8hd_inv_1 top_width_0_height_0__pin_8_ ltile_clb_0.mux_fle_0_in_1.INVTX1_8_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XPHY_838 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_11_515 vgnd vpwr scs8hd_fill_1
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
+ _620_/Y vgnd vpwr scs8hd_diode_2
XFILLER_2_202 vgnd vpwr scs8hd_decap_12
XFILLER_78_504 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_5_.TGATE_0_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_10_.scs8hd_inv_1/Y
+ _629_/Y ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_5_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_76_44 vgnd vpwr scs8hd_decap_12
XFILLER_65_209 vpwr vgnd scs8hd_fill_2
XANTENNA__559__A _559_/A vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_0_in_0.INVTX1_11_.scs8hd_inv_1 left_width_0_height_0__pin_11_
+ ltile_clb_0.mux_fle_0_in_0.INVTX1_11_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XFILLER_58_272 vgnd vpwr scs8hd_decap_3
XANTENNA_ltile_clb_0.mux_fle_2_in_1.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_2_in_1.LATCH_6_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_3_in_0.INVTX1_10_.scs8hd_inv_1 bottom_width_0_height_0__pin_10_
+ ltile_clb_0.mux_fle_3_in_0.INVTX1_10_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XFILLER_73_286 vpwr vgnd scs8hd_fill_2
XFILLER_73_297 vpwr vgnd scs8hd_fill_2
X_405_ _394_/A _398_/A _405_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_14_364 vgnd vpwr scs8hd_decap_3
XANTENNA__294__A _293_/X vgnd vpwr scs8hd_diode_2
XPHY_70 vgnd vpwr scs8hd_decap_3
XPHY_81 vgnd vpwr scs8hd_decap_3
XPHY_92 vgnd vpwr scs8hd_decap_3
X_336_ _263_/X _421_/A vgnd vpwr scs8hd_buf_1
X_267_ _304_/A _267_/X vgnd vpwr scs8hd_buf_1
Xltile_clb_0.mem_fle_1_in_3.LATCH_7_.latch data_in ltile_clb_0.mem_fle_1_in_3.LATCH_7_.latch/Q
+ _441_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA__460__C _384_/A vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mem_fle_1_in_0.LATCH_5_.latch_SLEEPB _476_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_2_in_1.mux_l1_in_3_.TGATE_2_.scs8hd_ebufn_2_A _649_/HI
+ vgnd vpwr scs8hd_diode_2
XANTENNA__469__A _436_/A vgnd vpwr scs8hd_diode_2
XFILLER_49_250 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.mem_fle_2_in_3.LATCH_6_.latch data_in ltile_clb_0.mem_fle_2_in_3.LATCH_6_.latch/Q
+ _389_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_37_412 vpwr vgnd scs8hd_fill_2
XFILLER_37_423 vgnd vpwr scs8hd_decap_4
XFILLER_37_434 vgnd vpwr scs8hd_decap_3
XFILLER_24_117 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.buf4_3_.scs8hd_buf_1
+ ltile_clb_0.mux_fle_0_in_3.INVTX1_14_.scs8hd_inv_1/Y _634_/A vgnd vpwr scs8hd_buf_1
Xltile_clb_0.mux_fle_0_in_1.INVTX1_13_.scs8hd_inv_1 right_width_0_height_0__pin_13_
+ ltile_clb_0.mux_fle_0_in_1.INVTX1_13_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
Xltile_clb_0.mux_fle_1_in_2.INVTX1_3_.scs8hd_inv_1 left_width_0_height_0__pin_3_ ltile_clb_0.mux_fle_1_in_2.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
Xltile_clb_0.mem_fle_3_in_3.LATCH_5_.latch data_in ltile_clb_0.mem_fle_3_in_3.LATCH_5_.latch/Q
+ _329_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
Xltile_clb_0.mux_fle_3_in_1.INVTX1_12_.scs8hd_inv_1 top_width_0_height_0__pin_12_
+ ltile_clb_0.mux_fle_3_in_1.INVTX1_12_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XFILLER_32_194 vgnd vpwr scs8hd_decap_4
XFILLER_21_39 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_11_.latch_D
+ data_in vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_1_in_1.INVTX1_9_.scs8hd_inv_1_A right_width_0_height_0__pin_9_
+ vgnd vpwr scs8hd_diode_2
XANTENNA__379__A _379_/A vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_2_in_2.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_2_in_2.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_28_401 vgnd vpwr scs8hd_decap_8
XANTENNA_ltile_clb_0.mux_fle_1_in_3.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_1_in_3.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_55_242 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.mux_fle_1_in_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_1_in_0.INVTX1_0_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_1_in_0.LATCH_0_.latch/Q ltile_clb_0.mux_fle_1_in_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_43_426 vgnd vpwr scs8hd_fill_1
XANTENNA_ltile_clb_0.mux_fle_2_in_1.INVTX1_10_.scs8hd_inv_1_A bottom_width_0_height_0__pin_10_
+ vgnd vpwr scs8hd_diode_2
XPHY_602 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_70_267 vgnd vpwr scs8hd_decap_8
XPHY_635 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_624 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_613 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_62_68 vgnd vpwr scs8hd_decap_12
XPHY_668 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_657 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_646 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_11_301 vpwr vgnd scs8hd_fill_2
XPHY_679 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_7_316 vpwr vgnd scs8hd_fill_2
XANTENNA__561__B _558_/B vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_3_in_2.INVTX1_14_.scs8hd_inv_1 ltile_clb_0.mux_fle_3_in_2.INVTX1_14_.scs8hd_inv_1/A
+ ltile_clb_0.mux_fle_3_in_2.INVTX1_14_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XANTENNA__289__A _267_/X vgnd vpwr scs8hd_diode_2
XFILLER_78_389 vgnd vpwr scs8hd_decap_8
XFILLER_19_423 vpwr vgnd scs8hd_fill_2
XFILLER_34_459 vgnd vpwr scs8hd_decap_6
XFILLER_36_80 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.mux_fle_0_in_3.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_0_in_3.INVTX1_6_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_0_in_3.LATCH_2_.latch/Q ltile_clb_0.mux_fle_0_in_3.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
Xltile_clb_0.mux_fle_2_in_3.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_2_in_3.INVTX1_1_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_2_in_3.LATCH_1_.latch/Q ltile_clb_0.mux_fle_2_in_3.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_ltile_clb_0.mux_fle_2_in_2.INVTX1_6_.scs8hd_inv_1_A bottom_width_0_height_0__pin_6_
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_3_in_0.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_3_in_0.INVTX1_12_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_3_in_0.LATCH_0_.latch/Q ltile_clb_0.mux_fle_3_in_0.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_42_492 vgnd vpwr scs8hd_decap_4
X_319_ _526_/D _358_/D vgnd vpwr scs8hd_buf_1
XANTENNA__471__B _226_/X vgnd vpwr scs8hd_diode_2
XFILLER_69_367 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.mux_fle_1_in_3.INVTX1_7_.scs8hd_inv_1 left_width_0_height_0__pin_7_ ltile_clb_0.mux_fle_1_in_3.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_25_437 vpwr vgnd scs8hd_fill_2
XFILLER_52_256 vgnd vpwr scs8hd_decap_3
XFILLER_32_27 vgnd vpwr scs8hd_decap_4
XFILLER_20_197 vgnd vpwr scs8hd_fill_1
XANTENNA_ltile_clb_0.mux_fle_3_in_3.INVTX1_3_.scs8hd_inv_1_A left_width_0_height_0__pin_3_
+ vgnd vpwr scs8hd_diode_2
XFILLER_75_315 vpwr vgnd scs8hd_fill_2
XFILLER_75_348 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2_TEB
+ _629_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_0_in_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_0_in_2.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__556__B _558_/B vgnd vpwr scs8hd_diode_2
XFILLER_16_426 vpwr vgnd scs8hd_fill_2
XFILLER_16_448 vgnd vpwr scs8hd_decap_8
XFILLER_28_297 vgnd vpwr scs8hd_decap_8
XFILLER_16_459 vgnd vpwr scs8hd_decap_4
XPHY_410 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_31_407 vgnd vpwr scs8hd_decap_3
XFILLER_43_256 vgnd vpwr scs8hd_fill_1
XPHY_421 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_432 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_443 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l4_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
+ _611_/Y vgnd vpwr scs8hd_diode_2
XPHY_454 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_465 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_476 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__572__A _546_/A vgnd vpwr scs8hd_diode_2
XPHY_487 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_498 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_7_135 vgnd vpwr scs8hd_decap_12
Xclkbuf_1_0_0_clk clkbuf_0_clk/X clkbuf_1_0_0_clk/X vgnd vpwr scs8hd_clkbuf_1
XFILLER_22_93 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.tap_buf4_0_.scs8hd_inv_1_A
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_3_352 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_0_in_1.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_0_in_1.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_3_396 vgnd vpwr scs8hd_fill_1
XFILLER_66_348 vgnd vpwr scs8hd_decap_6
XFILLER_81_318 vgnd vpwr scs8hd_decap_12
XFILLER_74_381 vgnd vpwr scs8hd_fill_1
XFILLER_19_297 vpwr vgnd scs8hd_fill_2
XANTENNA__466__B _462_/X vgnd vpwr scs8hd_diode_2
XFILLER_34_267 vgnd vpwr scs8hd_decap_8
Xltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_4_.scs8hd_inv_1/Y
+ _605_/Y ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA__482__A _380_/X vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_2_in_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_2_in_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ ltile_clb_0.mem_fle_2_in_0.LATCH_5_.latch/Q ltile_clb_0.mux_fle_2_in_0.INVTX1_14_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_30_484 vgnd vpwr scs8hd_decap_8
XFILLER_6_190 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mux_fle_2_in_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_2_in_2.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_1_in_0.INVTX1_14_.scs8hd_inv_1_A ltile_clb_0.mux_fle_1_in_0.INVTX1_14_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_57_326 vgnd vpwr scs8hd_fill_1
Xltile_clb_0.mux_fle_0_in_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_0_in_1.INVTX1_0_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_0_in_1.LATCH_0_.latch/Q ltile_clb_0.mux_fle_0_in_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_27_27 vgnd vpwr scs8hd_decap_12
XANTENNA__376__B _377_/B vgnd vpwr scs8hd_diode_2
XFILLER_25_267 vgnd vpwr scs8hd_decap_4
XFILLER_13_418 vgnd vpwr scs8hd_decap_6
XFILLER_40_215 vgnd vpwr scs8hd_decap_8
XFILLER_43_15 vgnd vpwr scs8hd_decap_12
XFILLER_40_237 vgnd vpwr scs8hd_decap_4
XFILLER_43_59 vpwr vgnd scs8hd_fill_2
XANTENNA__392__A _392_/A vgnd vpwr scs8hd_diode_2
XFILLER_21_484 vgnd vpwr scs8hd_decap_4
XFILLER_21_495 vpwr vgnd scs8hd_fill_2
XFILLER_4_105 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.mux_fle_3_in_0.INVTX1_4_.scs8hd_inv_1 top_width_0_height_0__pin_4_ ltile_clb_0.mux_fle_3_in_0.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
Xltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_6_.TGATE_1_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_13_.scs8hd_inv_1/Y
+ _604_/Y ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_3_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
Xltile_clb_0.mux_fle_3_in_3.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_3_in_3.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2/Z
+ ltile_clb_0.mem_fle_3_in_3.LATCH_6_.latch/Q ltile_clb_0.mux_fle_3_in_3.INVTX1_14_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
Xltile_clb_0.mux_fle_2_in_3.INVTX1_10_.scs8hd_inv_1 bottom_width_0_height_0__pin_10_
+ ltile_clb_0.mux_fle_2_in_3.INVTX1_10_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XFILLER_68_56 vgnd vpwr scs8hd_decap_12
XFILLER_0_366 vgnd vpwr scs8hd_decap_4
XFILLER_0_388 vgnd vpwr scs8hd_decap_4
XFILLER_75_123 vgnd vpwr scs8hd_decap_12
XFILLER_0_399 vpwr vgnd scs8hd_fill_2
XANTENNA__567__A _541_/A vgnd vpwr scs8hd_diode_2
X_653_ _653_/HI _653_/LO vgnd vpwr scs8hd_conb_1
XFILLER_56_370 vgnd vpwr scs8hd_fill_1
XANTENNA__286__B _286_/B vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_2_in_1.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_2_in_1.INVTX1_12_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_2_in_1.LATCH_0_.latch/Q ltile_clb_0.mux_fle_2_in_1.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
X_584_ _250_/X _585_/B _584_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_16_234 vgnd vpwr scs8hd_decap_3
XFILLER_16_245 vpwr vgnd scs8hd_fill_2
XFILLER_71_362 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_1_in_2.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_1_in_2.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XPHY_251 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_240 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_273 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_262 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_284 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_295 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_3_171 vgnd vpwr scs8hd_decap_12
XFILLER_79_484 vgnd vpwr scs8hd_decap_4
XFILLER_39_315 vpwr vgnd scs8hd_fill_2
XFILLER_39_326 vpwr vgnd scs8hd_fill_2
XFILLER_66_145 vgnd vpwr scs8hd_decap_3
XFILLER_12_3 vgnd vpwr scs8hd_decap_12
XFILLER_54_318 vpwr vgnd scs8hd_fill_2
XANTENNA__477__A _433_/A vgnd vpwr scs8hd_diode_2
XFILLER_54_329 vgnd vpwr scs8hd_fill_1
XFILLER_81_159 vgnd vpwr scs8hd_decap_12
XFILLER_62_362 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mux_fle_0_in_3.INVTX1_1_.scs8hd_inv_1_A right_width_0_height_0__pin_1_
+ vgnd vpwr scs8hd_diode_2
XFILLER_50_513 vgnd vpwr scs8hd_decap_3
XANTENNA_ltile_clb_0.mux_fle_1_in_1.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_1_in_1.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mem_fle_0_in_0.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
+ _607_/Y vgnd vpwr scs8hd_diode_2
XFILLER_30_292 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.mem_fle_0_in_2.LATCH_1_.latch data_in ltile_clb_0.mem_fle_0_in_2.LATCH_1_.latch/Q
+ _502_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_38_15 vgnd vpwr scs8hd_decap_12
XFILLER_57_123 vgnd vpwr scs8hd_decap_12
XANTENNA__387__A _387_/A vgnd vpwr scs8hd_diode_2
XFILLER_57_167 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.mem_fle_1_in_2.LATCH_0_.latch data_in ltile_clb_0.mem_fle_1_in_2.LATCH_0_.latch/Q
+ _459_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_72_159 vpwr vgnd scs8hd_fill_2
XFILLER_53_340 vpwr vgnd scs8hd_fill_2
XFILLER_38_392 vgnd vpwr scs8hd_decap_4
XFILLER_53_384 vpwr vgnd scs8hd_fill_2
XFILLER_53_362 vgnd vpwr scs8hd_fill_1
XFILLER_13_204 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.mux_fle_3_in_1.INVTX1_8_.scs8hd_inv_1 top_width_0_height_0__pin_8_ ltile_clb_0.mux_fle_3_in_1.INVTX1_8_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_13_259 vgnd vpwr scs8hd_decap_6
XFILLER_70_68 vgnd vpwr scs8hd_decap_12
XFILLER_21_270 vgnd vpwr scs8hd_decap_3
XANTENNA_ltile_clb_0.mux_fle_2_in_3.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_2_in_3.LATCH_5_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_21_292 vgnd vpwr scs8hd_decap_4
Xltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_11_.latch
+ data_in ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_11_.latch/Q
+ _534_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_76_443 vgnd vpwr scs8hd_decap_4
XFILLER_48_134 vpwr vgnd scs8hd_fill_2
XFILLER_76_454 vgnd vpwr scs8hd_decap_4
XANTENNA__297__A _296_/X vgnd vpwr scs8hd_diode_2
XFILLER_48_145 vgnd vpwr scs8hd_decap_4
XFILLER_48_189 vpwr vgnd scs8hd_fill_2
X_636_ _636_/HI _636_/LO vgnd vpwr scs8hd_conb_1
XFILLER_29_392 vpwr vgnd scs8hd_fill_2
X_567_ _541_/A _564_/B _567_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_71_192 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.mux_fle_1_in_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_1_in_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ ltile_clb_0.mem_fle_1_in_1.LATCH_5_.latch/Q ltile_clb_0.mux_fle_1_in_1.INVTX1_14_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_44_80 vgnd vpwr scs8hd_decap_12
X_498_ _328_/A _495_/X _498_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_12_270 vgnd vpwr scs8hd_decap_3
XANTENNA_ltile_clb_0.mux_fle_1_in_2.mux_l1_in_3_.TGATE_2_.scs8hd_ebufn_2_A _646_/HI
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_1_.latch_D
+ data_in vgnd vpwr scs8hd_diode_2
XFILLER_5_74 vgnd vpwr scs8hd_decap_12
XFILLER_67_443 vgnd vpwr scs8hd_decap_4
XFILLER_67_432 vpwr vgnd scs8hd_fill_2
XFILLER_39_123 vgnd vpwr scs8hd_decap_12
XFILLER_67_487 vgnd vpwr scs8hd_fill_1
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_35_340 vpwr vgnd scs8hd_fill_2
XFILLER_35_362 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.buf4_1_.scs8hd_buf_1
+ ltile_clb_0.mux_fle_3_in_1.INVTX1_14_.scs8hd_inv_1/Y _606_/A vgnd vpwr scs8hd_buf_1
XFILLER_50_321 vpwr vgnd scs8hd_fill_2
XFILLER_50_332 vpwr vgnd scs8hd_fill_2
XFILLER_50_398 vpwr vgnd scs8hd_fill_2
XFILLER_40_27 vgnd vpwr scs8hd_decap_4
XANTENNA_ltile_clb_0.mux_fle_1_in_3.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_1_in_3.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_0_in_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_0_in_0.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_2_417 vgnd vpwr scs8hd_decap_4
XFILLER_58_421 vgnd vpwr scs8hd_fill_1
XFILLER_58_498 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.mux_fle_1_in_2.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_1_in_2.INVTX1_12_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_1_in_2.LATCH_0_.latch/Q ltile_clb_0.mux_fle_1_in_2.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_6_.scs8hd_inv_1_A
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_6_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_26_362 vgnd vpwr scs8hd_decap_4
X_421_ _421_/A _435_/A vgnd vpwr scs8hd_buf_1
X_352_ _391_/A _353_/B _352_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_60_129 vpwr vgnd scs8hd_fill_2
XFILLER_53_170 vgnd vpwr scs8hd_fill_1
XANTENNA__564__B _564_/B vgnd vpwr scs8hd_diode_2
XFILLER_41_310 vpwr vgnd scs8hd_fill_2
XFILLER_41_376 vpwr vgnd scs8hd_fill_2
X_283_ _278_/X _324_/A _284_/A vgnd vpwr scs8hd_or2_4
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
+ _625_/Y vgnd vpwr scs8hd_diode_2
XANTENNA__580__A _579_/X vgnd vpwr scs8hd_diode_2
XFILLER_5_288 vpwr vgnd scs8hd_fill_2
XFILLER_30_93 vgnd vpwr scs8hd_decap_12
XFILLER_49_410 vpwr vgnd scs8hd_fill_2
XFILLER_49_443 vpwr vgnd scs8hd_fill_2
XFILLER_49_465 vgnd vpwr scs8hd_decap_4
XFILLER_64_402 vpwr vgnd scs8hd_fill_2
X_619_ _619_/A _619_/Y vgnd vpwr scs8hd_inv_8
XFILLER_32_310 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_1_in_1.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_1_in_1.LATCH_7_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__474__B _479_/B vgnd vpwr scs8hd_diode_2
XFILLER_20_505 vgnd vpwr scs8hd_decap_8
XFILLER_32_365 vpwr vgnd scs8hd_fill_2
XFILLER_32_398 vgnd vpwr scs8hd_decap_6
XANTENNA__490__A _421_/A vgnd vpwr scs8hd_diode_2
XFILLER_19_39 vgnd vpwr scs8hd_decap_12
XFILLER_67_273 vgnd vpwr scs8hd_decap_4
XFILLER_27_159 vgnd vpwr scs8hd_decap_8
XFILLER_55_479 vpwr vgnd scs8hd_fill_2
XFILLER_35_27 vgnd vpwr scs8hd_decap_12
XPHY_817 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_806 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_70_438 vgnd vpwr scs8hd_fill_1
XFILLER_23_332 vgnd vpwr scs8hd_decap_4
XFILLER_42_129 vgnd vpwr scs8hd_decap_12
XPHY_839 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_828 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mem_fle_0_in_2.LATCH_7_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_16_.scs8hd_inv_1_A
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_16_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_23_376 vpwr vgnd scs8hd_fill_2
XFILLER_23_398 vpwr vgnd scs8hd_fill_2
XFILLER_50_173 vpwr vgnd scs8hd_fill_2
XFILLER_51_15 vgnd vpwr scs8hd_decap_12
XFILLER_50_195 vgnd vpwr scs8hd_decap_8
XFILLER_51_59 vpwr vgnd scs8hd_fill_2
XFILLER_2_225 vgnd vpwr scs8hd_fill_1
XFILLER_76_56 vgnd vpwr scs8hd_decap_12
XFILLER_58_251 vgnd vpwr scs8hd_decap_4
XANTENNA__559__B _558_/B vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mem_fle_0_in_3.LATCH_5_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_46_402 vgnd vpwr scs8hd_fill_1
XFILLER_73_243 vgnd vpwr scs8hd_fill_1
Xltile_clb_0.mux_fle_0_in_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_0_in_2.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ ltile_clb_0.mem_fle_0_in_2.LATCH_5_.latch/Q ltile_clb_0.mux_fle_0_in_2.INVTX1_14_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA__575__A _575_/A vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_0_in_3.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_0_in_3.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_61_449 vgnd vpwr scs8hd_decap_8
Xltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_3_.TGATE_1_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_7_.TGATE_1_.scs8hd_ebufn_2/Z
+ _622_/Y ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_3_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
X_404_ _338_/A _399_/B _404_/Y vgnd vpwr scs8hd_nor2_4
XPHY_60 vgnd vpwr scs8hd_decap_3
XPHY_71 vgnd vpwr scs8hd_decap_3
XPHY_82 vgnd vpwr scs8hd_decap_3
X_335_ _392_/A _338_/B _335_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_14_376 vgnd vpwr scs8hd_decap_4
XFILLER_14_387 vgnd vpwr scs8hd_decap_8
XFILLER_14_398 vpwr vgnd scs8hd_fill_2
XFILLER_41_184 vgnd vpwr scs8hd_decap_3
XPHY_93 vgnd vpwr scs8hd_decap_3
XANTENNA_ltile_clb_0.mux_fle_1_in_3.INVTX1_7_.scs8hd_inv_1_A left_width_0_height_0__pin_7_
+ vgnd vpwr scs8hd_diode_2
X_266_ _248_/A _535_/A _266_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_1_.latch_SLEEPB
+ _545_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mem_fle_1_in_0.LATCH_7_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA__460__D _358_/D vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_2_in_0.INVTX1_3_.scs8hd_inv_1_A left_width_0_height_0__pin_3_
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_7_.TGATE_1_.scs8hd_ebufn_2_TEB
+ _628_/Y vgnd vpwr scs8hd_diode_2
XANTENNA__469__B _461_/X vgnd vpwr scs8hd_diode_2
XFILLER_49_240 vpwr vgnd scs8hd_fill_2
XFILLER_49_262 vgnd vpwr scs8hd_decap_4
XANTENNA__485__A _314_/A vgnd vpwr scs8hd_diode_2
XFILLER_37_468 vgnd vpwr scs8hd_decap_4
XFILLER_37_479 vpwr vgnd scs8hd_fill_2
XFILLER_64_287 vgnd vpwr scs8hd_fill_1
XFILLER_24_129 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mem_fle_1_in_1.LATCH_5_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_32_173 vgnd vpwr scs8hd_decap_6
XFILLER_20_335 vgnd vpwr scs8hd_fill_1
XFILLER_20_357 vgnd vpwr scs8hd_decap_4
XANTENNA_ltile_clb_0.mux_fle_1_in_3.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_1_in_3.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
+ _621_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l4_in_0_.TGATE_0_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mem_fle_1_in_2.LATCH_3_.latch_D data_in vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_0_in_3.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_0_in_3.INVTX1_12_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_0_in_3.LATCH_0_.latch/Q ltile_clb_0.mux_fle_0_in_3.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA__379__B _379_/B vgnd vpwr scs8hd_diode_2
XFILLER_28_424 vgnd vpwr scs8hd_decap_4
XFILLER_46_15 vgnd vpwr scs8hd_decap_12
XFILLER_55_232 vpwr vgnd scs8hd_fill_2
XANTENNA__395__A _379_/A vgnd vpwr scs8hd_diode_2
XFILLER_43_416 vpwr vgnd scs8hd_fill_2
XFILLER_70_213 vgnd vpwr scs8hd_fill_1
XANTENNA_ltile_clb_0.mux_fle_3_in_1.INVTX1_0_.scs8hd_inv_1_A top_width_0_height_0__pin_0_
+ vgnd vpwr scs8hd_diode_2
XPHY_625 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_614 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_603 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_669 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_658 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_647 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_636 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_ltile_clb_0.mem_fle_1_in_3.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_51_493 vpwr vgnd scs8hd_fill_2
XFILLER_11_324 vpwr vgnd scs8hd_fill_2
XFILLER_23_184 vpwr vgnd scs8hd_fill_2
XFILLER_7_339 vgnd vpwr scs8hd_decap_3
XFILLER_11_51 vgnd vpwr scs8hd_decap_8
XFILLER_3_501 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_8_.scs8hd_inv_1
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_8_.latch/Q
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_8_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_11_62 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_8_.scs8hd_inv_1_A
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_8_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_78_335 vgnd vpwr scs8hd_fill_1
XFILLER_78_346 vgnd vpwr scs8hd_decap_8
XANTENNA__289__B _541_/A vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_0_in_3.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_0_in_3.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_3_in_3.INVTX1_13_.scs8hd_inv_1_A right_width_0_height_0__pin_13_
+ vgnd vpwr scs8hd_diode_2
XFILLER_19_402 vgnd vpwr scs8hd_decap_4
XANTENNA_ltile_clb_0.mem_fle_2_in_0.LATCH_3_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_46_232 vgnd vpwr scs8hd_fill_1
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_34_449 vgnd vpwr scs8hd_decap_8
XANTENNA_ltile_clb_0.mux_fle_3_in_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_3_in_1.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_52_80 vgnd vpwr scs8hd_decap_12
X_318_ enable address[5] _526_/D vgnd vpwr scs8hd_nand2_4
XANTENNA__471__C _384_/A vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_7_.latch_D
+ data_in vgnd vpwr scs8hd_diode_2
X_249_ _246_/A _286_/A _286_/B address[1] _250_/A vgnd vpwr scs8hd_or4_4
Xltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l4_in_0_.TGATE_1_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l4_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ _618_/Y ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_16_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
Xltile_clb_0.mux_fle_0_in_0.mux_l1_in_2_.TGATE_3_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_0_in_0.INVTX1_11_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_0_in_0.LATCH_3_.latch/Q ltile_clb_0.mux_fle_0_in_0.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
Xltile_clb_0.mux_fle_2_in_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_2_in_0.INVTX1_6_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_2_in_0.LATCH_2_.latch/Q ltile_clb_0.mux_fle_2_in_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_ltile_clb_0.mem_fle_2_in_1.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_42_3 vgnd vpwr scs8hd_decap_12
XFILLER_69_379 vpwr vgnd scs8hd_fill_2
XFILLER_25_416 vpwr vgnd scs8hd_fill_2
XFILLER_37_276 vpwr vgnd scs8hd_fill_2
XFILLER_52_224 vgnd vpwr scs8hd_decap_12
XFILLER_20_154 vgnd vpwr scs8hd_decap_8
Xltile_clb_0.mux_fle_3_in_3.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_3_in_3.INVTX1_7_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_3_in_3.LATCH_3_.latch/Q ltile_clb_0.mux_fle_3_in_3.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_0_515 vgnd vpwr scs8hd_fill_1
XFILLER_68_390 vgnd vpwr scs8hd_decap_6
Xltile_clb_0.mux_fle_1_in_0.INVTX1_3_.scs8hd_inv_1 left_width_0_height_0__pin_3_ ltile_clb_0.mux_fle_1_in_0.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_16_416 vgnd vpwr scs8hd_decap_8
XPHY_400 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_43_235 vpwr vgnd scs8hd_fill_2
XPHY_411 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_422 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_31_419 vpwr vgnd scs8hd_fill_2
XPHY_433 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_444 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_11_110 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_9_.latch
+ data_in ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_9_.latch/Q
+ _273_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XPHY_455 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_466 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_477 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_ltile_clb_0.mem_fle_0_in_0.LATCH_0_.latch_SLEEPB _525_/Y vgnd vpwr scs8hd_diode_2
XANTENNA__572__B _554_/X vgnd vpwr scs8hd_diode_2
XPHY_488 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_499 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_7_147 vgnd vpwr scs8hd_decap_12
XFILLER_39_508 vgnd vpwr scs8hd_decap_8
XFILLER_78_154 vgnd vpwr scs8hd_decap_12
XFILLER_34_213 vgnd vpwr scs8hd_fill_1
XANTENNA_ltile_clb_0.mux_fle_0_in_3.mux_l1_in_3_.TGATE_2_.scs8hd_ebufn_2_A _643_/HI
+ vgnd vpwr scs8hd_diode_2
XFILLER_34_279 vgnd vpwr scs8hd_decap_8
XFILLER_30_430 vgnd vpwr scs8hd_fill_1
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_30_463 vgnd vpwr scs8hd_fill_1
XANTENNA__482__B _427_/B vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_3_in_1.mux_l1_in_3_.TGATE_2_.scs8hd_ebufn_2_A _653_/HI
+ vgnd vpwr scs8hd_diode_2
XFILLER_69_110 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_3_.latch_D
+ data_in vgnd vpwr scs8hd_diode_2
XFILLER_69_154 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_0_in_2.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_0_in_2.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_53_500 vgnd vpwr scs8hd_decap_12
XFILLER_27_39 vgnd vpwr scs8hd_decap_12
XFILLER_65_371 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_6_.latch_SLEEPB
+ _592_/Y vgnd vpwr scs8hd_diode_2
XFILLER_25_235 vpwr vgnd scs8hd_fill_2
XFILLER_40_205 vpwr vgnd scs8hd_fill_2
XFILLER_43_27 vgnd vpwr scs8hd_decap_12
XANTENNA__392__B _388_/B vgnd vpwr scs8hd_diode_2
XFILLER_4_117 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mux_fle_1_in_2.INVTX1_12_.scs8hd_inv_1_A top_width_0_height_0__pin_12_
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_3_in_2.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_3_in_2.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_0_in_1.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_0_in_1.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_68_68 vgnd vpwr scs8hd_decap_12
XFILLER_0_345 vgnd vpwr scs8hd_decap_4
Xltile_clb_0.mux_fle_1_in_1.INVTX1_7_.scs8hd_inv_1 left_width_0_height_0__pin_7_ ltile_clb_0.mux_fle_1_in_1.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_ltile_clb_0.mux_fle_3_in_0.INVTX1_9_.scs8hd_inv_1_A right_width_0_height_0__pin_9_
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_3_in_2.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_3_in_2.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_75_135 vgnd vpwr scs8hd_decap_12
X_652_ _652_/HI _652_/LO vgnd vpwr scs8hd_conb_1
XFILLER_63_319 vpwr vgnd scs8hd_fill_2
XANTENNA__567__B _564_/B vgnd vpwr scs8hd_diode_2
X_583_ _247_/X _585_/B _583_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA__286__C address[1] vgnd vpwr scs8hd_diode_2
XFILLER_71_385 vgnd vpwr scs8hd_decap_6
XANTENNA__583__A _247_/X vgnd vpwr scs8hd_diode_2
XPHY_252 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_241 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_230 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_0_.scs8hd_inv_1_A
+ ltile_clb_0.mux_fle_2_in_0.INVTX1_14_.scs8hd_inv_1/Y vgnd vpwr scs8hd_diode_2
XPHY_274 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_263 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_8_401 vgnd vpwr scs8hd_decap_4
XPHY_285 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xltile_clb_0.mux_fle_1_in_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_1_in_1.INVTX1_6_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_1_in_1.LATCH_2_.latch/Q ltile_clb_0.mux_fle_1_in_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
Xltile_clb_0.mux_fle_3_in_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_3_in_1.INVTX1_1_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_3_in_1.LATCH_1_.latch/Q ltile_clb_0.mux_fle_3_in_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XPHY_296 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_8_456 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_1_in_3.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_1_in_3.LATCH_6_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_2_in_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_2_in_0.LATCH_4_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l4_in_0_.TGATE_0_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l4_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_66_168 vpwr vgnd scs8hd_fill_2
XANTENNA__477__B _479_/B vgnd vpwr scs8hd_diode_2
XFILLER_62_341 vgnd vpwr scs8hd_fill_1
Xltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_4_.TGATE_0_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_8_.scs8hd_inv_1/Y
+ _613_/Y ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_4_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_62_374 vgnd vpwr scs8hd_decap_3
XFILLER_22_205 vpwr vgnd scs8hd_fill_2
XFILLER_22_249 vgnd vpwr scs8hd_decap_8
XANTENNA__493__A _380_/X vgnd vpwr scs8hd_diode_2
XFILLER_30_271 vgnd vpwr scs8hd_fill_1
XANTENNA_ltile_clb_0.mem_fle_2_in_3.LATCH_7_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_38_27 vgnd vpwr scs8hd_decap_4
Xltile_clb_0.mux_fle_2_in_2.INVTX1_2_.scs8hd_inv_1 bottom_width_0_height_0__pin_2_
+ ltile_clb_0.mux_fle_2_in_2.INVTX1_2_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XFILLER_57_135 vgnd vpwr scs8hd_decap_8
XFILLER_57_146 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_9_.latch
+ data_in ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_9_.latch/Q
+ _589_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_72_105 vgnd vpwr scs8hd_decap_12
XFILLER_57_179 vpwr vgnd scs8hd_fill_2
XFILLER_38_382 vgnd vpwr scs8hd_decap_3
XFILLER_45_319 vpwr vgnd scs8hd_fill_2
XFILLER_54_15 vgnd vpwr scs8hd_decap_12
XFILLER_53_374 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_1_.scs8hd_inv_1
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_1_.latch/Q
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_5_415 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mem_fle_3_in_1.LATCH_7_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA__578__A address[6] vgnd vpwr scs8hd_diode_2
XFILLER_48_168 vgnd vpwr scs8hd_decap_8
XFILLER_17_511 vgnd vpwr scs8hd_decap_4
XFILLER_28_93 vgnd vpwr scs8hd_decap_12
X_635_ _635_/A _635_/Y vgnd vpwr scs8hd_inv_8
XFILLER_44_341 vpwr vgnd scs8hd_fill_2
X_566_ _540_/A _564_/B _566_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_32_514 vpwr vgnd scs8hd_fill_2
XFILLER_44_352 vgnd vpwr scs8hd_decap_4
XFILLER_44_396 vgnd vpwr scs8hd_fill_1
X_497_ _325_/A _495_/X _497_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA_ltile_clb_0.mem_fle_3_in_2.LATCH_5_.latch_D data_in vgnd vpwr scs8hd_diode_2
Xltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.INVTX1_0_.scs8hd_inv_1
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.INVTX1_0_.scs8hd_inv_1/A
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_60_80 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mem_fle_3_in_3.LATCH_5_.latch_SLEEPB _329_/Y vgnd vpwr scs8hd_diode_2
XFILLER_5_86 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.tap_buf4_0_.scs8hd_inv_1
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.tap_buf4_0_.scs8hd_inv_1/A
+ left_width_0_height_0__pin_11_ vgnd vpwr scs8hd_inv_1
XFILLER_79_271 vgnd vpwr scs8hd_decap_8
XANTENNA__488__A _331_/A vgnd vpwr scs8hd_diode_2
XFILLER_39_135 vgnd vpwr scs8hd_decap_6
XANTENNA_ltile_clb_0.mem_fle_3_in_3.LATCH_3_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_54_105 vgnd vpwr scs8hd_decap_12
XFILLER_27_319 vpwr vgnd scs8hd_fill_2
XFILLER_39_179 vpwr vgnd scs8hd_fill_2
XFILLER_54_149 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_1_.scs8hd_inv_1/Y
+ _620_/Y ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_ltile_clb_0.mux_fle_0_in_0.INVTX1_7_.scs8hd_inv_1_A left_width_0_height_0__pin_7_
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_1_.TGATE_0_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_1_.TGATE_0_.scs8hd_ebufn_2/A
+ _609_/Y ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l4_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_ltile_clb_0.mux_fle_3_in_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_3_in_2.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_2_in_3.INVTX1_6_.scs8hd_inv_1 bottom_width_0_height_0__pin_6_
+ ltile_clb_0.mux_fle_2_in_3.INVTX1_6_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XFILLER_49_15 vgnd vpwr scs8hd_decap_12
XFILLER_49_59 vpwr vgnd scs8hd_fill_2
XANTENNA__398__A _398_/A vgnd vpwr scs8hd_diode_2
XFILLER_58_411 vpwr vgnd scs8hd_fill_2
XFILLER_58_455 vgnd vpwr scs8hd_fill_1
XFILLER_18_308 vgnd vpwr scs8hd_decap_4
X_420_ _434_/A _412_/B _420_/Y vgnd vpwr scs8hd_nor2_4
Xltile_clb_0.mux_fle_2_in_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_2_in_2.INVTX1_1_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_2_in_2.LATCH_1_.latch/Q ltile_clb_0.mux_fle_2_in_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
X_351_ _374_/A _353_/B _351_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_53_193 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.mux_fle_0_in_2.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_0_in_2.INVTX1_6_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_0_in_2.LATCH_2_.latch/Q ltile_clb_0.mux_fle_0_in_2.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_41_344 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.mux_fle_2_in_0.INVTX1_12_.scs8hd_inv_1 top_width_0_height_0__pin_12_
+ ltile_clb_0.mux_fle_2_in_0.INVTX1_12_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_5_.TGATE_1_.scs8hd_ebufn_2_TEB
+ _620_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.mem_ble4_out_0.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
X_282_ _286_/A _282_/B _282_/C _324_/A vgnd vpwr scs8hd_or3_4
XFILLER_5_223 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_1_in_1.INVTX1_4_.scs8hd_inv_1_A top_width_0_height_0__pin_4_
+ vgnd vpwr scs8hd_diode_2
XFILLER_1_473 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_2_in_2.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_2_in_2.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_36_105 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mux_fle_3_in_1.INVTX1_10_.scs8hd_inv_1_A bottom_width_0_height_0__pin_10_
+ vgnd vpwr scs8hd_diode_2
X_618_ _618_/A _618_/Y vgnd vpwr scs8hd_inv_8
XFILLER_17_385 vgnd vpwr scs8hd_fill_1
X_549_ _575_/A _548_/X _549_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA_ltile_clb_0.mux_fle_0_in_0.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_0_in_0.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_72_3 vgnd vpwr scs8hd_decap_12
XANTENNA__490__B _484_/X vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_0_in_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_0_in_0.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_2_in_1.INVTX1_14_.scs8hd_inv_1 ltile_clb_0.mux_fle_2_in_1.INVTX1_14_.scs8hd_inv_1/A
+ ltile_clb_0.mux_fle_2_in_1.INVTX1_14_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
Xltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_9_.latch
+ data_in ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_9_.latch/Q
+ _563_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_ltile_clb_0.mux_fle_3_in_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_3_in_1.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_9_.latch_D
+ data_in vgnd vpwr scs8hd_diode_2
XFILLER_82_211 vgnd vpwr scs8hd_decap_6
XFILLER_55_447 vgnd vpwr scs8hd_decap_4
XFILLER_35_39 vgnd vpwr scs8hd_decap_12
XPHY_818 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_807 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_63_480 vpwr vgnd scs8hd_fill_2
XFILLER_35_160 vgnd vpwr scs8hd_fill_1
XPHY_829 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_ltile_clb_0.mux_fle_2_in_2.INVTX1_1_.scs8hd_inv_1_A right_width_0_height_0__pin_1_
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_3_in_0.mux_l1_in_2_.TGATE_3_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_3_in_0.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_23_388 vgnd vpwr scs8hd_fill_1
XFILLER_51_27 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mem_fle_1_in_3.LATCH_6_.latch_SLEEPB _442_/Y vgnd vpwr scs8hd_diode_2
XFILLER_2_215 vgnd vpwr scs8hd_decap_3
XFILLER_76_68 vgnd vpwr scs8hd_decap_12
XFILLER_58_285 vpwr vgnd scs8hd_fill_2
XFILLER_18_105 vgnd vpwr scs8hd_decap_12
XFILLER_46_425 vgnd vpwr scs8hd_decap_3
XFILLER_73_222 vpwr vgnd scs8hd_fill_2
XFILLER_73_211 vpwr vgnd scs8hd_fill_2
XFILLER_46_436 vgnd vpwr scs8hd_decap_4
XFILLER_61_406 vpwr vgnd scs8hd_fill_2
XANTENNA__575__B _575_/B vgnd vpwr scs8hd_diode_2
X_403_ _392_/A _399_/B _403_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_61_439 vgnd vpwr scs8hd_fill_1
XFILLER_54_491 vpwr vgnd scs8hd_fill_2
XPHY_50 vgnd vpwr scs8hd_decap_3
XFILLER_26_193 vpwr vgnd scs8hd_fill_2
XPHY_61 vgnd vpwr scs8hd_decap_3
XPHY_72 vgnd vpwr scs8hd_decap_3
XPHY_83 vgnd vpwr scs8hd_decap_3
XPHY_94 vgnd vpwr scs8hd_decap_3
X_334_ _334_/A _392_/A vgnd vpwr scs8hd_buf_1
XANTENNA__591__A _539_/A vgnd vpwr scs8hd_diode_2
X_265_ _264_/X _535_/A vgnd vpwr scs8hd_buf_1
XFILLER_41_196 vpwr vgnd scs8hd_fill_2
XFILLER_1_270 vgnd vpwr scs8hd_decap_6
XFILLER_2_32 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.mux_fle_0_in_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_0_in_0.INVTX1_0_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_0_in_0.LATCH_0_.latch/Q ltile_clb_0.mux_fle_0_in_0.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_49_230 vgnd vpwr scs8hd_fill_1
XFILLER_49_285 vgnd vpwr scs8hd_decap_6
XFILLER_64_266 vpwr vgnd scs8hd_fill_2
XFILLER_64_255 vgnd vpwr scs8hd_decap_3
XFILLER_64_244 vpwr vgnd scs8hd_fill_2
XANTENNA__485__B _484_/X vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_2_in_2.mux_l1_in_3_.TGATE_2_.scs8hd_ebufn_2_A _650_/HI
+ vgnd vpwr scs8hd_diode_2
XFILLER_17_171 vgnd vpwr scs8hd_decap_3
XFILLER_17_182 vgnd vpwr scs8hd_fill_1
XFILLER_45_480 vpwr vgnd scs8hd_fill_2
XFILLER_32_141 vgnd vpwr scs8hd_decap_12
XFILLER_60_472 vgnd vpwr scs8hd_decap_4
XFILLER_20_325 vpwr vgnd scs8hd_fill_2
XFILLER_9_392 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.mux_fle_3_in_2.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_3_in_2.mux_l1_in_2_.TGATE_3_.scs8hd_ebufn_2/Z
+ ltile_clb_0.mem_fle_3_in_2.LATCH_6_.latch/Q ltile_clb_0.mux_fle_3_in_2.INVTX1_14_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_ltile_clb_0.mux_fle_0_in_0.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_0_in_0.INVTX1_10_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_1_.TGATE_0_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_1_.TGATE_0_.scs8hd_ebufn_2/A
+ _631_/Y ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_ltile_clb_0.mem_fle_2_in_2.LATCH_6_.latch_SLEEPB _400_/Y vgnd vpwr scs8hd_diode_2
XFILLER_46_27 vgnd vpwr scs8hd_decap_4
XANTENNA__395__B _387_/A vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_1_in_3.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_1_in_3.INVTX1_1_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_1_in_3.LATCH_1_.latch/Q ltile_clb_0.mux_fle_1_in_3.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_55_277 vpwr vgnd scs8hd_fill_2
XFILLER_55_266 vgnd vpwr scs8hd_decap_6
XANTENNA_ltile_clb_0.mux_fle_0_in_3.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_0_in_3.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_2_in_0.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_2_in_0.INVTX1_12_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_2_in_0.LATCH_0_.latch/Q ltile_clb_0.mux_fle_2_in_0.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_70_225 vpwr vgnd scs8hd_fill_2
XFILLER_55_299 vgnd vpwr scs8hd_decap_4
XFILLER_43_428 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_2_in_3.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_2_in_3.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_62_15 vgnd vpwr scs8hd_decap_12
XPHY_626 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_615 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_604 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_659 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_648 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_637 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_51_461 vpwr vgnd scs8hd_fill_2
XFILLER_23_196 vpwr vgnd scs8hd_fill_2
XFILLER_11_358 vgnd vpwr scs8hd_decap_4
XFILLER_11_74 vgnd vpwr scs8hd_decap_12
XFILLER_3_513 vgnd vpwr scs8hd_decap_3
XANTENNA_ltile_clb_0.mux_fle_2_in_0.INVTX1_14_.scs8hd_inv_1_A ltile_clb_0.mux_fle_2_in_0.INVTX1_14_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_2_3 vgnd vpwr scs8hd_decap_12
XANTENNA__586__A _261_/X vgnd vpwr scs8hd_diode_2
XFILLER_19_458 vpwr vgnd scs8hd_fill_2
XFILLER_46_244 vpwr vgnd scs8hd_fill_2
XFILLER_61_214 vpwr vgnd scs8hd_fill_2
XFILLER_27_480 vpwr vgnd scs8hd_fill_2
XFILLER_36_93 vgnd vpwr scs8hd_decap_12
XFILLER_14_141 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.mux_fle_3_in_3.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_3_in_3.INVTX1_13_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_3_in_3.LATCH_1_.latch/Q ltile_clb_0.mux_fle_3_in_3.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
X_317_ _380_/A address[7] _346_/C vgnd vpwr scs8hd_or2_4
Xltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_9_.latch
+ data_in ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_9_.latch/Q
+ _537_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA__471__D _346_/D vgnd vpwr scs8hd_diode_2
XFILLER_10_380 vpwr vgnd scs8hd_fill_2
X_248_ _248_/A _247_/X _248_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_6_351 vgnd vpwr scs8hd_decap_8
XFILLER_6_384 vgnd vpwr scs8hd_decap_4
XFILLER_6_373 vpwr vgnd scs8hd_fill_2
XFILLER_69_314 vgnd vpwr scs8hd_fill_1
XFILLER_35_3 vgnd vpwr scs8hd_decap_12
XFILLER_69_358 vpwr vgnd scs8hd_fill_2
XFILLER_69_336 vgnd vpwr scs8hd_fill_1
Xltile_clb_0.mux_fle_1_in_2.INVTX1_10_.scs8hd_inv_1 bottom_width_0_height_0__pin_10_
+ ltile_clb_0.mux_fle_1_in_2.INVTX1_10_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XFILLER_77_380 vpwr vgnd scs8hd_fill_2
XANTENNA__496__A _314_/A vgnd vpwr scs8hd_diode_2
XFILLER_37_222 vgnd vpwr scs8hd_decap_3
XFILLER_37_255 vpwr vgnd scs8hd_fill_2
XFILLER_37_299 vgnd vpwr scs8hd_decap_4
XFILLER_52_236 vpwr vgnd scs8hd_fill_2
XFILLER_40_409 vgnd vpwr scs8hd_decap_8
XFILLER_33_472 vgnd vpwr scs8hd_decap_3
XFILLER_60_280 vgnd vpwr scs8hd_decap_4
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_11_.latch_D
+ data_in vgnd vpwr scs8hd_diode_2
Xltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_13_.latch
+ data_in ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_13_.latch/Q
+ _558_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_ltile_clb_0.mem_fle_3_in_1.LATCH_6_.latch_SLEEPB _362_/Y vgnd vpwr scs8hd_diode_2
XFILLER_57_15 vgnd vpwr scs8hd_decap_12
XFILLER_57_59 vpwr vgnd scs8hd_fill_2
XFILLER_71_501 vgnd vpwr scs8hd_decap_12
XFILLER_16_406 vgnd vpwr scs8hd_fill_1
Xltile_clb_0.mux_fle_1_in_3.INVTX1_12_.scs8hd_inv_1 top_width_0_height_0__pin_12_
+ ltile_clb_0.mux_fle_1_in_3.INVTX1_12_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XFILLER_43_214 vpwr vgnd scs8hd_fill_2
XPHY_401 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_412 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_423 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_434 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xltile_clb_0.mux_fle_1_in_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_1_in_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ ltile_clb_0.mem_fle_1_in_0.LATCH_5_.latch/Q ltile_clb_0.mux_fle_1_in_0.INVTX1_14_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_24_494 vpwr vgnd scs8hd_fill_2
XPHY_445 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_456 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_467 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_478 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_489 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_11_188 vgnd vpwr scs8hd_fill_1
Xltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_3_.scs8hd_inv_1
+ ltile_clb_0.mux_fle_3_in_3.INVTX1_14_.scs8hd_inv_1/Y _611_/A vgnd vpwr scs8hd_inv_1
XFILLER_7_159 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mem_fle_0_in_2.LATCH_7_.latch_SLEEPB _496_/Y vgnd vpwr scs8hd_diode_2
XFILLER_78_166 vgnd vpwr scs8hd_decap_12
XFILLER_66_317 vpwr vgnd scs8hd_fill_2
XFILLER_66_328 vpwr vgnd scs8hd_fill_2
XFILLER_34_203 vpwr vgnd scs8hd_fill_2
XFILLER_34_247 vgnd vpwr scs8hd_decap_3
XFILLER_15_461 vpwr vgnd scs8hd_fill_2
XFILLER_30_420 vgnd vpwr scs8hd_decap_8
XFILLER_30_442 vpwr vgnd scs8hd_fill_2
XANTENNA__482__C _228_/X vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_2_in_3.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_2_in_3.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2/Z
+ ltile_clb_0.mem_fle_2_in_3.LATCH_6_.latch/Q ltile_clb_0.mux_fle_2_in_3.INVTX1_14_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_ltile_clb_0.mux_fle_3_in_2.INVTX1_7_.scs8hd_inv_1_A left_width_0_height_0__pin_7_
+ vgnd vpwr scs8hd_diode_2
XFILLER_57_306 vgnd vpwr scs8hd_decap_3
XANTENNA_ltile_clb_0.mux_fle_0_in_3.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_0_in_3.LATCH_7_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_69_188 vgnd vpwr scs8hd_fill_1
Xltile_clb_0.mux_fle_1_in_1.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_1_in_1.INVTX1_12_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_1_in_1.LATCH_0_.latch/Q ltile_clb_0.mux_fle_1_in_1.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_ltile_clb_0.mux_fle_1_in_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_1_in_0.LATCH_5_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_53_512 vgnd vpwr scs8hd_decap_4
XFILLER_25_203 vgnd vpwr scs8hd_decap_4
XANTENNA_ltile_clb_0.mux_fle_2_in_3.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_2_in_3.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_65_394 vgnd vpwr scs8hd_fill_1
XFILLER_25_225 vpwr vgnd scs8hd_fill_2
XFILLER_21_420 vpwr vgnd scs8hd_fill_2
XFILLER_21_431 vpwr vgnd scs8hd_fill_2
XFILLER_33_280 vpwr vgnd scs8hd_fill_2
XFILLER_43_39 vgnd vpwr scs8hd_decap_12
XFILLER_21_453 vgnd vpwr scs8hd_decap_3
Xltile_clb_0.mux_fle_0_in_2.INVTX1_1_.scs8hd_inv_1 right_width_0_height_0__pin_1_
+ ltile_clb_0.mux_fle_0_in_2.INVTX1_1_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.buf4_0_.scs8hd_buf_1_A
+ ltile_clb_0.mux_fle_1_in_0.INVTX1_14_.scs8hd_inv_1/Y vgnd vpwr scs8hd_diode_2
XFILLER_21_475 vgnd vpwr scs8hd_decap_3
XFILLER_4_129 vgnd vpwr scs8hd_decap_12
XFILLER_0_302 vpwr vgnd scs8hd_fill_2
XFILLER_0_324 vpwr vgnd scs8hd_fill_2
XFILLER_48_317 vpwr vgnd scs8hd_fill_2
XFILLER_48_328 vpwr vgnd scs8hd_fill_2
X_651_ _651_/HI _651_/LO vgnd vpwr scs8hd_conb_1
XFILLER_75_147 vgnd vpwr scs8hd_decap_12
XFILLER_56_350 vgnd vpwr scs8hd_fill_1
X_582_ _556_/A _585_/B _582_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_56_394 vgnd vpwr scs8hd_decap_3
XFILLER_17_51 vgnd vpwr scs8hd_decap_8
XFILLER_17_62 vgnd vpwr scs8hd_decap_12
XFILLER_71_375 vgnd vpwr scs8hd_fill_1
XPHY_242 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_231 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_220 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__583__B _585_/B vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mem_fle_1_in_1.LATCH_7_.latch_SLEEPB _463_/Y vgnd vpwr scs8hd_diode_2
XPHY_286 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_275 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_264 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_253 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_297 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_8_468 vgnd vpwr scs8hd_decap_3
XANTENNA_ltile_clb_0.mux_fle_1_in_3.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_1_in_3.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_3_184 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_1_.TGATE_0_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_1_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_58_80 vgnd vpwr scs8hd_decap_12
XFILLER_39_339 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_1_.scs8hd_inv_1_A
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_3_in_3.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_3_in_3.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_22_228 vgnd vpwr scs8hd_decap_12
XANTENNA__493__B _427_/B vgnd vpwr scs8hd_diode_2
Xltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_2_.TGATE_1_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_2_.TGATE_1_.scs8hd_ebufn_2/A
+ _606_/Y ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_1_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_9_.latch_SLEEPB
+ _537_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_3_in_2.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_3_in_2.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2_TEB
+ _612_/Y vgnd vpwr scs8hd_diode_2
XFILLER_72_117 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.mux_fle_0_in_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_0_in_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ ltile_clb_0.mem_fle_0_in_1.LATCH_5_.latch/Q ltile_clb_0.mux_fle_0_in_1.INVTX1_14_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_38_350 vgnd vpwr scs8hd_decap_4
XFILLER_65_191 vpwr vgnd scs8hd_fill_2
XFILLER_65_180 vgnd vpwr scs8hd_fill_1
XFILLER_54_27 vgnd vpwr scs8hd_decap_4
XFILLER_53_320 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.mux_fle_0_in_3.INVTX1_5_.scs8hd_inv_1 right_width_0_height_0__pin_5_
+ ltile_clb_0.mux_fle_0_in_3.INVTX1_5_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XFILLER_53_397 vgnd vpwr scs8hd_decap_4
XFILLER_13_228 vgnd vpwr scs8hd_decap_3
XFILLER_13_217 vgnd vpwr scs8hd_decap_4
XFILLER_70_15 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.buf4_2_.scs8hd_buf_1_A
+ ltile_clb_0.mux_fle_3_in_2.INVTX1_14_.scs8hd_inv_1/Y vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mem_fle_2_in_0.LATCH_7_.latch_SLEEPB _430_/Y vgnd vpwr scs8hd_diode_2
XANTENNA__578__B address[7] vgnd vpwr scs8hd_diode_2
XFILLER_0_187 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mux_fle_0_in_2.INVTX1_5_.scs8hd_inv_1_A right_width_0_height_0__pin_5_
+ vgnd vpwr scs8hd_diode_2
XFILLER_48_158 vgnd vpwr scs8hd_fill_1
X_634_ _634_/A _634_/Y vgnd vpwr scs8hd_inv_8
XFILLER_29_361 vpwr vgnd scs8hd_fill_2
XFILLER_63_139 vgnd vpwr scs8hd_fill_1
XFILLER_56_180 vpwr vgnd scs8hd_fill_2
XANTENNA__594__A _542_/A vgnd vpwr scs8hd_diode_2
X_565_ _539_/A _564_/B _565_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_11_.scs8hd_inv_1_A
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_11_.latch/Q
+ vgnd vpwr scs8hd_diode_2
X_496_ _314_/A _495_/X _496_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_44_93 vgnd vpwr scs8hd_decap_12
XFILLER_8_254 vgnd vpwr scs8hd_decap_8
XFILLER_8_243 vpwr vgnd scs8hd_fill_2
XFILLER_8_276 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.mem_ble4_out_0.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_5_98 vgnd vpwr scs8hd_decap_12
XFILLER_4_482 vgnd vpwr scs8hd_decap_12
XFILLER_4_471 vgnd vpwr scs8hd_decap_8
Xltile_clb_0.mux_fle_0_in_2.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_0_in_2.INVTX1_12_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_0_in_2.LATCH_0_.latch/Q ltile_clb_0.mux_fle_0_in_2.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_ltile_clb_0.mux_fle_1_in_3.mux_l1_in_3_.TGATE_2_.scs8hd_ebufn_2_A _647_/HI
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_6_.TGATE_0_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_12_.scs8hd_inv_1/Y
+ _621_/Y ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_3_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA__488__B _484_/X vgnd vpwr scs8hd_diode_2
XFILLER_67_467 vpwr vgnd scs8hd_fill_2
XFILLER_39_158 vpwr vgnd scs8hd_fill_2
XFILLER_82_404 vgnd vpwr scs8hd_decap_12
XFILLER_67_489 vgnd vpwr scs8hd_decap_12
XFILLER_54_117 vgnd vpwr scs8hd_decap_12
XFILLER_47_191 vpwr vgnd scs8hd_fill_2
XFILLER_23_504 vgnd vpwr scs8hd_decap_12
XFILLER_35_397 vgnd vpwr scs8hd_decap_4
XFILLER_50_312 vpwr vgnd scs8hd_fill_2
XFILLER_50_356 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_1_in_3.INVTX1_2_.scs8hd_inv_1_A bottom_width_0_height_0__pin_2_
+ vgnd vpwr scs8hd_diode_2
XFILLER_50_378 vpwr vgnd scs8hd_fill_2
XFILLER_50_389 vpwr vgnd scs8hd_fill_2
XFILLER_49_27 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mux_fle_2_in_1.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_2_in_1.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_65_15 vgnd vpwr scs8hd_decap_12
XFILLER_73_404 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_0_in_3.INVTX1_14_.scs8hd_inv_1_A ltile_clb_0.mux_fle_0_in_3.INVTX1_14_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_65_59 vpwr vgnd scs8hd_fill_2
XFILLER_45_139 vpwr vgnd scs8hd_fill_2
X_350_ _326_/A _353_/B _350_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_14_515 vgnd vpwr scs8hd_fill_1
XFILLER_26_386 vpwr vgnd scs8hd_fill_2
XFILLER_41_323 vpwr vgnd scs8hd_fill_2
X_281_ _267_/X _539_/A _281_/Y vgnd vpwr scs8hd_nor2_4
Xltile_clb_0.mux_fle_2_in_0.INVTX1_2_.scs8hd_inv_1 bottom_width_0_height_0__pin_2_
+ ltile_clb_0.mux_fle_2_in_0.INVTX1_2_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XANTENNA__589__A _272_/X vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB
+ _630_/Y vgnd vpwr scs8hd_diode_2
XFILLER_1_485 vgnd vpwr scs8hd_decap_3
XFILLER_49_423 vpwr vgnd scs8hd_fill_2
XFILLER_49_456 vgnd vpwr scs8hd_decap_3
XFILLER_36_117 vgnd vpwr scs8hd_decap_12
XFILLER_49_489 vgnd vpwr scs8hd_decap_4
XFILLER_64_459 vgnd vpwr scs8hd_decap_6
XFILLER_17_353 vpwr vgnd scs8hd_fill_2
X_617_ _617_/A _617_/Y vgnd vpwr scs8hd_inv_8
XFILLER_72_470 vgnd vpwr scs8hd_decap_12
X_548_ _547_/X _548_/X vgnd vpwr scs8hd_buf_1
XFILLER_44_183 vgnd vpwr scs8hd_fill_1
X_479_ _435_/A _479_/B _479_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_32_378 vpwr vgnd scs8hd_fill_2
XFILLER_32_389 vgnd vpwr scs8hd_decap_8
XFILLER_65_3 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_6_.TGATE_0_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_12_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_3_in_2.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_3_in_2.INVTX1_7_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_3_in_2.LATCH_3_.latch/Q ltile_clb_0.mux_fle_3_in_2.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_3_.scs8hd_inv_1_A
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_59_209 vpwr vgnd scs8hd_fill_2
XANTENNA__499__A _331_/A vgnd vpwr scs8hd_diode_2
Xltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_5_.scs8hd_inv_1/Y
+ _628_/Y ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_1_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_67_297 vpwr vgnd scs8hd_fill_2
XPHY_808 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_63_492 vpwr vgnd scs8hd_fill_2
XFILLER_23_301 vpwr vgnd scs8hd_fill_2
XPHY_819 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_6_.TGATE_0_.scs8hd_ebufn_2_TEB
+ _621_/Y vgnd vpwr scs8hd_diode_2
XFILLER_23_345 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_11_.latch
+ data_in ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_11_.latch/Q
+ _262_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_51_39 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.mem_fle_0_in_0.LATCH_4_.latch data_in ltile_clb_0.mem_fle_0_in_0.LATCH_4_.latch/Q
+ _521_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_1_.TGATE_0_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_1_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_58_264 vgnd vpwr scs8hd_decap_8
XFILLER_18_117 vgnd vpwr scs8hd_decap_12
XFILLER_73_256 vpwr vgnd scs8hd_fill_2
XFILLER_73_245 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_4_.scs8hd_inv_1
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_4_.latch/Q
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_ltile_clb_0.mem_fle_2_in_3.LATCH_0_.latch_SLEEPB _395_/Y vgnd vpwr scs8hd_diode_2
X_402_ _391_/A _399_/B _402_/Y vgnd vpwr scs8hd_nor2_4
Xltile_clb_0.mem_fle_1_in_0.LATCH_3_.latch data_in ltile_clb_0.mem_fle_1_in_0.LATCH_3_.latch/Q
+ _478_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XPHY_40 vgnd vpwr scs8hd_decap_3
XFILLER_26_172 vgnd vpwr scs8hd_decap_8
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__ff_0.DFFSRQ_0_.dff_SETB
+ set vgnd vpwr scs8hd_diode_2
XFILLER_25_51 vgnd vpwr scs8hd_decap_8
XFILLER_25_62 vgnd vpwr scs8hd_decap_12
XPHY_51 vgnd vpwr scs8hd_decap_3
XPHY_62 vgnd vpwr scs8hd_decap_3
XPHY_73 vgnd vpwr scs8hd_decap_3
X_333_ _333_/A _334_/A vgnd vpwr scs8hd_buf_1
XFILLER_41_175 vpwr vgnd scs8hd_fill_2
XPHY_84 vgnd vpwr scs8hd_decap_3
XPHY_95 vgnd vpwr scs8hd_decap_3
Xltile_clb_0.mux_fle_2_in_1.INVTX1_6_.scs8hd_inv_1 bottom_width_0_height_0__pin_6_
+ ltile_clb_0.mux_fle_2_in_1.INVTX1_6_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XANTENNA__591__B _588_/X vgnd vpwr scs8hd_diode_2
X_264_ _236_/X _263_/X _264_/X vgnd vpwr scs8hd_or2_4
XANTENNA_ltile_clb_0.mux_fle_3_in_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_3_in_1.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mem_fle_2_in_0.LATCH_2_.latch data_in ltile_clb_0.mem_fle_2_in_0.LATCH_2_.latch/Q
+ _435_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_1_282 vpwr vgnd scs8hd_fill_2
XFILLER_2_44 vgnd vpwr scs8hd_decap_12
XFILLER_37_404 vgnd vpwr scs8hd_decap_6
XFILLER_66_80 vgnd vpwr scs8hd_decap_12
XFILLER_49_297 vpwr vgnd scs8hd_fill_2
XFILLER_52_407 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.mem_fle_3_in_0.LATCH_1_.latch data_in ltile_clb_0.mem_fle_3_in_0.LATCH_1_.latch/Q
+ _378_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_45_470 vpwr vgnd scs8hd_fill_2
XFILLER_60_440 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_3_in_0.mux_l1_in_3_.TGATE_2_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_3_in_0.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_15_.scs8hd_inv_1
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_15_.latch/Q
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_15_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_20_315 vgnd vpwr scs8hd_fill_1
XFILLER_20_337 vgnd vpwr scs8hd_decap_4
XFILLER_9_360 vgnd vpwr scs8hd_decap_4
XANTENNA_ltile_clb_0.mux_fle_1_in_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_1_in_2.LATCH_4_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_9_371 vgnd vpwr scs8hd_decap_3
XFILLER_55_245 vpwr vgnd scs8hd_fill_2
XFILLER_70_215 vgnd vpwr scs8hd_decap_3
XFILLER_62_27 vgnd vpwr scs8hd_decap_4
XPHY_616 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_605 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
+ _608_/Y vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mem_fle_0_in_2.LATCH_7_.latch data_in ltile_clb_0.mem_fle_0_in_2.LATCH_7_.latch/Q
+ _496_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XPHY_649 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_638 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_627 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xltile_clb_0.mux_fle_1_in_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_1_in_0.INVTX1_6_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_1_in_0.LATCH_2_.latch/Q ltile_clb_0.mux_fle_1_in_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_51_484 vgnd vpwr scs8hd_decap_4
XFILLER_11_337 vgnd vpwr scs8hd_decap_4
Xltile_clb_0.mux_fle_3_in_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_3_in_0.INVTX1_1_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_3_in_0.LATCH_1_.latch/Q ltile_clb_0.mux_fle_3_in_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
Xltile_clb_0.mux_fle_3_in_2.INVTX1_1_.scs8hd_inv_1 right_width_0_height_0__pin_1_
+ ltile_clb_0.mux_fle_3_in_2.INVTX1_1_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XANTENNA_ltile_clb_0.mem_fle_3_in_2.LATCH_0_.latch_SLEEPB _356_/Y vgnd vpwr scs8hd_diode_2
XFILLER_11_86 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.mem_fle_1_in_2.LATCH_6_.latch data_in ltile_clb_0.mem_fle_1_in_2.LATCH_6_.latch/Q
+ _453_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_78_304 vpwr vgnd scs8hd_fill_2
XANTENNA__586__B _585_/B vgnd vpwr scs8hd_diode_2
XFILLER_19_437 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_2_.latch_SLEEPB
+ _570_/Y vgnd vpwr scs8hd_diode_2
XFILLER_34_407 vgnd vpwr scs8hd_decap_3
XFILLER_46_267 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.mem_fle_2_in_2.LATCH_5_.latch data_in ltile_clb_0.mem_fle_2_in_2.LATCH_5_.latch/Q
+ _401_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_61_248 vpwr vgnd scs8hd_fill_2
XFILLER_61_237 vgnd vpwr scs8hd_fill_1
XFILLER_27_492 vpwr vgnd scs8hd_fill_2
XFILLER_42_473 vgnd vpwr scs8hd_decap_6
X_316_ address[6] _380_/A vgnd vpwr scs8hd_inv_8
XFILLER_52_93 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.mux_fle_2_in_3.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_2_in_3.INVTX1_7_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_2_in_3.LATCH_3_.latch/Q ltile_clb_0.mux_fle_2_in_3.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
X_247_ _246_/X _247_/X vgnd vpwr scs8hd_buf_1
XANTENNA_ltile_clb_0.mux_fle_2_in_3.INVTX1_8_.scs8hd_inv_1_A top_width_0_height_0__pin_8_
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_2_in_2.INVTX1_12_.scs8hd_inv_1_A top_width_0_height_0__pin_12_
+ vgnd vpwr scs8hd_diode_2
XFILLER_6_330 vgnd vpwr scs8hd_decap_6
Xltile_clb_0.mem_fle_3_in_2.LATCH_4_.latch data_in ltile_clb_0.mem_fle_3_in_2.LATCH_4_.latch/Q
+ _352_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_ltile_clb_0.mux_fle_3_in_2.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_3_in_2.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_69_304 vgnd vpwr scs8hd_fill_1
Xltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_9_.scs8hd_inv_1
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_9_.latch/Q
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_9_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_ltile_clb_0.mux_fle_3_in_0.INVTX1_4_.scs8hd_inv_1_A top_width_0_height_0__pin_4_
+ vgnd vpwr scs8hd_diode_2
XFILLER_28_3 vgnd vpwr scs8hd_decap_12
XANTENNA__496__B _495_/X vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mem_fle_0_in_3.LATCH_1_.latch_SLEEPB _491_/Y vgnd vpwr scs8hd_diode_2
XFILLER_37_245 vgnd vpwr scs8hd_fill_1
XFILLER_18_470 vgnd vpwr scs8hd_decap_8
XFILLER_37_289 vgnd vpwr scs8hd_decap_8
XANTENNA_ltile_clb_0.mux_fle_1_in_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_1_in_0.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_5_.scs8hd_inv_1_A
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_5_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_33_484 vpwr vgnd scs8hd_fill_2
XFILLER_20_189 vpwr vgnd scs8hd_fill_2
XFILLER_57_27 vgnd vpwr scs8hd_decap_12
XFILLER_28_245 vgnd vpwr scs8hd_decap_8
XFILLER_28_256 vgnd vpwr scs8hd_decap_8
XFILLER_73_15 vgnd vpwr scs8hd_decap_12
XFILLER_71_513 vgnd vpwr scs8hd_decap_3
XFILLER_28_267 vpwr vgnd scs8hd_fill_2
XFILLER_28_289 vgnd vpwr scs8hd_decap_4
XFILLER_73_59 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_0_in_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_0_in_0.LATCH_6_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_43_248 vpwr vgnd scs8hd_fill_2
XFILLER_43_259 vgnd vpwr scs8hd_decap_4
XPHY_402 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_413 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_424 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_435 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xltile_clb_0.mux_fle_3_in_3.INVTX1_5_.scs8hd_inv_1 right_width_0_height_0__pin_5_
+ ltile_clb_0.mux_fle_3_in_3.INVTX1_5_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XFILLER_11_123 vgnd vpwr scs8hd_decap_12
XFILLER_24_484 vgnd vpwr scs8hd_fill_1
XPHY_446 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_457 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_468 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_479 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_6_.TGATE_0_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_12_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_3_322 vpwr vgnd scs8hd_fill_2
XFILLER_3_377 vpwr vgnd scs8hd_fill_2
XFILLER_3_399 vpwr vgnd scs8hd_fill_2
XFILLER_78_178 vgnd vpwr scs8hd_decap_12
XANTENNA__597__A _545_/A vgnd vpwr scs8hd_diode_2
XFILLER_19_234 vpwr vgnd scs8hd_fill_2
XFILLER_74_373 vpwr vgnd scs8hd_fill_2
XFILLER_19_267 vgnd vpwr scs8hd_fill_1
XFILLER_34_215 vgnd vpwr scs8hd_decap_4
XFILLER_34_237 vgnd vpwr scs8hd_decap_6
XFILLER_15_484 vpwr vgnd scs8hd_fill_2
XFILLER_8_32 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
+ _604_/Y vgnd vpwr scs8hd_diode_2
XANTENNA__482__D _526_/D vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mem_fle_1_in_2.LATCH_1_.latch_SLEEPB _458_/Y vgnd vpwr scs8hd_diode_2
XFILLER_69_123 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mux_fle_3_in_2.mux_l1_in_3_.TGATE_2_.scs8hd_ebufn_2_A _654_/HI
+ vgnd vpwr scs8hd_diode_2
XFILLER_69_178 vpwr vgnd scs8hd_fill_2
XFILLER_57_329 vpwr vgnd scs8hd_fill_2
XANTENNA__300__A _300_/A vgnd vpwr scs8hd_diode_2
XFILLER_65_351 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.buf4_3_.scs8hd_buf_1
+ ltile_clb_0.mux_fle_1_in_3.INVTX1_14_.scs8hd_inv_1/Y _626_/A vgnd vpwr scs8hd_buf_1
XFILLER_80_343 vgnd vpwr scs8hd_fill_1
XFILLER_25_248 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.mux_fle_0_in_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_0_in_1.INVTX1_6_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_0_in_1.LATCH_2_.latch/Q ltile_clb_0.mux_fle_0_in_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_80_354 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.mux_fle_2_in_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_2_in_1.INVTX1_1_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_2_in_1.LATCH_1_.latch/Q ltile_clb_0.mux_fle_2_in_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_80_398 vgnd vpwr scs8hd_decap_3
XFILLER_80_387 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_2_in_3.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_2_in_3.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_1_in_0.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_1_in_0.INVTX1_10_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_3_in_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_3_in_0.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_68_15 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l4_in_0_.TGATE_0_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l4_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ _635_/Y ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_16_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_75_159 vgnd vpwr scs8hd_decap_4
XANTENNA_ltile_clb_0.mux_fle_3_in_3.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_3_in_3.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_2_in_2.mux_l1_in_2_.TGATE_3_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_2_in_2.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
X_650_ _650_/HI _650_/LO vgnd vpwr scs8hd_conb_1
X_581_ _580_/X _585_/B vgnd vpwr scs8hd_buf_1
XFILLER_16_204 vgnd vpwr scs8hd_decap_4
XFILLER_16_215 vpwr vgnd scs8hd_fill_2
XFILLER_71_310 vpwr vgnd scs8hd_fill_2
XFILLER_17_74 vgnd vpwr scs8hd_decap_12
XFILLER_71_354 vpwr vgnd scs8hd_fill_2
XPHY_210 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_ltile_clb_0.mux_fle_0_in_1.INVTX1_11_.scs8hd_inv_1_A left_width_0_height_0__pin_11_
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_0_in_0.INVTX1_2_.scs8hd_inv_1_A bottom_width_0_height_0__pin_2_
+ vgnd vpwr scs8hd_diode_2
XPHY_243 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_232 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_221 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_31_229 vpwr vgnd scs8hd_fill_2
XFILLER_12_454 vgnd vpwr scs8hd_decap_4
XPHY_276 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_265 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_254 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_33_51 vgnd vpwr scs8hd_decap_8
XPHY_287 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_298 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_33_62 vgnd vpwr scs8hd_decap_12
XFILLER_79_443 vgnd vpwr scs8hd_decap_3
XFILLER_79_410 vgnd vpwr scs8hd_decap_8
XFILLER_3_196 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mem_fle_2_in_1.LATCH_1_.latch_SLEEPB _424_/Y vgnd vpwr scs8hd_diode_2
Xltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_15_.scs8hd_inv_1
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_15_.latch/Q
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_15_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_74_80 vgnd vpwr scs8hd_decap_12
XFILLER_50_505 vgnd vpwr scs8hd_decap_8
XFILLER_15_270 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.mem_ble4_out_0.LATCH_1_.latch_D
+ data_in vgnd vpwr scs8hd_diode_2
XANTENNA__493__C _228_/X vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_7_.latch_SLEEPB
+ _281_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.mem_ble4_out_0.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_7_.scs8hd_inv_1_A
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_7_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_72_129 vgnd vpwr scs8hd_decap_12
XFILLER_65_170 vgnd vpwr scs8hd_decap_4
XFILLER_53_365 vgnd vpwr scs8hd_fill_1
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
+ _622_/Y vgnd vpwr scs8hd_diode_2
XFILLER_70_27 vgnd vpwr scs8hd_decap_4
XFILLER_21_262 vpwr vgnd scs8hd_fill_2
XFILLER_5_428 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.mux_fle_1_in_0.INVTX1_14_.scs8hd_inv_1 ltile_clb_0.mux_fle_1_in_0.INVTX1_14_.scs8hd_inv_1/A
+ ltile_clb_0.mux_fle_1_in_0.INVTX1_14_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XANTENNA__578__C _227_/X vgnd vpwr scs8hd_diode_2
XFILLER_76_468 vgnd vpwr scs8hd_decap_12
XFILLER_0_199 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mux_fle_3_in_3.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_3_in_3.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
X_633_ _633_/A _633_/Y vgnd vpwr scs8hd_inv_8
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_0_.scs8hd_inv_1_A
+ ltile_clb_0.mux_fle_1_in_0.INVTX1_14_.scs8hd_inv_1/Y vgnd vpwr scs8hd_diode_2
Xltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ _615_/Y ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
Xltile_clb_0.mux_fle_0_in_0.INVTX1_1_.scs8hd_inv_1 right_width_0_height_0__pin_1_
+ ltile_clb_0.mux_fle_0_in_0.INVTX1_1_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XFILLER_44_310 vgnd vpwr scs8hd_decap_4
XFILLER_44_321 vpwr vgnd scs8hd_fill_2
XANTENNA__594__B _588_/X vgnd vpwr scs8hd_diode_2
X_564_ _564_/A _564_/B _564_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_71_184 vgnd vpwr scs8hd_decap_6
XFILLER_71_162 vpwr vgnd scs8hd_fill_2
X_495_ _502_/B _495_/X vgnd vpwr scs8hd_buf_1
XFILLER_44_398 vpwr vgnd scs8hd_fill_2
XFILLER_12_295 vgnd vpwr scs8hd_decap_6
XANTENNA_ltile_clb_0.mem_fle_3_in_0.LATCH_1_.latch_SLEEPB _378_/Y vgnd vpwr scs8hd_diode_2
XFILLER_60_93 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.mux_fle_3_in_1.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_3_in_1.mux_l1_in_2_.TGATE_3_.scs8hd_ebufn_2/Z
+ ltile_clb_0.mem_fle_3_in_1.LATCH_6_.latch/Q ltile_clb_0.mux_fle_3_in_1.INVTX1_14_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
Xltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_2_.scs8hd_inv_1
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_2_.latch/Q
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_ltile_clb_0.mux_fle_3_in_2.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_3_in_2.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_4_494 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_4_.TGATE_0_.scs8hd_ebufn_2_TEB
+ _613_/Y vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mem_fle_0_in_1.LATCH_0_.latch data_in ltile_clb_0.mem_fle_0_in_1.LATCH_0_.latch/Q
+ _514_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_79_284 vpwr vgnd scs8hd_fill_2
XFILLER_67_402 vpwr vgnd scs8hd_fill_2
XFILLER_67_457 vpwr vgnd scs8hd_fill_2
XFILLER_10_3 vgnd vpwr scs8hd_decap_12
XFILLER_82_416 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.mux_fle_1_in_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_1_in_2.INVTX1_1_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_1_in_2.LATCH_1_.latch/Q ltile_clb_0.mux_fle_1_in_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_82_438 vgnd vpwr scs8hd_decap_12
XFILLER_54_129 vgnd vpwr scs8hd_decap_6
XFILLER_35_321 vpwr vgnd scs8hd_fill_2
XFILLER_62_195 vgnd vpwr scs8hd_fill_1
XFILLER_49_39 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mux_fle_3_in_3.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_3_in_3.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_14_.latch_D
+ data_in vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mem_fle_0_in_1.LATCH_2_.latch_SLEEPB _512_/Y vgnd vpwr scs8hd_diode_2
XFILLER_65_27 vgnd vpwr scs8hd_decap_12
XFILLER_26_332 vpwr vgnd scs8hd_fill_2
XFILLER_81_471 vgnd vpwr scs8hd_decap_12
XFILLER_81_15 vgnd vpwr scs8hd_decap_12
XFILLER_53_173 vgnd vpwr scs8hd_decap_4
XFILLER_26_398 vgnd vpwr scs8hd_fill_1
XFILLER_41_302 vgnd vpwr scs8hd_decap_3
XFILLER_81_59 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.mux_fle_3_in_2.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_3_in_2.INVTX1_13_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_3_in_2.LATCH_1_.latch/Q ltile_clb_0.mux_fle_3_in_2.mux_l1_in_3_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
X_280_ _279_/X _539_/A vgnd vpwr scs8hd_buf_1
XFILLER_41_357 vpwr vgnd scs8hd_fill_2
XFILLER_5_236 vpwr vgnd scs8hd_fill_2
XFILLER_5_258 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_0_in_0.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_0_in_0.INVTX1_12_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__589__B _588_/X vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_0_in_1.INVTX1_5_.scs8hd_inv_1 right_width_0_height_0__pin_5_
+ ltile_clb_0.mux_fle_0_in_1.INVTX1_5_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XFILLER_76_276 vgnd vpwr scs8hd_decap_4
XFILLER_76_265 vpwr vgnd scs8hd_fill_2
XFILLER_76_287 vpwr vgnd scs8hd_fill_2
XFILLER_17_310 vgnd vpwr scs8hd_fill_1
XFILLER_36_129 vgnd vpwr scs8hd_decap_12
XFILLER_17_343 vgnd vpwr scs8hd_decap_3
X_616_ _616_/A _616_/Y vgnd vpwr scs8hd_inv_8
XFILLER_72_482 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_15_.latch
+ data_in ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_15_.latch/Q
+ _582_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
X_547_ _599_/A _526_/X _547_/X vgnd vpwr scs8hd_or2_4
XFILLER_32_302 vgnd vpwr scs8hd_fill_1
XANTENNA_ltile_clb_0.mux_fle_2_in_3.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_2_in_3.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mem_fle_0_in_3.LATCH_3_.latch data_in ltile_clb_0.mem_fle_0_in_3.LATCH_3_.latch/Q
+ _489_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
X_478_ _434_/A _479_/B _478_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA_ltile_clb_0.mux_fle_3_in_0.INVTX1_14_.scs8hd_inv_1_A ltile_clb_0.mux_fle_3_in_0.INVTX1_14_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_58_3 vgnd vpwr scs8hd_decap_12
XANTENNA__499__B _495_/X vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_0_in_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_0_in_1.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_2_in_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_2_in_1.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mem_fle_1_in_3.LATCH_2_.latch data_in ltile_clb_0.mem_fle_1_in_3.LATCH_2_.latch/Q
+ _446_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_67_243 vgnd vpwr scs8hd_fill_1
XFILLER_67_254 vpwr vgnd scs8hd_fill_2
XFILLER_55_416 vgnd vpwr scs8hd_decap_4
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XPHY_809 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xltile_clb_0.mem_fle_2_in_3.LATCH_1_.latch data_in ltile_clb_0.mem_fle_2_in_3.LATCH_1_.latch/Q
+ _394_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_35_195 vpwr vgnd scs8hd_fill_2
XFILLER_50_165 vgnd vpwr scs8hd_decap_8
XANTENNA_ltile_clb_0.mem_fle_1_in_0.LATCH_2_.latch_SLEEPB _479_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_1_in_0.INVTX1_8_.scs8hd_inv_1_A top_width_0_height_0__pin_8_
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_0_in_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_0_in_2.LATCH_5_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_3_.TGATE_0_.scs8hd_ebufn_2_TEB
+ _631_/Y vgnd vpwr scs8hd_diode_2
XFILLER_2_228 vgnd vpwr scs8hd_fill_1
Xltile_clb_0.mem_fle_3_in_3.LATCH_0_.latch data_in ltile_clb_0.mem_fle_3_in_3.LATCH_0_.latch/Q
+ _344_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_76_15 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.buf4_0_.scs8hd_buf_1
+ ltile_clb_0.mux_fle_0_in_0.INVTX1_14_.scs8hd_inv_1/Y _628_/A vgnd vpwr scs8hd_buf_1
Xltile_clb_0.mux_fle_0_in_1.INVTX1_10_.scs8hd_inv_1 bottom_width_0_height_0__pin_10_
+ ltile_clb_0.mux_fle_0_in_1.INVTX1_10_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_2_.TGATE_0_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_2_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_1_in_2.INVTX1_0_.scs8hd_inv_1 top_width_0_height_0__pin_0_ ltile_clb_0.mux_fle_1_in_2.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_73_235 vpwr vgnd scs8hd_fill_2
XFILLER_18_129 vgnd vpwr scs8hd_decap_12
X_401_ _374_/A _399_/B _401_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_61_419 vpwr vgnd scs8hd_fill_2
XPHY_30 vgnd vpwr scs8hd_decap_3
XFILLER_14_335 vgnd vpwr scs8hd_fill_1
XPHY_41 vgnd vpwr scs8hd_decap_3
XPHY_52 vgnd vpwr scs8hd_decap_3
XPHY_63 vgnd vpwr scs8hd_decap_3
XPHY_74 vgnd vpwr scs8hd_decap_3
XFILLER_41_110 vgnd vpwr scs8hd_decap_12
X_332_ _391_/A _338_/B _332_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_25_74 vgnd vpwr scs8hd_decap_12
XFILLER_41_154 vpwr vgnd scs8hd_fill_2
XPHY_85 vgnd vpwr scs8hd_decap_3
XPHY_96 vgnd vpwr scs8hd_decap_3
Xltile_clb_0.mux_fle_2_in_2.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_2_in_2.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2/A
+ ltile_clb_0.mem_fle_2_in_2.LATCH_6_.latch/Q ltile_clb_0.mux_fle_2_in_2.INVTX1_14_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
X_263_ _258_/X _282_/B _282_/C _263_/X vgnd vpwr scs8hd_or3_4
XFILLER_41_51 vgnd vpwr scs8hd_decap_8
XFILLER_41_62 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.mux_fle_0_in_2.INVTX1_9_.scs8hd_inv_1 right_width_0_height_0__pin_9_
+ ltile_clb_0.mux_fle_0_in_2.INVTX1_9_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
Xltile_clb_0.mux_fle_0_in_3.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_0_in_3.INVTX1_1_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_0_in_3.LATCH_1_.latch/Q ltile_clb_0.mux_fle_0_in_3.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_ltile_clb_0.mux_fle_2_in_1.INVTX1_5_.scs8hd_inv_1_A right_width_0_height_0__pin_5_
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_1_in_0.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_1_in_0.INVTX1_12_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_1_in_0.LATCH_0_.latch/Q ltile_clb_0.mux_fle_1_in_0.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_2_56 vgnd vpwr scs8hd_decap_12
XFILLER_49_254 vpwr vgnd scs8hd_fill_2
XFILLER_64_224 vgnd vpwr scs8hd_decap_3
Xltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_15_.scs8hd_inv_1
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_15_.latch/Q
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_15_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
Xltile_clb_0.mux_fle_0_in_2.INVTX1_12_.scs8hd_inv_1 top_width_0_height_0__pin_12_
+ ltile_clb_0.mux_fle_0_in_2.INVTX1_12_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XFILLER_64_279 vgnd vpwr scs8hd_decap_8
XFILLER_17_184 vgnd vpwr scs8hd_decap_4
Xltile_clb_0.mux_fle_3_in_2.INVTX1_11_.scs8hd_inv_1 left_width_0_height_0__pin_11_
+ ltile_clb_0.mux_fle_3_in_2.INVTX1_11_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XFILLER_32_154 vgnd vpwr scs8hd_decap_12
XFILLER_60_496 vgnd vpwr scs8hd_decap_12
XFILLER_60_485 vgnd vpwr scs8hd_decap_8
XFILLER_20_349 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_2_in_3.mux_l1_in_3_.TGATE_2_.scs8hd_ebufn_2_A _651_/HI
+ vgnd vpwr scs8hd_diode_2
XFILLER_9_383 vpwr vgnd scs8hd_fill_2
XANTENNA__303__A _302_/X vgnd vpwr scs8hd_diode_2
XFILLER_55_213 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_0_in_1.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_0_in_1.INVTX1_10_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_2_in_3.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_2_in_3.INVTX1_13_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_2_in_3.LATCH_1_.latch/Q ltile_clb_0.mux_fle_2_in_3.mux_l1_in_3_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_70_205 vgnd vpwr scs8hd_decap_8
XFILLER_70_249 vgnd vpwr scs8hd_decap_3
XFILLER_70_238 vgnd vpwr scs8hd_decap_8
XPHY_617 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_606 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_23_110 vgnd vpwr scs8hd_decap_12
XPHY_639 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_628 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xltile_clb_0.mux_fle_0_in_3.INVTX1_14_.scs8hd_inv_1 ltile_clb_0.mux_fle_0_in_3.INVTX1_14_.scs8hd_inv_1/A
+ ltile_clb_0.mux_fle_0_in_3.INVTX1_14_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XANTENNA_ltile_clb_0.mux_fle_3_in_2.INVTX1_2_.scs8hd_inv_1_A bottom_width_0_height_0__pin_2_
+ vgnd vpwr scs8hd_diode_2
XFILLER_7_309 vgnd vpwr scs8hd_decap_4
Xltile_clb_0.mux_fle_3_in_3.INVTX1_13_.scs8hd_inv_1 right_width_0_height_0__pin_13_
+ ltile_clb_0.mux_fle_3_in_3.INVTX1_13_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XANTENNA_ltile_clb_0.mux_fle_3_in_1.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_3_in_1.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_1_in_3.INVTX1_4_.scs8hd_inv_1 top_width_0_height_0__pin_4_ ltile_clb_0.mux_fle_1_in_3.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_11_98 vgnd vpwr scs8hd_decap_12
XFILLER_78_327 vpwr vgnd scs8hd_fill_2
XFILLER_78_316 vpwr vgnd scs8hd_fill_2
XFILLER_61_205 vpwr vgnd scs8hd_fill_2
XFILLER_61_227 vpwr vgnd scs8hd_fill_2
XFILLER_14_154 vgnd vpwr scs8hd_decap_12
X_315_ address[9] _369_/B vgnd vpwr scs8hd_inv_8
X_246_ _246_/A _286_/A _282_/C _282_/B _246_/X vgnd vpwr scs8hd_or4_4
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.mem_ble4_out_0.LATCH_1_.latch_SLEEPB
+ _550_/Y vgnd vpwr scs8hd_diode_2
XFILLER_77_393 vgnd vpwr scs8hd_decap_4
Xltile_clb_0.mux_fle_0_in_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_0_in_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ ltile_clb_0.mem_fle_0_in_0.LATCH_5_.latch/Q ltile_clb_0.mux_fle_0_in_0.INVTX1_14_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
+ _609_/Y vgnd vpwr scs8hd_diode_2
XFILLER_60_271 vgnd vpwr scs8hd_decap_4
XANTENNA_ltile_clb_0.mem_fle_0_in_0.LATCH_4_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_75_319 vpwr vgnd scs8hd_fill_2
XFILLER_57_39 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_1_.TGATE_1_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_1_.TGATE_1_.scs8hd_ebufn_2/A
+ _632_/Y ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l4_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_68_382 vpwr vgnd scs8hd_fill_2
XFILLER_28_224 vgnd vpwr scs8hd_decap_12
XFILLER_73_27 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mem_fle_0_in_1.LATCH_2_.latch_D data_in vgnd vpwr scs8hd_diode_2
Xltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_5_.TGATE_0_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_10_.scs8hd_inv_1/Y
+ _605_/Y ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_2_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_24_430 vgnd vpwr scs8hd_decap_4
Xltile_clb_0.mux_fle_1_in_3.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_1_in_3.mux_l1_in_2_.TGATE_3_.scs8hd_ebufn_2/Z
+ ltile_clb_0.mem_fle_1_in_3.LATCH_6_.latch/Q ltile_clb_0.mux_fle_1_in_3.INVTX1_14_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XPHY_403 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_414 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_425 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_36_290 vgnd vpwr scs8hd_decap_8
XPHY_436 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_447 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_458 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_11_135 vgnd vpwr scs8hd_decap_12
XPHY_469 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_ltile_clb_0.mux_fle_1_in_3.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_1_in_3.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_3_301 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_2_in_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_2_in_0.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_3_367 vgnd vpwr scs8hd_decap_3
XFILLER_3_356 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.mux_fle_0_in_1.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_0_in_1.INVTX1_12_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_0_in_1.LATCH_0_.latch/Q ltile_clb_0.mux_fle_0_in_1.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_ltile_clb_0.mem_fle_0_in_2.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA__597__B _580_/X vgnd vpwr scs8hd_diode_2
XFILLER_59_382 vpwr vgnd scs8hd_fill_2
XFILLER_74_341 vpwr vgnd scs8hd_fill_2
XFILLER_19_279 vpwr vgnd scs8hd_fill_2
XFILLER_74_385 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.mux_fle_3_in_0.INVTX1_1_.scs8hd_inv_1 right_width_0_height_0__pin_1_
+ ltile_clb_0.mux_fle_3_in_0.INVTX1_1_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XFILLER_27_290 vgnd vpwr scs8hd_decap_4
XFILLER_15_474 vpwr vgnd scs8hd_fill_2
XFILLER_42_271 vgnd vpwr scs8hd_decap_4
XFILLER_8_44 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_2_.scs8hd_inv_1
+ ltile_clb_0.mux_fle_2_in_2.INVTX1_14_.scs8hd_inv_1/Y _617_/A vgnd vpwr scs8hd_inv_1
X_229_ enable _229_/Y vgnd vpwr scs8hd_inv_8
XFILLER_10_190 vgnd vpwr scs8hd_decap_4
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_4_.latch_D
+ data_in vgnd vpwr scs8hd_diode_2
XFILLER_40_3 vgnd vpwr scs8hd_decap_12
XFILLER_69_135 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mux_fle_0_in_2.INVTX1_0_.scs8hd_inv_1_A top_width_0_height_0__pin_0_
+ vgnd vpwr scs8hd_diode_2
XFILLER_77_190 vgnd vpwr scs8hd_fill_1
XANTENNA_ltile_clb_0.mem_fle_1_in_0.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_65_363 vgnd vpwr scs8hd_fill_1
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_2_.TGATE_0_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_2_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_11_.latch_D
+ data_in vgnd vpwr scs8hd_diode_2
XFILLER_21_499 vpwr vgnd scs8hd_fill_2
XFILLER_68_27 vgnd vpwr scs8hd_decap_4
XFILLER_0_337 vpwr vgnd scs8hd_fill_2
XFILLER_48_308 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l4_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
+ _627_/Y vgnd vpwr scs8hd_diode_2
XFILLER_56_363 vgnd vpwr scs8hd_decap_4
X_580_ _579_/X _580_/X vgnd vpwr scs8hd_buf_1
XFILLER_71_333 vgnd vpwr scs8hd_decap_4
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.mem_ble4_out_0.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_3_.scs8hd_inv_1/Y
+ _612_/Y ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XPHY_200 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_16_249 vgnd vpwr scs8hd_decap_6
XFILLER_17_86 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.tap_buf4_0_.scs8hd_inv_1
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.tap_buf4_0_.scs8hd_inv_1/A
+ bottom_width_0_height_0__pin_10_ vgnd vpwr scs8hd_inv_1
XPHY_233 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_222 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_211 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB
+ _605_/Y vgnd vpwr scs8hd_diode_2
XFILLER_24_260 vpwr vgnd scs8hd_fill_2
XPHY_277 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_266 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_255 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_244 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_288 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_8_437 vpwr vgnd scs8hd_fill_2
XPHY_299 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_33_74 vgnd vpwr scs8hd_decap_12
XFILLER_8_448 vgnd vpwr scs8hd_decap_8
Xltile_clb_0.mux_fle_3_in_1.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_3_in_1.INVTX1_7_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_3_in_1.LATCH_3_.latch/Q ltile_clb_0.mux_fle_3_in_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA__401__A _374_/A vgnd vpwr scs8hd_diode_2
XFILLER_66_105 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_15_.scs8hd_inv_1
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_15_.latch/Q
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_15_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_39_319 vgnd vpwr scs8hd_decap_4
XFILLER_58_93 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mux_fle_1_in_3.INVTX1_14_.scs8hd_inv_1_A ltile_clb_0.mux_fle_1_in_3.INVTX1_14_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_3_in_1.INVTX1_5_.scs8hd_inv_1 right_width_0_height_0__pin_5_
+ ltile_clb_0.mux_fle_3_in_1.INVTX1_5_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XFILLER_35_503 vpwr vgnd scs8hd_fill_2
XFILLER_47_341 vpwr vgnd scs8hd_fill_2
XFILLER_47_352 vgnd vpwr scs8hd_decap_4
XFILLER_47_363 vgnd vpwr scs8hd_decap_3
XFILLER_47_374 vpwr vgnd scs8hd_fill_2
XFILLER_62_333 vgnd vpwr scs8hd_decap_3
XFILLER_47_385 vpwr vgnd scs8hd_fill_2
XFILLER_47_396 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_2_in_3.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_2_in_3.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__493__D _345_/A vgnd vpwr scs8hd_diode_2
XFILLER_15_282 vpwr vgnd scs8hd_fill_2
XFILLER_30_274 vgnd vpwr scs8hd_fill_1
XFILLER_30_285 vgnd vpwr scs8hd_decap_4
XFILLER_7_481 vpwr vgnd scs8hd_fill_2
XFILLER_7_470 vpwr vgnd scs8hd_fill_2
XANTENNA__311__A _270_/B vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_2_in_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_2_in_0.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_2_in_2.mux_l1_in_3_.TGATE_2_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_2_in_2.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_3_.scs8hd_inv_1
+ ltile_clb_0.mux_fle_0_in_3.INVTX1_14_.scs8hd_inv_1/Y _635_/A vgnd vpwr scs8hd_inv_1
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_0_.latch_D
+ data_in vgnd vpwr scs8hd_diode_2
XFILLER_38_396 vgnd vpwr scs8hd_fill_1
XFILLER_80_141 vgnd vpwr scs8hd_decap_12
XFILLER_53_344 vgnd vpwr scs8hd_decap_3
XFILLER_79_15 vgnd vpwr scs8hd_decap_12
XFILLER_79_59 vpwr vgnd scs8hd_fill_2
XFILLER_0_156 vgnd vpwr scs8hd_decap_12
XFILLER_48_105 vgnd vpwr scs8hd_decap_12
XANTENNA__578__D _526_/D vgnd vpwr scs8hd_diode_2
XFILLER_48_138 vgnd vpwr scs8hd_decap_4
X_632_ _632_/A _632_/Y vgnd vpwr scs8hd_inv_8
XFILLER_29_374 vpwr vgnd scs8hd_fill_2
XFILLER_29_396 vpwr vgnd scs8hd_fill_2
XFILLER_56_193 vpwr vgnd scs8hd_fill_2
X_563_ _272_/X _564_/B _563_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_32_506 vgnd vpwr scs8hd_decap_8
X_494_ _493_/X _502_/B vgnd vpwr scs8hd_buf_1
XFILLER_44_377 vpwr vgnd scs8hd_fill_2
XFILLER_44_388 vgnd vpwr scs8hd_decap_8
XFILLER_71_196 vgnd vpwr scs8hd_decap_4
XFILLER_12_252 vgnd vpwr scs8hd_decap_4
XFILLER_8_212 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_13_.scs8hd_inv_1_A
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_13_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_8_267 vgnd vpwr scs8hd_decap_8
Xltile_clb_0.mux_fle_3_in_2.INVTX1_9_.scs8hd_inv_1 right_width_0_height_0__pin_9_
+ ltile_clb_0.mux_fle_3_in_2.INVTX1_9_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XFILLER_67_436 vpwr vgnd scs8hd_fill_2
XFILLER_82_428 vgnd vpwr scs8hd_decap_6
XFILLER_35_344 vgnd vpwr scs8hd_decap_3
XFILLER_62_174 vgnd vpwr scs8hd_decap_6
XFILLER_62_163 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
+ _623_/Y vgnd vpwr scs8hd_diode_2
XFILLER_35_377 vpwr vgnd scs8hd_fill_2
XANTENNA__306__A _305_/X vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_0_in_1.INVTX1_9_.scs8hd_inv_1_A right_width_0_height_0__pin_9_
+ vgnd vpwr scs8hd_diode_2
XFILLER_58_425 vgnd vpwr scs8hd_decap_4
XANTENNA_ltile_clb_0.mem_fle_1_in_2.LATCH_6_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_65_39 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mux_fle_1_in_1.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_1_in_1.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_73_439 vpwr vgnd scs8hd_fill_2
XFILLER_73_428 vpwr vgnd scs8hd_fill_2
XFILLER_26_322 vgnd vpwr scs8hd_decap_3
XFILLER_38_171 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mux_fle_2_in_0.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_2_in_0.INVTX1_10_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_38_193 vgnd vpwr scs8hd_decap_3
XFILLER_81_483 vgnd vpwr scs8hd_decap_4
XFILLER_81_27 vgnd vpwr scs8hd_decap_12
XFILLER_26_366 vgnd vpwr scs8hd_fill_1
XFILLER_14_32 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.mux_fle_2_in_2.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_2_in_2.INVTX1_7_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_2_in_2.LATCH_3_.latch/Q ltile_clb_0.mux_fle_2_in_2.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_ltile_clb_0.mem_fle_1_in_3.LATCH_4_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_0_.TGATE_1_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.mem_ble4_out_0.LATCH_1_.latch_D
+ data_in vgnd vpwr scs8hd_diode_2
XFILLER_1_443 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_2_.TGATE_0_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_2_.TGATE_0_.scs8hd_ebufn_2/A
+ _623_/Y ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_1_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_39_51 vgnd vpwr scs8hd_decap_8
XFILLER_39_62 vgnd vpwr scs8hd_decap_12
XFILLER_64_406 vgnd vpwr scs8hd_decap_4
XFILLER_17_322 vpwr vgnd scs8hd_fill_2
XFILLER_29_171 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_1_in_2.INVTX1_6_.scs8hd_inv_1_A bottom_width_0_height_0__pin_6_
+ vgnd vpwr scs8hd_diode_2
XFILLER_72_450 vgnd vpwr scs8hd_decap_8
XANTENNA_ltile_clb_0.mem_fle_2_in_0.LATCH_6_.latch_D data_in vgnd vpwr scs8hd_diode_2
X_615_ _615_/A _615_/Y vgnd vpwr scs8hd_inv_8
XFILLER_29_193 vgnd vpwr scs8hd_decap_4
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.mem_ble4_out_0.LATCH_1_.latch_SLEEPB
+ _576_/Y vgnd vpwr scs8hd_diode_2
XFILLER_44_141 vpwr vgnd scs8hd_fill_2
XFILLER_17_377 vpwr vgnd scs8hd_fill_2
XFILLER_17_388 vpwr vgnd scs8hd_fill_2
X_546_ _546_/A _528_/X _546_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_32_314 vgnd vpwr scs8hd_decap_4
XFILLER_72_494 vgnd vpwr scs8hd_decap_12
XFILLER_44_196 vpwr vgnd scs8hd_fill_2
XFILLER_32_369 vpwr vgnd scs8hd_fill_2
X_477_ _433_/A _479_/B _477_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA_ltile_clb_0.mem_fle_2_in_1.LATCH_4_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_67_211 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.buf4_2_.scs8hd_buf_1_A
+ ltile_clb_0.mux_fle_0_in_2.INVTX1_14_.scs8hd_inv_1/Y vgnd vpwr scs8hd_diode_2
XFILLER_55_428 vgnd vpwr scs8hd_decap_4
XFILLER_48_491 vgnd vpwr scs8hd_decap_3
XFILLER_23_358 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mem_fle_2_in_2.LATCH_2_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_3_in_2.INVTX1_12_.scs8hd_inv_1_A top_width_0_height_0__pin_12_
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_2_in_3.INVTX1_3_.scs8hd_inv_1_A left_width_0_height_0__pin_3_
+ vgnd vpwr scs8hd_diode_2
XFILLER_76_27 vgnd vpwr scs8hd_decap_4
XFILLER_58_244 vgnd vpwr scs8hd_decap_4
XFILLER_46_406 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mem_fle_2_in_3.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_73_269 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_2_in_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_2_in_2.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
X_400_ _326_/A _399_/B _400_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_54_472 vgnd vpwr scs8hd_fill_1
XPHY_20 vgnd vpwr scs8hd_decap_3
XPHY_31 vgnd vpwr scs8hd_decap_3
XFILLER_26_141 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_0_.scs8hd_inv_1_A
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_14_325 vpwr vgnd scs8hd_fill_2
XPHY_42 vgnd vpwr scs8hd_decap_3
XPHY_53 vgnd vpwr scs8hd_decap_3
XPHY_64 vgnd vpwr scs8hd_decap_3
X_331_ _331_/A _391_/A vgnd vpwr scs8hd_buf_1
XFILLER_25_86 vgnd vpwr scs8hd_decap_12
XPHY_75 vgnd vpwr scs8hd_decap_3
XPHY_86 vgnd vpwr scs8hd_decap_3
XPHY_97 vgnd vpwr scs8hd_decap_3
X_262_ _248_/A _261_/X _262_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_22_391 vgnd vpwr scs8hd_decap_6
XFILLER_41_74 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mem_fle_3_in_0.LATCH_2_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_2_in_1.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_2_in_1.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_1_251 vpwr vgnd scs8hd_fill_2
XFILLER_1_240 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.mem_ble4_out_0.LATCH_1_.latch
+ data_in ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.mem_ble4_out_0.LATCH_1_.latch/Q
+ _550_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_49_222 vpwr vgnd scs8hd_fill_2
XFILLER_2_68 vgnd vpwr scs8hd_decap_12
XFILLER_37_428 vgnd vpwr scs8hd_decap_4
XFILLER_49_277 vpwr vgnd scs8hd_fill_2
XFILLER_66_93 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.mux_fle_2_in_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_2_in_0.INVTX1_1_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_2_in_0.LATCH_1_.latch/Q ltile_clb_0.mux_fle_2_in_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
Xltile_clb_0.mux_fle_0_in_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_0_in_0.INVTX1_6_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_0_in_0.LATCH_2_.latch/Q ltile_clb_0.mux_fle_0_in_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_ltile_clb_0.mem_fle_3_in_1.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
Xltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_5_.scs8hd_inv_1
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_5_.latch/Q
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
X_529_ _528_/X _529_/X vgnd vpwr scs8hd_buf_1
XFILLER_32_166 vgnd vpwr scs8hd_decap_4
XFILLER_70_3 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_6_.latch_D
+ data_in vgnd vpwr scs8hd_diode_2
XFILLER_55_203 vgnd vpwr scs8hd_decap_3
XFILLER_28_428 vgnd vpwr scs8hd_fill_1
XFILLER_55_236 vgnd vpwr scs8hd_decap_4
XPHY_607 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_51_420 vgnd vpwr scs8hd_decap_4
XPHY_629 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xltile_clb_0.mux_fle_1_in_3.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_1_in_3.INVTX1_7_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_1_in_3.LATCH_3_.latch/Q ltile_clb_0.mux_fle_1_in_3.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XPHY_618 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xltile_clb_0.mux_fle_3_in_3.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_3_in_3.INVTX1_2_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_3_in_3.LATCH_2_.latch/Q ltile_clb_0.mux_fle_3_in_3.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_11_306 vgnd vpwr scs8hd_decap_3
XFILLER_23_188 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
+ _636_/HI ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.mem_ble4_out_0.LATCH_2_.latch/Q
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_15_.latch_SLEEPB
+ _582_/Y vgnd vpwr scs8hd_diode_2
XFILLER_46_225 vgnd vpwr scs8hd_decap_4
XFILLER_42_431 vpwr vgnd scs8hd_fill_2
XFILLER_54_291 vgnd vpwr scs8hd_decap_4
XFILLER_14_166 vgnd vpwr scs8hd_decap_12
X_314_ _314_/A _388_/A vgnd vpwr scs8hd_buf_1
XANTENNA_ltile_clb_0.mux_fle_1_in_0.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_1_in_0.INVTX1_12_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
X_245_ address[0] _282_/C vgnd vpwr scs8hd_buf_1
XFILLER_10_361 vpwr vgnd scs8hd_fill_2
XANTENNA__404__A _338_/A vgnd vpwr scs8hd_diode_2
Xltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_4_.latch
+ data_in ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_4_.latch/Q
+ _292_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
Xltile_clb_0.mux_fle_1_in_0.INVTX1_0_.scs8hd_inv_1 top_width_0_height_0__pin_0_ ltile_clb_0.mux_fle_1_in_0.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_69_317 vpwr vgnd scs8hd_fill_2
XFILLER_69_306 vgnd vpwr scs8hd_decap_8
XFILLER_69_339 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_1_in_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_1_in_0.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_3_in_3.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_3_in_3.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__ff_0.DFFSRQ_0_.dff
+ clkbuf_1_0_0_clk/X ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.INVTX1_1_.scs8hd_inv_1/A
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.INVTX1_0_.scs8hd_inv_1/A
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__ff_0.DFFSRQ_0_.dff/QN
+ reset set vgnd vpwr scs8hd_dfbbp_1
XFILLER_37_203 vpwr vgnd scs8hd_fill_2
XFILLER_37_214 vgnd vpwr scs8hd_decap_6
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_6_.TGATE_1_.scs8hd_ebufn_2_TEB
+ _604_/Y vgnd vpwr scs8hd_diode_2
XFILLER_37_236 vpwr vgnd scs8hd_fill_2
XFILLER_80_515 vgnd vpwr scs8hd_fill_1
XFILLER_52_206 vgnd vpwr scs8hd_decap_3
XANTENNA_ltile_clb_0.mux_fle_1_in_1.INVTX1_11_.scs8hd_inv_1_A left_width_0_height_0__pin_11_
+ vgnd vpwr scs8hd_diode_2
XFILLER_45_280 vpwr vgnd scs8hd_fill_2
XFILLER_33_464 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.mux_fle_0_in_0.INVTX1_9_.scs8hd_inv_1 right_width_0_height_0__pin_9_
+ ltile_clb_0.mux_fle_0_in_0.INVTX1_9_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XANTENNA_ltile_clb_0.mux_fle_1_in_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_1_in_1.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_0_.TGATE_1_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XANTENNA__314__A _314_/A vgnd vpwr scs8hd_diode_2
XFILLER_73_39 vgnd vpwr scs8hd_decap_12
XFILLER_43_239 vgnd vpwr scs8hd_decap_4
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_2_.latch_D
+ data_in vgnd vpwr scs8hd_diode_2
XPHY_404 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_415 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_426 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_51_261 vgnd vpwr scs8hd_decap_6
XPHY_437 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_448 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_459 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_11_147 vgnd vpwr scs8hd_decap_12
XFILLER_22_32 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.mux_fle_3_in_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_3_in_0.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2/Z
+ ltile_clb_0.mem_fle_3_in_0.LATCH_6_.latch/Q ltile_clb_0.mux_fle_3_in_0.INVTX1_14_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_3_335 vpwr vgnd scs8hd_fill_2
XFILLER_0_3 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_3_.latch_SLEEPB
+ _595_/Y vgnd vpwr scs8hd_diode_2
XFILLER_66_309 vgnd vpwr scs8hd_decap_8
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_2_.scs8hd_inv_1_A
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_19_203 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.mux_fle_1_in_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_1_in_1.INVTX1_1_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_1_in_1.LATCH_1_.latch/Q ltile_clb_0.mux_fle_1_in_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_47_51 vgnd vpwr scs8hd_decap_8
XFILLER_47_62 vgnd vpwr scs8hd_decap_12
XFILLER_62_515 vgnd vpwr scs8hd_fill_1
XFILLER_30_456 vpwr vgnd scs8hd_fill_2
XFILLER_8_56 vgnd vpwr scs8hd_decap_12
XFILLER_30_467 vgnd vpwr scs8hd_decap_8
Xltile_clb_0.mux_fle_1_in_1.INVTX1_4_.scs8hd_inv_1 top_width_0_height_0__pin_4_ ltile_clb_0.mux_fle_1_in_1.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
X_228_ _227_/X _228_/X vgnd vpwr scs8hd_buf_1
XANTENNA_ltile_clb_0.mux_fle_3_in_3.INVTX1_9_.scs8hd_inv_1_A right_width_0_height_0__pin_9_
+ vgnd vpwr scs8hd_diode_2
XFILLER_33_3 vgnd vpwr scs8hd_decap_12
XFILLER_69_158 vgnd vpwr scs8hd_decap_3
XFILLER_69_147 vgnd vpwr scs8hd_decap_4
XFILLER_80_312 vgnd vpwr scs8hd_decap_3
XANTENNA_ltile_clb_0.mem_fle_3_in_3.LATCH_6_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_65_397 vpwr vgnd scs8hd_fill_2
XFILLER_65_386 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_25_239 vpwr vgnd scs8hd_fill_2
XFILLER_80_367 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mux_fle_3_in_3.mux_l1_in_3_.TGATE_2_.scs8hd_ebufn_2_A _655_/HI
+ vgnd vpwr scs8hd_diode_2
XFILLER_18_280 vpwr vgnd scs8hd_fill_2
XFILLER_18_291 vgnd vpwr scs8hd_decap_4
XANTENNA__309__A _308_/X vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_3_in_1.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_3_in_1.INVTX1_13_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_3_in_1.LATCH_1_.latch/Q ltile_clb_0.mux_fle_3_in_1.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_21_401 vpwr vgnd scs8hd_fill_2
XFILLER_21_412 vpwr vgnd scs8hd_fill_2
XFILLER_40_209 vgnd vpwr scs8hd_decap_4
XANTENNA_ltile_clb_0.mux_fle_1_in_3.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_1_in_3.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_21_489 vgnd vpwr scs8hd_decap_3
XANTENNA_ltile_clb_0.mux_fle_2_in_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_2_in_0.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_1_in_1.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_1_in_1.INVTX1_10_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_7_.TGATE_0_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_14_.scs8hd_inv_1/Y
+ _613_/Y ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_3_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_56_353 vgnd vpwr scs8hd_fill_1
XFILLER_44_504 vgnd vpwr scs8hd_decap_12
XFILLER_71_301 vpwr vgnd scs8hd_fill_2
XFILLER_56_386 vpwr vgnd scs8hd_fill_2
XFILLER_16_239 vgnd vpwr scs8hd_decap_3
XFILLER_71_367 vpwr vgnd scs8hd_fill_2
XPHY_201 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_17_98 vgnd vpwr scs8hd_decap_12
XPHY_234 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_223 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_212 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_272 vgnd vpwr scs8hd_decap_3
XPHY_267 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_256 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_245 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_4_.latch
+ data_in ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_4_.latch/Q
+ _594_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XPHY_289 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_278 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_8_405 vgnd vpwr scs8hd_fill_1
XFILLER_33_86 vgnd vpwr scs8hd_decap_12
XFILLER_3_110 vgnd vpwr scs8hd_decap_12
XFILLER_79_423 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.mem_ble4_out_0.LATCH_1_.latch_SLEEPB
+ _602_/Y vgnd vpwr scs8hd_diode_2
XANTENNA__401__B _399_/B vgnd vpwr scs8hd_diode_2
XFILLER_79_489 vgnd vpwr scs8hd_decap_12
XFILLER_66_117 vgnd vpwr scs8hd_decap_12
XFILLER_74_183 vgnd vpwr scs8hd_fill_1
XFILLER_62_312 vgnd vpwr scs8hd_decap_4
XFILLER_35_515 vgnd vpwr scs8hd_fill_1
XFILLER_74_93 vgnd vpwr scs8hd_decap_12
XFILLER_62_345 vpwr vgnd scs8hd_fill_2
XFILLER_62_389 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_3_in_1.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_3_in_1.LATCH_6_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_22_209 vgnd vpwr scs8hd_decap_3
Xltile_clb_0.mux_fle_1_in_2.INVTX1_8_.scs8hd_inv_1 top_width_0_height_0__pin_8_ ltile_clb_0.mux_fle_1_in_2.INVTX1_8_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XPHY_790 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_30_297 vgnd vpwr scs8hd_decap_6
Xltile_clb_0.mem_fle_3_in_0.LATCH_7_.latch data_in ltile_clb_0.mem_fle_3_in_0.LATCH_7_.latch/Q
+ _372_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA__311__B _309_/X vgnd vpwr scs8hd_diode_2
Xltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.mem_ble4_out_0.LATCH_1_.latch
+ data_in ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.mem_ble4_out_0.LATCH_1_.latch/Q
+ _602_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_26_504 vgnd vpwr scs8hd_decap_12
XFILLER_38_364 vgnd vpwr scs8hd_decap_3
XFILLER_53_301 vpwr vgnd scs8hd_fill_2
XFILLER_38_375 vgnd vpwr scs8hd_decap_4
XANTENNA_ltile_clb_0.mem_fle_3_in_3.LATCH_2_.latch_SLEEPB _338_/Y vgnd vpwr scs8hd_diode_2
XFILLER_53_378 vgnd vpwr scs8hd_decap_4
Xltile_clb_0.mux_fle_2_in_1.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_2_in_1.mux_l1_in_2_.TGATE_3_.scs8hd_ebufn_2/Z
+ ltile_clb_0.mem_fle_2_in_1.LATCH_6_.latch/Q ltile_clb_0.mux_fle_2_in_1.INVTX1_14_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_5_.TGATE_1_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_11_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_21_242 vpwr vgnd scs8hd_fill_2
XFILLER_21_275 vpwr vgnd scs8hd_fill_2
XFILLER_5_419 vpwr vgnd scs8hd_fill_2
XFILLER_79_27 vgnd vpwr scs8hd_decap_12
XANTENNA__502__A _423_/A vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_0_in_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_0_in_2.INVTX1_1_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_0_in_2.LATCH_1_.latch/Q ltile_clb_0.mux_fle_0_in_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_76_426 vgnd vpwr scs8hd_decap_8
XFILLER_76_415 vpwr vgnd scs8hd_fill_2
XFILLER_0_168 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_7_.scs8hd_inv_1/Y
+ _620_/Y ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_1_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_48_117 vgnd vpwr scs8hd_decap_12
XFILLER_76_437 vgnd vpwr scs8hd_decap_4
X_631_ _631_/A _631_/Y vgnd vpwr scs8hd_inv_8
XFILLER_29_331 vpwr vgnd scs8hd_fill_2
XFILLER_29_342 vpwr vgnd scs8hd_fill_2
XFILLER_17_515 vgnd vpwr scs8hd_fill_1
X_562_ _554_/X _564_/B vgnd vpwr scs8hd_buf_1
XANTENNA_ltile_clb_0.mux_fle_0_in_3.INVTX1_7_.scs8hd_inv_1_A left_width_0_height_0__pin_7_
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_2_in_3.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_2_in_3.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_44_345 vgnd vpwr scs8hd_decap_4
XFILLER_71_175 vpwr vgnd scs8hd_fill_2
X_493_ _380_/X _427_/B _228_/X _345_/A _493_/X vgnd vpwr scs8hd_or4_4
Xltile_clb_0.mux_fle_2_in_3.INVTX1_3_.scs8hd_inv_1 left_width_0_height_0__pin_3_ ltile_clb_0.mux_fle_2_in_3.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_ltile_clb_0.mux_fle_1_in_0.INVTX1_3_.scs8hd_inv_1_A left_width_0_height_0__pin_3_
+ vgnd vpwr scs8hd_diode_2
XFILLER_8_224 vgnd vpwr scs8hd_decap_6
XANTENNA__412__A _430_/A vgnd vpwr scs8hd_diode_2
XFILLER_79_220 vgnd vpwr scs8hd_decap_12
XFILLER_79_297 vpwr vgnd scs8hd_fill_2
XFILLER_75_481 vgnd vpwr scs8hd_decap_6
Xltile_clb_0.mux_fle_2_in_2.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_2_in_2.INVTX1_13_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_2_in_2.LATCH_1_.latch/Q ltile_clb_0.mux_fle_2_in_2.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_35_301 vpwr vgnd scs8hd_fill_2
XFILLER_47_161 vgnd vpwr scs8hd_decap_3
XFILLER_35_367 vgnd vpwr scs8hd_fill_1
XFILLER_50_337 vpwr vgnd scs8hd_fill_2
XANTENNA__322__A _341_/B vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_2_in_1.INVTX1_0_.scs8hd_inv_1_A top_width_0_height_0__pin_0_
+ vgnd vpwr scs8hd_diode_2
XFILLER_58_415 vgnd vpwr scs8hd_decap_6
XFILLER_58_448 vgnd vpwr scs8hd_fill_1
XFILLER_58_459 vgnd vpwr scs8hd_decap_3
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_15_.scs8hd_inv_1_A
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_15_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_4_.latch
+ data_in ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_4_.latch/Q
+ _568_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_53_131 vpwr vgnd scs8hd_fill_2
XFILLER_38_183 vgnd vpwr scs8hd_fill_1
XFILLER_53_153 vpwr vgnd scs8hd_fill_2
XFILLER_53_142 vpwr vgnd scs8hd_fill_2
XFILLER_14_507 vgnd vpwr scs8hd_decap_8
XFILLER_81_39 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.mux_fle_2_in_1.INVTX1_11_.scs8hd_inv_1 left_width_0_height_0__pin_11_
+ ltile_clb_0.mux_fle_2_in_1.INVTX1_11_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XFILLER_53_197 vgnd vpwr scs8hd_decap_3
XFILLER_14_44 vgnd vpwr scs8hd_decap_12
XFILLER_30_32 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_0_.scs8hd_inv_1_A
+ ltile_clb_0.mux_fle_0_in_0.INVTX1_14_.scs8hd_inv_1/Y vgnd vpwr scs8hd_diode_2
XFILLER_1_400 vpwr vgnd scs8hd_fill_2
XANTENNA__232__A address[4] vgnd vpwr scs8hd_diode_2
XFILLER_1_477 vgnd vpwr scs8hd_decap_8
XFILLER_76_234 vgnd vpwr scs8hd_decap_12
XFILLER_76_223 vpwr vgnd scs8hd_fill_2
XFILLER_76_212 vpwr vgnd scs8hd_fill_2
XFILLER_39_74 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mem_fle_1_in_3.LATCH_3_.latch_SLEEPB _445_/Y vgnd vpwr scs8hd_diode_2
XFILLER_17_301 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_0_in_1.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_0_in_1.INVTX1_12_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_72_440 vgnd vpwr scs8hd_fill_1
XFILLER_55_62 vgnd vpwr scs8hd_decap_12
XFILLER_55_51 vgnd vpwr scs8hd_decap_8
X_614_ _614_/A _614_/Y vgnd vpwr scs8hd_inv_8
XFILLER_72_462 vpwr vgnd scs8hd_fill_2
XFILLER_17_367 vgnd vpwr scs8hd_fill_1
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
X_545_ _545_/A _528_/X _545_/Y vgnd vpwr scs8hd_nor2_4
Xltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_0_.TGATE_1_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ _616_/Y ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l4_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_ltile_clb_0.mux_fle_1_in_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_1_in_2.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_44_175 vgnd vpwr scs8hd_fill_1
XFILLER_44_186 vgnd vpwr scs8hd_fill_1
X_476_ _432_/A _479_/B _476_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_32_359 vgnd vpwr scs8hd_decap_3
XANTENNA__407__A _314_/A vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_2_in_2.INVTX1_13_.scs8hd_inv_1 right_width_0_height_0__pin_13_
+ ltile_clb_0.mux_fle_2_in_2.INVTX1_13_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__ff_0.DFFSRQ_0_.dff_D
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.INVTX1_1_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_4_293 vgnd vpwr scs8hd_fill_1
XFILLER_67_245 vgnd vpwr scs8hd_decap_4
XANTENNA_ltile_clb_0.mux_fle_1_in_1.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_1_in_1.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_48_470 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_0_in_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_0_in_2.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_35_153 vgnd vpwr scs8hd_fill_1
XFILLER_35_164 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.mux_fle_1_in_2.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_1_in_2.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2/Z
+ ltile_clb_0.mem_fle_1_in_2.LATCH_6_.latch/Q ltile_clb_0.mux_fle_1_in_2.INVTX1_14_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_63_484 vpwr vgnd scs8hd_fill_2
XFILLER_35_175 vpwr vgnd scs8hd_fill_2
XANTENNA__317__A _380_/A vgnd vpwr scs8hd_diode_2
XFILLER_50_145 vgnd vpwr scs8hd_decap_6
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_14_.latch_SLEEPB
+ _557_/Y vgnd vpwr scs8hd_diode_2
XFILLER_50_178 vgnd vpwr scs8hd_decap_6
Xltile_clb_0.mux_fle_3_in_0.INVTX1_9_.scs8hd_inv_1 right_width_0_height_0__pin_9_
+ ltile_clb_0.mux_fle_3_in_0.INVTX1_9_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XANTENNA_ltile_clb_0.mux_fle_3_in_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_3_in_0.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_14_.latch_D
+ data_in vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_0_in_0.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_0_in_0.INVTX1_12_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_0_in_0.LATCH_0_.latch/Q ltile_clb_0.mux_fle_0_in_0.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_58_223 vgnd vpwr scs8hd_decap_12
XFILLER_58_289 vgnd vpwr scs8hd_decap_4
XFILLER_39_481 vgnd vpwr scs8hd_decap_4
XFILLER_39_492 vpwr vgnd scs8hd_fill_2
XPHY_21 vgnd vpwr scs8hd_decap_3
XPHY_10 vgnd vpwr scs8hd_decap_3
XFILLER_81_281 vgnd vpwr scs8hd_decap_8
XFILLER_14_337 vpwr vgnd scs8hd_fill_2
XPHY_32 vgnd vpwr scs8hd_decap_3
XPHY_43 vgnd vpwr scs8hd_decap_3
XPHY_54 vgnd vpwr scs8hd_decap_3
X_330_ _330_/A _331_/A vgnd vpwr scs8hd_buf_1
XPHY_65 vgnd vpwr scs8hd_decap_3
XFILLER_41_123 vgnd vpwr scs8hd_decap_12
XANTENNA__227__A address[8] vgnd vpwr scs8hd_diode_2
XPHY_76 vgnd vpwr scs8hd_decap_3
XPHY_87 vgnd vpwr scs8hd_decap_3
XPHY_98 vgnd vpwr scs8hd_decap_3
X_261_ _260_/X _261_/X vgnd vpwr scs8hd_buf_1
XFILLER_25_98 vgnd vpwr scs8hd_decap_12
XFILLER_6_503 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mem_fle_2_in_2.LATCH_3_.latch_SLEEPB _403_/Y vgnd vpwr scs8hd_diode_2
XFILLER_41_86 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.mux_fle_1_in_3.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_1_in_3.INVTX1_13_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_1_in_3.LATCH_1_.latch/Q ltile_clb_0.mux_fle_1_in_3.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
Xltile_clb_0.mux_fle_3_in_3.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_3_in_3.INVTX1_8_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_3_in_3.LATCH_0_.latch/Q ltile_clb_0.mux_fle_3_in_3.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_49_245 vpwr vgnd scs8hd_fill_2
XFILLER_64_248 vpwr vgnd scs8hd_fill_2
XFILLER_45_484 vpwr vgnd scs8hd_fill_2
X_528_ _528_/A _528_/X vgnd vpwr scs8hd_buf_1
XFILLER_20_307 vpwr vgnd scs8hd_fill_2
XFILLER_20_329 vgnd vpwr scs8hd_decap_6
X_459_ _437_/A _450_/X _459_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_9_352 vpwr vgnd scs8hd_fill_2
XFILLER_13_392 vgnd vpwr scs8hd_decap_4
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_5_.TGATE_1_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_11_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_63_3 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_4_.latch
+ data_in ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_4_.latch/Q
+ _542_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA__600__A _599_/X vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_0_in_0.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_0_in_0.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_63_281 vgnd vpwr scs8hd_decap_8
XPHY_608 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_36_473 vgnd vpwr scs8hd_decap_6
XPHY_619 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_51_465 vgnd vpwr scs8hd_decap_4
XFILLER_51_443 vpwr vgnd scs8hd_fill_2
XFILLER_23_123 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mux_fle_0_in_2.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_0_in_2.INVTX1_10_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_2_in_0.INVTX1_9_.scs8hd_inv_1_A right_width_0_height_0__pin_9_
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_3_in_0.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_3_in_0.INVTX1_7_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_3_in_0.LATCH_3_.latch/Q ltile_clb_0.mux_fle_3_in_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_ltile_clb_0.mux_fle_2_in_1.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_2_in_1.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_3_in_0.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_3_in_0.INVTX1_10_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__510__A _331_/A vgnd vpwr scs8hd_diode_2
XFILLER_46_215 vgnd vpwr scs8hd_fill_1
XFILLER_46_248 vgnd vpwr scs8hd_decap_8
XANTENNA_ltile_clb_0.mem_fle_3_in_1.LATCH_3_.latch_SLEEPB _365_/Y vgnd vpwr scs8hd_diode_2
XFILLER_27_473 vgnd vpwr scs8hd_fill_1
XFILLER_27_484 vgnd vpwr scs8hd_decap_4
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.mem_ble4_out_0.LATCH_1_.latch_SLEEPB
+ _311_/Y vgnd vpwr scs8hd_diode_2
X_313_ _313_/A _314_/A vgnd vpwr scs8hd_buf_1
X_244_ _248_/A _556_/A _244_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_1_.scs8hd_inv_1_A
+ ltile_clb_0.mux_fle_3_in_1.INVTX1_14_.scs8hd_inv_1/Y vgnd vpwr scs8hd_diode_2
XFILLER_10_384 vgnd vpwr scs8hd_decap_3
XANTENNA__404__B _399_/B vgnd vpwr scs8hd_diode_2
XFILLER_6_377 vgnd vpwr scs8hd_decap_4
XANTENNA_ltile_clb_0.mux_fle_3_in_3.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_3_in_3.LATCH_5_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_6_388 vgnd vpwr scs8hd_fill_1
XANTENNA__420__A _434_/A vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_0_in_3.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_0_in_3.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2/Z
+ ltile_clb_0.mem_fle_0_in_3.LATCH_6_.latch/Q ltile_clb_0.mux_fle_0_in_3.INVTX1_14_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_ltile_clb_0.mux_fle_3_in_1.INVTX1_6_.scs8hd_inv_1_A bottom_width_0_height_0__pin_6_
+ vgnd vpwr scs8hd_diode_2
XFILLER_18_462 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_0_.scs8hd_inv_1
+ ltile_clb_0.mux_fle_3_in_0.INVTX1_14_.scs8hd_inv_1/Y _605_/A vgnd vpwr scs8hd_inv_1
XFILLER_37_259 vpwr vgnd scs8hd_fill_2
XFILLER_60_240 vgnd vpwr scs8hd_decap_8
XFILLER_33_443 vpwr vgnd scs8hd_fill_2
XFILLER_33_498 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mem_fle_0_in_2.LATCH_4_.latch_SLEEPB _499_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_3_.TGATE_1_.scs8hd_ebufn_2_TEB
+ _614_/Y vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mem_fle_0_in_1.LATCH_6_.latch data_in ltile_clb_0.mem_fle_0_in_1.LATCH_6_.latch/Q
+ _508_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_9_171 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_1_.TGATE_1_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_1_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_0_509 vgnd vpwr scs8hd_decap_6
XANTENNA__330__A _330_/A vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_2_in_3.INVTX1_14_.scs8hd_inv_1_A ltile_clb_0.mux_fle_2_in_3.INVTX1_14_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mem_fle_1_in_1.LATCH_5_.latch data_in ltile_clb_0.mem_fle_1_in_1.LATCH_5_.latch/Q
+ _465_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_68_351 vgnd vpwr scs8hd_decap_3
XFILLER_56_513 vgnd vpwr scs8hd_decap_3
XFILLER_43_218 vpwr vgnd scs8hd_fill_2
XPHY_405 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_416 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_427 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_438 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_449 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xltile_clb_0.mem_fle_2_in_1.LATCH_4_.latch data_in ltile_clb_0.mem_fle_2_in_1.LATCH_4_.latch/Q
+ _418_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_51_295 vpwr vgnd scs8hd_fill_2
XFILLER_51_284 vpwr vgnd scs8hd_fill_2
XFILLER_24_498 vgnd vpwr scs8hd_decap_4
XFILLER_11_159 vgnd vpwr scs8hd_decap_12
XFILLER_22_44 vgnd vpwr scs8hd_decap_12
XANTENNA__505__A _504_/X vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_0_in_3.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_0_in_3.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_1_in_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_1_in_0.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__240__A address[0] vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mem_fle_3_in_1.LATCH_3_.latch data_in ltile_clb_0.mem_fle_3_in_1.LATCH_3_.latch/Q
+ _365_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_59_362 vpwr vgnd scs8hd_fill_2
XFILLER_47_502 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_7_.TGATE_0_.scs8hd_ebufn_2_TEB
+ _605_/Y vgnd vpwr scs8hd_diode_2
XFILLER_74_354 vgnd vpwr scs8hd_decap_8
XFILLER_19_248 vpwr vgnd scs8hd_fill_2
XFILLER_19_259 vpwr vgnd scs8hd_fill_2
XFILLER_34_207 vgnd vpwr scs8hd_decap_6
XFILLER_47_74 vgnd vpwr scs8hd_decap_12
XFILLER_15_410 vpwr vgnd scs8hd_fill_2
XFILLER_63_51 vgnd vpwr scs8hd_decap_8
XFILLER_15_443 vgnd vpwr scs8hd_decap_6
XFILLER_15_454 vgnd vpwr scs8hd_decap_4
XFILLER_63_62 vgnd vpwr scs8hd_decap_12
XFILLER_15_498 vgnd vpwr scs8hd_decap_12
XFILLER_30_446 vgnd vpwr scs8hd_decap_8
X_227_ address[8] address[9] _227_/X vgnd vpwr scs8hd_or2_4
XFILLER_8_68 vgnd vpwr scs8hd_decap_12
XANTENNA__415__A _328_/A vgnd vpwr scs8hd_diode_2
XFILLER_6_141 vgnd vpwr scs8hd_decap_12
XFILLER_26_3 vgnd vpwr scs8hd_decap_12
XFILLER_38_502 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mem_fle_1_in_1.LATCH_4_.latch_SLEEPB _466_/Y vgnd vpwr scs8hd_diode_2
XFILLER_65_332 vgnd vpwr scs8hd_decap_4
XFILLER_80_324 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_1_.TGATE_0_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2/Z
+ _607_/Y ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_25_207 vgnd vpwr scs8hd_fill_1
XFILLER_25_229 vgnd vpwr scs8hd_decap_3
XFILLER_80_346 vgnd vpwr scs8hd_decap_8
XFILLER_80_379 vgnd vpwr scs8hd_fill_1
XFILLER_21_424 vgnd vpwr scs8hd_decap_3
XFILLER_21_435 vgnd vpwr scs8hd_decap_3
XFILLER_33_284 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.mux_fle_2_in_1.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_2_in_1.INVTX1_7_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_2_in_1.LATCH_3_.latch/Q ltile_clb_0.mux_fle_2_in_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_ltile_clb_0.mux_fle_2_in_1.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_2_in_1.LATCH_7_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__325__A _325_/A vgnd vpwr scs8hd_diode_2
Xltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_1_.scs8hd_inv_1
+ ltile_clb_0.mux_fle_1_in_1.INVTX1_14_.scs8hd_inv_1/Y _623_/A vgnd vpwr scs8hd_inv_1
XFILLER_0_306 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.mem_fle_2_in_3.LATCH_7_.latch data_in ltile_clb_0.mem_fle_2_in_3.LATCH_7_.latch/Q
+ _388_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_29_502 vgnd vpwr scs8hd_decap_12
XFILLER_56_332 vpwr vgnd scs8hd_fill_2
XFILLER_68_192 vgnd vpwr scs8hd_decap_3
XPHY_224 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_213 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_202 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_268 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_257 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_246 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_235 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_6_.latch_SLEEPB
+ _540_/Y vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mem_fle_3_in_3.LATCH_6_.latch data_in ltile_clb_0.mem_fle_3_in_3.LATCH_6_.latch/Q
+ _326_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XPHY_279 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_12_468 vpwr vgnd scs8hd_fill_2
XANTENNA__235__A address[3] vgnd vpwr scs8hd_diode_2
XFILLER_33_98 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mux_fle_0_in_1.INVTX1_4_.scs8hd_inv_1_A top_width_0_height_0__pin_4_
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_0_in_3.INVTX1_2_.scs8hd_inv_1 bottom_width_0_height_0__pin_2_
+ ltile_clb_0.mux_fle_0_in_3.INVTX1_2_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XFILLER_79_457 vpwr vgnd scs8hd_fill_2
XFILLER_79_468 vpwr vgnd scs8hd_fill_2
XFILLER_66_129 vpwr vgnd scs8hd_fill_2
XFILLER_59_192 vpwr vgnd scs8hd_fill_2
XFILLER_74_162 vgnd vpwr scs8hd_decap_4
XANTENNA_ltile_clb_0.mux_fle_2_in_0.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_2_in_0.INVTX1_12_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_62_379 vgnd vpwr scs8hd_fill_1
XFILLER_15_251 vpwr vgnd scs8hd_fill_2
XPHY_780 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_30_243 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_1_in_3.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_1_in_3.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XPHY_791 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_ltile_clb_0.mem_fle_2_in_0.LATCH_4_.latch_SLEEPB _433_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_0_in_2.INVTX1_13_.scs8hd_inv_1_A right_width_0_height_0__pin_13_
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_11_.latch_D
+ data_in vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_1_in_2.INVTX1_1_.scs8hd_inv_1_A right_width_0_height_0__pin_1_
+ vgnd vpwr scs8hd_diode_2
XFILLER_38_354 vgnd vpwr scs8hd_fill_1
XFILLER_53_324 vgnd vpwr scs8hd_decap_4
XFILLER_65_195 vgnd vpwr scs8hd_decap_3
XFILLER_80_154 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mux_fle_2_in_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_2_in_1.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_21_210 vgnd vpwr scs8hd_decap_4
XFILLER_21_221 vpwr vgnd scs8hd_fill_2
XFILLER_21_298 vpwr vgnd scs8hd_fill_2
XFILLER_79_39 vgnd vpwr scs8hd_decap_12
XANTENNA__502__B _502_/B vgnd vpwr scs8hd_diode_2
XFILLER_0_125 vgnd vpwr scs8hd_decap_12
XFILLER_28_32 vgnd vpwr scs8hd_decap_12
XFILLER_48_129 vgnd vpwr scs8hd_decap_3
X_630_ _630_/A _630_/Y vgnd vpwr scs8hd_inv_8
X_561_ _535_/A _558_/B _561_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_29_365 vgnd vpwr scs8hd_fill_1
XFILLER_71_110 vgnd vpwr scs8hd_decap_12
XFILLER_56_184 vgnd vpwr scs8hd_decap_3
X_492_ _343_/A _492_/B _492_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_52_390 vgnd vpwr scs8hd_decap_6
XFILLER_12_287 vpwr vgnd scs8hd_fill_2
XFILLER_8_247 vgnd vpwr scs8hd_decap_4
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_15_.scs8hd_inv_1_A
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_15_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__412__B _412_/B vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_13_.latch_SLEEPB
+ _532_/Y vgnd vpwr scs8hd_diode_2
XFILLER_79_232 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_1_.TGATE_1_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_1_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_67_449 vgnd vpwr scs8hd_decap_6
XFILLER_47_151 vgnd vpwr scs8hd_decap_4
XFILLER_47_195 vpwr vgnd scs8hd_fill_2
XFILLER_62_198 vgnd vpwr scs8hd_fill_1
Xltile_clb_0.mux_fle_1_in_2.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_1_in_2.INVTX1_7_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_1_in_2.LATCH_3_.latch/Q ltile_clb_0.mux_fle_1_in_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_50_316 vgnd vpwr scs8hd_decap_3
Xltile_clb_0.mux_fle_3_in_2.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_3_in_2.INVTX1_2_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_3_in_2.LATCH_2_.latch/Q ltile_clb_0.mux_fle_3_in_2.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_43_390 vgnd vpwr scs8hd_decap_6
Xltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_2_.scs8hd_inv_1/Y
+ _629_/Y ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_ltile_clb_0.mux_fle_0_in_2.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_0_in_2.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2_TEB
+ _628_/Y vgnd vpwr scs8hd_diode_2
XANTENNA__603__A _603_/A vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l4_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
+ _610_/Y vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_1_in_0.INVTX1_8_.scs8hd_inv_1 top_width_0_height_0__pin_8_ ltile_clb_0.mux_fle_1_in_0.INVTX1_8_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
Xltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.buf4_3_.scs8hd_buf_1
+ ltile_clb_0.mux_fle_2_in_3.INVTX1_14_.scs8hd_inv_1/Y _618_/A vgnd vpwr scs8hd_buf_1
XFILLER_73_419 vpwr vgnd scs8hd_fill_2
XFILLER_26_302 vgnd vpwr scs8hd_fill_1
XFILLER_53_110 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mux_fle_0_in_1.mux_l1_in_2_.TGATE_3_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_0_in_1.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_26_357 vpwr vgnd scs8hd_fill_2
XFILLER_26_379 vgnd vpwr scs8hd_decap_4
XANTENNA_ltile_clb_0.mem_fle_0_in_0.LATCH_5_.latch_SLEEPB _520_/Y vgnd vpwr scs8hd_diode_2
XFILLER_41_327 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_2_in_1.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_2_in_1.INVTX1_10_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_14_56 vgnd vpwr scs8hd_decap_12
XFILLER_30_44 vgnd vpwr scs8hd_decap_12
XANTENNA__513__A _423_/A vgnd vpwr scs8hd_diode_2
Xltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_5_.TGATE_1_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_11_.scs8hd_inv_1/Y
+ _628_/Y ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_5_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA__232__B _231_/X vgnd vpwr scs8hd_diode_2
XFILLER_1_423 vpwr vgnd scs8hd_fill_2
XFILLER_1_456 vpwr vgnd scs8hd_fill_2
XFILLER_1_489 vgnd vpwr scs8hd_decap_12
XFILLER_76_246 vgnd vpwr scs8hd_decap_12
XFILLER_39_86 vgnd vpwr scs8hd_decap_12
XFILLER_57_460 vpwr vgnd scs8hd_fill_2
X_613_ _613_/A _613_/Y vgnd vpwr scs8hd_inv_8
XFILLER_57_482 vgnd vpwr scs8hd_fill_1
XFILLER_55_74 vgnd vpwr scs8hd_decap_12
XFILLER_17_357 vpwr vgnd scs8hd_fill_2
X_544_ _544_/A _528_/X _544_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_44_165 vpwr vgnd scs8hd_fill_2
X_475_ _431_/A _479_/B _475_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_71_62 vgnd vpwr scs8hd_decap_12
XFILLER_71_51 vgnd vpwr scs8hd_decap_8
XFILLER_40_393 vgnd vpwr scs8hd_decap_4
XANTENNA__423__A _423_/A vgnd vpwr scs8hd_diode_2
XFILLER_4_261 vgnd vpwr scs8hd_decap_3
Xltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_1_.scs8hd_inv_1
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_1_.latch/Q
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_67_224 vpwr vgnd scs8hd_fill_2
XFILLER_67_202 vgnd vpwr scs8hd_decap_6
XFILLER_67_235 vpwr vgnd scs8hd_fill_2
XFILLER_67_279 vpwr vgnd scs8hd_fill_2
XFILLER_82_249 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.mux_fle_2_in_1.INVTX1_3_.scs8hd_inv_1 left_width_0_height_0__pin_3_ ltile_clb_0.mux_fle_2_in_1.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_35_110 vgnd vpwr scs8hd_decap_12
XFILLER_63_463 vpwr vgnd scs8hd_fill_2
XFILLER_63_452 vpwr vgnd scs8hd_fill_2
XFILLER_63_441 vpwr vgnd scs8hd_fill_2
XFILLER_63_496 vgnd vpwr scs8hd_decap_12
XFILLER_35_187 vpwr vgnd scs8hd_fill_2
XFILLER_50_135 vgnd vpwr scs8hd_fill_1
XANTENNA__317__B address[7] vgnd vpwr scs8hd_diode_2
XFILLER_31_382 vgnd vpwr scs8hd_decap_4
XANTENNA__333__A _333_/A vgnd vpwr scs8hd_diode_2
XFILLER_58_202 vgnd vpwr scs8hd_fill_1
Xltile_clb_0.mux_fle_1_in_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_1_in_0.INVTX1_1_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_1_in_0.LATCH_1_.latch/Q ltile_clb_0.mux_fle_1_in_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
Xltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_12_.scs8hd_inv_1
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_12_.latch/Q
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_12_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_ltile_clb_0.mux_fle_2_in_1.INVTX1_11_.scs8hd_inv_1_A left_width_0_height_0__pin_11_
+ vgnd vpwr scs8hd_diode_2
XFILLER_39_471 vgnd vpwr scs8hd_decap_3
XFILLER_66_290 vgnd vpwr scs8hd_decap_4
XFILLER_54_452 vgnd vpwr scs8hd_fill_1
XPHY_22 vgnd vpwr scs8hd_decap_3
XPHY_11 vgnd vpwr scs8hd_decap_3
XFILLER_26_154 vgnd vpwr scs8hd_decap_12
XFILLER_54_496 vgnd vpwr scs8hd_decap_12
XFILLER_54_485 vgnd vpwr scs8hd_decap_4
XPHY_33 vgnd vpwr scs8hd_decap_3
XPHY_44 vgnd vpwr scs8hd_decap_3
XANTENNA__508__A _325_/A vgnd vpwr scs8hd_diode_2
XPHY_55 vgnd vpwr scs8hd_decap_3
XANTENNA_ltile_clb_0.mux_fle_1_in_2.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_1_in_2.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XPHY_66 vgnd vpwr scs8hd_decap_3
XPHY_77 vgnd vpwr scs8hd_decap_3
XFILLER_41_135 vgnd vpwr scs8hd_decap_12
XPHY_88 vgnd vpwr scs8hd_decap_3
XANTENNA__227__B address[9] vgnd vpwr scs8hd_diode_2
X_260_ _236_/X _333_/A _260_/X vgnd vpwr scs8hd_or2_4
XFILLER_22_360 vpwr vgnd scs8hd_fill_2
XFILLER_22_371 vpwr vgnd scs8hd_fill_2
XFILLER_41_179 vpwr vgnd scs8hd_fill_2
XPHY_99 vgnd vpwr scs8hd_decap_3
XFILLER_22_382 vpwr vgnd scs8hd_fill_2
XFILLER_6_515 vgnd vpwr scs8hd_fill_1
XANTENNA__243__A _242_/X vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mem_fle_0_in_2.LATCH_2_.latch data_in ltile_clb_0.mem_fle_0_in_2.LATCH_2_.latch/Q
+ _501_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_41_98 vgnd vpwr scs8hd_decap_12
XFILLER_2_15 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mux_fle_1_in_1.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_1_in_1.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_1_297 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
+ _606_/Y vgnd vpwr scs8hd_diode_2
XFILLER_37_419 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.mem_fle_1_in_2.LATCH_1_.latch data_in ltile_clb_0.mem_fle_1_in_2.LATCH_1_.latch/Q
+ _458_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_17_110 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.mux_fle_0_in_3.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_0_in_3.INVTX1_7_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_0_in_3.LATCH_3_.latch/Q ltile_clb_0.mux_fle_0_in_3.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
Xltile_clb_0.mux_fle_2_in_3.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_2_in_3.INVTX1_2_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_2_in_3.LATCH_2_.latch/Q ltile_clb_0.mux_fle_2_in_3.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_ltile_clb_0.mux_fle_2_in_2.INVTX1_7_.scs8hd_inv_1_A left_width_0_height_0__pin_7_
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_3_in_0.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_3_in_0.INVTX1_13_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_3_in_0.LATCH_1_.latch/Q ltile_clb_0.mux_fle_3_in_0.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_72_271 vgnd vpwr scs8hd_decap_4
XANTENNA__418__A _433_/A vgnd vpwr scs8hd_diode_2
XFILLER_17_176 vgnd vpwr scs8hd_decap_6
X_527_ address[4] _526_/X _528_/A vgnd vpwr scs8hd_or2_4
XFILLER_45_474 vgnd vpwr scs8hd_decap_3
XFILLER_60_444 vgnd vpwr scs8hd_decap_12
XFILLER_82_94 vgnd vpwr scs8hd_decap_12
X_458_ _436_/A _450_/X _458_/Y vgnd vpwr scs8hd_nor2_4
X_389_ _326_/A _388_/B _389_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_9_331 vgnd vpwr scs8hd_decap_6
XFILLER_13_371 vgnd vpwr scs8hd_decap_4
Xltile_clb_0.mem_fle_2_in_2.LATCH_0_.latch data_in ltile_clb_0.mem_fle_2_in_2.LATCH_0_.latch/Q
+ _406_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_56_3 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_12_.latch
+ data_in ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_12_.latch/Q
+ _533_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
Xltile_clb_0.mux_fle_2_in_2.INVTX1_7_.scs8hd_inv_1 left_width_0_height_0__pin_7_ ltile_clb_0.mux_fle_2_in_2.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_ltile_clb_0.mux_fle_2_in_3.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_2_in_3.LATCH_6_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_3_in_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_3_in_0.LATCH_4_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_55_249 vpwr vgnd scs8hd_fill_2
XANTENNA__328__A _328_/A vgnd vpwr scs8hd_diode_2
XPHY_609 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_23_135 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_6_.scs8hd_inv_1
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_6_.latch/Q
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_ltile_clb_0.mux_fle_3_in_3.INVTX1_4_.scs8hd_inv_1_A top_width_0_height_0__pin_4_
+ vgnd vpwr scs8hd_diode_2
XFILLER_78_308 vgnd vpwr scs8hd_decap_8
XFILLER_59_500 vgnd vpwr scs8hd_decap_12
XANTENNA__510__B _511_/B vgnd vpwr scs8hd_diode_2
XFILLER_19_419 vpwr vgnd scs8hd_fill_2
XFILLER_27_452 vpwr vgnd scs8hd_fill_2
XFILLER_36_32 vgnd vpwr scs8hd_decap_12
XANTENNA__238__A address[1] vgnd vpwr scs8hd_diode_2
XFILLER_27_496 vgnd vpwr scs8hd_decap_12
X_312_ _603_/A _309_/X _312_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_42_488 vpwr vgnd scs8hd_fill_2
X_243_ _242_/X _556_/A vgnd vpwr scs8hd_buf_1
XFILLER_42_499 vgnd vpwr scs8hd_decap_12
XFILLER_10_330 vgnd vpwr scs8hd_decap_6
XANTENNA_ltile_clb_0.mux_fle_1_in_1.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_1_in_1.INVTX1_12_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__420__B _412_/B vgnd vpwr scs8hd_diode_2
XFILLER_77_363 vgnd vpwr scs8hd_decap_3
Xltile_clb_0.mux_fle_3_in_3.INVTX1_2_.scs8hd_inv_1 bottom_width_0_height_0__pin_2_
+ ltile_clb_0.mux_fle_3_in_3.INVTX1_2_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XANTENNA_ltile_clb_0.mux_fle_0_in_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_0_in_0.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_33_400 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_5_.scs8hd_inv_1/Y
+ _604_/Y ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
Xltile_clb_0.mux_fle_2_in_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_2_in_0.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2/Z
+ ltile_clb_0.mem_fle_2_in_0.LATCH_6_.latch/Q ltile_clb_0.mux_fle_2_in_0.INVTX1_14_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_20_105 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mux_fle_0_in_0.INVTX1_10_.scs8hd_inv_1_A bottom_width_0_height_0__pin_10_
+ vgnd vpwr scs8hd_diode_2
XANTENNA__611__A _611_/A vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_0_in_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_0_in_1.INVTX1_1_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_0_in_1.LATCH_1_.latch/Q ltile_clb_0.mux_fle_0_in_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_ltile_clb_0.mux_fle_1_in_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_1_in_2.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
+ _624_/Y vgnd vpwr scs8hd_diode_2
XFILLER_68_396 vgnd vpwr scs8hd_fill_1
XFILLER_24_411 vgnd vpwr scs8hd_decap_8
XPHY_406 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_417 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_428 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_439 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xltile_clb_0.mux_fle_3_in_3.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_3_in_3.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2/Z
+ ltile_clb_0.mem_fle_3_in_3.LATCH_7_.latch/Q ltile_clb_0.mux_fle_3_in_3.INVTX1_14_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_22_56 vgnd vpwr scs8hd_decap_12
XFILLER_3_315 vgnd vpwr scs8hd_decap_4
Xltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.buf4_0_.scs8hd_buf_1
+ ltile_clb_0.mux_fle_1_in_0.INVTX1_14_.scs8hd_inv_1/Y _620_/A vgnd vpwr scs8hd_buf_1
XANTENNA__521__A _331_/A vgnd vpwr scs8hd_diode_2
XFILLER_78_105 vgnd vpwr scs8hd_decap_12
XFILLER_59_352 vpwr vgnd scs8hd_fill_2
XFILLER_47_514 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.mux_fle_2_in_1.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_2_in_1.INVTX1_13_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_2_in_1.LATCH_1_.latch/Q ltile_clb_0.mux_fle_2_in_1.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_19_238 vgnd vpwr scs8hd_decap_6
XFILLER_47_86 vgnd vpwr scs8hd_decap_12
XFILLER_74_377 vgnd vpwr scs8hd_decap_4
XFILLER_63_74 vgnd vpwr scs8hd_decap_12
X_226_ address[7] _226_/X vgnd vpwr scs8hd_buf_1
XANTENNA__431__A _431_/A vgnd vpwr scs8hd_diode_2
XFILLER_77_171 vgnd vpwr scs8hd_decap_12
XFILLER_19_3 vgnd vpwr scs8hd_decap_12
XFILLER_38_514 vpwr vgnd scs8hd_fill_2
XFILLER_65_355 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_0_in_3.INVTX1_2_.scs8hd_inv_1_A bottom_width_0_height_0__pin_2_
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_0_in_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_0_in_0.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_33_252 vgnd vpwr scs8hd_decap_8
XFILLER_33_263 vpwr vgnd scs8hd_fill_2
XANTENNA__606__A _606_/A vgnd vpwr scs8hd_diode_2
XFILLER_21_458 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_0_in_3.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_0_in_3.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__341__A _394_/A vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_1_in_0.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_1_in_0.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_12_.scs8hd_inv_1
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_12_.latch/Q
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_12_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_29_514 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_1_in_2.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_1_in_2.INVTX1_10_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_71_314 vpwr vgnd scs8hd_fill_2
XFILLER_16_208 vgnd vpwr scs8hd_fill_1
XFILLER_16_219 vpwr vgnd scs8hd_fill_2
XFILLER_71_358 vpwr vgnd scs8hd_fill_2
XPHY_225 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_214 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_203 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_12_436 vgnd vpwr scs8hd_decap_3
XPHY_258 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_247 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_236 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_285 vpwr vgnd scs8hd_fill_2
XANTENNA__516__A _516_/A vgnd vpwr scs8hd_diode_2
XPHY_269 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_4_.latch_SLEEPB
+ _292_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__251__A _248_/A vgnd vpwr scs8hd_diode_2
XFILLER_3_123 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_10_.scs8hd_inv_1_A
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_10_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_59_160 vpwr vgnd scs8hd_fill_2
XFILLER_47_322 vpwr vgnd scs8hd_fill_2
XFILLER_74_141 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
+ _620_/Y vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_1_in_1.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_1_in_1.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2/A
+ ltile_clb_0.mem_fle_1_in_1.LATCH_6_.latch/Q ltile_clb_0.mux_fle_1_in_1.INVTX1_14_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_62_325 vgnd vpwr scs8hd_decap_8
Xltile_clb_0.mux_fle_1_in_0.INVTX1_11_.scs8hd_inv_1 left_width_0_height_0__pin_11_
+ ltile_clb_0.mux_fle_1_in_0.INVTX1_11_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XFILLER_70_380 vgnd vpwr scs8hd_decap_4
XFILLER_30_200 vgnd vpwr scs8hd_decap_3
XPHY_781 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_770 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__426__A _437_/A vgnd vpwr scs8hd_diode_2
XFILLER_30_233 vgnd vpwr scs8hd_fill_1
XFILLER_30_255 vgnd vpwr scs8hd_decap_3
XPHY_792 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_3_.TGATE_0_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_6_.TGATE_1_.scs8hd_ebufn_2/Z
+ _615_/Y ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_1_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_78_480 vgnd vpwr scs8hd_decap_12
XFILLER_38_300 vgnd vpwr scs8hd_decap_6
XFILLER_38_388 vpwr vgnd scs8hd_fill_2
XFILLER_80_166 vgnd vpwr scs8hd_decap_12
XFILLER_53_358 vgnd vpwr scs8hd_decap_4
XFILLER_61_380 vpwr vgnd scs8hd_fill_2
XANTENNA__336__A _263_/X vgnd vpwr scs8hd_diode_2
XFILLER_21_266 vpwr vgnd scs8hd_fill_2
XFILLER_21_288 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.mux_fle_1_in_1.INVTX1_13_.scs8hd_inv_1 right_width_0_height_0__pin_13_
+ ltile_clb_0.mux_fle_1_in_1.INVTX1_13_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XFILLER_0_137 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.mux_fle_1_in_2.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_1_in_2.INVTX1_13_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_1_in_2.LATCH_1_.latch/Q ltile_clb_0.mux_fle_1_in_2.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
Xltile_clb_0.mux_fle_3_in_2.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_3_in_2.INVTX1_8_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_3_in_2.LATCH_0_.latch/Q ltile_clb_0.mux_fle_3_in_2.mux_l1_in_2_.TGATE_3_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_7_.scs8hd_inv_1_A
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_7_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_28_44 vgnd vpwr scs8hd_decap_12
XFILLER_56_163 vgnd vpwr scs8hd_decap_8
X_560_ _261_/X _558_/B _560_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_71_155 vgnd vpwr scs8hd_fill_1
XFILLER_44_32 vgnd vpwr scs8hd_decap_12
XFILLER_44_358 vpwr vgnd scs8hd_fill_2
X_491_ _423_/A _492_/B _491_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA_ltile_clb_0.mux_fle_1_in_3.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_1_in_3.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__246__A _246_/A vgnd vpwr scs8hd_diode_2
XFILLER_8_204 vgnd vpwr scs8hd_decap_8
XFILLER_5_15 vgnd vpwr scs8hd_decap_12
XFILLER_4_410 vpwr vgnd scs8hd_fill_2
XFILLER_5_59 vpwr vgnd scs8hd_fill_2
XFILLER_69_62 vgnd vpwr scs8hd_decap_12
XFILLER_69_51 vgnd vpwr scs8hd_decap_8
XFILLER_67_406 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_67_428 vgnd vpwr scs8hd_fill_1
XFILLER_75_461 vpwr vgnd scs8hd_fill_2
XFILLER_75_450 vpwr vgnd scs8hd_fill_2
XFILLER_35_325 vgnd vpwr scs8hd_decap_4
XFILLER_35_358 vpwr vgnd scs8hd_fill_2
XFILLER_50_328 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.mux_fle_0_in_1.INVTX1_2_.scs8hd_inv_1 bottom_width_0_height_0__pin_2_
+ ltile_clb_0.mux_fle_0_in_1.INVTX1_2_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
Xltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_10_.latch
+ data_in ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_10_.latch/Q
+ _587_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_7_292 vgnd vpwr scs8hd_decap_4
XANTENNA__603__B _600_/X vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__ff_0.DFFSRQ_0_.dff_SETB
+ set vgnd vpwr scs8hd_diode_2
XFILLER_66_450 vgnd vpwr scs8hd_decap_8
XFILLER_38_141 vgnd vpwr scs8hd_fill_1
XFILLER_26_314 vgnd vpwr scs8hd_decap_8
XFILLER_53_166 vgnd vpwr scs8hd_decap_4
Xltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l4_in_0_.TGATE_0_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l4_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ _611_/Y ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_16_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_26_369 vgnd vpwr scs8hd_fill_1
XFILLER_41_306 vpwr vgnd scs8hd_fill_2
XFILLER_14_68 vgnd vpwr scs8hd_decap_12
XFILLER_30_56 vgnd vpwr scs8hd_decap_12
XANTENNA__513__B _514_/B vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
+ _636_/HI vgnd vpwr scs8hd_diode_2
XFILLER_49_406 vpwr vgnd scs8hd_fill_2
XFILLER_49_417 vgnd vpwr scs8hd_decap_4
XFILLER_49_439 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.mux_fle_0_in_2.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_0_in_2.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2/Z
+ ltile_clb_0.mem_fle_0_in_2.LATCH_6_.latch/Q ltile_clb_0.mux_fle_0_in_2.INVTX1_14_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_39_98 vgnd vpwr scs8hd_decap_12
XFILLER_76_269 vgnd vpwr scs8hd_decap_6
X_612_ _612_/A _612_/Y vgnd vpwr scs8hd_inv_8
XFILLER_72_420 vgnd vpwr scs8hd_fill_1
XFILLER_55_86 vgnd vpwr scs8hd_decap_12
X_543_ _569_/A _528_/X _543_/Y vgnd vpwr scs8hd_nor2_4
X_474_ _430_/A _479_/B _474_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_32_328 vgnd vpwr scs8hd_decap_8
XANTENNA_ltile_clb_0.mux_fle_1_in_3.INVTX1_8_.scs8hd_inv_1_A top_width_0_height_0__pin_8_
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_0_in_2.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_0_in_2.INVTX1_12_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_71_74 vgnd vpwr scs8hd_decap_12
XFILLER_9_502 vpwr vgnd scs8hd_fill_2
XFILLER_40_350 vgnd vpwr scs8hd_decap_8
XFILLER_40_372 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_0_in_2.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_0_in_2.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_4_.TGATE_0_.scs8hd_ebufn_2_TEB
+ _629_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_2_in_0.INVTX1_4_.scs8hd_inv_1_A top_width_0_height_0__pin_4_
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_3_in_0.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_3_in_0.INVTX1_12_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_67_258 vpwr vgnd scs8hd_fill_2
XFILLER_63_420 vgnd vpwr scs8hd_decap_4
XANTENNA_ltile_clb_0.mux_fle_0_in_1.mux_l1_in_3_.TGATE_2_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_0_in_1.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_23_317 vgnd vpwr scs8hd_decap_6
XFILLER_23_328 vpwr vgnd scs8hd_fill_2
XFILLER_35_199 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.mux_fle_0_in_2.INVTX1_6_.scs8hd_inv_1 bottom_width_0_height_0__pin_6_
+ ltile_clb_0.mux_fle_0_in_2.INVTX1_6_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XFILLER_31_350 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_0_in_3.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_0_in_3.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__614__A _614_/A vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mem_fle_0_in_0.LATCH_7_.latch_D data_in vgnd vpwr scs8hd_diode_2
Xltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_12_.scs8hd_inv_1
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_12_.latch/Q
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_12_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
Xltile_clb_0.mux_fle_0_in_3.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_0_in_3.INVTX1_13_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_0_in_3.LATCH_1_.latch/Q ltile_clb_0.mux_fle_0_in_3.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
Xltile_clb_0.mux_fle_2_in_3.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_2_in_3.INVTX1_8_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_2_in_3.LATCH_0_.latch/Q ltile_clb_0.mux_fle_2_in_3.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_6_80 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_3_in_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_3_in_1.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_3_in_1.INVTX1_1_.scs8hd_inv_1_A right_width_0_height_0__pin_1_
+ vgnd vpwr scs8hd_diode_2
XFILLER_73_239 vpwr vgnd scs8hd_fill_2
XFILLER_54_431 vgnd vpwr scs8hd_decap_3
XPHY_12 vgnd vpwr scs8hd_decap_3
XANTENNA_ltile_clb_0.mux_fle_1_in_3.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_1_in_3.LATCH_7_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_2_in_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_2_in_0.LATCH_5_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_54_475 vgnd vpwr scs8hd_fill_1
XPHY_23 vgnd vpwr scs8hd_decap_3
XPHY_34 vgnd vpwr scs8hd_decap_3
XPHY_45 vgnd vpwr scs8hd_decap_3
XFILLER_26_166 vgnd vpwr scs8hd_decap_3
XANTENNA__508__B _511_/B vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mem_fle_0_in_1.LATCH_5_.latch_D data_in vgnd vpwr scs8hd_diode_2
XPHY_56 vgnd vpwr scs8hd_decap_3
XFILLER_81_294 vpwr vgnd scs8hd_fill_2
XPHY_67 vgnd vpwr scs8hd_decap_3
XPHY_78 vgnd vpwr scs8hd_decap_3
XFILLER_41_147 vpwr vgnd scs8hd_fill_2
XPHY_89 vgnd vpwr scs8hd_decap_3
XFILLER_41_158 vpwr vgnd scs8hd_fill_2
XANTENNA__524__A _423_/A vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_9_.scs8hd_inv_1_A
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_9_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_3_in_3.INVTX1_14_.scs8hd_inv_1_A ltile_clb_0.mux_fle_3_in_3.INVTX1_14_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_1_221 vpwr vgnd scs8hd_fill_2
XFILLER_77_501 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mem_fle_0_in_2.LATCH_3_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_2_27 vgnd vpwr scs8hd_decap_4
XFILLER_49_236 vpwr vgnd scs8hd_fill_2
XFILLER_64_206 vgnd vpwr scs8hd_decap_8
Xltile_clb_0.mux_fle_0_in_3.INVTX1_11_.scs8hd_inv_1 left_width_0_height_0__pin_11_
+ ltile_clb_0.mux_fle_0_in_3.INVTX1_11_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XFILLER_49_258 vpwr vgnd scs8hd_fill_2
XFILLER_45_420 vgnd vpwr scs8hd_decap_4
XFILLER_57_291 vpwr vgnd scs8hd_fill_2
XFILLER_45_453 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.mux_fle_3_in_3.INVTX1_10_.scs8hd_inv_1 bottom_width_0_height_0__pin_10_
+ ltile_clb_0.mux_fle_3_in_3.INVTX1_10_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XANTENNA__418__B _412_/B vgnd vpwr scs8hd_diode_2
XFILLER_60_412 vpwr vgnd scs8hd_fill_2
X_526_ _380_/A address[7] _228_/X _526_/D _526_/X vgnd vpwr scs8hd_or4_4
XFILLER_72_283 vgnd vpwr scs8hd_decap_3
XFILLER_60_456 vpwr vgnd scs8hd_fill_2
X_457_ _435_/A _451_/X _457_/Y vgnd vpwr scs8hd_nor2_4
X_388_ _388_/A _388_/B _388_/Y vgnd vpwr scs8hd_nor2_4
Xltile_clb_0.mux_fle_2_in_0.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_2_in_0.INVTX1_7_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_2_in_0.LATCH_3_.latch/Q ltile_clb_0.mux_fle_2_in_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
Xltile_clb_0.mux_fle_1_in_3.INVTX1_1_.scs8hd_inv_1 right_width_0_height_0__pin_1_
+ ltile_clb_0.mux_fle_1_in_3.INVTX1_1_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XANTENNA__434__A _434_/A vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mem_fle_0_in_3.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_9_387 vgnd vpwr scs8hd_decap_3
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_7_.latch_D
+ data_in vgnd vpwr scs8hd_diode_2
XFILLER_49_3 vgnd vpwr scs8hd_decap_12
XFILLER_28_409 vpwr vgnd scs8hd_fill_2
XFILLER_55_228 vpwr vgnd scs8hd_fill_2
XANTENNA__609__A _609_/A vgnd vpwr scs8hd_diode_2
XFILLER_36_453 vpwr vgnd scs8hd_fill_2
XFILLER_48_291 vgnd vpwr scs8hd_decap_3
XANTENNA_ltile_clb_0.mem_fle_1_in_0.LATCH_3_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_63_294 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_14_.latch_D
+ data_in vgnd vpwr scs8hd_diode_2
XFILLER_23_147 vgnd vpwr scs8hd_decap_12
XFILLER_51_489 vpwr vgnd scs8hd_fill_2
XANTENNA__344__A _379_/A vgnd vpwr scs8hd_diode_2
Xltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_0_.TGATE_0_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ _633_/Y ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l4_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_ltile_clb_0.mux_fle_0_in_3.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_0_in_3.INVTX1_10_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mem_fle_1_in_1.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_59_512 vgnd vpwr scs8hd_decap_4
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB
+ _607_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_74_504 vgnd vpwr scs8hd_decap_12
XFILLER_46_206 vgnd vpwr scs8hd_decap_8
XFILLER_27_431 vpwr vgnd scs8hd_fill_2
XFILLER_36_44 vgnd vpwr scs8hd_decap_12
XANTENNA__519__A _325_/A vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_3_in_1.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_3_in_1.INVTX1_10_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_61_209 vgnd vpwr scs8hd_decap_3
XFILLER_42_401 vpwr vgnd scs8hd_fill_2
XFILLER_42_423 vgnd vpwr scs8hd_decap_8
XFILLER_52_32 vgnd vpwr scs8hd_decap_12
X_311_ _270_/B _309_/X _311_/Y vgnd vpwr scs8hd_nor2_4
X_242_ _236_/X _313_/A _242_/X vgnd vpwr scs8hd_or2_4
XFILLER_10_342 vpwr vgnd scs8hd_fill_2
XANTENNA__254__A _286_/A vgnd vpwr scs8hd_diode_2
XFILLER_6_346 vgnd vpwr scs8hd_decap_3
XFILLER_77_62 vgnd vpwr scs8hd_decap_12
XFILLER_77_51 vgnd vpwr scs8hd_decap_8
XFILLER_77_397 vgnd vpwr scs8hd_fill_1
XFILLER_80_507 vgnd vpwr scs8hd_decap_8
XANTENNA__429__A _428_/X vgnd vpwr scs8hd_diode_2
XFILLER_18_453 vgnd vpwr scs8hd_decap_4
XFILLER_33_423 vpwr vgnd scs8hd_fill_2
X_509_ _328_/A _511_/B _509_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_20_117 vgnd vpwr scs8hd_decap_12
XFILLER_13_180 vgnd vpwr scs8hd_decap_3
XFILLER_9_184 vgnd vpwr scs8hd_decap_12
XFILLER_68_386 vpwr vgnd scs8hd_fill_2
XFILLER_28_206 vgnd vpwr scs8hd_decap_8
XANTENNA__339__A _339_/A vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_3_.latch_D
+ data_in vgnd vpwr scs8hd_diode_2
XFILLER_24_434 vgnd vpwr scs8hd_fill_1
XPHY_407 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_36_283 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_0_in_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_0_in_1.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_51_242 vpwr vgnd scs8hd_fill_2
XPHY_418 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_429 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_13_.latch_SLEEPB
+ _251_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_1_in_2.INVTX1_13_.scs8hd_inv_1_A right_width_0_height_0__pin_13_
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_2_in_0.INVTX1_7_.scs8hd_inv_1 left_width_0_height_0__pin_7_ ltile_clb_0.mux_fle_2_in_0.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_22_68 vgnd vpwr scs8hd_decap_12
XANTENNA__521__B _517_/X vgnd vpwr scs8hd_diode_2
XFILLER_78_117 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_0_.scs8hd_inv_1/Y
+ _613_/Y ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_59_331 vpwr vgnd scs8hd_fill_2
XFILLER_59_320 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_0_in_0.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_0_in_0.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_59_386 vgnd vpwr scs8hd_decap_3
XFILLER_19_217 vgnd vpwr scs8hd_decap_6
XFILLER_62_507 vgnd vpwr scs8hd_decap_8
XANTENNA__249__A _246_/A vgnd vpwr scs8hd_diode_2
XFILLER_47_98 vgnd vpwr scs8hd_decap_12
XFILLER_74_389 vgnd vpwr scs8hd_decap_8
XANTENNA_ltile_clb_0.mux_fle_3_in_1.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_3_in_1.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_1_.scs8hd_inv_1_A
+ ltile_clb_0.mux_fle_2_in_1.INVTX1_14_.scs8hd_inv_1/Y vgnd vpwr scs8hd_diode_2
XFILLER_15_423 vpwr vgnd scs8hd_fill_2
XFILLER_27_294 vgnd vpwr scs8hd_fill_1
Xltile_clb_0.mux_fle_1_in_1.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_1_in_1.INVTX1_7_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_1_in_1.LATCH_3_.latch/Q ltile_clb_0.mux_fle_1_in_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_15_478 vgnd vpwr scs8hd_decap_4
XFILLER_42_242 vgnd vpwr scs8hd_decap_3
Xltile_clb_0.mux_fle_3_in_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_3_in_1.INVTX1_2_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_3_in_1.LATCH_2_.latch/Q ltile_clb_0.mux_fle_3_in_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_63_86 vgnd vpwr scs8hd_decap_12
XFILLER_8_15 vgnd vpwr scs8hd_decap_12
XFILLER_30_459 vpwr vgnd scs8hd_fill_2
XFILLER_10_194 vgnd vpwr scs8hd_fill_1
XFILLER_6_154 vgnd vpwr scs8hd_decap_12
XANTENNA__431__B _429_/X vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
+ _625_/Y vgnd vpwr scs8hd_diode_2
XFILLER_2_382 vpwr vgnd scs8hd_fill_2
XFILLER_2_393 vgnd vpwr scs8hd_decap_4
XFILLER_65_301 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_4_.TGATE_1_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_9_.scs8hd_inv_1/Y
+ _612_/Y ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_4_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_77_194 vpwr vgnd scs8hd_fill_2
XFILLER_80_304 vgnd vpwr scs8hd_decap_8
XFILLER_65_367 vpwr vgnd scs8hd_fill_2
XFILLER_80_337 vgnd vpwr scs8hd_decap_6
XFILLER_18_272 vgnd vpwr scs8hd_decap_3
XFILLER_33_231 vpwr vgnd scs8hd_fill_2
XFILLER_33_297 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_12_.scs8hd_inv_1
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_12_.latch/Q
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_12_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA__622__A _622_/A vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_10_.scs8hd_inv_1_A
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_10_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__341__B _341_/B vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_3_in_1.INVTX1_2_.scs8hd_inv_1 bottom_width_0_height_0__pin_2_
+ ltile_clb_0.mux_fle_3_in_1.INVTX1_2_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XFILLER_56_323 vgnd vpwr scs8hd_decap_3
XFILLER_56_312 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_9_.scs8hd_inv_1
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_9_.latch/Q
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_9_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_ltile_clb_0.mem_fle_2_in_3.LATCH_5_.latch_SLEEPB _390_/Y vgnd vpwr scs8hd_diode_2
XFILLER_56_367 vgnd vpwr scs8hd_fill_1
XPHY_215 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_204 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_259 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_248 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_237 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_226 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_264 vgnd vpwr scs8hd_decap_8
XFILLER_8_408 vgnd vpwr scs8hd_decap_3
XFILLER_20_492 vgnd vpwr scs8hd_decap_4
XANTENNA__532__A _250_/X vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mem_fle_1_in_3.LATCH_7_.latch_D data_in vgnd vpwr scs8hd_diode_2
Xltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_0_.scs8hd_inv_1
+ ltile_clb_0.mux_fle_0_in_0.INVTX1_14_.scs8hd_inv_1/Y _629_/A vgnd vpwr scs8hd_inv_1
XFILLER_3_135 vgnd vpwr scs8hd_decap_12
XANTENNA__251__B _250_/X vgnd vpwr scs8hd_diode_2
XFILLER_79_437 vgnd vpwr scs8hd_decap_4
XFILLER_47_301 vpwr vgnd scs8hd_fill_2
XFILLER_47_345 vpwr vgnd scs8hd_fill_2
XFILLER_47_356 vgnd vpwr scs8hd_fill_1
XFILLER_74_175 vgnd vpwr scs8hd_decap_8
XFILLER_35_507 vgnd vpwr scs8hd_decap_8
XFILLER_47_367 vpwr vgnd scs8hd_fill_2
XFILLER_47_378 vpwr vgnd scs8hd_fill_2
XFILLER_47_389 vpwr vgnd scs8hd_fill_2
XFILLER_62_337 vpwr vgnd scs8hd_fill_2
XFILLER_15_220 vpwr vgnd scs8hd_fill_2
XFILLER_30_212 vpwr vgnd scs8hd_fill_2
XPHY_771 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_760 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__426__B _410_/X vgnd vpwr scs8hd_diode_2
XFILLER_15_297 vpwr vgnd scs8hd_fill_2
XPHY_793 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_782 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_ltile_clb_0.mux_fle_2_in_1.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_2_in_1.INVTX1_12_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_30_267 vgnd vpwr scs8hd_decap_4
XFILLER_30_289 vgnd vpwr scs8hd_fill_1
XANTENNA_ltile_clb_0.mux_fle_0_in_3.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_0_in_3.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_7_485 vgnd vpwr scs8hd_decap_3
XANTENNA__442__A _431_/A vgnd vpwr scs8hd_diode_2
XFILLER_31_3 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mem_fle_2_in_1.LATCH_7_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_2_190 vgnd vpwr scs8hd_decap_12
XFILLER_78_492 vgnd vpwr scs8hd_decap_12
XFILLER_65_153 vpwr vgnd scs8hd_fill_2
XFILLER_53_315 vgnd vpwr scs8hd_decap_3
Xltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.INVTX1_0_.scs8hd_inv_1
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.INVTX1_0_.scs8hd_inv_1/A
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_ltile_clb_0.mux_fle_0_in_0.INVTX1_8_.scs8hd_inv_1_A top_width_0_height_0__pin_8_
+ vgnd vpwr scs8hd_diode_2
XANTENNA__617__A _617_/A vgnd vpwr scs8hd_diode_2
XFILLER_80_178 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_1_.TGATE_1_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_1_.TGATE_1_.scs8hd_ebufn_2/A
+ _608_/Y ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l4_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_21_245 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.mux_fle_3_in_2.INVTX1_6_.scs8hd_inv_1 bottom_width_0_height_0__pin_6_
+ ltile_clb_0.mux_fle_3_in_2.INVTX1_6_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XANTENNA_ltile_clb_0.mem_fle_2_in_2.LATCH_5_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_2_in_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_2_in_2.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__352__A _391_/A vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_2_in_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_2_in_2.LATCH_4_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mem_fle_3_in_2.LATCH_5_.latch_SLEEPB _351_/Y vgnd vpwr scs8hd_diode_2
XFILLER_0_149 vgnd vpwr scs8hd_decap_6
XFILLER_29_301 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB
+ _621_/Y vgnd vpwr scs8hd_diode_2
XFILLER_28_56 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.mux_fle_2_in_2.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_2_in_2.INVTX1_2_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_2_in_2.LATCH_2_.latch/Q ltile_clb_0.mux_fle_2_in_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_7_.latch_SLEEPB
+ _565_/Y vgnd vpwr scs8hd_diode_2
XFILLER_29_378 vgnd vpwr scs8hd_decap_3
Xltile_clb_0.mux_fle_0_in_2.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_0_in_2.INVTX1_7_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_0_in_2.LATCH_3_.latch/Q ltile_clb_0.mux_fle_0_in_2.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_ltile_clb_0.mem_fle_2_in_3.LATCH_3_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_71_123 vgnd vpwr scs8hd_decap_12
XFILLER_44_337 vgnd vpwr scs8hd_fill_1
XANTENNA__527__A address[4] vgnd vpwr scs8hd_diode_2
X_490_ _421_/A _484_/X _490_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_44_44 vgnd vpwr scs8hd_decap_12
XANTENNA__246__B _286_/A vgnd vpwr scs8hd_diode_2
XFILLER_12_267 vgnd vpwr scs8hd_fill_1
XFILLER_60_32 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_14_.latch
+ data_in ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_14_.latch/Q
+ _557_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA__262__A _248_/A vgnd vpwr scs8hd_diode_2
XFILLER_5_27 vgnd vpwr scs8hd_decap_12
XFILLER_4_433 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_1_in_1.INVTX1_5_.scs8hd_inv_1_A right_width_0_height_0__pin_5_
+ vgnd vpwr scs8hd_diode_2
XFILLER_4_455 vgnd vpwr scs8hd_fill_1
XFILLER_4_444 vpwr vgnd scs8hd_fill_2
XFILLER_69_74 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mem_fle_3_in_0.LATCH_5_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_79_245 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mem_fle_0_in_3.LATCH_6_.latch_SLEEPB _486_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_3_in_1.INVTX1_11_.scs8hd_inv_1_A left_width_0_height_0__pin_11_
+ vgnd vpwr scs8hd_diode_2
XFILLER_47_131 vgnd vpwr scs8hd_fill_1
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__ff_0.DFFSRQ_0_.dff_D
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.INVTX1_1_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_47_175 vpwr vgnd scs8hd_fill_2
XANTENNA__437__A _437_/A vgnd vpwr scs8hd_diode_2
XFILLER_62_145 vpwr vgnd scs8hd_fill_2
XFILLER_43_370 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mem_fle_3_in_1.LATCH_3_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_43_381 vpwr vgnd scs8hd_fill_2
XFILLER_79_3 vgnd vpwr scs8hd_decap_12
XPHY_590 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_7_271 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_1_in_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_1_in_0.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mem_fle_3_in_2.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_66_440 vgnd vpwr scs8hd_fill_1
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_9_.latch_D
+ data_in vgnd vpwr scs8hd_diode_2
XFILLER_81_410 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mux_fle_2_in_2.INVTX1_2_.scs8hd_inv_1_A bottom_width_0_height_0__pin_2_
+ vgnd vpwr scs8hd_diode_2
XFILLER_53_123 vgnd vpwr scs8hd_decap_8
XFILLER_26_337 vgnd vpwr scs8hd_decap_3
XFILLER_81_487 vgnd vpwr scs8hd_fill_1
XANTENNA__347__A _347_/A vgnd vpwr scs8hd_diode_2
XFILLER_22_510 vgnd vpwr scs8hd_decap_6
XFILLER_5_219 vpwr vgnd scs8hd_fill_2
XFILLER_30_68 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mux_fle_2_in_2.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_2_in_2.INVTX1_10_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_76_215 vgnd vpwr scs8hd_decap_8
XFILLER_76_204 vgnd vpwr scs8hd_decap_8
X_611_ _611_/A _611_/Y vgnd vpwr scs8hd_inv_8
XFILLER_17_326 vgnd vpwr scs8hd_decap_3
XFILLER_29_175 vpwr vgnd scs8hd_fill_2
XFILLER_72_432 vpwr vgnd scs8hd_fill_2
X_542_ _542_/A _541_/B _542_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_44_145 vgnd vpwr scs8hd_decap_6
XFILLER_55_98 vgnd vpwr scs8hd_decap_12
XANTENNA__257__A _248_/A vgnd vpwr scs8hd_diode_2
XFILLER_32_318 vgnd vpwr scs8hd_fill_1
XANTENNA_ltile_clb_0.mux_fle_0_in_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_0_in_0.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
X_473_ _481_/B _479_/B vgnd vpwr scs8hd_buf_1
XFILLER_25_392 vpwr vgnd scs8hd_fill_2
XFILLER_9_514 vpwr vgnd scs8hd_fill_2
XFILLER_71_86 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mem_fle_1_in_2.LATCH_6_.latch_SLEEPB _453_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_1_in_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_1_in_0.LATCH_6_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_4_285 vgnd vpwr scs8hd_decap_8
Xltile_clb_0.mux_fle_0_in_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_0_in_0.INVTX1_1_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_0_in_0.LATCH_1_.latch/Q ltile_clb_0.mux_fle_0_in_0.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_4_296 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
+ _637_/HI vgnd vpwr scs8hd_diode_2
XFILLER_48_462 vgnd vpwr scs8hd_decap_8
XFILLER_82_218 vgnd vpwr scs8hd_decap_12
XFILLER_35_123 vgnd vpwr scs8hd_decap_12
XFILLER_35_156 vgnd vpwr scs8hd_decap_4
Xltile_clb_0.mux_fle_3_in_2.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_3_in_2.mux_l1_in_3_.TGATE_2_.scs8hd_ebufn_2/Z
+ ltile_clb_0.mem_fle_3_in_2.LATCH_7_.latch/Q ltile_clb_0.mux_fle_3_in_2.INVTX1_14_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
Xltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_1_.TGATE_1_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_1_.TGATE_1_.scs8hd_ebufn_2/A
+ _630_/Y ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA__630__A _630_/A vgnd vpwr scs8hd_diode_2
XFILLER_58_248 vgnd vpwr scs8hd_fill_1
Xltile_clb_0.mux_fle_1_in_3.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_1_in_3.INVTX1_2_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_1_in_3.LATCH_2_.latch/Q ltile_clb_0.mux_fle_1_in_3.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
Xltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_2_.scs8hd_inv_1
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_2_.latch/Q
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_73_207 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.mux_fle_2_in_0.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_2_in_0.INVTX1_13_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_2_in_0.LATCH_1_.latch/Q ltile_clb_0.mux_fle_2_in_0.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_73_218 vpwr vgnd scs8hd_fill_2
XPHY_13 vgnd vpwr scs8hd_decap_3
XPHY_24 vgnd vpwr scs8hd_decap_3
XFILLER_14_329 vgnd vpwr scs8hd_decap_6
XPHY_35 vgnd vpwr scs8hd_decap_3
XPHY_46 vgnd vpwr scs8hd_decap_3
XFILLER_26_189 vpwr vgnd scs8hd_fill_2
XPHY_57 vgnd vpwr scs8hd_decap_3
XPHY_68 vgnd vpwr scs8hd_decap_3
XPHY_79 vgnd vpwr scs8hd_decap_3
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_5_.latch_D
+ data_in vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_0_in_2.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_0_in_2.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__524__B _516_/X vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_3_in_3.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_3_in_3.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_1_in_0.INVTX1_10_.scs8hd_inv_1_A bottom_width_0_height_0__pin_10_
+ vgnd vpwr scs8hd_diode_2
XANTENNA__540__A _540_/A vgnd vpwr scs8hd_diode_2
XFILLER_9_3 vgnd vpwr scs8hd_decap_12
XFILLER_77_513 vgnd vpwr scs8hd_decap_3
XFILLER_1_255 vpwr vgnd scs8hd_fill_2
XFILLER_49_226 vgnd vpwr scs8hd_decap_4
XFILLER_64_229 vgnd vpwr scs8hd_decap_6
XANTENNA_ltile_clb_0.mem_fle_2_in_1.LATCH_6_.latch_SLEEPB _414_/Y vgnd vpwr scs8hd_diode_2
XFILLER_17_123 vgnd vpwr scs8hd_decap_12
XFILLER_45_443 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.mux_fle_3_in_3.mux_l1_in_3_.TGATE_2_.scs8hd_ebufn_2 _655_/HI ltile_clb_0.mem_fle_3_in_3.LATCH_2_.latch/Q
+ ltile_clb_0.mux_fle_3_in_3.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
X_525_ _343_/A _516_/X _525_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_82_63 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mux_fle_3_in_2.mux_l1_in_2_.TGATE_3_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_3_in_2.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_45_498 vpwr vgnd scs8hd_fill_2
XFILLER_60_468 vpwr vgnd scs8hd_fill_2
XFILLER_9_300 vpwr vgnd scs8hd_fill_2
X_456_ _434_/A _451_/X _456_/Y vgnd vpwr scs8hd_nor2_4
X_387_ _387_/A _388_/B vgnd vpwr scs8hd_buf_1
XANTENNA__434__B _429_/X vgnd vpwr scs8hd_diode_2
XFILLER_40_192 vgnd vpwr scs8hd_decap_4
XANTENNA__450__A _449_/X vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_12_.latch_SLEEPB
+ _585_/Y vgnd vpwr scs8hd_diode_2
XFILLER_48_270 vgnd vpwr scs8hd_decap_4
XFILLER_63_262 vgnd vpwr scs8hd_fill_1
XFILLER_63_240 vpwr vgnd scs8hd_fill_2
XFILLER_51_424 vgnd vpwr scs8hd_fill_1
XFILLER_23_159 vgnd vpwr scs8hd_decap_12
XANTENNA__625__A _625_/A vgnd vpwr scs8hd_diode_2
XANTENNA__344__B _341_/B vgnd vpwr scs8hd_diode_2
XFILLER_11_15 vgnd vpwr scs8hd_decap_12
XFILLER_11_59 vpwr vgnd scs8hd_fill_2
XANTENNA__360__A _368_/B vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_0_in_0.INVTX1_6_.scs8hd_inv_1 bottom_width_0_height_0__pin_6_
+ ltile_clb_0.mux_fle_0_in_0.INVTX1_6_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XFILLER_46_229 vgnd vpwr scs8hd_fill_1
XFILLER_39_281 vgnd vpwr scs8hd_decap_4
XANTENNA__519__B _517_/X vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_1_in_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_1_in_0.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2/Z
+ ltile_clb_0.mem_fle_1_in_0.LATCH_6_.latch/Q ltile_clb_0.mux_fle_1_in_0.INVTX1_14_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_27_476 vgnd vpwr scs8hd_fill_1
XFILLER_36_56 vgnd vpwr scs8hd_decap_12
XFILLER_42_413 vgnd vpwr scs8hd_fill_1
X_310_ _575_/A _309_/X _310_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_42_435 vgnd vpwr scs8hd_decap_3
XFILLER_42_457 vgnd vpwr scs8hd_fill_1
XFILLER_42_468 vgnd vpwr scs8hd_decap_3
XFILLER_52_44 vgnd vpwr scs8hd_decap_12
XANTENNA__535__A _535_/A vgnd vpwr scs8hd_diode_2
X_241_ _286_/A _282_/B _286_/B _313_/A vgnd vpwr scs8hd_or3_4
XFILLER_10_321 vpwr vgnd scs8hd_fill_2
XANTENNA__254__B _603_/A vgnd vpwr scs8hd_diode_2
XFILLER_10_365 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mem_fle_3_in_0.LATCH_6_.latch_SLEEPB _373_/Y vgnd vpwr scs8hd_diode_2
XFILLER_10_398 vgnd vpwr scs8hd_decap_6
Xltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_7_.scs8hd_inv_1
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_7_.latch/Q
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA__270__A _258_/X vgnd vpwr scs8hd_diode_2
XFILLER_77_74 vgnd vpwr scs8hd_decap_12
XFILLER_77_376 vpwr vgnd scs8hd_fill_2
XFILLER_18_410 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_1_in_2.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_1_in_2.INVTX1_12_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_45_240 vpwr vgnd scs8hd_fill_2
XFILLER_45_273 vpwr vgnd scs8hd_fill_2
XFILLER_45_284 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.mux_fle_2_in_3.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_2_in_3.mux_l1_in_3_.TGATE_2_.scs8hd_ebufn_2/Z
+ ltile_clb_0.mem_fle_2_in_3.LATCH_7_.latch/Q ltile_clb_0.mux_fle_2_in_3.INVTX1_14_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_ltile_clb_0.mux_fle_3_in_2.INVTX1_8_.scs8hd_inv_1_A top_width_0_height_0__pin_8_
+ vgnd vpwr scs8hd_diode_2
X_508_ _325_/A _511_/B _508_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_33_468 vpwr vgnd scs8hd_fill_2
XFILLER_60_287 vgnd vpwr scs8hd_decap_8
XFILLER_60_276 vpwr vgnd scs8hd_fill_2
XANTENNA__445__A _434_/A vgnd vpwr scs8hd_diode_2
XFILLER_20_129 vgnd vpwr scs8hd_decap_12
X_439_ _438_/X _447_/B vgnd vpwr scs8hd_buf_1
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_0_.latch_SLEEPB
+ _598_/Y vgnd vpwr scs8hd_diode_2
XFILLER_61_3 vgnd vpwr scs8hd_decap_12
XFILLER_9_196 vgnd vpwr scs8hd_decap_3
XANTENNA_ltile_clb_0.mem_fle_0_in_1.LATCH_7_.latch_SLEEPB _507_/Y vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_1_in_1.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_1_in_1.INVTX1_13_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_1_in_1.LATCH_1_.latch/Q ltile_clb_0.mux_fle_1_in_1.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_68_321 vpwr vgnd scs8hd_fill_2
XFILLER_68_310 vgnd vpwr scs8hd_decap_8
Xltile_clb_0.mux_fle_3_in_1.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_3_in_1.INVTX1_8_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_3_in_1.LATCH_0_.latch/Q ltile_clb_0.mux_fle_3_in_1.mux_l1_in_2_.TGATE_3_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_68_365 vgnd vpwr scs8hd_decap_8
XFILLER_56_505 vgnd vpwr scs8hd_decap_8
XANTENNA_ltile_clb_0.mux_fle_1_in_3.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_1_in_3.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_1_in_1.INVTX1_1_.scs8hd_inv_1 right_width_0_height_0__pin_1_
+ ltile_clb_0.mux_fle_1_in_1.INVTX1_1_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XFILLER_51_221 vpwr vgnd scs8hd_fill_2
XPHY_408 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_51_232 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.buf4_1_.scs8hd_buf_1_A
+ ltile_clb_0.mux_fle_1_in_1.INVTX1_14_.scs8hd_inv_1/Y vgnd vpwr scs8hd_diode_2
XFILLER_24_457 vgnd vpwr scs8hd_fill_1
XFILLER_24_468 vgnd vpwr scs8hd_decap_12
XPHY_419 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__355__A _394_/A vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_0_.TGATE_0_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_32_490 vpwr vgnd scs8hd_fill_2
XFILLER_3_339 vpwr vgnd scs8hd_fill_2
XFILLER_78_129 vgnd vpwr scs8hd_decap_12
XFILLER_74_335 vgnd vpwr scs8hd_fill_1
XANTENNA__249__B _286_/A vgnd vpwr scs8hd_diode_2
XFILLER_27_240 vpwr vgnd scs8hd_fill_2
XFILLER_27_262 vpwr vgnd scs8hd_fill_2
XFILLER_27_273 vpwr vgnd scs8hd_fill_2
XFILLER_42_221 vgnd vpwr scs8hd_fill_1
Xltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_12_.latch
+ data_in ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_12_.latch/Q
+ _257_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_63_98 vgnd vpwr scs8hd_decap_12
XANTENNA__265__A _264_/X vgnd vpwr scs8hd_diode_2
XFILLER_42_287 vgnd vpwr scs8hd_decap_12
XFILLER_8_27 vgnd vpwr scs8hd_decap_4
Xltile_clb_0.mux_fle_0_in_0.INVTX1_13_.scs8hd_inv_1 right_width_0_height_0__pin_13_
+ ltile_clb_0.mux_fle_0_in_0.INVTX1_13_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XFILLER_12_80 vgnd vpwr scs8hd_decap_12
XFILLER_6_166 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.mem_fle_0_in_0.LATCH_5_.latch data_in ltile_clb_0.mem_fle_0_in_0.LATCH_5_.latch/Q
+ _520_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
Xltile_clb_0.mux_fle_3_in_0.INVTX1_12_.scs8hd_inv_1 top_width_0_height_0__pin_12_
+ ltile_clb_0.mux_fle_3_in_0.INVTX1_12_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_6_.TGATE_1_.scs8hd_ebufn_2_TEB
+ _620_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_2_.scs8hd_inv_1_A
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_77_184 vgnd vpwr scs8hd_decap_6
Xltile_clb_0.mem_fle_1_in_0.LATCH_4_.latch data_in ltile_clb_0.mem_fle_1_in_0.LATCH_4_.latch/Q
+ _477_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_18_295 vgnd vpwr scs8hd_fill_1
XFILLER_33_243 vgnd vpwr scs8hd_fill_1
XFILLER_21_405 vpwr vgnd scs8hd_fill_2
XFILLER_21_416 vpwr vgnd scs8hd_fill_2
XFILLER_21_449 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_0_in_1.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_0_in_1.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mem_fle_1_in_0.LATCH_7_.latch_SLEEPB _474_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
+ _613_/Y vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mem_fle_2_in_0.LATCH_3_.latch data_in ltile_clb_0.mem_fle_2_in_0.LATCH_3_.latch/Q
+ _434_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_ltile_clb_0.mux_fle_0_in_0.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_0_in_0.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_0_in_1.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_0_in_1.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2/Z
+ ltile_clb_0.mem_fle_0_in_1.LATCH_6_.latch/Q ltile_clb_0.mux_fle_0_in_1.INVTX1_14_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
Xltile_clb_0.mux_fle_1_in_2.INVTX1_5_.scs8hd_inv_1 right_width_0_height_0__pin_5_
+ ltile_clb_0.mux_fle_1_in_2.INVTX1_5_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XFILLER_68_162 vpwr vgnd scs8hd_fill_2
XFILLER_56_346 vgnd vpwr scs8hd_decap_4
Xltile_clb_0.mux_fle_3_in_1.INVTX1_14_.scs8hd_inv_1 ltile_clb_0.mux_fle_3_in_1.INVTX1_14_.scs8hd_inv_1/A
+ ltile_clb_0.mux_fle_3_in_1.INVTX1_14_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XANTENNA_ltile_clb_0.mux_fle_3_in_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_3_in_1.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mem_fle_3_in_0.LATCH_2_.latch data_in ltile_clb_0.mem_fle_3_in_0.LATCH_2_.latch/Q
+ _377_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.buf4_3_.scs8hd_buf_1_A
+ ltile_clb_0.mux_fle_3_in_3.INVTX1_14_.scs8hd_inv_1/Y vgnd vpwr scs8hd_diode_2
XPHY_216 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_205 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_243 vpwr vgnd scs8hd_fill_2
XPHY_249 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_238 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_227 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_ltile_clb_0.mux_fle_1_in_3.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_1_in_3.INVTX1_10_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_4_.scs8hd_inv_1/Y
+ _621_/Y ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_1_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_20_471 vgnd vpwr scs8hd_decap_8
XANTENNA__532__B _529_/X vgnd vpwr scs8hd_diode_2
XFILLER_3_147 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mux_fle_0_in_2.INVTX1_6_.scs8hd_inv_1_A bottom_width_0_height_0__pin_6_
+ vgnd vpwr scs8hd_diode_2
XFILLER_58_32 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mux_fle_1_in_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_1_in_2.LATCH_5_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_47_313 vpwr vgnd scs8hd_fill_2
XFILLER_59_184 vgnd vpwr scs8hd_fill_1
XFILLER_74_154 vgnd vpwr scs8hd_fill_1
XFILLER_62_305 vgnd vpwr scs8hd_decap_4
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_12_.scs8hd_inv_1_A
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_12_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_74_187 vgnd vpwr scs8hd_decap_6
XFILLER_62_349 vgnd vpwr scs8hd_decap_4
XPHY_772 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_761 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_750 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_794 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_783 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_11_460 vpwr vgnd scs8hd_fill_2
XFILLER_11_482 vpwr vgnd scs8hd_fill_2
XFILLER_7_442 vgnd vpwr scs8hd_decap_3
XFILLER_7_453 vpwr vgnd scs8hd_fill_2
XANTENNA__442__B _446_/B vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_2_in_2.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_2_in_2.INVTX1_8_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_2_in_2.LATCH_0_.latch/Q ltile_clb_0.mux_fle_2_in_2.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
Xltile_clb_0.mux_fle_0_in_2.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_0_in_2.INVTX1_13_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_0_in_2.LATCH_1_.latch/Q ltile_clb_0.mux_fle_0_in_2.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
Xltile_clb_0.mem_fle_1_in_2.LATCH_7_.latch data_in ltile_clb_0.mem_fle_1_in_2.LATCH_7_.latch/Q
+ _452_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
Xltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_6_.TGATE_1_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_13_.scs8hd_inv_1/Y
+ _620_/Y ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_3_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_24_3 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.mux_fle_2_in_3.INVTX1_0_.scs8hd_inv_1 top_width_0_height_0__pin_0_ ltile_clb_0.mux_fle_2_in_3.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_65_110 vgnd vpwr scs8hd_decap_12
XFILLER_38_346 vpwr vgnd scs8hd_fill_2
XFILLER_38_379 vgnd vpwr scs8hd_fill_1
Xltile_clb_0.mem_fle_2_in_2.LATCH_6_.latch data_in ltile_clb_0.mem_fle_2_in_2.LATCH_6_.latch/Q
+ _400_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_65_187 vpwr vgnd scs8hd_fill_2
XFILLER_65_176 vgnd vpwr scs8hd_decap_4
XANTENNA_ltile_clb_0.mux_fle_1_in_3.INVTX1_3_.scs8hd_inv_1_A left_width_0_height_0__pin_3_
+ vgnd vpwr scs8hd_diode_2
XFILLER_0_94 vgnd vpwr scs8hd_decap_12
XFILLER_61_360 vpwr vgnd scs8hd_fill_2
XANTENNA__633__A _633_/A vgnd vpwr scs8hd_diode_2
XANTENNA__352__B _353_/B vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mem_fle_3_in_2.LATCH_5_.latch data_in ltile_clb_0.mem_fle_3_in_2.LATCH_5_.latch/Q
+ _351_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
Xltile_clb_0.mux_fle_1_in_3.INVTX1_9_.scs8hd_inv_1 right_width_0_height_0__pin_9_
+ ltile_clb_0.mux_fle_1_in_3.INVTX1_9_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XFILLER_0_106 vgnd vpwr scs8hd_decap_12
XFILLER_76_419 vgnd vpwr scs8hd_decap_4
XFILLER_29_313 vgnd vpwr scs8hd_decap_4
XFILLER_29_346 vpwr vgnd scs8hd_fill_2
XFILLER_28_68 vgnd vpwr scs8hd_decap_12
XFILLER_29_357 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_5_.TGATE_0_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_10_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_71_135 vgnd vpwr scs8hd_decap_12
XFILLER_71_179 vgnd vpwr scs8hd_decap_4
XANTENNA__527__B _526_/X vgnd vpwr scs8hd_diode_2
XFILLER_44_56 vgnd vpwr scs8hd_decap_12
XFILLER_12_224 vgnd vpwr scs8hd_decap_12
XFILLER_12_213 vgnd vpwr scs8hd_fill_1
XANTENNA__246__C _282_/C vgnd vpwr scs8hd_diode_2
XFILLER_60_44 vgnd vpwr scs8hd_decap_12
XANTENNA__543__A _569_/A vgnd vpwr scs8hd_diode_2
XANTENNA__262__B _261_/X vgnd vpwr scs8hd_diode_2
XFILLER_20_290 vgnd vpwr scs8hd_decap_6
XFILLER_5_39 vgnd vpwr scs8hd_decap_12
XFILLER_79_257 vgnd vpwr scs8hd_decap_3
XFILLER_69_86 vgnd vpwr scs8hd_decap_12
XFILLER_79_279 vgnd vpwr scs8hd_decap_3
XFILLER_67_419 vgnd vpwr scs8hd_decap_6
XFILLER_47_110 vgnd vpwr scs8hd_decap_12
XFILLER_47_187 vpwr vgnd scs8hd_fill_2
XFILLER_62_157 vgnd vpwr scs8hd_decap_4
XFILLER_62_135 vgnd vpwr scs8hd_fill_1
XANTENNA__437__B _428_/X vgnd vpwr scs8hd_diode_2
XFILLER_50_308 vpwr vgnd scs8hd_fill_2
XPHY_580 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_591 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_0_.TGATE_0_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XANTENNA__453__A _431_/A vgnd vpwr scs8hd_diode_2
XFILLER_11_290 vgnd vpwr scs8hd_decap_4
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_4_.scs8hd_inv_1_A
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_4_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mem_fle_1_in_3.LATCH_0_.latch_SLEEPB _448_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_0_in_0.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_0_in_0.LATCH_7_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_78_290 vgnd vpwr scs8hd_decap_4
XFILLER_38_154 vgnd vpwr scs8hd_decap_4
XFILLER_81_422 vgnd vpwr scs8hd_decap_4
XFILLER_66_474 vgnd vpwr scs8hd_decap_12
XANTENNA__628__A _628_/A vgnd vpwr scs8hd_diode_2
XFILLER_81_433 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.mux_fle_2_in_2.INVTX1_10_.scs8hd_inv_1 bottom_width_0_height_0__pin_10_
+ ltile_clb_0.mux_fle_2_in_2.INVTX1_10_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XFILLER_26_349 vgnd vpwr scs8hd_decap_8
XFILLER_38_198 vgnd vpwr scs8hd_decap_3
XFILLER_53_179 vpwr vgnd scs8hd_fill_2
XFILLER_14_15 vgnd vpwr scs8hd_decap_12
XFILLER_34_371 vgnd vpwr scs8hd_decap_6
XANTENNA__363__A _374_/A vgnd vpwr scs8hd_diode_2
XFILLER_1_404 vpwr vgnd scs8hd_fill_2
XFILLER_29_110 vgnd vpwr scs8hd_decap_12
XFILLER_57_441 vgnd vpwr scs8hd_fill_1
X_610_ _610_/A _610_/Y vgnd vpwr scs8hd_inv_8
XFILLER_57_485 vgnd vpwr scs8hd_decap_3
XFILLER_57_474 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_11_.latch_SLEEPB
+ _560_/Y vgnd vpwr scs8hd_diode_2
XANTENNA__538__A _564_/A vgnd vpwr scs8hd_diode_2
X_541_ _541_/A _541_/B _541_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_17_338 vgnd vpwr scs8hd_decap_3
Xltile_clb_0.mux_fle_3_in_0.INVTX1_6_.scs8hd_inv_1 bottom_width_0_height_0__pin_6_
+ ltile_clb_0.mux_fle_3_in_0.INVTX1_6_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XFILLER_72_466 vpwr vgnd scs8hd_fill_2
XANTENNA__257__B _559_/A vgnd vpwr scs8hd_diode_2
XFILLER_44_179 vgnd vpwr scs8hd_decap_4
X_472_ _471_/X _481_/B vgnd vpwr scs8hd_buf_1
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_7_.TGATE_1_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_15_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_25_371 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.mux_fle_2_in_3.INVTX1_12_.scs8hd_inv_1 top_width_0_height_0__pin_12_
+ ltile_clb_0.mux_fle_2_in_3.INVTX1_12_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XFILLER_71_98 vgnd vpwr scs8hd_decap_12
XANTENNA__273__A _267_/X vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_1_in_3.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_1_in_3.INVTX1_8_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_1_in_3.LATCH_0_.latch/Q ltile_clb_0.mux_fle_1_in_3.mux_l1_in_2_.TGATE_3_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_ltile_clb_0.mux_fle_0_in_3.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_0_in_3.INVTX1_12_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_4_253 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_2_in_3.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_2_in_3.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_20_80 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mux_fle_3_in_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_3_in_0.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_75_282 vpwr vgnd scs8hd_fill_2
XFILLER_75_271 vgnd vpwr scs8hd_decap_4
XANTENNA__448__A _437_/A vgnd vpwr scs8hd_diode_2
XFILLER_75_293 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_3_in_1.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_3_in_1.INVTX1_12_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_35_135 vgnd vpwr scs8hd_decap_12
XFILLER_35_168 vpwr vgnd scs8hd_fill_2
XFILLER_35_179 vgnd vpwr scs8hd_decap_4
XFILLER_50_105 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mem_fle_2_in_2.LATCH_0_.latch_SLEEPB _406_/Y vgnd vpwr scs8hd_diode_2
XFILLER_6_93 vgnd vpwr scs8hd_decap_12
XFILLER_39_441 vpwr vgnd scs8hd_fill_2
XFILLER_66_271 vgnd vpwr scs8hd_decap_4
XANTENNA__358__A address[8] vgnd vpwr scs8hd_diode_2
XFILLER_39_485 vgnd vpwr scs8hd_fill_1
XFILLER_39_496 vgnd vpwr scs8hd_decap_12
XFILLER_54_455 vgnd vpwr scs8hd_decap_3
XANTENNA_ltile_clb_0.mux_fle_3_in_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_3_in_2.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_1_in_0.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_1_in_0.INVTX1_7_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_1_in_0.LATCH_3_.latch/Q ltile_clb_0.mux_fle_1_in_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XPHY_25 vgnd vpwr scs8hd_decap_3
XPHY_14 vgnd vpwr scs8hd_decap_3
XFILLER_14_308 vgnd vpwr scs8hd_decap_6
XPHY_36 vgnd vpwr scs8hd_decap_3
XPHY_47 vgnd vpwr scs8hd_decap_3
Xltile_clb_0.mux_fle_3_in_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_3_in_0.INVTX1_2_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_3_in_0.LATCH_2_.latch/Q ltile_clb_0.mux_fle_3_in_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XPHY_58 vgnd vpwr scs8hd_decap_3
XPHY_69 vgnd vpwr scs8hd_decap_3
XFILLER_22_352 vpwr vgnd scs8hd_fill_2
XFILLER_10_514 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
+ _638_/HI vgnd vpwr scs8hd_diode_2
XANTENNA__540__B _541_/B vgnd vpwr scs8hd_diode_2
XFILLER_1_245 vgnd vpwr scs8hd_decap_3
XFILLER_49_205 vpwr vgnd scs8hd_fill_2
XFILLER_1_278 vpwr vgnd scs8hd_fill_2
XFILLER_66_32 vgnd vpwr scs8hd_decap_12
XFILLER_72_230 vpwr vgnd scs8hd_fill_2
XFILLER_17_135 vgnd vpwr scs8hd_decap_12
XANTENNA__268__A _286_/B vgnd vpwr scs8hd_diode_2
XFILLER_32_105 vgnd vpwr scs8hd_decap_12
XFILLER_45_466 vpwr vgnd scs8hd_fill_2
X_524_ _423_/A _516_/X _524_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_82_75 vgnd vpwr scs8hd_decap_12
X_455_ _433_/A _451_/X _455_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_13_330 vgnd vpwr scs8hd_decap_4
XFILLER_13_341 vpwr vgnd scs8hd_fill_2
XFILLER_13_352 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_2_in_3.INVTX1_9_.scs8hd_inv_1_A right_width_0_height_0__pin_9_
+ vgnd vpwr scs8hd_diode_2
X_386_ _385_/X _387_/A vgnd vpwr scs8hd_buf_1
XANTENNA_ltile_clb_0.mux_fle_2_in_2.INVTX1_13_.scs8hd_inv_1_A right_width_0_height_0__pin_13_
+ vgnd vpwr scs8hd_diode_2
XFILLER_40_171 vgnd vpwr scs8hd_decap_12
XFILLER_9_367 vpwr vgnd scs8hd_fill_2
XFILLER_9_356 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_3_in_0.INVTX1_5_.scs8hd_inv_1_A right_width_0_height_0__pin_5_
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mem_fle_3_in_1.LATCH_0_.latch_SLEEPB _368_/Y vgnd vpwr scs8hd_diode_2
XFILLER_51_403 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_5_.TGATE_0_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_10_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_6_.scs8hd_inv_1_A
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_6_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_36_488 vgnd vpwr scs8hd_decap_8
XFILLER_51_447 vgnd vpwr scs8hd_decap_3
XFILLER_36_499 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mux_fle_3_in_3.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_3_in_3.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_31_193 vgnd vpwr scs8hd_decap_4
XANTENNA_ltile_clb_0.mux_fle_2_in_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_2_in_0.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_11_27 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.mem_fle_0_in_1.LATCH_1_.latch data_in ltile_clb_0.mem_fle_0_in_1.LATCH_1_.latch/Q
+ _513_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
Xltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.buf4_3_.scs8hd_buf_1
+ ltile_clb_0.mux_fle_3_in_3.INVTX1_14_.scs8hd_inv_1/Y _610_/A vgnd vpwr scs8hd_buf_1
XFILLER_27_400 vgnd vpwr scs8hd_decap_4
XANTENNA_ltile_clb_0.mem_fle_0_in_2.LATCH_1_.latch_SLEEPB _502_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_3_in_2.mux_l1_in_3_.TGATE_2_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_3_in_2.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_54_252 vgnd vpwr scs8hd_fill_1
XFILLER_36_68 vgnd vpwr scs8hd_decap_12
XFILLER_14_105 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_4_.TGATE_1_.scs8hd_ebufn_2_TEB
+ _612_/Y vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mem_fle_1_in_1.LATCH_0_.latch data_in ltile_clb_0.mem_fle_1_in_1.LATCH_0_.latch/Q
+ _470_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_52_56 vgnd vpwr scs8hd_decap_12
XANTENNA__535__B _529_/X vgnd vpwr scs8hd_diode_2
X_240_ address[0] _286_/B vgnd vpwr scs8hd_inv_8
XANTENNA_ltile_clb_0.mux_fle_3_in_2.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_3_in_2.INVTX1_10_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_6_326 vpwr vgnd scs8hd_fill_2
XFILLER_6_359 vgnd vpwr scs8hd_decap_3
XANTENNA__551__A _603_/A vgnd vpwr scs8hd_diode_2
XANTENNA__270__B _270_/B vgnd vpwr scs8hd_diode_2
XFILLER_77_355 vpwr vgnd scs8hd_fill_2
XFILLER_77_344 vpwr vgnd scs8hd_fill_2
XFILLER_77_333 vgnd vpwr scs8hd_decap_4
XFILLER_77_86 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mux_fle_1_in_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_1_in_0.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_18_422 vgnd vpwr scs8hd_decap_3
XFILLER_18_466 vpwr vgnd scs8hd_fill_2
XFILLER_45_252 vpwr vgnd scs8hd_fill_2
XFILLER_60_200 vgnd vpwr scs8hd_decap_12
X_507_ _314_/A _511_/B _507_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_33_447 vgnd vpwr scs8hd_decap_6
XANTENNA__445__B _446_/B vgnd vpwr scs8hd_diode_2
X_438_ _380_/X _226_/X _384_/X _358_/D _438_/X vgnd vpwr scs8hd_or4_4
X_369_ address[8] _369_/B _369_/C _346_/D _370_/A vgnd vpwr scs8hd_or4_4
XFILLER_13_193 vgnd vpwr scs8hd_decap_4
XFILLER_41_480 vpwr vgnd scs8hd_fill_2
XANTENNA__461__A _460_/X vgnd vpwr scs8hd_diode_2
XFILLER_54_3 vgnd vpwr scs8hd_decap_12
XFILLER_5_381 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_14_.latch_D
+ data_in vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_0_in_1.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_0_in_1.INVTX1_7_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_0_in_1.LATCH_3_.latch/Q ltile_clb_0.mux_fle_0_in_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
Xltile_clb_0.mux_fle_2_in_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_2_in_1.INVTX1_2_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_2_in_1.LATCH_2_.latch/Q ltile_clb_0.mux_fle_2_in_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XPHY_409 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xltile_clb_0.mem_fle_0_in_3.LATCH_4_.latch data_in ltile_clb_0.mem_fle_0_in_3.LATCH_4_.latch/Q
+ _488_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA__355__B _355_/B vgnd vpwr scs8hd_diode_2
XFILLER_51_288 vgnd vpwr scs8hd_decap_4
XFILLER_51_299 vgnd vpwr scs8hd_decap_4
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_7_.TGATE_1_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_15_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_22_15 vgnd vpwr scs8hd_decap_12
XANTENNA__371__A _379_/B vgnd vpwr scs8hd_diode_2
Xltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l4_in_0_.TGATE_1_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l4_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ _634_/Y ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_16_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_ltile_clb_0.mem_fle_1_in_1.LATCH_1_.latch_SLEEPB _469_/Y vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mem_fle_1_in_3.LATCH_3_.latch data_in ltile_clb_0.mem_fle_1_in_3.LATCH_3_.latch/Q
+ _445_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_59_377 vgnd vpwr scs8hd_decap_3
XANTENNA_ltile_clb_0.mux_fle_0_in_1.INVTX1_12_.scs8hd_inv_1_A top_width_0_height_0__pin_12_
+ vgnd vpwr scs8hd_diode_2
XANTENNA__249__C _286_/B vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_0_in_0.INVTX1_3_.scs8hd_inv_1_A left_width_0_height_0__pin_3_
+ vgnd vpwr scs8hd_diode_2
XFILLER_15_414 vpwr vgnd scs8hd_fill_2
XFILLER_42_211 vgnd vpwr scs8hd_decap_3
Xltile_clb_0.mem_fle_2_in_3.LATCH_2_.latch data_in ltile_clb_0.mem_fle_2_in_3.LATCH_2_.latch/Q
+ _393_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_ltile_clb_0.mux_fle_2_in_1.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_2_in_1.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_15_458 vgnd vpwr scs8hd_fill_1
XANTENNA__546__A _546_/A vgnd vpwr scs8hd_diode_2
XFILLER_42_255 vgnd vpwr scs8hd_fill_1
XFILLER_23_480 vgnd vpwr scs8hd_decap_4
XFILLER_42_299 vgnd vpwr scs8hd_fill_1
XFILLER_10_141 vgnd vpwr scs8hd_decap_12
XANTENNA__281__A _267_/X vgnd vpwr scs8hd_diode_2
XFILLER_6_178 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.mem_fle_3_in_3.LATCH_1_.latch data_in ltile_clb_0.mem_fle_3_in_3.LATCH_1_.latch/Q
+ _341_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_2_340 vgnd vpwr scs8hd_decap_3
XFILLER_65_336 vgnd vpwr scs8hd_fill_1
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_3_.latch_SLEEPB
+ _543_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_3_.TGATE_1_.scs8hd_ebufn_2_TEB
+ _630_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_0_in_2.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_0_in_2.LATCH_6_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_73_380 vpwr vgnd scs8hd_fill_2
XFILLER_18_263 vpwr vgnd scs8hd_fill_2
XANTENNA__456__A _434_/A vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_1_in_1.INVTX1_0_.scs8hd_inv_1_A top_width_0_height_0__pin_0_
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_8_.scs8hd_inv_1_A
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_8_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_68_141 vgnd vpwr scs8hd_decap_12
XFILLER_71_306 vpwr vgnd scs8hd_fill_2
XFILLER_17_15 vgnd vpwr scs8hd_decap_12
XFILLER_71_339 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mem_fle_2_in_0.LATCH_1_.latch_SLEEPB _436_/Y vgnd vpwr scs8hd_diode_2
XFILLER_17_59 vpwr vgnd scs8hd_fill_2
XANTENNA__366__A _338_/A vgnd vpwr scs8hd_diode_2
XPHY_206 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_233 vgnd vpwr scs8hd_fill_1
XFILLER_12_428 vgnd vpwr scs8hd_decap_8
XPHY_239 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_228 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_217 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_20_450 vgnd vpwr scs8hd_decap_8
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_7_.TGATE_0_.scs8hd_ebufn_2_TEB
+ _621_/Y vgnd vpwr scs8hd_diode_2
XFILLER_3_159 vgnd vpwr scs8hd_decap_12
XFILLER_58_44 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_1_.scs8hd_inv_1_A
+ ltile_clb_0.mux_fle_1_in_1.INVTX1_14_.scs8hd_inv_1/Y vgnd vpwr scs8hd_diode_2
Xltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ _614_/Y ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_59_141 vgnd vpwr scs8hd_decap_6
XFILLER_74_32 vgnd vpwr scs8hd_decap_12
XFILLER_55_380 vpwr vgnd scs8hd_fill_2
XANTENNA__276__A _276_/A vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_3_in_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_3_in_2.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_15_266 vpwr vgnd scs8hd_fill_2
XFILLER_15_277 vgnd vpwr scs8hd_decap_3
XPHY_762 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_751 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_740 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_30_225 vgnd vpwr scs8hd_decap_8
XPHY_795 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_784 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_773 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xltile_clb_0.mux_fle_3_in_1.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_3_in_1.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2/Z
+ ltile_clb_0.mem_fle_3_in_1.LATCH_7_.latch/Q ltile_clb_0.mux_fle_3_in_1.INVTX1_14_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_30_247 vgnd vpwr scs8hd_decap_8
XFILLER_7_498 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_2_in_2.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_2_in_2.INVTX1_12_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_1_in_2.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_1_in_2.INVTX1_2_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_1_in_2.LATCH_2_.latch/Q ltile_clb_0.mux_fle_1_in_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_78_450 vgnd vpwr scs8hd_decap_8
Xltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.INVTX1_1_.scs8hd_inv_1
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.INVTX1_1_.scs8hd_inv_1/A
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_ltile_clb_0.mux_fle_3_in_1.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_3_in_1.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_17_3 vgnd vpwr scs8hd_decap_12
XFILLER_38_369 vgnd vpwr scs8hd_decap_3
XFILLER_53_328 vgnd vpwr scs8hd_fill_1
XANTENNA_ltile_clb_0.mux_fle_0_in_0.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_0_in_0.INVTX1_8_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_10_.latch_SLEEPB
+ _535_/Y vgnd vpwr scs8hd_diode_2
XFILLER_21_214 vgnd vpwr scs8hd_fill_1
XFILLER_21_236 vgnd vpwr scs8hd_decap_4
XFILLER_0_118 vgnd vpwr scs8hd_decap_6
XANTENNA_ltile_clb_0.mux_fle_2_in_3.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_2_in_3.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_69_461 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.mux_fle_3_in_2.mux_l1_in_3_.TGATE_2_.scs8hd_ebufn_2 _654_/HI ltile_clb_0.mem_fle_3_in_2.LATCH_2_.latch/Q
+ ltile_clb_0.mux_fle_3_in_2.mux_l1_in_3_.TGATE_2_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XFILLER_44_306 vpwr vgnd scs8hd_fill_2
XFILLER_44_317 vpwr vgnd scs8hd_fill_2
XFILLER_44_328 vgnd vpwr scs8hd_decap_8
XFILLER_71_158 vpwr vgnd scs8hd_fill_2
XFILLER_71_147 vgnd vpwr scs8hd_decap_8
XFILLER_37_380 vgnd vpwr scs8hd_decap_4
Xltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_4_.TGATE_0_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_8_.scs8hd_inv_1/Y
+ _629_/Y ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_2_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_44_68 vgnd vpwr scs8hd_decap_12
XFILLER_52_383 vgnd vpwr scs8hd_decap_4
XFILLER_52_372 vpwr vgnd scs8hd_fill_2
XFILLER_12_236 vgnd vpwr scs8hd_decap_3
XANTENNA__246__D _282_/B vgnd vpwr scs8hd_diode_2
XANTENNA__543__B _528_/X vgnd vpwr scs8hd_diode_2
XFILLER_60_56 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
+ _608_/Y vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_1_in_0.INVTX1_5_.scs8hd_inv_1 right_width_0_height_0__pin_5_
+ ltile_clb_0.mux_fle_1_in_0.INVTX1_5_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
Xltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.buf4_0_.scs8hd_buf_1
+ ltile_clb_0.mux_fle_2_in_0.INVTX1_14_.scs8hd_inv_1/Y _612_/A vgnd vpwr scs8hd_buf_1
XFILLER_69_98 vgnd vpwr scs8hd_decap_12
XFILLER_75_431 vgnd vpwr scs8hd_decap_3
XANTENNA_ltile_clb_0.mem_fle_0_in_0.LATCH_2_.latch_SLEEPB _523_/Y vgnd vpwr scs8hd_diode_2
XFILLER_18_80 vgnd vpwr scs8hd_decap_12
XFILLER_35_317 vpwr vgnd scs8hd_fill_2
XFILLER_47_199 vgnd vpwr scs8hd_decap_3
XPHY_570 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_592 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__453__B _451_/X vgnd vpwr scs8hd_diode_2
XPHY_581 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_ltile_clb_0.mux_fle_2_in_0.INVTX1_10_.scs8hd_inv_1_A bottom_width_0_height_0__pin_10_
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_1_.TGATE_0_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_1_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_7_240 vpwr vgnd scs8hd_fill_2
XFILLER_78_280 vgnd vpwr scs8hd_fill_1
XANTENNA_ltile_clb_0.mux_fle_2_in_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_2_in_0.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_66_486 vgnd vpwr scs8hd_decap_12
XFILLER_26_328 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_1_in_1.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_1_in_1.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_19_380 vpwr vgnd scs8hd_fill_2
XFILLER_19_391 vpwr vgnd scs8hd_fill_2
XFILLER_81_489 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mux_fle_1_in_0.INVTX1_9_.scs8hd_inv_1_A right_width_0_height_0__pin_9_
+ vgnd vpwr scs8hd_diode_2
XFILLER_14_27 vgnd vpwr scs8hd_decap_4
XFILLER_34_394 vgnd vpwr scs8hd_fill_1
XANTENNA__363__B _365_/B vgnd vpwr scs8hd_diode_2
XFILLER_30_15 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.mux_fle_2_in_1.INVTX1_0_.scs8hd_inv_1 top_width_0_height_0__pin_0_ ltile_clb_0.mux_fle_2_in_1.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_8_.latch_SLEEPB
+ _590_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_2_in_3.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_2_in_3.INVTX1_10_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_57_464 vpwr vgnd scs8hd_fill_2
XANTENNA__538__B _541_/B vgnd vpwr scs8hd_diode_2
XFILLER_17_306 vgnd vpwr scs8hd_decap_4
X_540_ _540_/A _541_/B _540_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_29_199 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.mux_fle_2_in_2.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_2_in_2.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2/Z
+ ltile_clb_0.mem_fle_2_in_2.LATCH_7_.latch/Q ltile_clb_0.mux_fle_2_in_2.INVTX1_14_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
X_471_ _409_/A _226_/X _384_/A _346_/D _471_/X vgnd vpwr scs8hd_or4_4
XFILLER_25_350 vpwr vgnd scs8hd_fill_2
XFILLER_44_169 vgnd vpwr scs8hd_decap_6
XFILLER_52_191 vgnd vpwr scs8hd_decap_12
XANTENNA__554__A _553_/X vgnd vpwr scs8hd_diode_2
XANTENNA__273__B _272_/X vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_1_in_1.INVTX1_9_.scs8hd_inv_1 right_width_0_height_0__pin_9_
+ ltile_clb_0.mux_fle_1_in_1.INVTX1_9_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_10_.latch_D
+ data_in vgnd vpwr scs8hd_diode_2
Xltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_1_.TGATE_0_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_1_.TGATE_0_.scs8hd_ebufn_2/A
+ _625_/Y ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_ltile_clb_0.mux_fle_0_in_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_0_in_1.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_0_in_3.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_0_in_3.INVTX1_2_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_0_in_3.LATCH_2_.latch/Q ltile_clb_0.mux_fle_0_in_3.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_ltile_clb_0.mux_fle_2_in_1.INVTX1_6_.scs8hd_inv_1_A bottom_width_0_height_0__pin_6_
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_1_in_0.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_1_in_0.INVTX1_13_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_1_in_0.LATCH_1_.latch/Q ltile_clb_0.mux_fle_1_in_0.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
Xltile_clb_0.mux_fle_3_in_0.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_3_in_0.INVTX1_8_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_3_in_0.LATCH_0_.latch/Q ltile_clb_0.mux_fle_3_in_0.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_67_239 vpwr vgnd scs8hd_fill_2
XFILLER_67_228 vpwr vgnd scs8hd_fill_2
XFILLER_0_493 vgnd vpwr scs8hd_decap_3
XFILLER_48_453 vgnd vpwr scs8hd_decap_4
XFILLER_75_250 vpwr vgnd scs8hd_fill_2
XFILLER_48_475 vpwr vgnd scs8hd_fill_2
XFILLER_48_486 vgnd vpwr scs8hd_decap_3
XFILLER_63_456 vpwr vgnd scs8hd_fill_2
XFILLER_63_445 vgnd vpwr scs8hd_decap_4
XANTENNA__448__B _447_/B vgnd vpwr scs8hd_diode_2
XFILLER_35_147 vgnd vpwr scs8hd_decap_6
XFILLER_48_497 vpwr vgnd scs8hd_fill_2
XFILLER_63_467 vpwr vgnd scs8hd_fill_2
XFILLER_16_394 vgnd vpwr scs8hd_decap_3
XFILLER_50_117 vgnd vpwr scs8hd_decap_12
XANTENNA__464__A _431_/A vgnd vpwr scs8hd_diode_2
XFILLER_31_364 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l4_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
+ _626_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_3_.TGATE_1_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_7_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB
+ _604_/Y vgnd vpwr scs8hd_diode_2
XFILLER_58_206 vgnd vpwr scs8hd_decap_8
Xltile_clb_0.mux_fle_2_in_3.mux_l1_in_3_.TGATE_2_.scs8hd_ebufn_2 _651_/HI ltile_clb_0.mem_fle_2_in_3.LATCH_2_.latch/Q
+ ltile_clb_0.mux_fle_2_in_3.mux_l1_in_3_.TGATE_2_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XFILLER_39_453 vpwr vgnd scs8hd_fill_2
XFILLER_54_412 vgnd vpwr scs8hd_decap_8
XFILLER_81_220 vgnd vpwr scs8hd_decap_12
XFILLER_66_294 vgnd vpwr scs8hd_fill_1
XANTENNA__358__B _369_/B vgnd vpwr scs8hd_diode_2
XPHY_26 vgnd vpwr scs8hd_decap_3
XPHY_15 vgnd vpwr scs8hd_decap_3
XPHY_37 vgnd vpwr scs8hd_decap_3
XFILLER_25_15 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mux_fle_3_in_2.INVTX1_3_.scs8hd_inv_1_A left_width_0_height_0__pin_3_
+ vgnd vpwr scs8hd_diode_2
XPHY_48 vgnd vpwr scs8hd_decap_3
XFILLER_25_59 vpwr vgnd scs8hd_fill_2
XPHY_59 vgnd vpwr scs8hd_decap_3
XANTENNA__374__A _374_/A vgnd vpwr scs8hd_diode_2
XFILLER_22_375 vgnd vpwr scs8hd_decap_4
XFILLER_22_386 vgnd vpwr scs8hd_decap_3
Xltile_clb_0.mux_fle_2_in_2.INVTX1_4_.scs8hd_inv_1 top_width_0_height_0__pin_4_ ltile_clb_0.mux_fle_2_in_2.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_ltile_clb_0.mux_fle_2_in_3.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_2_in_3.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_3_in_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_3_in_0.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_66_44 vgnd vpwr scs8hd_decap_12
XANTENNA__549__A _575_/A vgnd vpwr scs8hd_diode_2
XFILLER_45_412 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_3_.scs8hd_inv_1
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_3_.latch/Q
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA__268__B address[1] vgnd vpwr scs8hd_diode_2
XFILLER_82_32 vgnd vpwr scs8hd_decap_12
XFILLER_17_147 vgnd vpwr scs8hd_decap_12
X_523_ _421_/A _517_/X _523_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_32_117 vgnd vpwr scs8hd_decap_12
X_454_ _432_/A _451_/X _454_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_82_87 vgnd vpwr scs8hd_decap_6
XANTENNA__284__A _284_/A vgnd vpwr scs8hd_diode_2
X_385_ _380_/X _427_/B _384_/X _358_/D _385_/X vgnd vpwr scs8hd_or4_4
XFILLER_68_504 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
+ _639_/HI vgnd vpwr scs8hd_diode_2
Xltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_2_.scs8hd_inv_1/Y
+ _605_/Y ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
Xltile_clb_0.mux_fle_0_in_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_0_in_0.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2/Z
+ ltile_clb_0.mem_fle_0_in_0.LATCH_6_.latch/Q ltile_clb_0.mux_fle_0_in_0.INVTX1_14_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA__459__A _437_/A vgnd vpwr scs8hd_diode_2
XFILLER_55_209 vpwr vgnd scs8hd_fill_2
XFILLER_36_434 vpwr vgnd scs8hd_fill_2
XFILLER_36_445 vgnd vpwr scs8hd_decap_8
XANTENNA_ltile_clb_0.mem_fle_3_in_3.LATCH_7_.latch_SLEEPB _323_/Y vgnd vpwr scs8hd_diode_2
XFILLER_11_39 vgnd vpwr scs8hd_decap_12
XANTENNA__369__A address[8] vgnd vpwr scs8hd_diode_2
Xltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_5_.TGATE_1_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_11_.scs8hd_inv_1/Y
+ _604_/Y ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_2_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_27_423 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.mux_fle_1_in_3.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_1_in_3.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2/Z
+ ltile_clb_0.mem_fle_1_in_3.LATCH_7_.latch/Q ltile_clb_0.mux_fle_1_in_3.INVTX1_14_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_27_456 vpwr vgnd scs8hd_fill_2
XFILLER_54_297 vpwr vgnd scs8hd_fill_2
XFILLER_14_117 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.mux_fle_2_in_3.INVTX1_8_.scs8hd_inv_1 top_width_0_height_0__pin_8_ ltile_clb_0.mux_fle_2_in_3.INVTX1_8_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_50_470 vpwr vgnd scs8hd_fill_2
XFILLER_52_68 vgnd vpwr scs8hd_decap_12
XFILLER_10_389 vgnd vpwr scs8hd_decap_8
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_1_.TGATE_0_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XANTENNA__551__B _548_/X vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_0_in_1.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_0_in_1.INVTX1_13_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_0_in_1.LATCH_1_.latch/Q ltile_clb_0.mux_fle_0_in_1.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
Xltile_clb_0.mux_fle_2_in_1.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_2_in_1.INVTX1_8_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_2_in_1.LATCH_0_.latch/Q ltile_clb_0.mux_fle_2_in_1.mux_l1_in_2_.TGATE_3_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
+ _622_/Y vgnd vpwr scs8hd_diode_2
XANTENNA__279__A _278_/X vgnd vpwr scs8hd_diode_2
XFILLER_77_98 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.mux_fle_2_in_0.INVTX1_14_.scs8hd_inv_1 ltile_clb_0.mux_fle_2_in_0.INVTX1_14_.scs8hd_inv_1/A
+ ltile_clb_0.mux_fle_2_in_0.INVTX1_14_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.tap_buf4_0_.scs8hd_inv_1_A
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_60_212 vpwr vgnd scs8hd_fill_2
XFILLER_18_489 vgnd vpwr scs8hd_decap_8
X_506_ _514_/B _511_/B vgnd vpwr scs8hd_buf_1
XFILLER_33_404 vgnd vpwr scs8hd_decap_4
XFILLER_45_297 vpwr vgnd scs8hd_fill_2
XFILLER_26_80 vgnd vpwr scs8hd_decap_12
X_437_ _437_/A _428_/X _437_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_60_267 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_1_in_3.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_1_in_3.INVTX1_12_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_3_in_3.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_3_in_3.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
X_368_ _379_/A _368_/B _368_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_13_172 vpwr vgnd scs8hd_fill_2
XFILLER_9_110 vgnd vpwr scs8hd_decap_12
X_299_ _286_/B address[1] address[3] _258_/X _300_/A vgnd vpwr scs8hd_or4_4
XFILLER_5_360 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_0_in_2.INVTX1_1_.scs8hd_inv_1_A right_width_0_height_0__pin_1_
+ vgnd vpwr scs8hd_diode_2
XFILLER_47_3 vgnd vpwr scs8hd_decap_12
XFILLER_3_51 vgnd vpwr scs8hd_decap_8
XFILLER_3_62 vgnd vpwr scs8hd_decap_12
XFILLER_36_242 vgnd vpwr scs8hd_decap_4
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_5_.TGATE_0_.scs8hd_ebufn_2_TEB
+ _613_/Y vgnd vpwr scs8hd_diode_2
XFILLER_24_437 vgnd vpwr scs8hd_decap_3
XFILLER_51_256 vgnd vpwr scs8hd_decap_3
XFILLER_22_27 vgnd vpwr scs8hd_decap_4
XFILLER_3_319 vgnd vpwr scs8hd_fill_1
XFILLER_59_367 vgnd vpwr scs8hd_fill_1
XFILLER_59_356 vgnd vpwr scs8hd_decap_4
XFILLER_74_337 vpwr vgnd scs8hd_fill_2
XANTENNA__249__D address[1] vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mem_fle_0_in_0.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_70_510 vgnd vpwr scs8hd_decap_6
XANTENNA__546__B _528_/X vgnd vpwr scs8hd_diode_2
XFILLER_27_297 vpwr vgnd scs8hd_fill_2
XFILLER_42_267 vpwr vgnd scs8hd_fill_2
XANTENNA__562__A _554_/X vgnd vpwr scs8hd_diode_2
XFILLER_10_197 vpwr vgnd scs8hd_fill_2
XANTENNA__281__B _539_/A vgnd vpwr scs8hd_diode_2
XFILLER_12_93 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_3_.TGATE_1_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_3_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_0_in_3.INVTX1_10_.scs8hd_inv_1_A bottom_width_0_height_0__pin_10_
+ vgnd vpwr scs8hd_diode_2
XFILLER_65_315 vpwr vgnd scs8hd_fill_2
XFILLER_65_359 vgnd vpwr scs8hd_decap_4
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_1_.latch_SLEEPB
+ _301_/Y vgnd vpwr scs8hd_diode_2
XFILLER_18_231 vgnd vpwr scs8hd_decap_6
XANTENNA__456__B _451_/X vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.mem_ble4_out_0.LATCH_2_.latch_D
+ data_in vgnd vpwr scs8hd_diode_2
XFILLER_33_267 vpwr vgnd scs8hd_fill_2
XANTENNA__472__A _471_/X vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_2_in_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_2_in_2.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_0_in_2.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_0_in_2.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.mem_ble4_out_0.LATCH_2_.latch
+ data_in ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.mem_ble4_out_0.LATCH_2_.latch/Q
+ _549_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_68_197 vgnd vpwr scs8hd_decap_3
XFILLER_68_175 vgnd vpwr scs8hd_decap_8
XFILLER_17_27 vgnd vpwr scs8hd_decap_12
XFILLER_71_329 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_2_in_1.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_2_in_1.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_3_in_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_3_in_0.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XANTENNA__366__B _365_/B vgnd vpwr scs8hd_diode_2
XPHY_207 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_212 vpwr vgnd scs8hd_fill_2
XPHY_229 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_218 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_0_.latch_D
+ data_in vgnd vpwr scs8hd_diode_2
XFILLER_33_15 vgnd vpwr scs8hd_decap_12
XFILLER_24_289 vgnd vpwr scs8hd_decap_12
XFILLER_33_59 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.mux_fle_1_in_2.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_1_in_2.INVTX1_8_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_1_in_2.LATCH_0_.latch/Q ltile_clb_0.mux_fle_1_in_2.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA__382__A _381_/Y vgnd vpwr scs8hd_diode_2
XFILLER_79_418 vgnd vpwr scs8hd_decap_3
XFILLER_58_56 vgnd vpwr scs8hd_decap_12
XFILLER_59_164 vpwr vgnd scs8hd_fill_2
XFILLER_59_175 vpwr vgnd scs8hd_fill_2
XFILLER_47_326 vpwr vgnd scs8hd_fill_2
XFILLER_47_359 vpwr vgnd scs8hd_fill_2
XFILLER_74_44 vgnd vpwr scs8hd_decap_12
XANTENNA__557__A _247_/X vgnd vpwr scs8hd_diode_2
XFILLER_15_212 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.mux_fle_1_in_1.INVTX1_10_.scs8hd_inv_1 bottom_width_0_height_0__pin_10_
+ ltile_clb_0.mux_fle_1_in_1.INVTX1_10_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XFILLER_15_245 vgnd vpwr scs8hd_decap_4
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_14_.scs8hd_inv_1_A
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_14_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XPHY_763 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_752 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_741 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_70_395 vpwr vgnd scs8hd_fill_2
XPHY_730 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_30_215 vgnd vpwr scs8hd_fill_1
XPHY_796 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_785 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_774 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_11_451 vgnd vpwr scs8hd_decap_4
XANTENNA__292__A _267_/X vgnd vpwr scs8hd_diode_2
XFILLER_7_400 vgnd vpwr scs8hd_decap_4
XFILLER_7_466 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_2_in_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_2_in_0.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_7_477 vpwr vgnd scs8hd_fill_2
XFILLER_65_123 vgnd vpwr scs8hd_decap_12
XANTENNA__467__A _434_/A vgnd vpwr scs8hd_diode_2
XFILLER_0_63 vgnd vpwr scs8hd_decap_12
XFILLER_61_384 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.mux_fle_1_in_2.INVTX1_12_.scs8hd_inv_1 top_width_0_height_0__pin_12_
+ ltile_clb_0.mux_fle_1_in_2.INVTX1_12_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
Xltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_5_.latch
+ data_in ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_5_.latch/Q
+ _289_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_28_15 vgnd vpwr scs8hd_decap_12
XFILLER_56_145 vgnd vpwr scs8hd_decap_8
XANTENNA__377__A _338_/A vgnd vpwr scs8hd_diode_2
XFILLER_56_189 vpwr vgnd scs8hd_fill_2
XFILLER_52_351 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_1_in_0.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_1_in_0.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_12_259 vgnd vpwr scs8hd_decap_8
XFILLER_12_248 vpwr vgnd scs8hd_fill_2
XFILLER_60_68 vgnd vpwr scs8hd_decap_12
XFILLER_4_414 vgnd vpwr scs8hd_decap_4
Xltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_2_.TGATE_1_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_2_.TGATE_1_.scs8hd_ebufn_2/A
+ _622_/Y ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_1_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
Xltile_clb_0.mux_fle_1_in_3.INVTX1_14_.scs8hd_inv_1 ltile_clb_0.mux_fle_1_in_3.INVTX1_14_.scs8hd_inv_1/A
+ ltile_clb_0.mux_fle_1_in_3.INVTX1_14_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XANTENNA_ltile_clb_0.mux_fle_3_in_1.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_3_in_1.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_1_in_2.INVTX1_7_.scs8hd_inv_1_A left_width_0_height_0__pin_7_
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mem_fle_0_in_2.LATCH_6_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_75_454 vpwr vgnd scs8hd_fill_2
XFILLER_47_123 vgnd vpwr scs8hd_decap_8
XFILLER_47_134 vpwr vgnd scs8hd_fill_2
XFILLER_75_487 vgnd vpwr scs8hd_fill_1
XFILLER_75_465 vpwr vgnd scs8hd_fill_2
XANTENNA__287__A _278_/X vgnd vpwr scs8hd_diode_2
XFILLER_43_351 vgnd vpwr scs8hd_decap_4
XFILLER_43_362 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.INVTX1_0_.scs8hd_inv_1/Y
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.mem_ble4_out_0.LATCH_0_.latch/Q
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_31_513 vgnd vpwr scs8hd_decap_3
XFILLER_70_192 vpwr vgnd scs8hd_fill_2
XFILLER_34_80 vgnd vpwr scs8hd_decap_12
XPHY_560 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_571 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_593 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_582 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_ltile_clb_0.mem_fle_0_in_3.LATCH_4_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_7_296 vgnd vpwr scs8hd_fill_1
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.buf4_3_.scs8hd_buf_1_A
+ ltile_clb_0.mux_fle_0_in_3.INVTX1_14_.scs8hd_inv_1/Y vgnd vpwr scs8hd_diode_2
XFILLER_66_421 vgnd vpwr scs8hd_decap_8
XFILLER_66_432 vpwr vgnd scs8hd_fill_2
XFILLER_38_145 vpwr vgnd scs8hd_fill_2
XFILLER_38_167 vpwr vgnd scs8hd_fill_2
XFILLER_66_498 vgnd vpwr scs8hd_decap_12
XFILLER_34_351 vgnd vpwr scs8hd_decap_6
Xltile_clb_0.mux_fle_0_in_3.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_0_in_3.INVTX1_8_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_0_in_3.LATCH_0_.latch/Q ltile_clb_0.mux_fle_0_in_3.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_ltile_clb_0.mem_fle_1_in_0.LATCH_6_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_3_in_2.INVTX1_13_.scs8hd_inv_1_A right_width_0_height_0__pin_13_
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_2_in_3.INVTX1_4_.scs8hd_inv_1_A top_width_0_height_0__pin_4_
+ vgnd vpwr scs8hd_diode_2
XFILLER_61_192 vpwr vgnd scs8hd_fill_2
XFILLER_30_27 vgnd vpwr scs8hd_decap_4
XANTENNA_ltile_clb_0.mux_fle_3_in_0.INVTX1_0_.scs8hd_inv_1_A top_width_0_height_0__pin_0_
+ vgnd vpwr scs8hd_diode_2
XFILLER_1_439 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mem_fle_1_in_1.LATCH_4_.latch_D data_in vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_0_in_2.INVTX1_3_.scs8hd_inv_1 left_width_0_height_0__pin_3_ ltile_clb_0.mux_fle_0_in_2.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_29_123 vgnd vpwr scs8hd_decap_12
XFILLER_72_413 vgnd vpwr scs8hd_fill_1
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_1_.scs8hd_inv_1_A
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
X_470_ _437_/A _461_/X _470_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_13_502 vpwr vgnd scs8hd_fill_2
XFILLER_25_362 vpwr vgnd scs8hd_fill_2
XFILLER_9_506 vgnd vpwr scs8hd_decap_8
XFILLER_40_321 vgnd vpwr scs8hd_decap_4
XFILLER_40_376 vpwr vgnd scs8hd_fill_2
XFILLER_40_398 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mem_fle_1_in_2.LATCH_2_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA__570__A _544_/A vgnd vpwr scs8hd_diode_2
XFILLER_20_93 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mux_fle_1_in_3.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_1_in_3.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_0_450 vpwr vgnd scs8hd_fill_2
XFILLER_0_461 vgnd vpwr scs8hd_decap_4
Xltile_clb_0.mux_fle_2_in_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_2_in_0.INVTX1_2_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_2_in_0.LATCH_2_.latch/Q ltile_clb_0.mux_fle_2_in_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_ltile_clb_0.mux_fle_2_in_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_2_in_0.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_0_in_0.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_0_in_0.INVTX1_7_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_0_in_0.LATCH_3_.latch/Q ltile_clb_0.mux_fle_0_in_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_48_421 vgnd vpwr scs8hd_decap_8
XFILLER_48_432 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mem_fle_1_in_3.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_63_424 vgnd vpwr scs8hd_fill_1
Xltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_5_.latch
+ data_in ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_5_.latch/Q
+ _593_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
X_599_ _599_/A _578_/X _599_/X vgnd vpwr scs8hd_or2_4
XFILLER_50_129 vgnd vpwr scs8hd_decap_6
XFILLER_31_321 vpwr vgnd scs8hd_fill_2
XFILLER_31_343 vpwr vgnd scs8hd_fill_2
XANTENNA__464__B _462_/X vgnd vpwr scs8hd_diode_2
XFILLER_31_354 vpwr vgnd scs8hd_fill_2
XFILLER_77_3 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mux_fle_3_in_2.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_3_in_2.INVTX1_12_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XPHY_390 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__480__A _436_/A vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mem_fle_2_in_0.LATCH_2_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_0_in_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_0_in_1.LATCH_4_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_58_218 vgnd vpwr scs8hd_decap_3
XANTENNA_ltile_clb_0.mux_fle_1_in_0.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_1_in_0.INVTX1_8_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__358__C _369_/C vgnd vpwr scs8hd_diode_2
XFILLER_81_232 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.mux_fle_3_in_3.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_3_in_3.INVTX1_3_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_3_in_3.LATCH_3_.latch/Q ltile_clb_0.mux_fle_3_in_3.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_54_468 vgnd vpwr scs8hd_decap_4
XPHY_16 vgnd vpwr scs8hd_decap_3
XPHY_27 vgnd vpwr scs8hd_decap_3
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_6_.latch_D
+ data_in vgnd vpwr scs8hd_diode_2
XPHY_38 vgnd vpwr scs8hd_decap_3
XFILLER_25_27 vgnd vpwr scs8hd_decap_12
XFILLER_81_298 vgnd vpwr scs8hd_decap_6
XPHY_49 vgnd vpwr scs8hd_decap_3
XANTENNA__374__B _377_/B vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mem_fle_2_in_1.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_34_192 vgnd vpwr scs8hd_decap_8
XFILLER_22_398 vgnd vpwr scs8hd_fill_1
XFILLER_41_15 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mux_fle_3_in_3.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_3_in_3.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_41_59 vpwr vgnd scs8hd_fill_2
XANTENNA__390__A _374_/A vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_3_in_1.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_3_in_1.LATCH_7_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_0_in_3.INVTX1_7_.scs8hd_inv_1 left_width_0_height_0__pin_7_ ltile_clb_0.mux_fle_0_in_3.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_1_236 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.mem_ble4_out_0.LATCH_2_.latch
+ data_in ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.mem_ble4_out_0.LATCH_2_.latch/Q
+ _601_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA__549__B _548_/X vgnd vpwr scs8hd_diode_2
XFILLER_66_56 vgnd vpwr scs8hd_decap_12
XFILLER_57_262 vpwr vgnd scs8hd_fill_2
XFILLER_57_295 vpwr vgnd scs8hd_fill_2
XFILLER_57_273 vgnd vpwr scs8hd_decap_3
XFILLER_45_424 vgnd vpwr scs8hd_fill_1
XFILLER_72_243 vgnd vpwr scs8hd_decap_12
XFILLER_17_159 vgnd vpwr scs8hd_decap_12
X_522_ _334_/A _517_/X _522_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_82_44 vgnd vpwr scs8hd_decap_12
XFILLER_60_416 vgnd vpwr scs8hd_decap_12
XANTENNA__565__A _539_/A vgnd vpwr scs8hd_diode_2
XFILLER_32_129 vgnd vpwr scs8hd_decap_12
X_453_ _431_/A _451_/X _453_/Y vgnd vpwr scs8hd_nor2_4
X_384_ _384_/A _384_/X vgnd vpwr scs8hd_buf_1
XFILLER_9_314 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2_TEB
+ _605_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_1_in_1.INVTX1_12_.scs8hd_inv_1_A top_width_0_height_0__pin_12_
+ vgnd vpwr scs8hd_diode_2
XANTENNA__459__B _450_/X vgnd vpwr scs8hd_diode_2
XFILLER_48_251 vgnd vpwr scs8hd_decap_3
XFILLER_63_221 vpwr vgnd scs8hd_fill_2
XFILLER_63_254 vpwr vgnd scs8hd_fill_2
XFILLER_63_232 vpwr vgnd scs8hd_fill_2
XFILLER_36_457 vgnd vpwr scs8hd_fill_1
XFILLER_36_468 vgnd vpwr scs8hd_decap_3
XFILLER_63_298 vpwr vgnd scs8hd_fill_2
XFILLER_63_265 vgnd vpwr scs8hd_decap_3
XFILLER_51_416 vpwr vgnd scs8hd_fill_2
XANTENNA__475__A _431_/A vgnd vpwr scs8hd_diode_2
XFILLER_16_192 vgnd vpwr scs8hd_decap_3
XANTENNA_ltile_clb_0.mux_fle_2_in_3.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_2_in_3.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_2_in_1.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_2_in_1.mux_l1_in_2_.TGATE_3_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XANTENNA__369__B _369_/B vgnd vpwr scs8hd_diode_2
XFILLER_39_240 vgnd vpwr scs8hd_fill_1
XFILLER_39_262 vpwr vgnd scs8hd_fill_2
XFILLER_27_435 vgnd vpwr scs8hd_decap_4
XFILLER_36_15 vgnd vpwr scs8hd_decap_12
XFILLER_39_273 vpwr vgnd scs8hd_fill_2
XANTENNA__385__A _380_/X vgnd vpwr scs8hd_diode_2
XFILLER_54_287 vpwr vgnd scs8hd_fill_2
XFILLER_54_276 vgnd vpwr scs8hd_decap_8
XFILLER_42_405 vpwr vgnd scs8hd_fill_2
XFILLER_14_129 vgnd vpwr scs8hd_decap_12
XFILLER_42_449 vgnd vpwr scs8hd_decap_8
Xltile_clb_0.mux_fle_3_in_0.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_3_in_0.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2/Z
+ ltile_clb_0.mem_fle_3_in_0.LATCH_7_.latch/Q ltile_clb_0.mux_fle_3_in_0.INVTX1_14_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_10_302 vgnd vpwr scs8hd_decap_8
XFILLER_10_346 vgnd vpwr scs8hd_decap_4
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_2_.latch_D
+ data_in vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_3_in_3.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_3_in_3.INVTX1_10_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_3_.scs8hd_inv_1_A
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_7_3 vgnd vpwr scs8hd_decap_12
XFILLER_77_313 vgnd vpwr scs8hd_decap_3
XFILLER_77_302 vgnd vpwr scs8hd_decap_3
Xltile_clb_0.mux_fle_1_in_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_1_in_1.INVTX1_2_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_1_in_1.LATCH_2_.latch/Q ltile_clb_0.mux_fle_1_in_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
Xltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_5_.latch
+ data_in ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_5_.latch/Q
+ _567_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_65_508 vgnd vpwr scs8hd_decap_8
XANTENNA__279__B _313_/A vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_10_.latch_SLEEPB
+ _266_/Y vgnd vpwr scs8hd_diode_2
XFILLER_18_457 vgnd vpwr scs8hd_fill_1
XANTENNA__295__A _304_/A vgnd vpwr scs8hd_diode_2
X_505_ _504_/X _514_/B vgnd vpwr scs8hd_buf_1
Xltile_clb_0.mux_fle_2_in_0.INVTX1_4_.scs8hd_inv_1 top_width_0_height_0__pin_4_ ltile_clb_0.mux_fle_2_in_0.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_ltile_clb_0.mux_fle_1_in_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_1_in_1.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
X_436_ _436_/A _428_/X _436_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_60_257 vgnd vpwr scs8hd_decap_8
X_367_ _394_/A _368_/B _367_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_13_184 vpwr vgnd scs8hd_fill_2
XFILLER_42_80 vgnd vpwr scs8hd_decap_12
X_298_ _304_/A _544_/A _298_/Y vgnd vpwr scs8hd_nor2_4
Xltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_6_.scs8hd_inv_1/Y
+ _613_/Y ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_1_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_68_346 vgnd vpwr scs8hd_decap_3
XFILLER_3_74 vgnd vpwr scs8hd_decap_12
XFILLER_36_210 vgnd vpwr scs8hd_decap_4
Xltile_clb_0.mux_fle_3_in_1.mux_l1_in_3_.TGATE_2_.scs8hd_ebufn_2 _653_/HI ltile_clb_0.mem_fle_3_in_1.LATCH_2_.latch/Q
+ ltile_clb_0.mux_fle_3_in_1.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XFILLER_36_221 vgnd vpwr scs8hd_fill_1
XFILLER_36_265 vpwr vgnd scs8hd_fill_2
XFILLER_24_449 vgnd vpwr scs8hd_decap_8
XFILLER_36_298 vgnd vpwr scs8hd_fill_1
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB
+ _623_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_1_in_2.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_1_in_2.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_59_313 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_7_.TGATE_1_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_15_.scs8hd_inv_1/Y
+ _612_/Y ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_3_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_59_335 vpwr vgnd scs8hd_fill_2
XFILLER_59_324 vpwr vgnd scs8hd_fill_2
XFILLER_74_327 vgnd vpwr scs8hd_decap_8
XFILLER_27_210 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mem_fle_2_in_3.LATCH_6_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_1_in_1.mux_l1_in_2_.TGATE_3_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_1_in_1.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_10_154 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_6_.scs8hd_inv_1
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_6_.latch/Q
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_ltile_clb_0.mem_fle_2_in_3.LATCH_2_.latch_SLEEPB _393_/Y vgnd vpwr scs8hd_diode_2
XFILLER_77_110 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_4_.TGATE_1_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_9_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_77_198 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.mux_fle_2_in_1.INVTX1_8_.scs8hd_inv_1 top_width_0_height_0__pin_8_ ltile_clb_0.mux_fle_2_in_1.INVTX1_8_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_73_360 vgnd vpwr scs8hd_decap_4
XFILLER_18_276 vpwr vgnd scs8hd_fill_2
XFILLER_73_393 vgnd vpwr scs8hd_decap_4
XFILLER_18_298 vgnd vpwr scs8hd_fill_1
XFILLER_33_235 vgnd vpwr scs8hd_decap_8
X_419_ _334_/A _434_/A vgnd vpwr scs8hd_buf_1
XANTENNA_ltile_clb_0.mem_fle_3_in_1.LATCH_6_.latch_D data_in vgnd vpwr scs8hd_diode_2
Xltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_0_.TGATE_0_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ _609_/Y ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l4_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_68_154 vgnd vpwr scs8hd_decap_8
XANTENNA_ltile_clb_0.mem_fle_3_in_2.LATCH_4_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_17_39 vgnd vpwr scs8hd_decap_12
XFILLER_64_393 vgnd vpwr scs8hd_decap_4
Xltile_clb_0.mux_fle_2_in_1.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_2_in_1.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2/Z
+ ltile_clb_0.mem_fle_2_in_1.LATCH_7_.latch/Q ltile_clb_0.mux_fle_2_in_1.INVTX1_14_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XPHY_219 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_208 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_33_27 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mux_fle_3_in_0.INVTX1_10_.scs8hd_inv_1_A bottom_width_0_height_0__pin_10_
+ vgnd vpwr scs8hd_diode_2
XFILLER_32_290 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_5_.latch
+ data_in ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_5_.latch/Q
+ _541_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
Xltile_clb_0.mux_fle_0_in_2.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_0_in_2.INVTX1_2_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_0_in_2.LATCH_2_.latch/Q ltile_clb_0.mux_fle_0_in_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_ltile_clb_0.mem_fle_3_in_3.LATCH_2_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_59_110 vgnd vpwr scs8hd_decap_12
XFILLER_58_68 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mux_fle_0_in_3.INVTX1_8_.scs8hd_inv_1_A top_width_0_height_0__pin_8_
+ vgnd vpwr scs8hd_diode_2
XFILLER_74_56 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.mux_fle_3_in_2.INVTX1_3_.scs8hd_inv_1 left_width_0_height_0__pin_3_ ltile_clb_0.mux_fle_3_in_2.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA__557__B _558_/B vgnd vpwr scs8hd_diode_2
XFILLER_43_511 vgnd vpwr scs8hd_decap_4
XANTENNA_ltile_clb_0.mux_fle_1_in_0.INVTX1_4_.scs8hd_inv_1_A top_width_0_height_0__pin_4_
+ vgnd vpwr scs8hd_diode_2
XFILLER_55_393 vpwr vgnd scs8hd_fill_2
XFILLER_15_235 vpwr vgnd scs8hd_fill_2
XPHY_720 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_753 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_742 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_731 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_ltile_clb_0.mem_fle_3_in_2.LATCH_2_.latch_SLEEPB _354_/Y vgnd vpwr scs8hd_diode_2
XANTENNA__573__A _599_/A vgnd vpwr scs8hd_diode_2
XPHY_786 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_775 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_764 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_ltile_clb_0.mux_fle_2_in_2.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_2_in_2.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XPHY_797 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__292__B _542_/A vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_4_.latch_SLEEPB
+ _568_/Y vgnd vpwr scs8hd_diode_2
XFILLER_78_430 vgnd vpwr scs8hd_decap_4
Xltile_clb_0.mux_fle_2_in_2.mux_l1_in_3_.TGATE_2_.scs8hd_ebufn_2 _650_/HI ltile_clb_0.mem_fle_2_in_2.LATCH_2_.latch/Q
+ ltile_clb_0.mux_fle_2_in_2.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XANTENNA_ltile_clb_0.mux_fle_2_in_3.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_2_in_3.INVTX1_12_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_65_135 vgnd vpwr scs8hd_decap_12
XFILLER_80_105 vgnd vpwr scs8hd_decap_12
XFILLER_65_157 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_2_in_1.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_2_in_1.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__467__B _462_/X vgnd vpwr scs8hd_diode_2
XFILLER_0_75 vgnd vpwr scs8hd_decap_12
XFILLER_73_190 vpwr vgnd scs8hd_fill_2
XFILLER_61_341 vpwr vgnd scs8hd_fill_2
XANTENNA__483__A _482_/X vgnd vpwr scs8hd_diode_2
XFILLER_9_62 vgnd vpwr scs8hd_decap_12
XFILLER_9_51 vgnd vpwr scs8hd_decap_8
XFILLER_21_249 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_0_in_1.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_0_in_1.INVTX1_8_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mem_fle_0_in_3.LATCH_3_.latch_SLEEPB _489_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_2_in_1.INVTX1_1_.scs8hd_inv_1_A right_width_0_height_0__pin_1_
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_16_.scs8hd_inv_1_A
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_16_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_69_485 vgnd vpwr scs8hd_decap_3
XFILLER_28_27 vgnd vpwr scs8hd_decap_4
XFILLER_29_327 vpwr vgnd scs8hd_fill_2
XFILLER_56_135 vgnd vpwr scs8hd_fill_1
XANTENNA__377__B _377_/B vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_3_in_3.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_3_in_3.LATCH_6_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_44_15 vgnd vpwr scs8hd_decap_12
XANTENNA__393__A _338_/A vgnd vpwr scs8hd_diode_2
XFILLER_52_396 vgnd vpwr scs8hd_fill_1
XFILLER_12_205 vgnd vpwr scs8hd_decap_8
Xltile_clb_0.mem_fle_0_in_1.LATCH_7_.latch data_in ltile_clb_0.mem_fle_0_in_1.LATCH_7_.latch/Q
+ _507_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_8_.latch_D
+ data_in vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_1_.scs8hd_inv_1_A
+ ltile_clb_0.mux_fle_0_in_1.INVTX1_14_.scs8hd_inv_1/Y vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.mem_ble4_out_0.LATCH_2_.latch_D
+ data_in vgnd vpwr scs8hd_diode_2
XFILLER_4_459 vgnd vpwr scs8hd_decap_3
Xltile_clb_0.mux_fle_3_in_3.INVTX1_7_.scs8hd_inv_1 left_width_0_height_0__pin_7_ ltile_clb_0.mux_fle_3_in_3.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
Xltile_clb_0.mem_fle_1_in_1.LATCH_6_.latch data_in ltile_clb_0.mem_fle_1_in_1.LATCH_6_.latch/Q
+ _464_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_75_422 vgnd vpwr scs8hd_decap_3
XANTENNA__568__A _542_/A vgnd vpwr scs8hd_diode_2
XFILLER_62_105 vgnd vpwr scs8hd_decap_12
XANTENNA__287__B _286_/X vgnd vpwr scs8hd_diode_2
XFILLER_47_157 vpwr vgnd scs8hd_fill_2
XFILLER_47_179 vpwr vgnd scs8hd_fill_2
XFILLER_18_93 vgnd vpwr scs8hd_decap_12
XFILLER_28_371 vgnd vpwr scs8hd_decap_3
XFILLER_28_382 vpwr vgnd scs8hd_fill_2
XFILLER_62_149 vpwr vgnd scs8hd_fill_2
XFILLER_43_330 vpwr vgnd scs8hd_fill_2
XFILLER_43_341 vpwr vgnd scs8hd_fill_2
XFILLER_70_171 vpwr vgnd scs8hd_fill_2
XFILLER_43_374 vgnd vpwr scs8hd_decap_4
Xltile_clb_0.mem_fle_2_in_1.LATCH_5_.latch data_in ltile_clb_0.mem_fle_2_in_1.LATCH_5_.latch/Q
+ _416_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XPHY_550 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_561 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_594 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_572 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_583 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_7_275 vpwr vgnd scs8hd_fill_2
XFILLER_50_80 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.mem_fle_3_in_1.LATCH_4_.latch data_in ltile_clb_0.mem_fle_3_in_1.LATCH_4_.latch/Q
+ _364_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_22_3 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.mux_fle_1_in_2.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_1_in_2.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2/Z
+ ltile_clb_0.mem_fle_1_in_2.LATCH_7_.latch/Q ltile_clb_0.mux_fle_1_in_2.INVTX1_14_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA__478__A _434_/A vgnd vpwr scs8hd_diode_2
XFILLER_81_447 vgnd vpwr scs8hd_decap_12
XFILLER_53_138 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mem_fle_1_in_2.LATCH_3_.latch_SLEEPB _456_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_1_in_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_1_in_0.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_53_149 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ _631_/Y ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_61_171 vgnd vpwr scs8hd_fill_1
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_7_.TGATE_1_.scs8hd_ebufn_2_TEB
+ _604_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_1_in_2.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_1_in_2.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_2_in_0.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_2_in_0.INVTX1_8_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_2_in_0.LATCH_0_.latch/Q ltile_clb_0.mux_fle_2_in_0.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
Xltile_clb_0.mux_fle_0_in_0.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_0_in_0.INVTX1_13_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_0_in_0.LATCH_1_.latch/Q ltile_clb_0.mux_fle_0_in_0.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_39_15 vgnd vpwr scs8hd_decap_12
XFILLER_69_260 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_4_.TGATE_1_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_9_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_39_59 vpwr vgnd scs8hd_fill_2
XANTENNA__388__A _388_/A vgnd vpwr scs8hd_diode_2
XFILLER_57_433 vpwr vgnd scs8hd_fill_2
XFILLER_29_135 vgnd vpwr scs8hd_decap_12
XFILLER_29_179 vpwr vgnd scs8hd_fill_2
XFILLER_72_436 vgnd vpwr scs8hd_decap_4
XFILLER_44_105 vgnd vpwr scs8hd_decap_12
XFILLER_13_514 vpwr vgnd scs8hd_fill_2
XFILLER_25_396 vpwr vgnd scs8hd_fill_2
XFILLER_40_333 vgnd vpwr scs8hd_decap_3
XFILLER_4_212 vpwr vgnd scs8hd_fill_2
XANTENNA__570__B _554_/X vgnd vpwr scs8hd_diode_2
XFILLER_4_267 vgnd vpwr scs8hd_decap_8
Xltile_clb_0.mux_fle_1_in_3.mux_l1_in_3_.TGATE_2_.scs8hd_ebufn_2 _647_/HI ltile_clb_0.mem_fle_1_in_3.LATCH_2_.latch/Q
+ ltile_clb_0.mux_fle_1_in_3.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
Xltile_clb_0.mux_fle_3_in_3.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_3_in_3.INVTX1_9_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_3_in_3.LATCH_1_.latch/Q ltile_clb_0.mux_fle_3_in_3.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_ltile_clb_0.mux_fle_0_in_2.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_0_in_2.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_67_208 vgnd vpwr scs8hd_fill_1
XFILLER_0_473 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.tap_buf4_0_.scs8hd_inv_1_A
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_48_411 vgnd vpwr scs8hd_fill_1
XANTENNA__298__A _304_/A vgnd vpwr scs8hd_diode_2
XFILLER_63_403 vpwr vgnd scs8hd_fill_2
X_598_ _546_/A _580_/X _598_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_16_352 vgnd vpwr scs8hd_decap_4
XFILLER_43_160 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.mem_fle_3_in_3.LATCH_7_.latch data_in ltile_clb_0.mem_fle_3_in_3.LATCH_7_.latch/Q
+ _323_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_ltile_clb_0.mux_fle_3_in_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_3_in_0.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_clkbuf_1_1_0_clk_A clkbuf_0_clk/X vgnd vpwr scs8hd_diode_2
XPHY_380 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_391 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_31_388 vgnd vpwr scs8hd_decap_4
XANTENNA__480__B _481_/B vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mem_fle_2_in_1.LATCH_3_.latch_SLEEPB _420_/Y vgnd vpwr scs8hd_diode_2
XFILLER_39_466 vgnd vpwr scs8hd_decap_3
XFILLER_39_477 vpwr vgnd scs8hd_fill_2
XFILLER_66_285 vgnd vpwr scs8hd_decap_3
XFILLER_54_436 vgnd vpwr scs8hd_decap_3
XANTENNA__358__D _358_/D vgnd vpwr scs8hd_diode_2
XFILLER_26_105 vgnd vpwr scs8hd_decap_12
XPHY_28 vgnd vpwr scs8hd_decap_3
XPHY_17 vgnd vpwr scs8hd_decap_3
XPHY_39 vgnd vpwr scs8hd_decap_3
XFILLER_25_39 vgnd vpwr scs8hd_decap_12
XFILLER_10_506 vgnd vpwr scs8hd_decap_8
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_9_.latch_SLEEPB
+ _273_/Y vgnd vpwr scs8hd_diode_2
XFILLER_41_27 vgnd vpwr scs8hd_decap_12
XANTENNA__390__B _388_/B vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_1_in_3.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_1_in_3.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_2_in_0.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_2_in_0.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_66_68 vgnd vpwr scs8hd_decap_12
XFILLER_57_241 vgnd vpwr scs8hd_decap_3
XFILLER_57_230 vgnd vpwr scs8hd_decap_4
XFILLER_72_255 vgnd vpwr scs8hd_fill_1
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_10_.latch_D
+ data_in vgnd vpwr scs8hd_diode_2
X_521_ _331_/A _517_/X _521_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_45_447 vgnd vpwr scs8hd_decap_4
XFILLER_82_56 vgnd vpwr scs8hd_decap_6
XFILLER_72_288 vpwr vgnd scs8hd_fill_2
XFILLER_60_428 vgnd vpwr scs8hd_fill_1
XANTENNA__565__B _564_/B vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
X_452_ _430_/A _451_/X _452_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_72_299 vpwr vgnd scs8hd_fill_2
X_383_ address[8] _369_/B _384_/A vgnd vpwr scs8hd_nand2_4
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_2_.scs8hd_inv_1_A
+ ltile_clb_0.mux_fle_3_in_2.INVTX1_14_.scs8hd_inv_1/Y vgnd vpwr scs8hd_diode_2
XFILLER_25_171 vgnd vpwr scs8hd_decap_6
XFILLER_25_193 vgnd vpwr scs8hd_decap_4
XFILLER_9_304 vgnd vpwr scs8hd_fill_1
XFILLER_40_141 vgnd vpwr scs8hd_fill_1
XANTENNA__581__A _580_/X vgnd vpwr scs8hd_diode_2
XFILLER_13_388 vpwr vgnd scs8hd_fill_2
XFILLER_13_399 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.mux_fle_0_in_0.INVTX1_3_.scs8hd_inv_1 left_width_0_height_0__pin_3_ ltile_clb_0.mux_fle_0_in_0.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
Xltile_clb_0.mux_fle_0_in_3.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_0_in_3.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2/Z
+ ltile_clb_0.mem_fle_0_in_3.LATCH_7_.latch/Q ltile_clb_0.mux_fle_0_in_3.INVTX1_14_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_ltile_clb_0.mux_fle_3_in_1.INVTX1_7_.scs8hd_inv_1_A left_width_0_height_0__pin_7_
+ vgnd vpwr scs8hd_diode_2
XFILLER_0_270 vpwr vgnd scs8hd_fill_2
XFILLER_63_200 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
+ _615_/Y vgnd vpwr scs8hd_diode_2
XFILLER_48_274 vgnd vpwr scs8hd_fill_1
XANTENNA_ltile_clb_0.mem_fle_3_in_0.LATCH_3_.latch_SLEEPB _376_/Y vgnd vpwr scs8hd_diode_2
XFILLER_63_277 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_4_.scs8hd_inv_1
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_4_.latch/Q
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA__475__B _479_/B vgnd vpwr scs8hd_diode_2
XFILLER_51_439 vpwr vgnd scs8hd_fill_2
XFILLER_31_163 vgnd vpwr scs8hd_fill_1
Xltile_clb_0.mux_fle_1_in_1.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_1_in_1.INVTX1_8_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_1_in_1.LATCH_0_.latch/Q ltile_clb_0.mux_fle_1_in_1.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA__491__A _423_/A vgnd vpwr scs8hd_diode_2
XFILLER_8_370 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_1_in_3.INVTX1_10_.scs8hd_inv_1_A bottom_width_0_height_0__pin_10_
+ vgnd vpwr scs8hd_diode_2
XANTENNA__369__C _369_/C vgnd vpwr scs8hd_diode_2
XFILLER_39_252 vgnd vpwr scs8hd_decap_4
XFILLER_54_211 vgnd vpwr scs8hd_decap_3
XFILLER_36_27 vgnd vpwr scs8hd_decap_4
XFILLER_39_285 vgnd vpwr scs8hd_fill_1
XFILLER_54_244 vgnd vpwr scs8hd_decap_8
XFILLER_27_469 vgnd vpwr scs8hd_decap_4
XANTENNA__385__B _427_/B vgnd vpwr scs8hd_diode_2
XFILLER_54_255 vgnd vpwr scs8hd_decap_3
XFILLER_52_15 vgnd vpwr scs8hd_decap_12
XFILLER_35_480 vpwr vgnd scs8hd_fill_2
XFILLER_22_141 vgnd vpwr scs8hd_decap_12
XFILLER_50_450 vpwr vgnd scs8hd_fill_2
XFILLER_10_325 vgnd vpwr scs8hd_decap_3
XFILLER_22_174 vgnd vpwr scs8hd_decap_3
XANTENNA_ltile_clb_0.mem_fle_0_in_1.LATCH_4_.latch_SLEEPB _510_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_0_in_2.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_0_in_2.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_18_414 vgnd vpwr scs8hd_decap_8
XANTENNA__576__A _270_/B vgnd vpwr scs8hd_diode_2
XFILLER_45_222 vgnd vpwr scs8hd_fill_1
X_504_ _409_/A _381_/Y _228_/X _526_/D _504_/X vgnd vpwr scs8hd_or4_4
XANTENNA__295__B _569_/A vgnd vpwr scs8hd_diode_2
XFILLER_26_93 vgnd vpwr scs8hd_decap_12
XFILLER_26_480 vgnd vpwr scs8hd_decap_4
XFILLER_33_439 vpwr vgnd scs8hd_fill_2
X_435_ _435_/A _429_/X _435_/Y vgnd vpwr scs8hd_nor2_4
X_366_ _338_/A _365_/B _366_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_9_123 vgnd vpwr scs8hd_decap_12
X_297_ _296_/X _544_/A vgnd vpwr scs8hd_buf_1
Xltile_clb_0.mux_fle_0_in_1.INVTX1_7_.scs8hd_inv_1 left_width_0_height_0__pin_7_ ltile_clb_0.mux_fle_0_in_1.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_ltile_clb_0.mux_fle_2_in_3.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_2_in_3.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_5_340 vgnd vpwr scs8hd_decap_4
XFILLER_3_86 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_1_.TGATE_1_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_1_.TGATE_1_.scs8hd_ebufn_2/A
+ _606_/Y ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
Xltile_clb_0.mem_fle_0_in_0.LATCH_0_.latch data_in ltile_clb_0.mem_fle_0_in_0.LATCH_0_.latch/Q
+ _525_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA__486__A _325_/A vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_0_in_0.INVTX1_10_.scs8hd_inv_1 bottom_width_0_height_0__pin_10_
+ ltile_clb_0.mux_fle_0_in_0.INVTX1_10_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XFILLER_51_236 vgnd vpwr scs8hd_decap_4
XFILLER_51_225 vpwr vgnd scs8hd_fill_2
XFILLER_51_269 vpwr vgnd scs8hd_fill_2
XFILLER_32_450 vgnd vpwr scs8hd_decap_4
XFILLER_32_483 vgnd vpwr scs8hd_fill_1
XFILLER_32_494 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mux_fle_2_in_0.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_2_in_0.INVTX1_8_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_59_303 vpwr vgnd scs8hd_fill_2
XFILLER_47_15 vgnd vpwr scs8hd_decap_12
XFILLER_47_59 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mem_fle_1_in_0.LATCH_4_.latch_SLEEPB _477_/Y vgnd vpwr scs8hd_diode_2
XFILLER_67_391 vpwr vgnd scs8hd_fill_2
XANTENNA__396__A _380_/X vgnd vpwr scs8hd_diode_2
XFILLER_27_277 vpwr vgnd scs8hd_fill_2
XFILLER_15_428 vpwr vgnd scs8hd_fill_2
XFILLER_42_225 vpwr vgnd scs8hd_fill_2
XFILLER_30_409 vgnd vpwr scs8hd_decap_8
XANTENNA_ltile_clb_0.mux_fle_0_in_1.INVTX1_5_.scs8hd_inv_1_A right_width_0_height_0__pin_5_
+ vgnd vpwr scs8hd_diode_2
XFILLER_42_247 vgnd vpwr scs8hd_decap_8
XFILLER_23_472 vgnd vpwr scs8hd_decap_3
Xltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.buf4_2_.scs8hd_buf_1
+ ltile_clb_0.mux_fle_0_in_2.INVTX1_14_.scs8hd_inv_1/Y _632_/A vgnd vpwr scs8hd_buf_1
Xltile_clb_0.mux_fle_0_in_1.INVTX1_12_.scs8hd_inv_1 top_width_0_height_0__pin_12_
+ ltile_clb_0.mux_fle_0_in_1.INVTX1_12_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XFILLER_10_166 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.mux_fle_1_in_2.INVTX1_2_.scs8hd_inv_1 bottom_width_0_height_0__pin_2_
+ ltile_clb_0.mux_fle_1_in_2.INVTX1_2_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
Xltile_clb_0.mux_fle_3_in_1.INVTX1_11_.scs8hd_inv_1 left_width_0_height_0__pin_11_
+ ltile_clb_0.mux_fle_3_in_1.INVTX1_11_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XFILLER_2_398 vgnd vpwr scs8hd_decap_4
XFILLER_65_339 vgnd vpwr scs8hd_decap_3
XFILLER_33_214 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.mux_fle_0_in_2.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_0_in_2.INVTX1_8_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_0_in_2.LATCH_0_.latch/Q ltile_clb_0.mux_fle_0_in_2.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
Xltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_5_.TGATE_0_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_10_.scs8hd_inv_1/Y
+ _621_/Y ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_2_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_14_450 vgnd vpwr scs8hd_decap_8
X_418_ _433_/A _412_/B _418_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA_ltile_clb_0.mux_fle_0_in_2.INVTX1_14_.scs8hd_inv_1_A ltile_clb_0.mux_fle_0_in_2.INVTX1_14_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_41_291 vpwr vgnd scs8hd_fill_2
X_349_ _388_/A _353_/B _349_/Y vgnd vpwr scs8hd_nor2_4
Xltile_clb_0.mem_fle_0_in_2.LATCH_3_.latch data_in ltile_clb_0.mem_fle_0_in_2.LATCH_3_.latch/Q
+ _500_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_52_3 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.mux_fle_0_in_2.INVTX1_14_.scs8hd_inv_1 ltile_clb_0.mux_fle_0_in_2.INVTX1_14_.scs8hd_inv_1/A
+ ltile_clb_0.mux_fle_0_in_2.INVTX1_14_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XANTENNA_ltile_clb_0.mux_fle_1_in_2.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_1_in_2.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_1_in_2.INVTX1_2_.scs8hd_inv_1_A bottom_width_0_height_0__pin_2_
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_3_in_2.INVTX1_13_.scs8hd_inv_1 right_width_0_height_0__pin_13_
+ ltile_clb_0.mux_fle_3_in_2.INVTX1_13_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XFILLER_56_328 vpwr vgnd scs8hd_fill_2
XFILLER_56_306 vgnd vpwr scs8hd_decap_4
XANTENNA_ltile_clb_0.mux_fle_0_in_3.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_0_in_3.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mem_fle_1_in_2.LATCH_2_.latch data_in ltile_clb_0.mem_fle_1_in_2.LATCH_2_.latch/Q
+ _457_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_64_361 vgnd vpwr scs8hd_decap_8
XFILLER_24_225 vgnd vpwr scs8hd_decap_8
XFILLER_12_409 vgnd vpwr scs8hd_decap_8
XPHY_209 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_247 vgnd vpwr scs8hd_decap_4
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_1_in_1.mux_l1_in_3_.TGATE_2_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_1_in_1.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_33_39 vgnd vpwr scs8hd_decap_12
XFILLER_20_420 vgnd vpwr scs8hd_decap_6
Xltile_clb_0.mem_fle_2_in_2.LATCH_1_.latch data_in ltile_clb_0.mem_fle_2_in_2.LATCH_1_.latch/Q
+ _405_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_ltile_clb_0.mux_fle_3_in_1.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_3_in_1.mux_l1_in_2_.TGATE_3_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_13_.latch
+ data_in ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_13_.latch/Q
+ _532_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
Xltile_clb_0.mem_fle_3_in_2.LATCH_0_.latch data_in ltile_clb_0.mem_fle_3_in_2.LATCH_0_.latch/Q
+ _356_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_59_188 vpwr vgnd scs8hd_fill_2
XFILLER_47_317 vpwr vgnd scs8hd_fill_2
XFILLER_74_158 vpwr vgnd scs8hd_fill_2
XFILLER_74_68 vgnd vpwr scs8hd_decap_12
XFILLER_62_309 vgnd vpwr scs8hd_fill_1
XFILLER_82_180 vgnd vpwr scs8hd_decap_6
XPHY_710 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_ltile_clb_0.mux_fle_2_in_3.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_2_in_3.LATCH_7_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XPHY_754 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_743 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_732 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_721 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xltile_clb_0.mux_fle_1_in_3.INVTX1_6_.scs8hd_inv_1 bottom_width_0_height_0__pin_6_
+ ltile_clb_0.mux_fle_1_in_3.INVTX1_6_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XFILLER_30_206 vgnd vpwr scs8hd_decap_4
XANTENNA__573__B _552_/X vgnd vpwr scs8hd_diode_2
XPHY_787 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_776 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_765 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_798 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_ltile_clb_0.mux_fle_3_in_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_3_in_0.LATCH_5_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_11_464 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_16_.scs8hd_inv_1_A
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_16_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_11_486 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_2_in_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_2_in_1.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_38_317 vgnd vpwr scs8hd_decap_8
XFILLER_38_328 vgnd vpwr scs8hd_decap_8
XFILLER_65_147 vgnd vpwr scs8hd_fill_1
XFILLER_48_80 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
+ _629_/Y vgnd vpwr scs8hd_diode_2
XFILLER_0_32 vgnd vpwr scs8hd_decap_12
XFILLER_80_117 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.mux_fle_3_in_2.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_3_in_2.INVTX1_3_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_3_in_2.LATCH_3_.latch/Q ltile_clb_0.mux_fle_3_in_2.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_0_87 vgnd vpwr scs8hd_decap_6
Xltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_3_.scs8hd_inv_1/Y
+ _628_/Y ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_61_364 vpwr vgnd scs8hd_fill_2
XFILLER_21_217 vpwr vgnd scs8hd_fill_2
XFILLER_9_74 vgnd vpwr scs8hd_decap_12
XFILLER_29_317 vgnd vpwr scs8hd_fill_1
XFILLER_37_361 vgnd vpwr scs8hd_decap_3
XFILLER_44_27 vgnd vpwr scs8hd_decap_4
XANTENNA__393__B _388_/B vgnd vpwr scs8hd_diode_2
XFILLER_40_515 vgnd vpwr scs8hd_fill_1
XFILLER_60_15 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mux_fle_0_in_0.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_0_in_0.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.buf4_0_.scs8hd_buf_1_A
+ ltile_clb_0.mux_fle_2_in_0.INVTX1_14_.scs8hd_inv_1/Y vgnd vpwr scs8hd_diode_2
XFILLER_4_449 vgnd vpwr scs8hd_decap_6
XFILLER_4_438 vgnd vpwr scs8hd_decap_4
XFILLER_4_427 vgnd vpwr scs8hd_decap_4
XFILLER_75_401 vpwr vgnd scs8hd_fill_2
XANTENNA__568__B _564_/B vgnd vpwr scs8hd_diode_2
XFILLER_75_489 vgnd vpwr scs8hd_decap_12
XFILLER_62_117 vgnd vpwr scs8hd_decap_12
XANTENNA__584__A _250_/X vgnd vpwr scs8hd_diode_2
XFILLER_28_394 vgnd vpwr scs8hd_decap_3
XFILLER_43_386 vpwr vgnd scs8hd_fill_2
XPHY_540 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_551 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_562 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_595 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_34_93 vgnd vpwr scs8hd_decap_12
XPHY_573 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_584 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_11_283 vpwr vgnd scs8hd_fill_2
XFILLER_11_261 vgnd vpwr scs8hd_decap_6
XFILLER_7_221 vgnd vpwr scs8hd_decap_4
XFILLER_11_294 vgnd vpwr scs8hd_fill_1
XFILLER_7_254 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.mux_fle_3_in_0.INVTX1_3_.scs8hd_inv_1 left_width_0_height_0__pin_3_ ltile_clb_0.mux_fle_3_in_0.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_78_250 vgnd vpwr scs8hd_decap_8
XFILLER_66_412 vpwr vgnd scs8hd_fill_2
XFILLER_78_294 vgnd vpwr scs8hd_fill_1
XFILLER_15_3 vgnd vpwr scs8hd_decap_12
XANTENNA__478__B _479_/B vgnd vpwr scs8hd_diode_2
XFILLER_81_437 vgnd vpwr scs8hd_fill_1
XFILLER_81_426 vgnd vpwr scs8hd_fill_1
XFILLER_19_361 vgnd vpwr scs8hd_decap_3
XFILLER_81_459 vgnd vpwr scs8hd_decap_12
XANTENNA__494__A _493_/X vgnd vpwr scs8hd_diode_2
XFILLER_34_386 vgnd vpwr scs8hd_decap_8
Xltile_clb_0.mux_fle_1_in_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_1_in_0.INVTX1_2_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_1_in_0.LATCH_2_.latch/Q ltile_clb_0.mux_fle_1_in_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_1_419 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_2_in_1.INVTX1_12_.scs8hd_inv_1_A top_width_0_height_0__pin_12_
+ vgnd vpwr scs8hd_diode_2
XFILLER_39_27 vgnd vpwr scs8hd_decap_12
XFILLER_57_412 vgnd vpwr scs8hd_decap_4
XANTENNA__388__B _388_/B vgnd vpwr scs8hd_diode_2
XFILLER_69_283 vpwr vgnd scs8hd_fill_2
XFILLER_69_272 vpwr vgnd scs8hd_fill_2
XFILLER_57_445 vpwr vgnd scs8hd_fill_2
XFILLER_57_423 vpwr vgnd scs8hd_fill_2
XFILLER_57_478 vgnd vpwr scs8hd_decap_4
XFILLER_57_456 vpwr vgnd scs8hd_fill_2
XFILLER_55_15 vgnd vpwr scs8hd_decap_12
XFILLER_29_147 vgnd vpwr scs8hd_decap_12
XFILLER_57_489 vgnd vpwr scs8hd_decap_12
XFILLER_55_59 vpwr vgnd scs8hd_fill_2
XFILLER_44_117 vgnd vpwr scs8hd_decap_12
XFILLER_25_320 vpwr vgnd scs8hd_fill_2
XFILLER_25_375 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_1_in_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_1_in_1.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_40_389 vpwr vgnd scs8hd_fill_2
XFILLER_4_202 vgnd vpwr scs8hd_decap_8
XFILLER_4_257 vpwr vgnd scs8hd_fill_2
XFILLER_0_430 vpwr vgnd scs8hd_fill_2
XANTENNA__579__A address[4] vgnd vpwr scs8hd_diode_2
XFILLER_48_401 vgnd vpwr scs8hd_decap_4
Xltile_clb_0.mux_fle_2_in_3.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_2_in_3.INVTX1_3_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_2_in_3.LATCH_3_.latch/Q ltile_clb_0.mux_fle_2_in_3.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_ltile_clb_0.mux_fle_2_in_2.INVTX1_8_.scs8hd_inv_1_A top_width_0_height_0__pin_8_
+ vgnd vpwr scs8hd_diode_2
XANTENNA__298__B _544_/A vgnd vpwr scs8hd_diode_2
XFILLER_0_485 vgnd vpwr scs8hd_decap_8
Xltile_clb_0.mux_fle_3_in_0.mux_l1_in_3_.TGATE_2_.scs8hd_ebufn_2 _652_/HI ltile_clb_0.mem_fle_3_in_0.LATCH_2_.latch/Q
+ ltile_clb_0.mux_fle_3_in_0.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XFILLER_75_242 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_0_in_3.mux_l1_in_2_.TGATE_3_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_0_in_3.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_75_297 vpwr vgnd scs8hd_fill_2
XFILLER_75_275 vgnd vpwr scs8hd_fill_1
XANTENNA_ltile_clb_0.mux_fle_1_in_0.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_1_in_0.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_28_191 vpwr vgnd scs8hd_fill_2
X_597_ _545_/A _580_/X _597_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_31_301 vpwr vgnd scs8hd_fill_2
XPHY_370 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_31_378 vpwr vgnd scs8hd_fill_2
XPHY_381 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_392 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xltile_clb_0.mux_fle_3_in_1.INVTX1_7_.scs8hd_inv_1 left_width_0_height_0__pin_7_ ltile_clb_0.mux_fle_3_in_1.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_ltile_clb_0.mux_fle_3_in_3.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_3_in_3.INVTX1_12_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__489__A _334_/A vgnd vpwr scs8hd_diode_2
XFILLER_39_423 vpwr vgnd scs8hd_fill_2
XFILLER_39_445 vpwr vgnd scs8hd_fill_2
XFILLER_66_297 vgnd vpwr scs8hd_fill_1
XFILLER_26_117 vgnd vpwr scs8hd_decap_12
XFILLER_81_245 vgnd vpwr scs8hd_decap_12
XFILLER_54_448 vgnd vpwr scs8hd_decap_4
XPHY_18 vgnd vpwr scs8hd_decap_3
XPHY_29 vgnd vpwr scs8hd_decap_3
XFILLER_81_289 vpwr vgnd scs8hd_fill_2
XFILLER_62_470 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_1_in_1.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_1_in_1.INVTX1_8_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_22_334 vpwr vgnd scs8hd_fill_2
XFILLER_22_356 vpwr vgnd scs8hd_fill_2
XFILLER_41_39 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mux_fle_3_in_3.INVTX1_5_.scs8hd_inv_1_A right_width_0_height_0__pin_5_
+ vgnd vpwr scs8hd_diode_2
XANTENNA__399__A _388_/A vgnd vpwr scs8hd_diode_2
XFILLER_49_209 vpwr vgnd scs8hd_fill_2
XFILLER_72_201 vpwr vgnd scs8hd_fill_2
X_520_ _328_/A _517_/X _520_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_72_267 vpwr vgnd scs8hd_fill_2
X_451_ _450_/X _451_/X vgnd vpwr scs8hd_buf_1
XFILLER_53_492 vpwr vgnd scs8hd_fill_2
X_382_ _381_/Y _427_/B vgnd vpwr scs8hd_buf_1
XFILLER_13_356 vgnd vpwr scs8hd_decap_8
XFILLER_13_367 vpwr vgnd scs8hd_fill_2
XFILLER_15_51 vgnd vpwr scs8hd_decap_8
XFILLER_15_62 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.buf4_0_.scs8hd_buf_1
+ ltile_clb_0.mux_fle_3_in_0.INVTX1_14_.scs8hd_inv_1/Y _604_/A vgnd vpwr scs8hd_buf_1
Xltile_clb_0.mux_fle_2_in_0.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_2_in_0.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2/Z
+ ltile_clb_0.mem_fle_2_in_0.LATCH_7_.latch/Q ltile_clb_0.mux_fle_2_in_0.INVTX1_14_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_56_80 vgnd vpwr scs8hd_decap_12
X_649_ _649_/HI _649_/LO vgnd vpwr scs8hd_conb_1
XFILLER_82_3 vgnd vpwr scs8hd_decap_12
XFILLER_31_175 vpwr vgnd scs8hd_fill_2
XFILLER_31_197 vgnd vpwr scs8hd_fill_1
XANTENNA_ltile_clb_0.mux_fle_0_in_0.INVTX1_11_.scs8hd_inv_1_A left_width_0_height_0__pin_11_
+ vgnd vpwr scs8hd_diode_2
XANTENNA__491__B _492_/B vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_0_in_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_0_in_1.INVTX1_2_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_0_in_1.LATCH_2_.latch/Q ltile_clb_0.mux_fle_0_in_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_ltile_clb_0.mux_fle_1_in_3.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_1_in_3.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__369__D _346_/D vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_2_in_2.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_2_in_2.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_54_234 vgnd vpwr scs8hd_fill_1
XFILLER_39_297 vpwr vgnd scs8hd_fill_2
XANTENNA__385__C _384_/X vgnd vpwr scs8hd_diode_2
XFILLER_54_267 vgnd vpwr scs8hd_decap_8
XFILLER_35_492 vpwr vgnd scs8hd_fill_2
XFILLER_52_27 vgnd vpwr scs8hd_decap_4
XFILLER_10_337 vpwr vgnd scs8hd_fill_2
XFILLER_50_495 vgnd vpwr scs8hd_fill_1
Xltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_11_.latch
+ data_in ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_11_.latch/Q
+ _586_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
Xltile_clb_0.mux_fle_2_in_1.mux_l1_in_3_.TGATE_2_.scs8hd_ebufn_2 _649_/HI ltile_clb_0.mem_fle_2_in_1.LATCH_2_.latch/Q
+ ltile_clb_0.mux_fle_2_in_1.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XANTENNA_ltile_clb_0.mux_fle_3_in_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_3_in_2.LATCH_4_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_77_359 vpwr vgnd scs8hd_fill_2
XFILLER_77_348 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__ff_0.DFFSRQ_0_.dff
+ clkbuf_1_1_0_clk/X ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.INVTX1_1_.scs8hd_inv_1/A
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.INVTX1_0_.scs8hd_inv_1/A
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__ff_0.DFFSRQ_0_.dff/QN
+ reset set vgnd vpwr scs8hd_dfbbp_1
XANTENNA__576__B _575_/B vgnd vpwr scs8hd_diode_2
XFILLER_45_245 vgnd vpwr scs8hd_decap_4
XFILLER_45_256 vpwr vgnd scs8hd_fill_2
X_503_ _343_/A _502_/B _503_/Y vgnd vpwr scs8hd_nor2_4
X_434_ _434_/A _429_/X _434_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_60_215 vgnd vpwr scs8hd_fill_1
XFILLER_26_470 vgnd vpwr scs8hd_decap_3
XANTENNA__592__A _540_/A vgnd vpwr scs8hd_diode_2
XFILLER_41_440 vpwr vgnd scs8hd_fill_2
X_365_ _392_/A _365_/B _365_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_41_484 vpwr vgnd scs8hd_fill_2
XFILLER_9_135 vgnd vpwr scs8hd_decap_12
X_296_ _282_/C _282_/B address[3] _258_/X _296_/X vgnd vpwr scs8hd_or4_4
XANTENNA_ltile_clb_0.mux_fle_1_in_2.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_1_in_2.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_42_93 vgnd vpwr scs8hd_decap_12
XFILLER_5_385 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_0_in_3.INVTX1_3_.scs8hd_inv_1_A left_width_0_height_0__pin_3_
+ vgnd vpwr scs8hd_diode_2
XFILLER_3_98 vgnd vpwr scs8hd_decap_12
XFILLER_76_392 vgnd vpwr scs8hd_decap_4
XANTENNA__486__B _484_/X vgnd vpwr scs8hd_diode_2
XFILLER_24_407 vpwr vgnd scs8hd_fill_2
XFILLER_51_204 vpwr vgnd scs8hd_fill_2
XFILLER_8_190 vgnd vpwr scs8hd_decap_6
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_0_.latch_SLEEPB
+ _546_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_4_.TGATE_1_.scs8hd_ebufn_2_TEB
+ _628_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_0_in_2.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_0_in_2.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_59_348 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.mem_ble4_out_0.LATCH_0_.latch_D
+ data_in vgnd vpwr scs8hd_diode_2
XFILLER_47_27 vgnd vpwr scs8hd_decap_12
XANTENNA__396__B _427_/B vgnd vpwr scs8hd_diode_2
XFILLER_63_15 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_7_.TGATE_0_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_14_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_15_418 vgnd vpwr scs8hd_decap_3
XFILLER_27_245 vpwr vgnd scs8hd_fill_2
XFILLER_82_373 vgnd vpwr scs8hd_decap_12
XFILLER_42_215 vgnd vpwr scs8hd_decap_6
XFILLER_63_59 vpwr vgnd scs8hd_fill_2
XFILLER_23_484 vgnd vpwr scs8hd_fill_1
XFILLER_6_105 vgnd vpwr scs8hd_decap_12
XFILLER_10_178 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_11_.scs8hd_inv_1_A
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_11_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_77_123 vgnd vpwr scs8hd_decap_12
XANTENNA__587__A _535_/A vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_1_in_1.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_1_in_1.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2/A
+ ltile_clb_0.mem_fle_1_in_1.LATCH_7_.latch/Q ltile_clb_0.mux_fle_1_in_1.INVTX1_14_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_58_392 vgnd vpwr scs8hd_decap_4
XFILLER_58_381 vpwr vgnd scs8hd_fill_2
XFILLER_18_267 vgnd vpwr scs8hd_decap_3
XFILLER_33_248 vpwr vgnd scs8hd_fill_2
XFILLER_14_473 vgnd vpwr scs8hd_decap_12
X_417_ _331_/A _433_/A vgnd vpwr scs8hd_buf_1
X_348_ _355_/B _353_/B vgnd vpwr scs8hd_buf_1
X_279_ _278_/X _313_/A _279_/X vgnd vpwr scs8hd_or2_4
XANTENNA_ltile_clb_0.mux_fle_2_in_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_2_in_0.LATCH_6_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_5_171 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_3_.TGATE_1_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_3_.TGATE_1_.scs8hd_ebufn_2/A
+ _614_/Y ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_1_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_45_3 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_7_.scs8hd_inv_1
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_7_.latch/Q
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA__497__A _325_/A vgnd vpwr scs8hd_diode_2
XFILLER_49_392 vgnd vpwr scs8hd_decap_3
XFILLER_24_215 vgnd vpwr scs8hd_fill_1
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_20_443 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.mux_fle_1_in_2.mux_l1_in_3_.TGATE_2_.scs8hd_ebufn_2 _646_/HI ltile_clb_0.mem_fle_1_in_2.LATCH_2_.latch/Q
+ ltile_clb_0.mux_fle_1_in_2.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
Xltile_clb_0.mux_fle_3_in_2.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_3_in_2.INVTX1_9_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_3_in_2.LATCH_1_.latch/Q ltile_clb_0.mux_fle_3_in_2.mux_l1_in_2_.TGATE_3_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_8_.scs8hd_inv_1_A
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_8_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_58_15 vgnd vpwr scs8hd_decap_12
XFILLER_59_123 vgnd vpwr scs8hd_decap_6
XFILLER_55_362 vpwr vgnd scs8hd_fill_2
XPHY_711 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_700 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_744 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_70_387 vgnd vpwr scs8hd_decap_6
XFILLER_70_376 vpwr vgnd scs8hd_fill_2
XPHY_733 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_722 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_777 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_766 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_755 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_70_398 vpwr vgnd scs8hd_fill_2
XFILLER_23_270 vpwr vgnd scs8hd_fill_2
XPHY_799 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_788 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_23_51 vgnd vpwr scs8hd_decap_8
XFILLER_23_62 vgnd vpwr scs8hd_decap_12
XFILLER_11_498 vgnd vpwr scs8hd_decap_3
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_13_.latch_D
+ data_in vgnd vpwr scs8hd_diode_2
XFILLER_7_447 vgnd vpwr scs8hd_decap_4
XANTENNA_ltile_clb_0.mux_fle_1_in_2.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_1_in_2.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_78_410 vgnd vpwr scs8hd_decap_4
XFILLER_2_141 vgnd vpwr scs8hd_decap_12
XFILLER_78_443 vgnd vpwr scs8hd_decap_4
Xltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_7_.TGATE_0_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_14_.scs8hd_inv_1/Y
+ _629_/Y ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_7_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_0_44 vgnd vpwr scs8hd_decap_12
XFILLER_80_129 vgnd vpwr scs8hd_decap_12
XFILLER_34_513 vgnd vpwr scs8hd_decap_3
XFILLER_46_373 vpwr vgnd scs8hd_fill_2
XFILLER_46_384 vpwr vgnd scs8hd_fill_2
XFILLER_64_80 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.mux_fle_1_in_0.INVTX1_2_.scs8hd_inv_1 bottom_width_0_height_0__pin_2_
+ ltile_clb_0.mux_fle_1_in_0.INVTX1_2_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB
+ _606_/Y vgnd vpwr scs8hd_diode_2
XFILLER_9_86 vgnd vpwr scs8hd_decap_12
XFILLER_6_491 vgnd vpwr scs8hd_decap_12
XFILLER_69_443 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_0_in_2.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_0_in_2.INVTX1_8_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_69_465 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l4_in_0_.TGATE_1_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l4_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ _610_/Y ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_16_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_64_170 vpwr vgnd scs8hd_fill_2
XFILLER_37_384 vgnd vpwr scs8hd_fill_1
XFILLER_52_387 vgnd vpwr scs8hd_fill_1
XFILLER_52_376 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_3_in_0.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_3_in_0.INVTX1_8_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_60_27 vgnd vpwr scs8hd_decap_4
XFILLER_20_240 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.mux_fle_0_in_2.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_0_in_2.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2/Z
+ ltile_clb_0.mem_fle_0_in_2.LATCH_7_.latch/Q ltile_clb_0.mux_fle_0_in_2.INVTX1_14_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_ltile_clb_0.mux_fle_1_in_3.INVTX1_9_.scs8hd_inv_1_A right_width_0_height_0__pin_9_
+ vgnd vpwr scs8hd_diode_2
XFILLER_62_129 vgnd vpwr scs8hd_decap_6
XANTENNA__584__B _585_/B vgnd vpwr scs8hd_diode_2
XFILLER_31_505 vgnd vpwr scs8hd_decap_8
XFILLER_70_184 vgnd vpwr scs8hd_decap_8
XANTENNA_ltile_clb_0.mux_fle_2_in_0.INVTX1_5_.scs8hd_inv_1_A right_width_0_height_0__pin_5_
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_1_in_0.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_1_in_0.INVTX1_8_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_1_in_0.LATCH_0_.latch/Q ltile_clb_0.mux_fle_1_in_0.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_5_.latch_SLEEPB
+ _593_/Y vgnd vpwr scs8hd_diode_2
XFILLER_43_398 vpwr vgnd scs8hd_fill_2
XPHY_530 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_541 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_552 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_596 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_585 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_11_240 vpwr vgnd scs8hd_fill_2
XPHY_563 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_574 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_7_211 vgnd vpwr scs8hd_decap_4
XFILLER_7_299 vpwr vgnd scs8hd_fill_2
XFILLER_7_288 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_0_in_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_0_in_1.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_50_93 vgnd vpwr scs8hd_decap_12
XFILLER_3_472 vpwr vgnd scs8hd_fill_2
XFILLER_3_483 vpwr vgnd scs8hd_fill_2
XFILLER_78_284 vgnd vpwr scs8hd_decap_4
Xltile_clb_0.mux_fle_1_in_1.INVTX1_6_.scs8hd_inv_1 bottom_width_0_height_0__pin_6_
+ ltile_clb_0.mux_fle_1_in_1.INVTX1_6_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_7_.TGATE_0_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_14_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_61_140 vpwr vgnd scs8hd_fill_2
XFILLER_61_184 vgnd vpwr scs8hd_fill_1
XANTENNA_ltile_clb_0.mux_fle_0_in_0.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_0_in_0.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_0_in_3.mux_l1_in_3_.TGATE_2_.scs8hd_ebufn_2 _643_/HI ltile_clb_0.mem_fle_0_in_3.LATCH_2_.latch/Q
+ ltile_clb_0.mux_fle_0_in_3.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
Xltile_clb_0.mux_fle_2_in_3.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_2_in_3.INVTX1_9_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_2_in_3.LATCH_1_.latch/Q ltile_clb_0.mux_fle_2_in_3.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_ltile_clb_0.mux_fle_1_in_3.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_1_in_3.mux_l1_in_2_.TGATE_3_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_39_39 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mux_fle_3_in_1.INVTX1_2_.scs8hd_inv_1_A bottom_width_0_height_0__pin_2_
+ vgnd vpwr scs8hd_diode_2
XFILLER_69_240 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l4_in_0_.TGATE_1_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_57_468 vgnd vpwr scs8hd_decap_3
XFILLER_29_159 vgnd vpwr scs8hd_decap_12
XFILLER_72_416 vgnd vpwr scs8hd_decap_4
XFILLER_55_27 vgnd vpwr scs8hd_decap_12
XFILLER_44_129 vgnd vpwr scs8hd_decap_12
XFILLER_80_471 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
+ _624_/Y vgnd vpwr scs8hd_diode_2
XFILLER_25_354 vgnd vpwr scs8hd_fill_1
XFILLER_71_15 vgnd vpwr scs8hd_decap_12
XFILLER_40_313 vgnd vpwr scs8hd_fill_1
XFILLER_71_59 vpwr vgnd scs8hd_fill_2
XFILLER_40_346 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_2_in_3.INVTX1_10_.scs8hd_inv_1_A bottom_width_0_height_0__pin_10_
+ vgnd vpwr scs8hd_diode_2
XFILLER_4_236 vgnd vpwr scs8hd_decap_8
XANTENNA__579__B _578_/X vgnd vpwr scs8hd_diode_2
XFILLER_75_221 vpwr vgnd scs8hd_fill_2
XFILLER_0_497 vgnd vpwr scs8hd_decap_12
XFILLER_75_254 vpwr vgnd scs8hd_fill_2
XFILLER_48_457 vgnd vpwr scs8hd_fill_1
XFILLER_63_416 vpwr vgnd scs8hd_fill_2
XANTENNA__595__A _569_/A vgnd vpwr scs8hd_diode_2
XFILLER_48_479 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.mux_fle_2_in_2.INVTX1_1_.scs8hd_inv_1 right_width_0_height_0__pin_1_
+ ltile_clb_0.mux_fle_2_in_2.INVTX1_1_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XANTENNA_ltile_clb_0.mux_fle_0_in_3.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_0_in_3.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
X_596_ _544_/A _580_/X _596_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_16_343 vpwr vgnd scs8hd_fill_2
XFILLER_16_398 vpwr vgnd scs8hd_fill_2
XFILLER_43_195 vpwr vgnd scs8hd_fill_2
XPHY_360 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XPHY_371 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_382 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_393 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_6_32 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mux_fle_3_in_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_3_in_1.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_0_.scs8hd_inv_1
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_0_.latch/Q
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_3_291 vgnd vpwr scs8hd_fill_1
XFILLER_39_402 vpwr vgnd scs8hd_fill_2
XANTENNA__489__B _484_/X vgnd vpwr scs8hd_diode_2
XPHY_19 vgnd vpwr scs8hd_decap_3
XFILLER_26_129 vgnd vpwr scs8hd_decap_12
XFILLER_81_257 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_0_.TGATE_1_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ _632_/Y ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l4_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_22_313 vgnd vpwr scs8hd_decap_4
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_3_.TGATE_0_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_6_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_4_.TGATE_0_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_8_.scs8hd_inv_1/Y
+ _605_/Y ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_2_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_1_217 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mem_fle_3_in_3.LATCH_4_.latch_SLEEPB _332_/Y vgnd vpwr scs8hd_diode_2
XANTENNA__399__B _399_/B vgnd vpwr scs8hd_diode_2
XFILLER_66_15 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mux_fle_0_in_3.mux_l1_in_3_.TGATE_2_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_0_in_3.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_72_213 vgnd vpwr scs8hd_fill_1
XFILLER_57_287 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_1_in_0.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_1_in_0.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_45_416 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.mux_fle_0_in_1.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_0_in_1.INVTX1_8_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_0_in_1.LATCH_0_.latch/Q ltile_clb_0.mux_fle_0_in_1.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_38_490 vgnd vpwr scs8hd_decap_12
XFILLER_72_279 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mem_fle_0_in_0.LATCH_3_.latch_D data_in vgnd vpwr scs8hd_diode_2
X_450_ _449_/X _450_/X vgnd vpwr scs8hd_buf_1
X_381_ _226_/X _381_/Y vgnd vpwr scs8hd_inv_8
XFILLER_9_306 vgnd vpwr scs8hd_decap_3
XFILLER_15_74 vgnd vpwr scs8hd_decap_12
XFILLER_9_339 vpwr vgnd scs8hd_fill_2
XFILLER_40_154 vgnd vpwr scs8hd_decap_6
XFILLER_5_501 vgnd vpwr scs8hd_decap_12
XFILLER_31_51 vgnd vpwr scs8hd_decap_8
XFILLER_31_62 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mem_fle_0_in_1.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_2_in_3.INVTX1_5_.scs8hd_inv_1 right_width_0_height_0__pin_5_
+ ltile_clb_0.mux_fle_2_in_3.INVTX1_5_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XFILLER_0_283 vgnd vpwr scs8hd_decap_4
XFILLER_48_265 vgnd vpwr scs8hd_decap_3
XANTENNA_ltile_clb_0.mux_fle_2_in_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_2_in_2.LATCH_5_.latch/Q
+ vgnd vpwr scs8hd_diode_2
X_648_ _648_/HI _648_/LO vgnd vpwr scs8hd_conb_1
XFILLER_31_110 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mux_fle_0_in_1.INVTX1_0_.scs8hd_inv_1_A top_width_0_height_0__pin_0_
+ vgnd vpwr scs8hd_diode_2
XFILLER_44_482 vpwr vgnd scs8hd_fill_2
XFILLER_44_493 vpwr vgnd scs8hd_fill_2
XFILLER_72_80 vgnd vpwr scs8hd_decap_12
X_579_ address[4] _578_/X _579_/X vgnd vpwr scs8hd_or2_4
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB
+ _620_/Y vgnd vpwr scs8hd_diode_2
Xltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_15_.latch
+ data_in ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_15_.latch/Q
+ _556_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_75_3 vgnd vpwr scs8hd_decap_12
XPHY_190 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xltile_clb_0.mux_fle_2_in_0.INVTX1_11_.scs8hd_inv_1 left_width_0_height_0__pin_11_
+ ltile_clb_0.mux_fle_2_in_0.INVTX1_11_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XFILLER_8_383 vpwr vgnd scs8hd_fill_2
XFILLER_39_210 vpwr vgnd scs8hd_fill_2
XFILLER_39_221 vpwr vgnd scs8hd_fill_2
XFILLER_39_232 vpwr vgnd scs8hd_fill_2
XFILLER_39_243 vgnd vpwr scs8hd_fill_1
XFILLER_54_224 vpwr vgnd scs8hd_fill_2
XANTENNA__385__D _358_/D vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_1_in_2.INVTX1_14_.scs8hd_inv_1_A ltile_clb_0.mux_fle_1_in_2.INVTX1_14_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_62_290 vgnd vpwr scs8hd_decap_6
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_3_.latch_D
+ data_in vgnd vpwr scs8hd_diode_2
XFILLER_22_154 vgnd vpwr scs8hd_decap_12
XFILLER_50_474 vpwr vgnd scs8hd_fill_2
XFILLER_6_309 vgnd vpwr scs8hd_decap_8
Xltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_1_.scs8hd_inv_1/Y
+ _612_/Y ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_10_.latch_D
+ data_in vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_2_in_1.INVTX1_13_.scs8hd_inv_1 right_width_0_height_0__pin_13_
+ ltile_clb_0.mux_fle_2_in_1.INVTX1_13_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_2_.scs8hd_inv_1_A
+ ltile_clb_0.mux_fle_2_in_2.INVTX1_14_.scs8hd_inv_1/Y vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mux_fle_3_in_1.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_3_in_1.INVTX1_3_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_3_in_1.LATCH_3_.latch/Q ltile_clb_0.mux_fle_3_in_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_18_438 vgnd vpwr scs8hd_decap_8
XFILLER_18_449 vpwr vgnd scs8hd_fill_2
XFILLER_33_419 vpwr vgnd scs8hd_fill_2
X_502_ _423_/A _502_/B _502_/Y vgnd vpwr scs8hd_nor2_4
X_433_ _433_/A _429_/X _433_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_60_227 vpwr vgnd scs8hd_fill_2
XFILLER_13_110 vgnd vpwr scs8hd_decap_12
XANTENNA__592__B _588_/X vgnd vpwr scs8hd_diode_2
XFILLER_26_493 vgnd vpwr scs8hd_decap_8
XFILLER_13_176 vpwr vgnd scs8hd_fill_2
XFILLER_41_463 vpwr vgnd scs8hd_fill_2
X_364_ _391_/A _365_/B _364_/Y vgnd vpwr scs8hd_nor2_4
X_295_ _304_/A _569_/A _295_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_9_147 vgnd vpwr scs8hd_decap_12
XFILLER_5_364 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mem_fle_1_in_3.LATCH_5_.latch_SLEEPB _443_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l4_in_0_.TGATE_1_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l4_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_17_482 vpwr vgnd scs8hd_fill_2
XFILLER_24_419 vpwr vgnd scs8hd_fill_2
XFILLER_36_279 vpwr vgnd scs8hd_fill_2
XFILLER_32_430 vgnd vpwr scs8hd_decap_6
XFILLER_44_290 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_11_.scs8hd_inv_1_A
+ ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_11_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_1_in_0.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_1_in_0.LATCH_7_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_74_308 vgnd vpwr scs8hd_decap_8
XFILLER_67_360 vgnd vpwr scs8hd_decap_4
XANTENNA_ltile_clb_0.mux_fle_2_in_1.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_2_in_1.INVTX1_8_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_47_39 vgnd vpwr scs8hd_decap_12
XANTENNA__396__C _384_/X vgnd vpwr scs8hd_diode_2
XFILLER_82_385 vgnd vpwr scs8hd_decap_12
XFILLER_63_27 vgnd vpwr scs8hd_decap_12
XFILLER_23_452 vgnd vpwr scs8hd_fill_1
XFILLER_50_260 vgnd vpwr scs8hd_decap_12
XFILLER_6_117 vgnd vpwr scs8hd_decap_12
XFILLER_5_3 vgnd vpwr scs8hd_decap_12
XFILLER_2_345 vgnd vpwr scs8hd_decap_3
XFILLER_2_378 vpwr vgnd scs8hd_fill_2
XFILLER_2_389 vpwr vgnd scs8hd_fill_2
XFILLER_77_135 vgnd vpwr scs8hd_decap_12
XFILLER_65_319 vpwr vgnd scs8hd_fill_2
XFILLER_58_360 vgnd vpwr scs8hd_decap_4
XANTENNA__587__B _585_/B vgnd vpwr scs8hd_diode_2
XFILLER_46_500 vgnd vpwr scs8hd_decap_12
XFILLER_18_213 vgnd vpwr scs8hd_fill_1
XFILLER_18_224 vgnd vpwr scs8hd_decap_4
XANTENNA_ltile_clb_0.mux_fle_0_in_3.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_0_in_3.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_18_246 vgnd vpwr scs8hd_decap_6
XANTENNA_ltile_clb_0.mem_fle_2_in_2.LATCH_5_.latch_SLEEPB _401_/Y vgnd vpwr scs8hd_diode_2
XFILLER_61_514 vpwr vgnd scs8hd_fill_2
X_416_ _432_/A _412_/B _416_/Y vgnd vpwr scs8hd_nor2_4
X_347_ _347_/A _355_/B vgnd vpwr scs8hd_buf_1
XFILLER_14_485 vpwr vgnd scs8hd_fill_2
XFILLER_14_496 vgnd vpwr scs8hd_decap_8
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_3_.TGATE_0_.scs8hd_ebufn_2_A
+ ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_6_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
X_278_ address[3] _278_/X vgnd vpwr scs8hd_buf_1
XANTENNA_ltile_clb_0.mem_fle_0_in_3.LATCH_7_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_0_in_2.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_0_in_2.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_5_.TGATE_0_.scs8hd_ebufn_2_TEB
+ _629_/Y vgnd vpwr scs8hd_diode_2
XFILLER_38_3 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mux_fle_3_in_3.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_3_in_3.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__497__B _495_/X vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_0_in_0.INVTX1_9_.scs8hd_inv_1_A right_width_0_height_0__pin_9_
+ vgnd vpwr scs8hd_diode_2
XFILLER_49_371 vpwr vgnd scs8hd_fill_2
XFILLER_64_341 vpwr vgnd scs8hd_fill_2
XFILLER_20_488 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_3_in_2.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_3_in_2.mux_l1_in_2_.TGATE_3_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_58_27 vgnd vpwr scs8hd_decap_4
Xltile_clb_0.mux_fle_2_in_2.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_2_in_2.INVTX1_3_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_2_in_2.LATCH_3_.latch/Q ltile_clb_0.mux_fle_2_in_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_74_105 vgnd vpwr scs8hd_decap_12
XFILLER_59_179 vpwr vgnd scs8hd_fill_2
XFILLER_59_168 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_0_.latch
+ data_in ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_0_.latch/Q
+ _304_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_ltile_clb_0.mem_fle_1_in_1.LATCH_7_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_74_15 vgnd vpwr scs8hd_decap_12
XFILLER_55_330 vpwr vgnd scs8hd_fill_2
XFILLER_15_216 vpwr vgnd scs8hd_fill_2
XFILLER_43_503 vpwr vgnd scs8hd_fill_2
XPHY_701 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_1_.TGATE_0_.scs8hd_ebufn_2
+ ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_1_.TGATE_0_.scs8hd_ebufn_2/A
+ _623_/Y ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XPHY_745 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_734 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_723 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_712 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_778 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_767 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_756 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_11_400 vpwr vgnd scs8hd_fill_2
XPHY_789 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_7_415 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_1_in_1.INVTX1_6_.scs8hd_inv_1_A bottom_width_0_height_0__pin_6_
+ vgnd vpwr scs8hd_diode_2
XFILLER_11_477 vgnd vpwr scs8hd_decap_3
XFILLER_23_74 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mem_fle_1_in_2.LATCH_5_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mem_fle_3_in_1.LATCH_5_.latch_SLEEPB _363_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_3_in_1.INVTX1_12_.scs8hd_inv_1_A top_width_0_height_0__pin_12_
+ vgnd vpwr scs8hd_diode_2
XANTENNA__598__A _546_/A vgnd vpwr scs8hd_diode_2
XFILLER_48_93 vgnd vpwr scs8hd_decap_12
XFILLER_58_190 vgnd vpwr scs8hd_decap_6
XFILLER_46_352 vgnd vpwr scs8hd_decap_4
XANTENNA_ltile_clb_0.mem_fle_1_in_3.LATCH_3_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_0_56 vgnd vpwr scs8hd_decap_6
XFILLER_73_182 vgnd vpwr scs8hd_fill_1
XFILLER_61_322 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_2_in_2.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_2_in_2.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.mem_ble4_out_0.LATCH_0_.latch_D
+ data_in vgnd vpwr scs8hd_diode_2
XFILLER_46_396 vgnd vpwr scs8hd_fill_1
Xltile_clb_0.mux_fle_1_in_3.INVTX1_11_.scs8hd_inv_1 left_width_0_height_0__pin_11_
+ ltile_clb_0.mux_fle_1_in_3.INVTX1_11_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
XFILLER_61_399 vgnd vpwr scs8hd_decap_4
XFILLER_80_80 vgnd vpwr scs8hd_decap_12
XFILLER_9_98 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_2_.scs8hd_inv_1
+ ltile_clb_0.mux_fle_3_in_2.INVTX1_14_.scs8hd_inv_1/Y _609_/A vgnd vpwr scs8hd_inv_1
XANTENNA_ltile_clb_0.mux_fle_0_in_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_0_in_0.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mem_fle_2_in_0.LATCH_5_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_69_477 vgnd vpwr scs8hd_decap_8
XANTENNA_ltile_clb_0.mux_fle_2_in_2.INVTX1_3_.scs8hd_inv_1_A left_width_0_height_0__pin_3_
+ vgnd vpwr scs8hd_diode_2
XANTENNA__301__A _304_/A vgnd vpwr scs8hd_diode_2
XFILLER_56_105 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mem_fle_0_in_2.LATCH_6_.latch_SLEEPB _497_/Y vgnd vpwr scs8hd_diode_2
XFILLER_37_330 vgnd vpwr scs8hd_decap_3
XFILLER_25_503 vgnd vpwr scs8hd_decap_12
XFILLER_64_193 vgnd vpwr scs8hd_decap_4
XFILLER_52_333 vgnd vpwr scs8hd_decap_3
XFILLER_52_322 vgnd vpwr scs8hd_fill_1
XFILLER_52_355 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_9_.latch_D
+ data_in vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mem_fle_2_in_1.LATCH_3_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_20_252 vgnd vpwr scs8hd_fill_1
XFILLER_20_285 vgnd vpwr scs8hd_decap_3
XFILLER_69_15 vgnd vpwr scs8hd_decap_12
XFILLER_79_208 vgnd vpwr scs8hd_decap_12
XFILLER_69_59 vpwr vgnd scs8hd_fill_2
XFILLER_75_436 vgnd vpwr scs8hd_decap_3
XFILLER_75_414 vgnd vpwr scs8hd_decap_8
XFILLER_75_469 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mem_fle_2_in_2.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_47_138 vpwr vgnd scs8hd_fill_2
XFILLER_28_352 vgnd vpwr scs8hd_decap_4
XFILLER_70_141 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_3_.TGATE_0_.scs8hd_ebufn_2_TEB
+ _607_/Y vgnd vpwr scs8hd_diode_2
XPHY_520 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_531 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_542 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_553 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_ltile_clb_0.mux_fle_3_in_3.INVTX1_0_.scs8hd_inv_1_A top_width_0_height_0__pin_0_
+ vgnd vpwr scs8hd_diode_2
XPHY_586 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_564 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_575 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_597 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xltile_clb_0.mux_fle_0_in_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_0_in_0.INVTX1_2_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_0_in_0.LATCH_2_.latch/Q ltile_clb_0.mux_fle_0_in_0.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
Xltile_clb_0.mux_fle_0_in_2.INVTX1_0_.scs8hd_inv_1 top_width_0_height_0__pin_0_ ltile_clb_0.mux_fle_0_in_2.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_3_451 vpwr vgnd scs8hd_fill_2
XFILLER_66_436 vpwr vgnd scs8hd_fill_2
XFILLER_38_105 vgnd vpwr scs8hd_decap_12
XFILLER_19_330 vgnd vpwr scs8hd_decap_6
XFILLER_38_149 vgnd vpwr scs8hd_decap_4
XFILLER_81_428 vgnd vpwr scs8hd_decap_3
XFILLER_34_300 vpwr vgnd scs8hd_fill_2
XFILLER_74_480 vgnd vpwr scs8hd_decap_12
XFILLER_34_333 vgnd vpwr scs8hd_fill_1
XFILLER_46_182 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_13_.latch
+ data_in ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_13_.latch/Q
+ _251_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_ltile_clb_0.mem_fle_3_in_0.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_61_163 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mem_fle_1_in_1.LATCH_6_.latch_SLEEPB _464_/Y vgnd vpwr scs8hd_diode_2
Xltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_0_.latch
+ data_in ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_0_.latch/Q
+ _598_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
Xltile_clb_0.mem_fle_0_in_0.LATCH_6_.latch data_in ltile_clb_0.mem_fle_0_in_0.LATCH_6_.latch/Q
+ _519_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
Xltile_clb_0.mux_fle_1_in_3.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_1_in_3.INVTX1_3_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_1_in_3.LATCH_3_.latch/Q ltile_clb_0.mux_fle_1_in_3.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
Xltile_clb_0.mux_fle_2_in_0.mux_l1_in_3_.TGATE_2_.scs8hd_ebufn_2 _648_/HI ltile_clb_0.mem_fle_2_in_0.LATCH_2_.latch/Q
+ ltile_clb_0.mux_fle_2_in_0.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XFILLER_69_252 vpwr vgnd scs8hd_fill_2
XFILLER_69_296 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_0_in_0.mux_l1_in_2_.TGATE_3_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_0_in_0.INVTX1_11_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_55_39 vgnd vpwr scs8hd_decap_12
Xltile_clb_0.mem_fle_1_in_0.LATCH_5_.latch data_in ltile_clb_0.mem_fle_1_in_0.LATCH_5_.latch/Q
+ _476_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_65_480 vgnd vpwr scs8hd_decap_8
Xltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_3_.scs8hd_inv_1
+ ltile_clb_0.mux_fle_1_in_3.INVTX1_14_.scs8hd_inv_1/Y _627_/A vgnd vpwr scs8hd_inv_1
XFILLER_25_333 vpwr vgnd scs8hd_fill_2
XFILLER_37_193 vpwr vgnd scs8hd_fill_2
XFILLER_80_450 vgnd vpwr scs8hd_decap_8
XFILLER_13_506 vgnd vpwr scs8hd_decap_8
XFILLER_80_483 vgnd vpwr scs8hd_decap_12
XFILLER_71_27 vgnd vpwr scs8hd_decap_12
XFILLER_40_358 vgnd vpwr scs8hd_fill_1
XANTENNA_ltile_clb_0.mux_fle_1_in_0.INVTX1_11_.scs8hd_inv_1_A left_width_0_height_0__pin_11_
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_0.mem_fle_2_in_0.LATCH_4_.latch data_in ltile_clb_0.mem_fle_2_in_0.LATCH_4_.latch/Q
+ _433_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_4_215 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_5_.latch_D
+ data_in vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_0_in_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_0_in_1.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_0_421 vpwr vgnd scs8hd_fill_2
XFILLER_0_454 vgnd vpwr scs8hd_decap_4
XANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
+ _612_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_8_.latch_SLEEPB
+ _538_/Y vgnd vpwr scs8hd_diode_2
XFILLER_29_51 vgnd vpwr scs8hd_decap_8
XFILLER_29_62 vgnd vpwr scs8hd_decap_12
XFILLER_48_436 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.mem_fle_3_in_0.LATCH_3_.latch data_in ltile_clb_0.mem_fle_3_in_0.LATCH_3_.latch/Q
+ _376_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_63_428 vpwr vgnd scs8hd_fill_2
XANTENNA__595__B _580_/X vgnd vpwr scs8hd_diode_2
XFILLER_16_333 vgnd vpwr scs8hd_decap_3
XFILLER_71_461 vgnd vpwr scs8hd_decap_12
X_595_ _569_/A _580_/X _595_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_16_366 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_0.mux_fle_0_in_0.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_0_in_0.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_16_377 vgnd vpwr scs8hd_decap_8
XFILLER_16_388 vgnd vpwr scs8hd_decap_4
XFILLER_31_325 vgnd vpwr scs8hd_decap_4
XPHY_350 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_361 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_31_358 vgnd vpwr scs8hd_decap_4
Xltile_clb_0.mux_fle_0_in_3.INVTX1_4_.scs8hd_inv_1 top_width_0_height_0__pin_4_ ltile_clb_0.mux_fle_0_in_3.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XPHY_372 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_383 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_394 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_ltile_clb_0.mux_fle_3_in_1.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_3_in_1.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_6_44 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mux_fle_0_in_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_0_in_0.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_20_3 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mem_fle_2_in_0.LATCH_6_.latch_SLEEPB _431_/Y vgnd vpwr scs8hd_diode_2
XFILLER_19_182 vgnd vpwr scs8hd_fill_1
XFILLER_81_269 vgnd vpwr scs8hd_decap_12
XFILLER_34_141 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.mux_fle_1_in_2.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB ltile_clb_0.mem_fle_1_in_2.LATCH_6_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_0.mux_fle_1_in_2.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A ltile_clb_0.mux_fle_1_in_2.INVTX1_8_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_66_27 vgnd vpwr scs8hd_decap_4
XFILLER_57_200 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.mux_fle_1_in_0.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_1_in_0.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2/Z
+ ltile_clb_0.mem_fle_1_in_0.LATCH_7_.latch/Q ltile_clb_0.mux_fle_1_in_0.INVTX1_14_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
Xltile_clb_0.mem_fle_2_in_2.LATCH_7_.latch data_in ltile_clb_0.mem_fle_2_in_2.LATCH_7_.latch/Q
+ _399_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_57_299 vgnd vpwr scs8hd_decap_4
XFILLER_45_439 vpwr vgnd scs8hd_fill_2
XFILLER_82_15 vgnd vpwr scs8hd_decap_12
X_380_ _380_/A _380_/X vgnd vpwr scs8hd_buf_1
XFILLER_53_483 vpwr vgnd scs8hd_fill_2
XFILLER_9_318 vpwr vgnd scs8hd_fill_2
XFILLER_15_86 vgnd vpwr scs8hd_decap_12
XFILLER_21_380 vpwr vgnd scs8hd_fill_2
XFILLER_40_188 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.mem_fle_3_in_2.LATCH_6_.latch data_in ltile_clb_0.mem_fle_3_in_2.LATCH_6_.latch/Q
+ _350_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_5_513 vgnd vpwr scs8hd_decap_3
XFILLER_31_74 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_1_.latch_D
+ data_in vgnd vpwr scs8hd_diode_2
XFILLER_48_222 vgnd vpwr scs8hd_decap_3
XANTENNA_ltile_clb_0.mux_fle_3_in_2.INVTX1_9_.scs8hd_inv_1_A right_width_0_height_0__pin_9_
+ vgnd vpwr scs8hd_diode_2
XFILLER_63_236 vpwr vgnd scs8hd_fill_2
XFILLER_63_225 vgnd vpwr scs8hd_decap_4
XFILLER_56_93 vgnd vpwr scs8hd_decap_12
XFILLER_36_428 vgnd vpwr scs8hd_decap_4
XFILLER_63_258 vgnd vpwr scs8hd_decap_4
XFILLER_16_141 vgnd vpwr scs8hd_decap_12
XFILLER_44_450 vgnd vpwr scs8hd_decap_8
X_647_ _647_/HI _647_/LO vgnd vpwr scs8hd_conb_1
X_578_ address[6] address[7] _227_/X _526_/D _578_/X vgnd vpwr scs8hd_or4_4
Xltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_0_.latch
+ data_in ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_0_.latch/Q
+ _572_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_15_.latch_SLEEPB
+ _530_/Y vgnd vpwr scs8hd_diode_2
XPHY_180 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_191 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_68_3 vgnd vpwr scs8hd_decap_12
XFILLER_8_395 vpwr vgnd scs8hd_fill_2
Xltile_clb_0.mux_fle_1_in_1.mux_l1_in_3_.TGATE_2_.scs8hd_ebufn_2 _645_/HI ltile_clb_0.mem_fle_1_in_1.LATCH_2_.latch/Q
+ ltile_clb_0.mux_fle_1_in_1.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2/A vgnd vpwr scs8hd_ebufn_2
Xltile_clb_0.mux_fle_3_in_1.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2 ltile_clb_0.mux_fle_3_in_1.INVTX1_9_.scs8hd_inv_1/Y
+ ltile_clb_0.mem_fle_3_in_1.LATCH_1_.latch/Q ltile_clb_0.mux_fle_3_in_1.mux_l1_in_2_.TGATE_3_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
Xltile_clb_0.mux_fle_2_in_0.INVTX1_1_.scs8hd_inv_1 right_width_0_height_0__pin_1_
+ ltile_clb_0.mux_fle_2_in_0.INVTX1_1_.scs8hd_inv_1/Y vgnd vpwr scs8hd_inv_1
.ends

