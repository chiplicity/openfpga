* NGSPICE file created from cby_0__1_.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_12 abstract view
.subckt sky130_fd_sc_hd__decap_12 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A X VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_1 abstract view
.subckt sky130_fd_sc_hd__dfxtp_1 D Q CLK VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A X VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A X VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
.subckt sky130_fd_sc_hd__conb_1 HI LO VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S X VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A X VGND VNB VPB VPWR
.ends

.subckt cby_0__1_ ccff_head ccff_tail chany_bottom_in[0] chany_bottom_in[10] chany_bottom_in[11]
+ chany_bottom_in[12] chany_bottom_in[13] chany_bottom_in[14] chany_bottom_in[15]
+ chany_bottom_in[16] chany_bottom_in[17] chany_bottom_in[18] chany_bottom_in[19]
+ chany_bottom_in[1] chany_bottom_in[2] chany_bottom_in[3] chany_bottom_in[4] chany_bottom_in[5]
+ chany_bottom_in[6] chany_bottom_in[7] chany_bottom_in[8] chany_bottom_in[9] chany_bottom_out[0]
+ chany_bottom_out[10] chany_bottom_out[11] chany_bottom_out[12] chany_bottom_out[13]
+ chany_bottom_out[14] chany_bottom_out[15] chany_bottom_out[16] chany_bottom_out[17]
+ chany_bottom_out[18] chany_bottom_out[19] chany_bottom_out[1] chany_bottom_out[2]
+ chany_bottom_out[3] chany_bottom_out[4] chany_bottom_out[5] chany_bottom_out[6]
+ chany_bottom_out[7] chany_bottom_out[8] chany_bottom_out[9] chany_top_in[0] chany_top_in[10]
+ chany_top_in[11] chany_top_in[12] chany_top_in[13] chany_top_in[14] chany_top_in[15]
+ chany_top_in[16] chany_top_in[17] chany_top_in[18] chany_top_in[19] chany_top_in[1]
+ chany_top_in[2] chany_top_in[3] chany_top_in[4] chany_top_in[5] chany_top_in[6]
+ chany_top_in[7] chany_top_in[8] chany_top_in[9] chany_top_out[0] chany_top_out[10]
+ chany_top_out[11] chany_top_out[12] chany_top_out[13] chany_top_out[14] chany_top_out[15]
+ chany_top_out[16] chany_top_out[17] chany_top_out[18] chany_top_out[19] chany_top_out[1]
+ chany_top_out[2] chany_top_out[3] chany_top_out[4] chany_top_out[5] chany_top_out[6]
+ chany_top_out[7] chany_top_out[8] chany_top_out[9] gfpga_pad_EMBEDDED_IO_SOC_DIR
+ gfpga_pad_EMBEDDED_IO_SOC_IN gfpga_pad_EMBEDDED_IO_SOC_OUT left_grid_pin_0_ prog_clk
+ right_width_0_height_0__pin_0_ right_width_0_height_0__pin_1_lower right_width_0_height_0__pin_1_upper
+ VPWR VGND
XFILLER_7_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_50_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mem_right_ipin_0.sky130_fd_sc_hd__dfxtp_1_2__CLK clkbuf_1_1_0_prog_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_mux_right_ipin_0.sky130_fd_sc_hd__buf_4_0__A mux_right_ipin_0.mux_l4_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_61_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mux_right_ipin_0.mux_l1_in_0__S mux_right_ipin_0.mux_l1_in_2_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_1_0_0_prog_clk_A clkbuf_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_ipin_0.mux_l1_in_1__A0 chany_top_in[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__04__A chany_bottom_in[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_mux_right_ipin_0.mux_l2_in_0__A0 mux_right_ipin_0.mux_l1_in_1_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_mem_right_ipin_0.sky130_fd_sc_hd__dfxtp_1_0__D ccff_head VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_7_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__12__A chany_bottom_in[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__07__A chany_bottom_in[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_right_ipin_0.mux_l1_in_1__A1 chany_bottom_in[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_29_ chany_top_in[11] chany_bottom_out[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_61_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mem_right_ipin_0.sky130_fd_sc_hd__dfxtp_1_3__D mux_right_ipin_0.mux_l3_in_1_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__20__A gfpga_pad_EMBEDDED_IO_SOC_IN VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_mux_right_ipin_0.mux_l2_in_0__A1 mux_right_ipin_0.mux_l1_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15__A chany_bottom_in[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_45_ chany_bottom_in[15] chany_top_out[15] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_61_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__23__A chany_top_in[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28_ chany_top_in[12] chany_bottom_out[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_61_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__18__A right_width_0_height_0__pin_0_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_right_ipin_0.mux_l2_in_1__S mux_right_ipin_0.mux_l2_in_3_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__31__A chany_top_in[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__26__A chany_top_in[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_44_ chany_bottom_in[16] chany_top_out[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_59_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_27_ chany_top_in[13] chany_bottom_out[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_1_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_right_ipin_0.mux_l2_in_3__A0 _01_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__34__A chany_top_in[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_56_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__29__A chany_top_in[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_0 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_ltile_io_mode_io__0.ltile_io_physical__iopad_0.EMBEDDED_IO_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_0__CLK
+ clkbuf_1_0_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__42__A chany_bottom_in[18] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__37__A chany_top_in[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_43_ chany_bottom_in[17] chany_top_out[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_55_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_26_ chany_top_in[14] chany_bottom_out[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XANTENNA_mux_right_ipin_0.mux_l2_in_3__A1 chany_top_in[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09_ chany_bottom_in[7] chany_top_out[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XPHY_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_56_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__45__A chany_bottom_in[15] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmem_right_ipin_0.sky130_fd_sc_hd__dfxtp_1_3_ mux_right_ipin_0.mux_l3_in_1_/S mux_right_ipin_0.mux_l4_in_0_/S
+ clkbuf_1_0_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_53_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_42_ chany_bottom_in[18] chany_top_out[18] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_55_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_25_ chany_top_in[15] chany_bottom_out[15] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_1_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08_ chany_bottom_in[8] chany_top_out[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_56_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmem_right_ipin_0.sky130_fd_sc_hd__dfxtp_1_2_ mux_right_ipin_0.mux_l2_in_3_/S mux_right_ipin_0.mux_l3_in_1_/S
+ clkbuf_1_1_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_16_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_41_ chany_bottom_in[19] chany_top_out[19] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_34_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24_ chany_top_in[16] chany_bottom_out[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_45_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07_ chany_bottom_in[9] chany_top_out[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XPHY_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_right_ipin_0.sky130_fd_sc_hd__dfxtp_1_1_ mux_right_ipin_0.mux_l1_in_2_/S mux_right_ipin_0.mux_l2_in_3_/S
+ clkbuf_1_1_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_42_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_40_ chany_top_in[0] chany_bottom_out[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_13_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23_ chany_top_in[17] chany_bottom_out[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_61_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_06_ chany_bottom_in[10] chany_top_out[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_25_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_56_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_right_ipin_0.sky130_fd_sc_hd__dfxtp_1_0_ ccff_head mux_right_ipin_0.mux_l1_in_2_/S
+ clkbuf_1_1_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XANTENNA_clkbuf_1_1_0_prog_clk_A clkbuf_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_right_ipin_0.mux_l4_in_0__S mux_right_ipin_0.mux_l4_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22_ chany_top_in[18] chany_bottom_out[18] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_60_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_05_ chany_bottom_in[11] chany_top_out[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XPHY_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_56_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_59_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21_ chany_top_in[19] chany_bottom_out[19] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_28_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_04_ chany_bottom_in[12] chany_top_out[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XPHY_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mem_right_ipin_0.sky130_fd_sc_hd__dfxtp_1_1__CLK clkbuf_1_1_0_prog_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_20_ gfpga_pad_EMBEDDED_IO_SOC_IN right_width_0_height_0__pin_1_upper VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__buf_2
XFILLER_37_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_0_prog_clk prog_clk clkbuf_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__clkbuf_16
XFILLER_28_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_03_ chany_bottom_in[13] chany_top_out[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XPHY_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_right_ipin_0.mux_l1_in_0__A0 chany_top_in[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_02_ chany_bottom_in[14] chany_top_out[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XPHY_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_right_ipin_0.mux_l1_in_1__S mux_right_ipin_0.mux_l1_in_2_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_right_ipin_0.sky130_fd_sc_hd__buf_4_0_ mux_right_ipin_0.mux_l4_in_0_/X left_grid_pin_0_
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_4
XFILLER_58_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__02__A chany_bottom_in[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_right_ipin_0.mux_l1_in_0__A1 chany_bottom_in[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_51_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_01_ _01_/HI _01_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XFILLER_33_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__10__A chany_bottom_in[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_57_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__05__A chany_bottom_in[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mem_right_ipin_0.sky130_fd_sc_hd__dfxtp_1_1__D mux_right_ipin_0.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_43_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__13__A chany_bottom_in[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__08__A chany_bottom_in[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_51_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__21__A chany_top_in[19] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__16__A chany_bottom_in[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_43_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_right_ipin_0.mux_l2_in_3_ _01_/HI chany_top_in[16] mux_right_ipin_0.mux_l2_in_3_/S
+ mux_right_ipin_0.mux_l2_in_3_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_4_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_clkbuf_0_prog_clk_A prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_right_ipin_0.mux_l4_in_0_ mux_right_ipin_0.mux_l3_in_1_/X mux_right_ipin_0.mux_l3_in_0_/X
+ mux_right_ipin_0.mux_l4_in_0_/S mux_right_ipin_0.mux_l4_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XFILLER_10_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_right_ipin_0.mux_l2_in_2__A0 chany_bottom_in[16] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_18_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24__A chany_top_in[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__19__A gfpga_pad_EMBEDDED_IO_SOC_IN VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_right_ipin_0.mux_l3_in_1_ mux_right_ipin_0.mux_l2_in_3_/X mux_right_ipin_0.mux_l2_in_2_/X
+ mux_right_ipin_0.mux_l3_in_1_/S mux_right_ipin_0.mux_l3_in_1_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XFILLER_23_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_ipin_0.mux_l3_in_1__A0 mux_right_ipin_0.mux_l2_in_3_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_right_ipin_0.mux_l2_in_2_ chany_bottom_in[16] chany_top_in[10] mux_right_ipin_0.mux_l2_in_3_/S
+ mux_right_ipin_0.mux_l2_in_2_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mux_right_ipin_0.mux_l2_in_2__S mux_right_ipin_0.mux_l2_in_3_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__32__A chany_top_in[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xltile_io_mode_io__0.ltile_io_physical__iopad_0.EMBEDDED_IO_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_0_
+ mux_right_ipin_0.mux_l4_in_0_/S ccff_tail clkbuf_1_0_0_prog_clk/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__dfxtp_1
XANTENNA_mux_right_ipin_0.mux_l4_in_0__A0 mux_right_ipin_0.mux_l3_in_1_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__27__A chany_top_in[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__40__A chany_top_in[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_right_ipin_0.mux_l2_in_2__A1 chany_top_in[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_62_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__35__A chany_top_in[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_right_ipin_0.mux_l3_in_0_ mux_right_ipin_0.mux_l2_in_1_/X mux_right_ipin_0.mux_l2_in_0_/X
+ mux_right_ipin_0.mux_l3_in_1_/S mux_right_ipin_0.mux_l3_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XFILLER_21_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_right_ipin_0.mux_l3_in_1__A1 mux_right_ipin_0.mux_l2_in_2_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_right_ipin_0.mux_l2_in_1_ chany_bottom_in[10] mux_right_ipin_0.mux_l1_in_2_/X
+ mux_right_ipin_0.mux_l2_in_3_/S mux_right_ipin_0.mux_l2_in_1_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XPHY_260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_mux_right_ipin_0.mux_l4_in_0__A1 mux_right_ipin_0.mux_l3_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_57_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__43__A chany_bottom_in[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmux_right_ipin_0.mux_l1_in_2_ chany_top_in[4] chany_bottom_in[4] mux_right_ipin_0.mux_l1_in_2_/S
+ mux_right_ipin_0.mux_l1_in_2_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_24_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__38__A chany_top_in[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_right_ipin_0.mux_l2_in_0_ mux_right_ipin_0.mux_l1_in_1_/X mux_right_ipin_0.mux_l1_in_0_/X
+ mux_right_ipin_0.mux_l2_in_3_/S mux_right_ipin_0.mux_l2_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XPHY_261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_right_ipin_0.mux_l3_in_0__S mux_right_ipin_0.mux_l3_in_1_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_right_ipin_0.mux_l1_in_1_ chany_top_in[2] chany_bottom_in[2] mux_right_ipin_0.mux_l1_in_2_/S
+ mux_right_ipin_0.mux_l1_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_36_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_39_ chany_top_in[1] chany_bottom_out[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_32_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_right_ipin_0.mux_l1_in_0_ chany_top_in[0] chany_bottom_in[0] mux_right_ipin_0.mux_l1_in_2_/S
+ mux_right_ipin_0.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_60_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_42_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_38_ chany_top_in[2] chany_bottom_out[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_11_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_37_ chany_top_in[3] chany_bottom_out[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_57_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_36_ chany_top_in[4] chany_bottom_out[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_20_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mem_right_ipin_0.sky130_fd_sc_hd__dfxtp_1_0__CLK clkbuf_1_1_0_prog_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_19_ gfpga_pad_EMBEDDED_IO_SOC_IN right_width_0_height_0__pin_1_lower VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__buf_2
XPHY_254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_35_ chany_top_in[5] chany_bottom_out[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_57_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18_ right_width_0_height_0__pin_0_ gfpga_pad_EMBEDDED_IO_SOC_OUT VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__buf_2
XFILLER_40_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_34_ chany_top_in[6] chany_bottom_out[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_11_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_17_ ccff_tail gfpga_pad_EMBEDDED_IO_SOC_DIR VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_8_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mem_right_ipin_0.sky130_fd_sc_hd__dfxtp_1_3__CLK clkbuf_1_0_0_prog_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_33_ chany_top_in[7] chany_bottom_out[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_14_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_16_ chany_bottom_in[0] chany_top_out[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_26_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_right_ipin_0.mux_l1_in_2__S mux_right_ipin_0.mux_l1_in_2_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__03__A chany_bottom_in[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_32_ chany_top_in[8] chany_bottom_out[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_47_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11__A chany_bottom_in[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15_ chany_bottom_in[1] chany_top_out[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_8_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06__A chany_bottom_in[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mem_right_ipin_0.sky130_fd_sc_hd__dfxtp_1_2__D mux_right_ipin_0.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_44_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_ipin_0.mux_l1_in_2__A0 chany_top_in[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__14__A chany_bottom_in[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mux_right_ipin_0.mux_l2_in_1__A0 chany_bottom_in[10] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XPHY_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__09__A chany_bottom_in[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_31_ chany_top_in[9] chany_bottom_out[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XANTENNA_mux_right_ipin_0.mux_l3_in_0__A0 mux_right_ipin_0.mux_l2_in_1_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14_ chany_bottom_in[2] chany_top_out[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XPHY_259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__22__A chany_top_in[18] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__17__A ccff_tail VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_right_ipin_0.mux_l1_in_2__A1 chany_bottom_in[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mux_right_ipin_0.mux_l2_in_0__S mux_right_ipin_0.mux_l2_in_3_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__30__A chany_top_in[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mux_right_ipin_0.mux_l2_in_1__A1 mux_right_ipin_0.mux_l1_in_2_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__25__A chany_top_in[15] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_30_ chany_top_in[10] chany_bottom_out[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_61_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_right_ipin_0.mux_l3_in_0__A1 mux_right_ipin_0.mux_l2_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13_ chany_bottom_in[3] chany_top_out[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XPHY_249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_right_ipin_0.mux_l2_in_3__S mux_right_ipin_0.mux_l2_in_3_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__33__A chany_top_in[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__28__A chany_top_in[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_50_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__41__A chany_bottom_in[19] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__36__A chany_top_in[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12_ chany_bottom_in[4] chany_top_out[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_6_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__44__A chany_bottom_in[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__39__A chany_top_in[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11_ chany_bottom_in[5] chany_top_out[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XPHY_229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_1_1_0_prog_clk clkbuf_0_prog_clk/X clkbuf_1_1_0_prog_clk/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_30_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_right_ipin_0.mux_l3_in_1__S mux_right_ipin_0.mux_l3_in_1_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_10_ chany_bottom_in[6] chany_top_out[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XPHY_219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_59_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_56_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_io_mode_io__0.ltile_io_physical__iopad_0.EMBEDDED_IO_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_0__D
+ mux_right_ipin_0.mux_l4_in_0_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_1_0_0_prog_clk clkbuf_0_prog_clk/X clkbuf_1_0_0_prog_clk/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_31_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_58_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
.ends

