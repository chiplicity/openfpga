* NGSPICE file created from decoder6to61.ext - technology: EFS8A

* Black-box entry subcircuit for scs8hd_decap_12 abstract view
.subckt scs8hd_decap_12 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_decap_3 abstract view
.subckt scs8hd_decap_3 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_diode_2 abstract view
.subckt scs8hd_diode_2 DIODE vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_inv_8 abstract view
.subckt scs8hd_inv_8 A Y vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_fill_2 abstract view
.subckt scs8hd_fill_2 vpwr vgnd
.ends

* Black-box entry subcircuit for scs8hd_buf_1 abstract view
.subckt scs8hd_buf_1 A X vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_decap_4 abstract view
.subckt scs8hd_decap_4 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_fill_1 abstract view
.subckt scs8hd_fill_1 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_decap_6 abstract view
.subckt scs8hd_decap_6 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_tapvpwrvgnd_1 abstract view
.subckt scs8hd_tapvpwrvgnd_1 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_nor2_4 abstract view
.subckt scs8hd_nor2_4 A B Y vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_decap_8 abstract view
.subckt scs8hd_decap_8 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_or4_4 abstract view
.subckt scs8hd_or4_4 A B C D X vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_or3_4 abstract view
.subckt scs8hd_or3_4 A B C X vgnd vpwr
.ends

.subckt decoder6to61 address[0] address[1] address[2] address[3] address[4] address[5]
+ data_out[0] data_out[10] data_out[11] data_out[12] data_out[13] data_out[14] data_out[15]
+ data_out[16] data_out[17] data_out[18] data_out[19] data_out[1] data_out[20] data_out[21]
+ data_out[22] data_out[23] data_out[24] data_out[25] data_out[26] data_out[27] data_out[28]
+ data_out[29] data_out[2] data_out[30] data_out[31] data_out[32] data_out[33] data_out[34]
+ data_out[35] data_out[36] data_out[37] data_out[38] data_out[39] data_out[3] data_out[40]
+ data_out[41] data_out[42] data_out[43] data_out[44] data_out[45] data_out[46] data_out[47]
+ data_out[48] data_out[49] data_out[4] data_out[50] data_out[51] data_out[52] data_out[53]
+ data_out[54] data_out[55] data_out[56] data_out[57] data_out[58] data_out[59] data_out[5]
+ data_out[60] data_out[6] data_out[7] data_out[8] data_out[9] enable vpwr vgnd
XFILLER_22_166 vgnd vpwr scs8hd_decap_12
XFILLER_26_41 vgnd vpwr scs8hd_decap_3
XANTENNA__113__B _112_/B vgnd vpwr scs8hd_diode_2
XFILLER_9_159 vgnd vpwr scs8hd_decap_12
XANTENNA__108__B _142_/B vgnd vpwr scs8hd_diode_2
XFILLER_6_129 vgnd vpwr scs8hd_decap_12
XANTENNA__124__A _092_/X vgnd vpwr scs8hd_diode_2
XFILLER_5_184 vgnd vpwr scs8hd_decap_12
X_062_ address[4] _063_/A vgnd vpwr scs8hd_inv_8
XFILLER_23_75 vgnd vpwr scs8hd_decap_12
XFILLER_23_53 vpwr vgnd scs8hd_fill_2
X_131_ _181_/A _151_/A vgnd vpwr scs8hd_buf_1
XANTENNA__119__A _089_/A vgnd vpwr scs8hd_diode_2
XFILLER_2_154 vgnd vpwr scs8hd_decap_12
XFILLER_9_33 vpwr vgnd scs8hd_fill_2
XFILLER_34_41 vpwr vgnd scs8hd_fill_2
X_114_ address[2] _154_/A vgnd vpwr scs8hd_buf_1
XFILLER_11_220 vgnd vpwr scs8hd_decap_12
XFILLER_29_117 vgnd vpwr scs8hd_decap_4
XFILLER_29_41 vgnd vpwr scs8hd_fill_1
XFILLER_20_32 vpwr vgnd scs8hd_fill_2
XFILLER_20_10 vpwr vgnd scs8hd_fill_2
XFILLER_4_227 vgnd vpwr scs8hd_decap_6
XFILLER_13_3 vgnd vpwr scs8hd_decap_3
XANTENNA__132__A _151_/A vgnd vpwr scs8hd_diode_2
XFILLER_6_23 vpwr vgnd scs8hd_fill_2
XFILLER_6_89 vgnd vpwr scs8hd_decap_3
XFILLER_31_31 vpwr vgnd scs8hd_fill_2
XFILLER_15_65 vpwr vgnd scs8hd_fill_2
XFILLER_1_208 vgnd vpwr scs8hd_decap_12
XPHY_192 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_31_123 vgnd vpwr scs8hd_decap_12
XPHY_181 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_170 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_0_230 vgnd vpwr scs8hd_decap_3
XANTENNA__127__A _090_/X vgnd vpwr scs8hd_diode_2
XFILLER_22_178 vgnd vpwr scs8hd_decap_12
XFILLER_26_64 vgnd vpwr scs8hd_decap_12
XFILLER_26_53 vpwr vgnd scs8hd_fill_2
XFILLER_13_123 vgnd vpwr scs8hd_decap_12
XFILLER_18_215 vgnd vpwr scs8hd_decap_12
XFILLER_12_22 vpwr vgnd scs8hd_fill_2
XANTENNA__140__A _147_/A vgnd vpwr scs8hd_diode_2
XANTENNA__108__C _107_/X vgnd vpwr scs8hd_diode_2
XANTENNA__124__B _124_/B vgnd vpwr scs8hd_diode_2
XFILLER_5_196 vgnd vpwr scs8hd_decap_12
X_130_ _092_/X _134_/B data_out[3] vgnd vpwr scs8hd_nor2_4
XFILLER_23_87 vgnd vpwr scs8hd_decap_12
XANTENNA__135__A _171_/A vgnd vpwr scs8hd_diode_2
XFILLER_2_166 vgnd vpwr scs8hd_decap_12
XANTENNA__119__B _116_/X vgnd vpwr scs8hd_diode_2
XFILLER_9_56 vgnd vpwr scs8hd_decap_3
XFILLER_34_20 vgnd vpwr scs8hd_fill_1
XFILLER_18_10 vpwr vgnd scs8hd_fill_2
XFILLER_11_232 vgnd vpwr scs8hd_fill_1
X_113_ _090_/X _112_/B data_out[12] vgnd vpwr scs8hd_nor2_4
XFILLER_29_53 vpwr vgnd scs8hd_fill_2
XFILLER_29_20 vpwr vgnd scs8hd_fill_2
XFILLER_20_77 vgnd vpwr scs8hd_decap_12
XFILLER_19_184 vgnd vpwr scs8hd_decap_12
XANTENNA__132__B _134_/B vgnd vpwr scs8hd_diode_2
XFILLER_34_154 vgnd vpwr scs8hd_decap_12
XFILLER_15_55 vpwr vgnd scs8hd_fill_2
XFILLER_15_33 vgnd vpwr scs8hd_decap_3
XPHY_193 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_31_135 vgnd vpwr scs8hd_decap_12
XFILLER_31_65 vpwr vgnd scs8hd_fill_2
XFILLER_31_54 vpwr vgnd scs8hd_fill_2
XPHY_182 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_171 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_160 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_16_154 vgnd vpwr scs8hd_decap_12
XFILLER_15_77 vgnd vpwr scs8hd_decap_12
XANTENNA__127__B _124_/B vgnd vpwr scs8hd_diode_2
XANTENNA__143__A _142_/X vgnd vpwr scs8hd_diode_2
XFILLER_30_190 vgnd vpwr scs8hd_decap_12
XFILLER_26_76 vgnd vpwr scs8hd_decap_12
XFILLER_13_135 vgnd vpwr scs8hd_decap_12
XANTENNA__138__A _138_/A vgnd vpwr scs8hd_diode_2
XFILLER_12_190 vgnd vpwr scs8hd_decap_12
XFILLER_3_14 vpwr vgnd scs8hd_fill_2
XFILLER_3_36 vpwr vgnd scs8hd_fill_2
XFILLER_3_47 vpwr vgnd scs8hd_fill_2
XFILLER_10_105 vgnd vpwr scs8hd_decap_12
XFILLER_33_208 vgnd vpwr scs8hd_decap_12
XANTENNA__140__B _139_/X vgnd vpwr scs8hd_diode_2
XFILLER_18_227 vgnd vpwr scs8hd_decap_6
XANTENNA__108__D _064_/X vgnd vpwr scs8hd_diode_2
XFILLER_15_208 vgnd vpwr scs8hd_decap_12
XFILLER_23_99 vgnd vpwr scs8hd_decap_12
XFILLER_23_33 vgnd vpwr scs8hd_decap_4
XFILLER_23_22 vpwr vgnd scs8hd_fill_2
XFILLER_0_15 vpwr vgnd scs8hd_fill_2
XFILLER_2_178 vgnd vpwr scs8hd_decap_12
XFILLER_3_3 vpwr vgnd scs8hd_fill_2
XFILLER_9_13 vpwr vgnd scs8hd_fill_2
XANTENNA__151__A _151_/A vgnd vpwr scs8hd_diode_2
X_112_ _089_/A _112_/B data_out[13] vgnd vpwr scs8hd_nor2_4
XANTENNA__146__A _146_/A vgnd vpwr scs8hd_diode_2
XFILLER_22_9 vgnd vpwr scs8hd_decap_3
XFILLER_20_89 vgnd vpwr scs8hd_decap_3
XFILLER_20_23 vpwr vgnd scs8hd_fill_2
XFILLER_29_65 vpwr vgnd scs8hd_fill_2
XFILLER_28_141 vgnd vpwr scs8hd_decap_12
XFILLER_20_6 vpwr vgnd scs8hd_fill_2
XFILLER_6_14 vpwr vgnd scs8hd_fill_2
XFILLER_34_166 vgnd vpwr scs8hd_decap_12
XFILLER_19_196 vgnd vpwr scs8hd_decap_12
XFILLER_31_11 vgnd vpwr scs8hd_decap_8
XFILLER_16_166 vgnd vpwr scs8hd_decap_12
XFILLER_15_89 vgnd vpwr scs8hd_decap_12
XFILLER_15_12 vpwr vgnd scs8hd_fill_2
XPHY_194 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_31_147 vgnd vpwr scs8hd_decap_12
XPHY_183 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_172 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_161 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_150 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_26_88 vgnd vpwr scs8hd_decap_4
XFILLER_13_147 vgnd vpwr scs8hd_decap_12
XFILLER_9_107 vgnd vpwr scs8hd_decap_12
XANTENNA__154__A _154_/A vgnd vpwr scs8hd_diode_2
XFILLER_3_59 vpwr vgnd scs8hd_fill_2
XANTENNA__064__A address[5] vgnd vpwr scs8hd_diode_2
XFILLER_12_35 vpwr vgnd scs8hd_fill_2
XFILLER_10_117 vgnd vpwr scs8hd_decap_12
XFILLER_5_110 vgnd vpwr scs8hd_decap_12
XANTENNA__149__A _149_/A vgnd vpwr scs8hd_diode_2
XFILLER_23_220 vgnd vpwr scs8hd_decap_12
XFILLER_0_27 vpwr vgnd scs8hd_fill_2
XANTENNA__151__B _149_/X vgnd vpwr scs8hd_diode_2
XFILLER_29_3 vpwr vgnd scs8hd_fill_2
XFILLER_18_67 vpwr vgnd scs8hd_fill_2
XFILLER_18_45 vpwr vgnd scs8hd_fill_2
XFILLER_18_23 vpwr vgnd scs8hd_fill_2
XANTENNA__146__B _147_/B vgnd vpwr scs8hd_diode_2
X_111_ _086_/X _112_/B data_out[14] vgnd vpwr scs8hd_nor2_4
XANTENNA__162__A _144_/A vgnd vpwr scs8hd_diode_2
XANTENNA__072__A _071_/X vgnd vpwr scs8hd_diode_2
XFILLER_29_33 vpwr vgnd scs8hd_fill_2
XFILLER_34_178 vgnd vpwr scs8hd_decap_12
XANTENNA__157__A _151_/A vgnd vpwr scs8hd_diode_2
XFILLER_25_123 vgnd vpwr scs8hd_decap_12
XANTENNA__067__A _063_/X vgnd vpwr scs8hd_diode_2
XFILLER_0_211 vgnd vpwr scs8hd_decap_6
XPHY_195 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_31_159 vgnd vpwr scs8hd_decap_12
XPHY_184 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_173 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_162 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_151 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_140 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_16_178 vgnd vpwr scs8hd_decap_12
XFILLER_11_3 vgnd vpwr scs8hd_fill_1
XFILLER_26_23 vpwr vgnd scs8hd_fill_2
XFILLER_13_159 vgnd vpwr scs8hd_decap_12
XFILLER_9_119 vgnd vpwr scs8hd_decap_3
XANTENNA__154__B _148_/B vgnd vpwr scs8hd_diode_2
XANTENNA__170__A _146_/A vgnd vpwr scs8hd_diode_2
XFILLER_12_14 vpwr vgnd scs8hd_fill_2
XFILLER_10_129 vgnd vpwr scs8hd_decap_12
XFILLER_8_141 vgnd vpwr scs8hd_decap_12
XANTENNA__080__A _068_/X vgnd vpwr scs8hd_diode_2
XANTENNA__165__A _147_/A vgnd vpwr scs8hd_diode_2
XFILLER_23_232 vgnd vpwr scs8hd_fill_1
XFILLER_23_57 vpwr vgnd scs8hd_fill_2
XANTENNA__075__A _071_/A vgnd vpwr scs8hd_diode_2
XFILLER_9_37 vgnd vpwr scs8hd_decap_4
XFILLER_20_202 vgnd vpwr scs8hd_decap_12
XFILLER_34_89 vgnd vpwr scs8hd_decap_3
XFILLER_34_45 vgnd vpwr scs8hd_decap_12
XFILLER_34_23 vgnd vpwr scs8hd_decap_8
XFILLER_34_12 vpwr vgnd scs8hd_fill_2
X_110_ _092_/X _112_/B data_out[15] vgnd vpwr scs8hd_nor2_4
XANTENNA__162__B _165_/B vgnd vpwr scs8hd_diode_2
XFILLER_1_60 vgnd vpwr scs8hd_fill_1
XFILLER_28_154 vgnd vpwr scs8hd_decap_12
XFILLER_20_36 vpwr vgnd scs8hd_fill_2
XANTENNA__157__B _155_/X vgnd vpwr scs8hd_diode_2
XANTENNA__173__A _172_/X vgnd vpwr scs8hd_diode_2
XFILLER_3_220 vgnd vpwr scs8hd_decap_12
XFILLER_6_27 vpwr vgnd scs8hd_fill_2
XFILLER_31_35 vpwr vgnd scs8hd_fill_2
XFILLER_25_135 vgnd vpwr scs8hd_decap_12
XFILLER_15_69 vpwr vgnd scs8hd_fill_2
XANTENNA__067__B _064_/X vgnd vpwr scs8hd_diode_2
XANTENNA__083__A _071_/A vgnd vpwr scs8hd_diode_2
XPHY_196 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_185 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_31_105 vgnd vpwr scs8hd_decap_12
XPHY_174 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_163 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_190 vgnd vpwr scs8hd_decap_12
XPHY_152 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_141 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_130 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__168__A _144_/A vgnd vpwr scs8hd_diode_2
XFILLER_22_105 vgnd vpwr scs8hd_decap_12
XFILLER_26_57 vgnd vpwr scs8hd_decap_4
XFILLER_26_35 vgnd vpwr scs8hd_decap_4
XFILLER_21_171 vgnd vpwr scs8hd_decap_12
XANTENNA__078__A _071_/A vgnd vpwr scs8hd_diode_2
XFILLER_35_230 vgnd vpwr scs8hd_decap_3
XANTENNA__154__C _063_/A vgnd vpwr scs8hd_diode_2
XFILLER_27_208 vgnd vpwr scs8hd_decap_12
XANTENNA__170__B _167_/X vgnd vpwr scs8hd_diode_2
XFILLER_16_90 vpwr vgnd scs8hd_fill_2
XANTENNA__080__B _171_/A vgnd vpwr scs8hd_diode_2
XFILLER_12_59 vgnd vpwr scs8hd_fill_1
XFILLER_12_26 vpwr vgnd scs8hd_fill_2
XANTENNA__165__B _165_/B vgnd vpwr scs8hd_diode_2
XFILLER_5_123 vgnd vpwr scs8hd_decap_12
XANTENNA__181__A _181_/A vgnd vpwr scs8hd_diode_2
XFILLER_4_93 vgnd vpwr scs8hd_decap_12
XANTENNA__075__B _074_/Y vgnd vpwr scs8hd_diode_2
XANTENNA__091__A _090_/X vgnd vpwr scs8hd_diode_2
XANTENNA__176__A _176_/A vgnd vpwr scs8hd_diode_2
XFILLER_34_57 vgnd vpwr scs8hd_decap_12
XANTENNA__086__A _181_/A vgnd vpwr scs8hd_diode_2
XFILLER_1_3 vpwr vgnd scs8hd_fill_2
X_169_ _151_/A _167_/X data_out[42] vgnd vpwr scs8hd_nor2_4
XFILLER_29_57 vpwr vgnd scs8hd_fill_2
XFILLER_28_166 vgnd vpwr scs8hd_decap_12
XFILLER_19_90 vgnd vpwr scs8hd_decap_12
XFILLER_10_81 vgnd vpwr scs8hd_decap_8
XFILLER_3_232 vgnd vpwr scs8hd_fill_1
XFILLER_31_58 vgnd vpwr scs8hd_decap_3
XFILLER_25_147 vgnd vpwr scs8hd_decap_12
XFILLER_15_59 vpwr vgnd scs8hd_fill_2
XANTENNA__067__C _065_/Y vgnd vpwr scs8hd_diode_2
XANTENNA__083__B _074_/Y vgnd vpwr scs8hd_diode_2
XPHY_197 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_186 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_31_117 vgnd vpwr scs8hd_decap_4
XFILLER_31_69 vgnd vpwr scs8hd_decap_12
XPHY_175 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_164 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_153 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_142 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_131 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_120 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__168__B _167_/X vgnd vpwr scs8hd_diode_2
XFILLER_22_117 vgnd vpwr scs8hd_decap_12
XANTENNA__184__A _068_/X vgnd vpwr scs8hd_diode_2
XPHY_0 vgnd vpwr scs8hd_decap_3
XFILLER_13_106 vgnd vpwr scs8hd_decap_12
XANTENNA__078__B address[0] vgnd vpwr scs8hd_diode_2
XFILLER_3_18 vpwr vgnd scs8hd_fill_2
XANTENNA__094__A _093_/X vgnd vpwr scs8hd_diode_2
XANTENNA__154__D _148_/D vgnd vpwr scs8hd_diode_2
XANTENNA__179__A _178_/X vgnd vpwr scs8hd_diode_2
XFILLER_8_154 vgnd vpwr scs8hd_decap_12
XANTENNA__089__A _089_/A vgnd vpwr scs8hd_diode_2
XFILLER_17_220 vgnd vpwr scs8hd_decap_12
XFILLER_5_135 vgnd vpwr scs8hd_decap_12
XFILLER_23_37 vgnd vpwr scs8hd_fill_1
XFILLER_23_26 vpwr vgnd scs8hd_fill_2
XANTENNA__181__B _179_/X vgnd vpwr scs8hd_diode_2
XANTENNA__075__C address[1] vgnd vpwr scs8hd_diode_2
XFILLER_4_190 vgnd vpwr scs8hd_decap_12
XFILLER_13_70 vgnd vpwr scs8hd_decap_12
XANTENNA__091__B _082_/X vgnd vpwr scs8hd_diode_2
XFILLER_0_19 vpwr vgnd scs8hd_fill_2
XFILLER_2_105 vgnd vpwr scs8hd_decap_12
XFILLER_9_17 vpwr vgnd scs8hd_fill_2
XFILLER_20_215 vgnd vpwr scs8hd_decap_12
XANTENNA__176__B _174_/B vgnd vpwr scs8hd_diode_2
XFILLER_1_171 vgnd vpwr scs8hd_decap_12
XFILLER_34_69 vgnd vpwr scs8hd_decap_12
XFILLER_7_208 vgnd vpwr scs8hd_decap_12
X_168_ _144_/A _167_/X data_out[43] vgnd vpwr scs8hd_nor2_4
X_099_ _063_/X _064_/X address[2] address[3] _099_/X vgnd vpwr scs8hd_or4_4
XFILLER_29_69 vgnd vpwr scs8hd_decap_12
XFILLER_20_49 vpwr vgnd scs8hd_fill_2
XFILLER_20_27 vpwr vgnd scs8hd_fill_2
XFILLER_1_62 vgnd vpwr scs8hd_decap_12
XFILLER_28_178 vgnd vpwr scs8hd_decap_12
XFILLER_19_123 vgnd vpwr scs8hd_decap_12
XFILLER_10_93 vgnd vpwr scs8hd_decap_12
XFILLER_6_18 vgnd vpwr scs8hd_decap_3
XANTENNA__097__A _089_/A vgnd vpwr scs8hd_diode_2
XFILLER_25_159 vgnd vpwr scs8hd_decap_12
XFILLER_25_104 vgnd vpwr scs8hd_decap_12
XFILLER_15_38 vpwr vgnd scs8hd_fill_2
XFILLER_15_16 vpwr vgnd scs8hd_fill_2
XANTENNA__067__D _066_/Y vgnd vpwr scs8hd_diode_2
XPHY_198 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_187 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_176 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_165 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_154 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_143 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_132 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_121 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__083__C _071_/C vgnd vpwr scs8hd_diode_2
XPHY_110 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_22_129 vgnd vpwr scs8hd_decap_12
XANTENNA__184__B _180_/A vgnd vpwr scs8hd_diode_2
XPHY_1 vgnd vpwr scs8hd_decap_3
XFILLER_21_184 vgnd vpwr scs8hd_decap_12
XFILLER_13_118 vgnd vpwr scs8hd_decap_4
XANTENNA__078__C address[1] vgnd vpwr scs8hd_diode_2
XFILLER_16_70 vpwr vgnd scs8hd_fill_2
XFILLER_8_166 vgnd vpwr scs8hd_decap_12
XANTENNA__089__B _082_/X vgnd vpwr scs8hd_diode_2
XFILLER_12_39 vgnd vpwr scs8hd_decap_3
XFILLER_5_147 vgnd vpwr scs8hd_decap_12
XFILLER_32_202 vgnd vpwr scs8hd_decap_12
XFILLER_17_232 vgnd vpwr scs8hd_fill_1
XFILLER_14_202 vgnd vpwr scs8hd_decap_12
XFILLER_2_117 vgnd vpwr scs8hd_decap_12
XFILLER_20_227 vgnd vpwr scs8hd_decap_6
X_184_ _068_/X _180_/A data_out[31] vgnd vpwr scs8hd_nor2_4
XFILLER_13_82 vgnd vpwr scs8hd_decap_12
XFILLER_13_60 vgnd vpwr scs8hd_fill_1
XFILLER_18_49 vgnd vpwr scs8hd_decap_3
XFILLER_18_27 vpwr vgnd scs8hd_fill_2
X_167_ _167_/A _167_/X vgnd vpwr scs8hd_buf_1
XFILLER_24_81 vgnd vpwr scs8hd_decap_8
X_098_ _090_/X _096_/B data_out[20] vgnd vpwr scs8hd_nor2_4
XFILLER_1_74 vgnd vpwr scs8hd_decap_12
XFILLER_1_52 vgnd vpwr scs8hd_decap_8
XFILLER_1_41 vpwr vgnd scs8hd_fill_2
XFILLER_29_37 vgnd vpwr scs8hd_decap_4
XFILLER_19_102 vgnd vpwr scs8hd_decap_12
XANTENNA__097__B _096_/B vgnd vpwr scs8hd_diode_2
XFILLER_10_50 vgnd vpwr scs8hd_decap_4
XFILLER_34_105 vgnd vpwr scs8hd_decap_12
XFILLER_19_135 vgnd vpwr scs8hd_decap_12
XFILLER_33_171 vgnd vpwr scs8hd_decap_12
XFILLER_25_116 vgnd vpwr scs8hd_decap_6
XFILLER_18_190 vgnd vpwr scs8hd_decap_12
XFILLER_16_105 vgnd vpwr scs8hd_decap_12
XPHY_100 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_199 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_188 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_177 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_166 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_155 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_21_71 vpwr vgnd scs8hd_fill_2
XPHY_144 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_133 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_15_171 vgnd vpwr scs8hd_decap_12
XPHY_122 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_111 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_2 vgnd vpwr scs8hd_decap_3
XFILLER_30_141 vgnd vpwr scs8hd_decap_12
XFILLER_26_27 vpwr vgnd scs8hd_fill_2
XFILLER_21_196 vgnd vpwr scs8hd_decap_12
XFILLER_7_51 vgnd vpwr scs8hd_decap_8
XFILLER_7_62 vgnd vpwr scs8hd_decap_12
XFILLER_32_81 vgnd vpwr scs8hd_decap_8
XFILLER_16_93 vgnd vpwr scs8hd_decap_12
XFILLER_12_141 vgnd vpwr scs8hd_decap_12
XFILLER_8_178 vgnd vpwr scs8hd_decap_12
XFILLER_35_211 vgnd vpwr scs8hd_decap_6
XFILLER_12_18 vpwr vgnd scs8hd_fill_2
XFILLER_5_159 vgnd vpwr scs8hd_decap_12
XFILLER_27_81 vgnd vpwr scs8hd_decap_12
XFILLER_4_41 vgnd vpwr scs8hd_decap_12
XFILLER_2_129 vgnd vpwr scs8hd_decap_12
X_183_ _171_/A _179_/X data_out[32] vgnd vpwr scs8hd_nor2_4
XFILLER_13_94 vgnd vpwr scs8hd_decap_12
XFILLER_1_184 vgnd vpwr scs8hd_decap_12
XFILLER_34_16 vgnd vpwr scs8hd_decap_4
XFILLER_24_93 vgnd vpwr scs8hd_decap_12
X_166_ _154_/A _142_/B _107_/X _148_/D _167_/A vgnd vpwr scs8hd_or4_4
X_097_ _089_/A _096_/B data_out[21] vgnd vpwr scs8hd_nor2_4
XFILLER_1_86 vgnd vpwr scs8hd_decap_12
XFILLER_29_16 vpwr vgnd scs8hd_fill_2
XFILLER_34_117 vgnd vpwr scs8hd_decap_12
X_149_ _149_/A _149_/X vgnd vpwr scs8hd_buf_1
XFILLER_32_3 vgnd vpwr scs8hd_fill_1
XFILLER_19_147 vgnd vpwr scs8hd_decap_12
XFILLER_19_114 vgnd vpwr scs8hd_decap_8
XFILLER_31_39 vpwr vgnd scs8hd_fill_2
XFILLER_15_29 vpwr vgnd scs8hd_fill_2
XPHY_189 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_178 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_167 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_156 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_145 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_134 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_16_117 vgnd vpwr scs8hd_decap_12
XPHY_123 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_112 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_101 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_3 vgnd vpwr scs8hd_decap_3
XFILLER_7_41 vgnd vpwr scs8hd_decap_8
XFILLER_7_74 vgnd vpwr scs8hd_decap_12
XFILLER_29_220 vgnd vpwr scs8hd_decap_12
XFILLER_32_93 vgnd vpwr scs8hd_decap_12
XFILLER_32_215 vgnd vpwr scs8hd_decap_12
XFILLER_27_93 vgnd vpwr scs8hd_decap_12
XFILLER_4_53 vgnd vpwr scs8hd_decap_12
X_182_ _176_/A _179_/X data_out[33] vgnd vpwr scs8hd_nor2_4
XFILLER_14_215 vgnd vpwr scs8hd_decap_12
XFILLER_13_62 vpwr vgnd scs8hd_fill_2
XFILLER_1_196 vgnd vpwr scs8hd_decap_12
XANTENNA__100__A _099_/X vgnd vpwr scs8hd_diode_2
X_165_ _147_/A _165_/B data_out[44] vgnd vpwr scs8hd_nor2_4
X_096_ _086_/X _096_/B data_out[22] vgnd vpwr scs8hd_nor2_4
XFILLER_1_98 vgnd vpwr scs8hd_decap_12
XFILLER_34_129 vgnd vpwr scs8hd_decap_12
X_148_ _148_/A _148_/B _063_/A _148_/D _149_/A vgnd vpwr scs8hd_or4_4
XFILLER_19_159 vgnd vpwr scs8hd_decap_12
XFILLER_19_50 vpwr vgnd scs8hd_fill_2
XFILLER_10_30 vgnd vpwr scs8hd_fill_1
XFILLER_33_184 vgnd vpwr scs8hd_decap_12
XFILLER_25_3 vpwr vgnd scs8hd_fill_2
X_079_ _079_/A _171_/A vgnd vpwr scs8hd_buf_1
XPHY_179 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_168 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_157 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_146 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_135 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_16_129 vgnd vpwr scs8hd_decap_12
XPHY_124 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_113 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_102 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_30_154 vgnd vpwr scs8hd_decap_12
XFILLER_15_184 vgnd vpwr scs8hd_decap_12
XPHY_4 vgnd vpwr scs8hd_decap_3
XFILLER_7_20 vpwr vgnd scs8hd_fill_2
XFILLER_7_86 vgnd vpwr scs8hd_decap_12
XFILLER_29_232 vgnd vpwr scs8hd_fill_1
XFILLER_12_154 vgnd vpwr scs8hd_decap_12
XANTENNA__103__A _089_/A vgnd vpwr scs8hd_diode_2
XFILLER_26_202 vgnd vpwr scs8hd_decap_12
XFILLER_32_227 vgnd vpwr scs8hd_decap_6
XFILLER_4_65 vgnd vpwr scs8hd_decap_12
X_181_ _181_/A _179_/X data_out[34] vgnd vpwr scs8hd_nor2_4
XFILLER_14_227 vgnd vpwr scs8hd_decap_6
XFILLER_13_52 vpwr vgnd scs8hd_fill_2
XFILLER_9_220 vgnd vpwr scs8hd_decap_12
XFILLER_11_208 vgnd vpwr scs8hd_decap_12
X_164_ _146_/A _165_/B data_out[45] vgnd vpwr scs8hd_nor2_4
X_095_ _092_/X _096_/B data_out[23] vgnd vpwr scs8hd_nor2_4
XFILLER_1_22 vgnd vpwr scs8hd_decap_4
XANTENNA__111__A _086_/X vgnd vpwr scs8hd_diode_2
XFILLER_28_105 vgnd vpwr scs8hd_decap_12
XFILLER_35_94 vgnd vpwr scs8hd_decap_12
XFILLER_27_171 vgnd vpwr scs8hd_decap_12
XFILLER_19_62 vgnd vpwr scs8hd_decap_3
XFILLER_33_196 vgnd vpwr scs8hd_decap_12
X_147_ _147_/A _147_/B data_out[56] vgnd vpwr scs8hd_nor2_4
XFILLER_31_19 vgnd vpwr scs8hd_fill_1
XANTENNA__106__A _066_/Y vgnd vpwr scs8hd_diode_2
X_078_ _071_/A address[0] address[1] _079_/A vgnd vpwr scs8hd_or3_4
XPHY_169 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_141 vgnd vpwr scs8hd_decap_12
XPHY_158 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_21_52 vpwr vgnd scs8hd_fill_2
XPHY_147 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_136 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_125 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_114 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_0_218 vgnd vpwr scs8hd_decap_12
XPHY_103 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_30_166 vgnd vpwr scs8hd_decap_12
XFILLER_15_196 vgnd vpwr scs8hd_decap_12
XPHY_5 vgnd vpwr scs8hd_decap_3
XFILLER_7_98 vgnd vpwr scs8hd_decap_12
XFILLER_26_19 vpwr vgnd scs8hd_fill_2
XFILLER_21_111 vgnd vpwr scs8hd_decap_8
XFILLER_16_74 vpwr vgnd scs8hd_fill_2
XFILLER_16_41 vgnd vpwr scs8hd_decap_3
XFILLER_12_166 vgnd vpwr scs8hd_decap_12
XANTENNA__103__B _100_/X vgnd vpwr scs8hd_diode_2
XFILLER_27_40 vpwr vgnd scs8hd_fill_2
XANTENNA__114__A address[2] vgnd vpwr scs8hd_diode_2
XFILLER_4_77 vgnd vpwr scs8hd_decap_12
X_180_ _180_/A _179_/X data_out[35] vgnd vpwr scs8hd_nor2_4
XFILLER_1_110 vgnd vpwr scs8hd_decap_12
XANTENNA__109__A _108_/X vgnd vpwr scs8hd_diode_2
XFILLER_9_232 vgnd vpwr scs8hd_fill_1
X_163_ _151_/A _165_/B data_out[46] vgnd vpwr scs8hd_nor2_4
XFILLER_24_52 vpwr vgnd scs8hd_fill_2
X_094_ _093_/X _096_/B vgnd vpwr scs8hd_buf_1
XANTENNA__111__B _112_/B vgnd vpwr scs8hd_diode_2
XFILLER_6_202 vgnd vpwr scs8hd_decap_12
XFILLER_28_117 vgnd vpwr scs8hd_decap_12
XFILLER_19_74 vpwr vgnd scs8hd_fill_2
XFILLER_10_21 vgnd vpwr scs8hd_decap_3
X_146_ _146_/A _147_/B data_out[57] vgnd vpwr scs8hd_nor2_4
XANTENNA__122__A _148_/A vgnd vpwr scs8hd_diode_2
X_077_ _068_/X _176_/A data_out[29] vgnd vpwr scs8hd_nor2_4
XPHY_159 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_148 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_137 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_126 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_115 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_104 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_30_178 vgnd vpwr scs8hd_decap_12
XFILLER_21_75 vgnd vpwr scs8hd_decap_12
XPHY_6 vgnd vpwr scs8hd_decap_3
XANTENNA__117__A _092_/X vgnd vpwr scs8hd_diode_2
XFILLER_30_3 vgnd vpwr scs8hd_decap_3
XFILLER_21_123 vgnd vpwr scs8hd_decap_12
X_129_ _128_/X _134_/B vgnd vpwr scs8hd_buf_1
XFILLER_16_64 vgnd vpwr scs8hd_decap_3
XFILLER_12_178 vgnd vpwr scs8hd_decap_12
XFILLER_8_105 vgnd vpwr scs8hd_decap_12
XFILLER_7_171 vgnd vpwr scs8hd_decap_12
XFILLER_26_215 vgnd vpwr scs8hd_decap_12
XFILLER_27_30 vgnd vpwr scs8hd_decap_4
XANTENNA__130__A _092_/X vgnd vpwr scs8hd_diode_2
XFILLER_4_23 vpwr vgnd scs8hd_fill_2
XFILLER_4_89 vgnd vpwr scs8hd_decap_3
XFILLER_4_141 vgnd vpwr scs8hd_decap_12
XFILLER_13_32 vgnd vpwr scs8hd_decap_4
XANTENNA__125__A _086_/X vgnd vpwr scs8hd_diode_2
X_162_ _144_/A _165_/B data_out[47] vgnd vpwr scs8hd_nor2_4
XFILLER_24_20 vpwr vgnd scs8hd_fill_2
X_093_ _063_/X _064_/X _065_/Y address[3] _093_/X vgnd vpwr scs8hd_or4_4
XFILLER_28_129 vgnd vpwr scs8hd_decap_12
XFILLER_35_63 vgnd vpwr scs8hd_decap_12
X_145_ _151_/A _147_/B data_out[58] vgnd vpwr scs8hd_nor2_4
XFILLER_27_184 vgnd vpwr scs8hd_decap_12
XANTENNA__122__B _148_/B vgnd vpwr scs8hd_diode_2
X_076_ _076_/A _176_/A vgnd vpwr scs8hd_buf_1
XFILLER_33_110 vgnd vpwr scs8hd_decap_12
XPHY_116 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_105 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_154 vgnd vpwr scs8hd_decap_12
XFILLER_21_87 vgnd vpwr scs8hd_decap_12
XPHY_149 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_138 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_15_121 vgnd vpwr scs8hd_fill_1
XPHY_127 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_7 vgnd vpwr scs8hd_decap_3
XFILLER_23_3 vgnd vpwr scs8hd_decap_4
X_128_ _154_/A _148_/B _107_/X address[5] _128_/X vgnd vpwr scs8hd_or4_4
XFILLER_21_135 vgnd vpwr scs8hd_decap_12
XANTENNA__133__A _176_/A vgnd vpwr scs8hd_diode_2
XANTENNA__117__B _116_/X vgnd vpwr scs8hd_diode_2
XFILLER_7_12 vpwr vgnd scs8hd_fill_2
XFILLER_20_190 vgnd vpwr scs8hd_decap_12
XFILLER_16_32 vpwr vgnd scs8hd_fill_2
XFILLER_8_117 vgnd vpwr scs8hd_decap_12
XANTENNA__128__A _154_/A vgnd vpwr scs8hd_diode_2
XFILLER_26_227 vgnd vpwr scs8hd_decap_6
XFILLER_27_53 vpwr vgnd scs8hd_fill_2
XANTENNA__130__B _134_/B vgnd vpwr scs8hd_diode_2
XFILLER_23_208 vgnd vpwr scs8hd_decap_12
XFILLER_13_66 vpwr vgnd scs8hd_fill_2
XFILLER_1_123 vgnd vpwr scs8hd_decap_12
XANTENNA__141__A _180_/A vgnd vpwr scs8hd_diode_2
XANTENNA__125__B _124_/B vgnd vpwr scs8hd_diode_2
X_161_ _161_/A _165_/B vgnd vpwr scs8hd_buf_1
XFILLER_24_32 vgnd vpwr scs8hd_decap_4
XFILLER_6_215 vgnd vpwr scs8hd_decap_12
XFILLER_1_14 vpwr vgnd scs8hd_fill_2
XANTENNA__136__A _147_/A vgnd vpwr scs8hd_diode_2
X_092_ _180_/A _092_/X vgnd vpwr scs8hd_buf_1
XFILLER_35_75 vgnd vpwr scs8hd_decap_12
X_144_ _144_/A _147_/B data_out[59] vgnd vpwr scs8hd_nor2_4
XFILLER_27_196 vgnd vpwr scs8hd_decap_12
XFILLER_19_54 vpwr vgnd scs8hd_fill_2
XANTENNA__122__C _107_/X vgnd vpwr scs8hd_diode_2
X_075_ _071_/A _074_/Y address[1] _076_/A vgnd vpwr scs8hd_or3_4
XFILLER_10_89 vgnd vpwr scs8hd_decap_3
XFILLER_18_141 vgnd vpwr scs8hd_decap_12
XFILLER_18_6 vpwr vgnd scs8hd_fill_2
XFILLER_24_166 vgnd vpwr scs8hd_decap_12
XFILLER_21_99 vgnd vpwr scs8hd_decap_12
XPHY_139 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_128 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_117 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_106 vgnd vpwr scs8hd_tapvpwrvgnd_1
X_127_ _090_/X _124_/B data_out[4] vgnd vpwr scs8hd_nor2_4
XPHY_8 vgnd vpwr scs8hd_decap_3
XFILLER_7_24 vpwr vgnd scs8hd_fill_2
XFILLER_21_147 vgnd vpwr scs8hd_decap_12
XFILLER_32_32 vpwr vgnd scs8hd_fill_2
XANTENNA__144__A _144_/A vgnd vpwr scs8hd_diode_2
XANTENNA__128__B _148_/B vgnd vpwr scs8hd_diode_2
XFILLER_8_129 vgnd vpwr scs8hd_decap_12
XFILLER_7_184 vgnd vpwr scs8hd_decap_12
XFILLER_27_65 vpwr vgnd scs8hd_fill_2
XFILLER_4_14 vpwr vgnd scs8hd_fill_2
XFILLER_4_154 vgnd vpwr scs8hd_decap_12
XFILLER_31_220 vgnd vpwr scs8hd_decap_12
XANTENNA__139__A _148_/A vgnd vpwr scs8hd_diode_2
XFILLER_13_56 vpwr vgnd scs8hd_fill_2
XFILLER_1_135 vgnd vpwr scs8hd_decap_12
XFILLER_13_220 vgnd vpwr scs8hd_decap_12
X_160_ _148_/A _142_/B _107_/X _148_/D _161_/A vgnd vpwr scs8hd_or4_4
X_091_ _090_/X _082_/X data_out[24] vgnd vpwr scs8hd_nor2_4
XFILLER_1_48 vpwr vgnd scs8hd_fill_2
XFILLER_1_37 vpwr vgnd scs8hd_fill_2
XANTENNA__136__B _134_/B vgnd vpwr scs8hd_diode_2
XFILLER_6_227 vgnd vpwr scs8hd_decap_6
XANTENNA__152__A _146_/A vgnd vpwr scs8hd_diode_2
XFILLER_35_87 vgnd vpwr scs8hd_decap_6
XFILLER_35_32 vgnd vpwr scs8hd_decap_12
X_143_ _142_/X _147_/B vgnd vpwr scs8hd_buf_1
XANTENNA__062__A address[4] vgnd vpwr scs8hd_diode_2
XFILLER_19_33 vpwr vgnd scs8hd_fill_2
XFILLER_19_11 vpwr vgnd scs8hd_fill_2
X_074_ address[0] _074_/Y vgnd vpwr scs8hd_inv_8
XFILLER_10_57 vgnd vpwr scs8hd_decap_12
XFILLER_10_46 vpwr vgnd scs8hd_fill_2
XFILLER_3_208 vgnd vpwr scs8hd_decap_12
XFILLER_10_13 vpwr vgnd scs8hd_fill_2
XFILLER_10_35 vpwr vgnd scs8hd_fill_2
XFILLER_33_123 vgnd vpwr scs8hd_decap_12
XANTENNA__147__A _147_/A vgnd vpwr scs8hd_diode_2
XANTENNA__122__D address[5] vgnd vpwr scs8hd_diode_2
XFILLER_24_178 vgnd vpwr scs8hd_decap_12
XFILLER_21_56 vgnd vpwr scs8hd_decap_3
XFILLER_21_12 vpwr vgnd scs8hd_fill_2
XPHY_129 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_118 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_107 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_15_123 vgnd vpwr scs8hd_decap_12
XFILLER_15_101 vgnd vpwr scs8hd_decap_12
X_126_ _089_/A _124_/B data_out[5] vgnd vpwr scs8hd_nor2_4
XPHY_9 vgnd vpwr scs8hd_decap_3
XFILLER_21_159 vgnd vpwr scs8hd_decap_12
XFILLER_16_23 vpwr vgnd scs8hd_fill_2
XFILLER_16_12 vpwr vgnd scs8hd_fill_2
XFILLER_35_218 vgnd vpwr scs8hd_decap_12
XANTENNA__128__C _107_/X vgnd vpwr scs8hd_diode_2
XFILLER_16_78 vgnd vpwr scs8hd_decap_12
XANTENNA__144__B _147_/B vgnd vpwr scs8hd_diode_2
XANTENNA__160__A _148_/A vgnd vpwr scs8hd_diode_2
X_109_ _108_/X _112_/B vgnd vpwr scs8hd_buf_1
XFILLER_7_196 vgnd vpwr scs8hd_decap_12
XANTENNA__070__A address[1] vgnd vpwr scs8hd_diode_2
XFILLER_31_232 vgnd vpwr scs8hd_fill_1
XANTENNA__155__A _155_/A vgnd vpwr scs8hd_diode_2
XANTENNA__139__B _142_/B vgnd vpwr scs8hd_diode_2
XFILLER_4_166 vgnd vpwr scs8hd_decap_12
XANTENNA__065__A address[2] vgnd vpwr scs8hd_diode_2
XFILLER_1_147 vgnd vpwr scs8hd_decap_12
XFILLER_13_232 vgnd vpwr scs8hd_fill_1
XFILLER_0_180 vgnd vpwr scs8hd_decap_6
XFILLER_24_89 vgnd vpwr scs8hd_decap_3
XFILLER_24_56 vpwr vgnd scs8hd_fill_2
X_090_ _171_/A _090_/X vgnd vpwr scs8hd_buf_1
XFILLER_10_202 vgnd vpwr scs8hd_decap_12
XFILLER_6_3 vpwr vgnd scs8hd_fill_2
XANTENNA__152__B _149_/X vgnd vpwr scs8hd_diode_2
XFILLER_35_44 vgnd vpwr scs8hd_decap_12
XFILLER_27_121 vgnd vpwr scs8hd_fill_1
X_142_ _154_/A _142_/B _063_/X _148_/D _142_/X vgnd vpwr scs8hd_or4_4
XFILLER_19_78 vgnd vpwr scs8hd_decap_12
XFILLER_10_69 vgnd vpwr scs8hd_decap_12
XFILLER_33_135 vgnd vpwr scs8hd_decap_12
XANTENNA__147__B _147_/B vgnd vpwr scs8hd_diode_2
XANTENNA__163__A _151_/A vgnd vpwr scs8hd_diode_2
XFILLER_18_154 vgnd vpwr scs8hd_decap_12
X_073_ _068_/X _181_/A data_out[30] vgnd vpwr scs8hd_nor2_4
XFILLER_32_190 vgnd vpwr scs8hd_decap_12
XFILLER_21_35 vpwr vgnd scs8hd_fill_2
XANTENNA__073__A _068_/X vgnd vpwr scs8hd_diode_2
XPHY_119 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_108 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_30_105 vgnd vpwr scs8hd_decap_12
XFILLER_15_135 vgnd vpwr scs8hd_decap_12
XFILLER_15_113 vgnd vpwr scs8hd_decap_8
X_125_ _086_/X _124_/B data_out[6] vgnd vpwr scs8hd_nor2_4
XFILLER_7_37 vpwr vgnd scs8hd_fill_2
XFILLER_7_59 vpwr vgnd scs8hd_fill_2
XANTENNA__158__A _146_/A vgnd vpwr scs8hd_diode_2
XFILLER_14_190 vgnd vpwr scs8hd_decap_12
XFILLER_32_89 vgnd vpwr scs8hd_decap_3
XFILLER_32_23 vgnd vpwr scs8hd_decap_8
XANTENNA__068__A _067_/X vgnd vpwr scs8hd_diode_2
XFILLER_16_46 vpwr vgnd scs8hd_fill_2
XFILLER_12_105 vgnd vpwr scs8hd_decap_12
XANTENNA__160__B _142_/B vgnd vpwr scs8hd_diode_2
XANTENNA__128__D address[5] vgnd vpwr scs8hd_diode_2
X_108_ _148_/A _142_/B _107_/X _064_/X _108_/X vgnd vpwr scs8hd_or4_4
XFILLER_11_171 vgnd vpwr scs8hd_decap_12
XFILLER_27_12 vpwr vgnd scs8hd_fill_2
XFILLER_17_208 vgnd vpwr scs8hd_decap_12
XANTENNA__139__C _063_/X vgnd vpwr scs8hd_diode_2
XFILLER_4_27 vpwr vgnd scs8hd_fill_2
XFILLER_4_178 vgnd vpwr scs8hd_decap_12
XANTENNA__171__A _171_/A vgnd vpwr scs8hd_diode_2
XFILLER_13_36 vgnd vpwr scs8hd_fill_1
XANTENNA__081__A _063_/X vgnd vpwr scs8hd_diode_2
XFILLER_1_159 vgnd vpwr scs8hd_decap_12
XANTENNA__166__A _154_/A vgnd vpwr scs8hd_diode_2
XFILLER_24_24 vgnd vpwr scs8hd_decap_4
XANTENNA__076__A _076_/A vgnd vpwr scs8hd_diode_2
XFILLER_35_56 vgnd vpwr scs8hd_decap_6
XFILLER_19_24 vpwr vgnd scs8hd_fill_2
XFILLER_10_26 vpwr vgnd scs8hd_fill_2
XFILLER_33_147 vgnd vpwr scs8hd_decap_12
X_141_ _180_/A _144_/A vgnd vpwr scs8hd_buf_1
XFILLER_18_166 vgnd vpwr scs8hd_decap_12
X_072_ _071_/X _181_/A vgnd vpwr scs8hd_buf_1
XANTENNA__163__B _165_/B vgnd vpwr scs8hd_diode_2
XFILLER_2_93 vgnd vpwr scs8hd_decap_12
XPHY_109 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_30_117 vgnd vpwr scs8hd_decap_12
XANTENNA__073__B _181_/A vgnd vpwr scs8hd_diode_2
XFILLER_15_147 vgnd vpwr scs8hd_decap_12
X_124_ _092_/X _124_/B data_out[7] vgnd vpwr scs8hd_nor2_4
XFILLER_7_16 vpwr vgnd scs8hd_fill_2
XANTENNA__158__B _155_/X vgnd vpwr scs8hd_diode_2
XANTENNA__174__A _144_/A vgnd vpwr scs8hd_diode_2
XFILLER_32_57 vgnd vpwr scs8hd_decap_12
XFILLER_32_46 vgnd vpwr scs8hd_decap_8
XFILLER_32_13 vgnd vpwr scs8hd_decap_8
XFILLER_16_36 vpwr vgnd scs8hd_fill_2
XFILLER_12_117 vgnd vpwr scs8hd_decap_12
XANTENNA__084__A _083_/X vgnd vpwr scs8hd_diode_2
X_107_ address[4] _107_/X vgnd vpwr scs8hd_buf_1
XANTENNA__160__C _107_/X vgnd vpwr scs8hd_diode_2
XFILLER_7_110 vgnd vpwr scs8hd_decap_12
XFILLER_27_57 vpwr vgnd scs8hd_fill_2
XANTENNA__169__A _151_/A vgnd vpwr scs8hd_diode_2
XANTENNA__079__A _079_/A vgnd vpwr scs8hd_diode_2
XANTENNA__139__D _148_/D vgnd vpwr scs8hd_diode_2
XFILLER_25_220 vgnd vpwr scs8hd_decap_12
XANTENNA__171__B _167_/X vgnd vpwr scs8hd_diode_2
XFILLER_13_15 vpwr vgnd scs8hd_fill_2
XANTENNA__081__B _064_/X vgnd vpwr scs8hd_diode_2
XANTENNA__166__B _142_/B vgnd vpwr scs8hd_diode_2
XANTENNA__182__A _176_/A vgnd vpwr scs8hd_diode_2
XFILLER_24_69 vgnd vpwr scs8hd_decap_12
XFILLER_24_36 vgnd vpwr scs8hd_fill_1
XFILLER_10_215 vgnd vpwr scs8hd_decap_12
XANTENNA__092__A _180_/A vgnd vpwr scs8hd_diode_2
XFILLER_1_18 vpwr vgnd scs8hd_fill_2
XFILLER_19_58 vgnd vpwr scs8hd_decap_3
XANTENNA__177__A _171_/A vgnd vpwr scs8hd_diode_2
X_140_ _147_/A _139_/X data_out[60] vgnd vpwr scs8hd_nor2_4
XFILLER_27_123 vgnd vpwr scs8hd_decap_12
X_071_ _071_/A address[0] _071_/C _071_/X vgnd vpwr scs8hd_or3_4
XANTENNA__087__A _086_/X vgnd vpwr scs8hd_diode_2
XFILLER_33_159 vgnd vpwr scs8hd_decap_12
XFILLER_18_178 vgnd vpwr scs8hd_decap_12
XPHY_90 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_30_129 vgnd vpwr scs8hd_decap_12
XFILLER_15_159 vgnd vpwr scs8hd_decap_12
XANTENNA__174__B _174_/B vgnd vpwr scs8hd_diode_2
X_123_ _122_/X _124_/B vgnd vpwr scs8hd_buf_1
XFILLER_32_69 vgnd vpwr scs8hd_decap_12
XFILLER_32_36 vgnd vpwr scs8hd_fill_1
XFILLER_16_59 vgnd vpwr scs8hd_decap_3
XFILLER_12_129 vgnd vpwr scs8hd_decap_12
XANTENNA__160__D _148_/D vgnd vpwr scs8hd_diode_2
XFILLER_22_91 vgnd vpwr scs8hd_fill_1
X_106_ _066_/Y _142_/B vgnd vpwr scs8hd_buf_1
XFILLER_11_184 vgnd vpwr scs8hd_decap_12
XANTENNA__169__B _167_/X vgnd vpwr scs8hd_diode_2
XFILLER_8_93 vgnd vpwr scs8hd_decap_12
XFILLER_27_69 vgnd vpwr scs8hd_decap_12
XFILLER_27_36 vpwr vgnd scs8hd_fill_2
XFILLER_25_232 vgnd vpwr scs8hd_fill_1
XANTENNA__095__A _092_/X vgnd vpwr scs8hd_diode_2
XFILLER_4_18 vgnd vpwr scs8hd_decap_3
XFILLER_22_202 vgnd vpwr scs8hd_decap_12
XANTENNA__081__C address[2] vgnd vpwr scs8hd_diode_2
XANTENNA__166__C _107_/X vgnd vpwr scs8hd_diode_2
XFILLER_24_48 vpwr vgnd scs8hd_fill_2
XANTENNA__182__B _179_/X vgnd vpwr scs8hd_diode_2
XFILLER_10_227 vgnd vpwr scs8hd_decap_6
XFILLER_14_81 vgnd vpwr scs8hd_decap_8
XFILLER_5_220 vgnd vpwr scs8hd_decap_12
XFILLER_30_80 vgnd vpwr scs8hd_decap_12
XANTENNA__177__B _174_/B vgnd vpwr scs8hd_diode_2
XFILLER_10_39 vpwr vgnd scs8hd_fill_2
XFILLER_10_17 vpwr vgnd scs8hd_fill_2
XFILLER_27_135 vgnd vpwr scs8hd_decap_12
XFILLER_19_37 vpwr vgnd scs8hd_fill_2
XANTENNA__087__B _082_/X vgnd vpwr scs8hd_diode_2
X_070_ address[1] _071_/C vgnd vpwr scs8hd_inv_8
XFILLER_4_3 vpwr vgnd scs8hd_fill_2
XFILLER_26_190 vgnd vpwr scs8hd_decap_12
XFILLER_25_80 vgnd vpwr scs8hd_decap_12
XPHY_80 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_91 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_105 vgnd vpwr scs8hd_decap_12
XFILLER_21_16 vpwr vgnd scs8hd_fill_2
XANTENNA__098__A _090_/X vgnd vpwr scs8hd_diode_2
XFILLER_23_171 vgnd vpwr scs8hd_decap_12
XFILLER_23_9 vpwr vgnd scs8hd_fill_2
X_122_ _148_/A _148_/B _107_/X address[5] _122_/X vgnd vpwr scs8hd_or4_4
XFILLER_29_208 vgnd vpwr scs8hd_decap_12
XFILLER_21_119 vgnd vpwr scs8hd_decap_3
XFILLER_20_141 vgnd vpwr scs8hd_decap_12
XFILLER_16_27 vpwr vgnd scs8hd_fill_2
XFILLER_16_16 vpwr vgnd scs8hd_fill_2
X_105_ _065_/Y _148_/A vgnd vpwr scs8hd_buf_1
XFILLER_11_196 vgnd vpwr scs8hd_decap_12
XFILLER_7_123 vgnd vpwr scs8hd_decap_12
XANTENNA__095__B _096_/B vgnd vpwr scs8hd_diode_2
XANTENNA__081__D _066_/Y vgnd vpwr scs8hd_diode_2
XFILLER_13_39 vpwr vgnd scs8hd_fill_2
XANTENNA__166__D _148_/D vgnd vpwr scs8hd_diode_2
XFILLER_24_16 vpwr vgnd scs8hd_fill_2
XFILLER_5_62 vgnd vpwr scs8hd_decap_12
XFILLER_14_93 vgnd vpwr scs8hd_decap_12
XFILLER_5_232 vgnd vpwr scs8hd_fill_1
XFILLER_35_180 vgnd vpwr scs8hd_decap_6
XFILLER_27_147 vgnd vpwr scs8hd_decap_12
XFILLER_2_202 vgnd vpwr scs8hd_decap_12
XPHY_70 vgnd vpwr scs8hd_decap_3
XFILLER_25_92 vgnd vpwr scs8hd_decap_12
XPHY_81 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_92 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_117 vgnd vpwr scs8hd_decap_12
XFILLER_21_39 vpwr vgnd scs8hd_fill_2
XFILLER_2_41 vgnd vpwr scs8hd_decap_12
X_121_ address[3] _148_/B vgnd vpwr scs8hd_buf_1
XFILLER_11_50 vpwr vgnd scs8hd_fill_2
XANTENNA__098__B _096_/B vgnd vpwr scs8hd_diode_2
XFILLER_22_93 vgnd vpwr scs8hd_decap_12
XFILLER_22_71 vgnd vpwr scs8hd_decap_12
XFILLER_19_220 vgnd vpwr scs8hd_decap_12
XFILLER_14_6 vpwr vgnd scs8hd_fill_2
X_104_ _090_/X _100_/X data_out[16] vgnd vpwr scs8hd_nor2_4
XFILLER_7_135 vgnd vpwr scs8hd_decap_12
XFILLER_27_16 vgnd vpwr scs8hd_decap_3
XFILLER_4_105 vgnd vpwr scs8hd_decap_12
XFILLER_6_190 vgnd vpwr scs8hd_decap_12
XFILLER_17_82 vpwr vgnd scs8hd_fill_2
XFILLER_17_71 vpwr vgnd scs8hd_fill_2
XFILLER_22_215 vgnd vpwr scs8hd_decap_12
XFILLER_12_3 vpwr vgnd scs8hd_fill_2
XFILLER_3_171 vgnd vpwr scs8hd_decap_12
XFILLER_9_208 vgnd vpwr scs8hd_decap_12
XFILLER_28_81 vgnd vpwr scs8hd_decap_8
XFILLER_5_30 vpwr vgnd scs8hd_fill_2
XFILLER_5_41 vpwr vgnd scs8hd_fill_2
XFILLER_5_74 vgnd vpwr scs8hd_decap_12
XFILLER_24_28 vgnd vpwr scs8hd_fill_1
XFILLER_30_93 vgnd vpwr scs8hd_decap_12
XFILLER_27_159 vgnd vpwr scs8hd_decap_12
XFILLER_19_28 vgnd vpwr scs8hd_decap_3
XPHY_71 vgnd vpwr scs8hd_decap_3
XPHY_60 vgnd vpwr scs8hd_decap_3
XFILLER_25_60 vgnd vpwr scs8hd_fill_1
XPHY_82 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_93 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_129 vgnd vpwr scs8hd_decap_12
XFILLER_21_29 vgnd vpwr scs8hd_decap_4
XFILLER_2_53 vgnd vpwr scs8hd_decap_12
XFILLER_23_184 vgnd vpwr scs8hd_decap_12
XFILLER_11_62 vgnd vpwr scs8hd_decap_12
X_120_ _090_/X _116_/X data_out[8] vgnd vpwr scs8hd_nor2_4
XFILLER_20_154 vgnd vpwr scs8hd_decap_12
XFILLER_34_202 vgnd vpwr scs8hd_decap_12
XFILLER_22_83 vgnd vpwr scs8hd_decap_8
XFILLER_19_232 vgnd vpwr scs8hd_fill_1
XFILLER_11_110 vgnd vpwr scs8hd_decap_12
XFILLER_7_147 vgnd vpwr scs8hd_decap_12
X_103_ _089_/A _100_/X data_out[17] vgnd vpwr scs8hd_nor2_4
XFILLER_8_30 vgnd vpwr scs8hd_fill_1
XFILLER_8_41 vgnd vpwr scs8hd_decap_8
XFILLER_8_52 vgnd vpwr scs8hd_decap_12
XFILLER_16_202 vgnd vpwr scs8hd_decap_12
XFILLER_4_117 vgnd vpwr scs8hd_decap_12
XFILLER_22_227 vgnd vpwr scs8hd_decap_6
XFILLER_13_19 vpwr vgnd scs8hd_fill_2
XFILLER_28_93 vgnd vpwr scs8hd_decap_12
XFILLER_5_86 vgnd vpwr scs8hd_decap_12
XANTENNA__101__A _092_/X vgnd vpwr scs8hd_diode_2
XFILLER_27_105 vgnd vpwr scs8hd_decap_12
XPHY_61 vgnd vpwr scs8hd_decap_3
XPHY_50 vgnd vpwr scs8hd_decap_3
XFILLER_18_105 vgnd vpwr scs8hd_decap_12
XPHY_83 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_72 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_2_215 vgnd vpwr scs8hd_decap_12
XPHY_94 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_32_141 vgnd vpwr scs8hd_decap_12
XFILLER_17_171 vgnd vpwr scs8hd_decap_12
XFILLER_2_65 vgnd vpwr scs8hd_decap_12
XFILLER_23_196 vgnd vpwr scs8hd_decap_12
X_179_ _178_/X _179_/X vgnd vpwr scs8hd_buf_1
XFILLER_14_141 vgnd vpwr scs8hd_decap_12
XFILLER_11_74 vgnd vpwr scs8hd_decap_12
XFILLER_2_3 vgnd vpwr scs8hd_decap_3
XFILLER_35_3 vpwr vgnd scs8hd_fill_2
XFILLER_20_166 vgnd vpwr scs8hd_decap_12
XFILLER_7_159 vgnd vpwr scs8hd_decap_12
X_102_ _086_/X _100_/X data_out[18] vgnd vpwr scs8hd_nor2_4
XFILLER_8_20 vgnd vpwr scs8hd_decap_4
XFILLER_8_64 vgnd vpwr scs8hd_decap_12
XFILLER_4_129 vgnd vpwr scs8hd_decap_12
XFILLER_3_184 vgnd vpwr scs8hd_decap_12
XANTENNA__104__A _090_/X vgnd vpwr scs8hd_diode_2
XFILLER_0_187 vgnd vpwr scs8hd_decap_12
XFILLER_5_98 vgnd vpwr scs8hd_decap_12
XFILLER_14_52 vpwr vgnd scs8hd_fill_2
XFILLER_27_117 vgnd vpwr scs8hd_decap_4
XANTENNA__101__B _100_/X vgnd vpwr scs8hd_diode_2
XFILLER_18_117 vgnd vpwr scs8hd_decap_12
XFILLER_2_227 vgnd vpwr scs8hd_decap_6
XPHY_62 vgnd vpwr scs8hd_decap_3
XPHY_51 vgnd vpwr scs8hd_decap_3
XPHY_40 vgnd vpwr scs8hd_decap_3
XFILLER_2_77 vgnd vpwr scs8hd_decap_12
XPHY_73 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_84 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_95 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__112__A _089_/A vgnd vpwr scs8hd_diode_2
XANTENNA__107__A address[4] vgnd vpwr scs8hd_diode_2
XFILLER_11_86 vgnd vpwr scs8hd_decap_12
X_178_ _154_/A _148_/B address[4] _138_/A _178_/X vgnd vpwr scs8hd_or4_4
XFILLER_20_178 vgnd vpwr scs8hd_decap_12
XFILLER_22_63 vpwr vgnd scs8hd_fill_2
XFILLER_22_52 vpwr vgnd scs8hd_fill_2
XFILLER_22_41 vpwr vgnd scs8hd_fill_2
XFILLER_11_123 vgnd vpwr scs8hd_decap_12
X_101_ _092_/X _100_/X data_out[19] vgnd vpwr scs8hd_nor2_4
XFILLER_34_215 vgnd vpwr scs8hd_decap_12
XFILLER_8_76 vgnd vpwr scs8hd_decap_12
XFILLER_33_62 vgnd vpwr scs8hd_decap_12
XFILLER_17_52 vpwr vgnd scs8hd_fill_2
XFILLER_17_41 vpwr vgnd scs8hd_fill_2
XFILLER_17_30 vpwr vgnd scs8hd_fill_2
XFILLER_16_215 vgnd vpwr scs8hd_decap_12
XANTENNA__120__A _090_/X vgnd vpwr scs8hd_diode_2
XFILLER_3_196 vgnd vpwr scs8hd_decap_12
XANTENNA__104__B _100_/X vgnd vpwr scs8hd_diode_2
XFILLER_0_199 vgnd vpwr scs8hd_decap_12
XANTENNA__115__A _154_/A vgnd vpwr scs8hd_diode_2
XFILLER_10_3 vgnd vpwr scs8hd_fill_1
XFILLER_30_52 vpwr vgnd scs8hd_fill_2
XFILLER_30_41 vgnd vpwr scs8hd_decap_3
XFILLER_35_19 vgnd vpwr scs8hd_decap_12
XPHY_63 vgnd vpwr scs8hd_decap_3
XPHY_52 vgnd vpwr scs8hd_decap_3
XFILLER_25_52 vpwr vgnd scs8hd_fill_2
XPHY_41 vgnd vpwr scs8hd_decap_3
XFILLER_18_129 vgnd vpwr scs8hd_decap_12
XPHY_30 vgnd vpwr scs8hd_decap_3
XFILLER_2_23 vpwr vgnd scs8hd_fill_2
XPHY_74 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_2_89 vgnd vpwr scs8hd_decap_3
XPHY_85 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__112__B _112_/B vgnd vpwr scs8hd_diode_2
XPHY_96 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_32_154 vgnd vpwr scs8hd_decap_12
XFILLER_17_184 vgnd vpwr scs8hd_decap_12
XFILLER_14_154 vgnd vpwr scs8hd_decap_12
XFILLER_11_98 vgnd vpwr scs8hd_decap_12
XFILLER_11_54 vpwr vgnd scs8hd_fill_2
XFILLER_11_21 vgnd vpwr scs8hd_decap_3
X_177_ _171_/A _174_/B data_out[36] vgnd vpwr scs8hd_nor2_4
XANTENNA__123__A _122_/X vgnd vpwr scs8hd_diode_2
XFILLER_28_202 vgnd vpwr scs8hd_decap_12
XFILLER_11_135 vgnd vpwr scs8hd_decap_12
X_100_ _099_/X _100_/X vgnd vpwr scs8hd_buf_1
XFILLER_34_227 vgnd vpwr scs8hd_decap_6
XFILLER_10_190 vgnd vpwr scs8hd_decap_12
XANTENNA__118__A _086_/X vgnd vpwr scs8hd_diode_2
XFILLER_8_88 vgnd vpwr scs8hd_decap_4
XPHY_200 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_33_74 vgnd vpwr scs8hd_decap_12
XFILLER_33_30 vpwr vgnd scs8hd_fill_2
XFILLER_31_208 vgnd vpwr scs8hd_decap_12
XFILLER_17_86 vgnd vpwr scs8hd_decap_12
XFILLER_17_75 vpwr vgnd scs8hd_fill_2
XFILLER_16_227 vgnd vpwr scs8hd_decap_6
XANTENNA__120__B _116_/X vgnd vpwr scs8hd_diode_2
XFILLER_28_52 vpwr vgnd scs8hd_fill_2
XFILLER_13_208 vgnd vpwr scs8hd_decap_12
XFILLER_0_156 vgnd vpwr scs8hd_decap_12
XANTENNA__115__B _142_/B vgnd vpwr scs8hd_diode_2
XANTENNA__131__A _181_/A vgnd vpwr scs8hd_diode_2
XFILLER_5_34 vpwr vgnd scs8hd_fill_2
XFILLER_5_45 vgnd vpwr scs8hd_decap_12
XFILLER_14_10 vpwr vgnd scs8hd_fill_2
XFILLER_29_171 vgnd vpwr scs8hd_decap_12
XANTENNA__126__A _089_/A vgnd vpwr scs8hd_diode_2
XPHY_64 vgnd vpwr scs8hd_decap_3
XPHY_53 vgnd vpwr scs8hd_decap_3
XFILLER_26_141 vgnd vpwr scs8hd_decap_12
XFILLER_25_31 vpwr vgnd scs8hd_fill_2
XPHY_42 vgnd vpwr scs8hd_decap_3
XPHY_31 vgnd vpwr scs8hd_decap_3
XPHY_75 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_86 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_97 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_20 vgnd vpwr scs8hd_decap_3
XFILLER_32_166 vgnd vpwr scs8hd_decap_12
XFILLER_17_196 vgnd vpwr scs8hd_decap_12
XFILLER_23_111 vgnd vpwr scs8hd_decap_8
XFILLER_11_33 vpwr vgnd scs8hd_fill_2
X_176_ _176_/A _174_/B data_out[37] vgnd vpwr scs8hd_nor2_4
XFILLER_14_166 vgnd vpwr scs8hd_decap_12
XFILLER_22_21 vpwr vgnd scs8hd_fill_2
XFILLER_11_147 vgnd vpwr scs8hd_decap_12
XFILLER_0_3 vgnd vpwr scs8hd_decap_3
XANTENNA__118__B _116_/X vgnd vpwr scs8hd_diode_2
XFILLER_8_12 vpwr vgnd scs8hd_fill_2
X_159_ _147_/A _155_/X data_out[48] vgnd vpwr scs8hd_nor2_4
XANTENNA__134__A _146_/A vgnd vpwr scs8hd_diode_2
XPHY_201 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_33_86 vgnd vpwr scs8hd_decap_12
XFILLER_33_20 vgnd vpwr scs8hd_fill_1
XFILLER_17_98 vgnd vpwr scs8hd_decap_12
XFILLER_3_110 vgnd vpwr scs8hd_decap_12
XANTENNA__129__A _128_/X vgnd vpwr scs8hd_diode_2
XFILLER_28_20 vgnd vpwr scs8hd_decap_4
XFILLER_21_220 vgnd vpwr scs8hd_decap_12
XFILLER_0_168 vgnd vpwr scs8hd_decap_12
XANTENNA__115__C _107_/X vgnd vpwr scs8hd_diode_2
XFILLER_5_13 vpwr vgnd scs8hd_fill_2
XFILLER_5_57 vgnd vpwr scs8hd_decap_4
XFILLER_8_202 vgnd vpwr scs8hd_decap_12
XANTENNA__142__A _154_/A vgnd vpwr scs8hd_diode_2
XANTENNA__126__B _124_/B vgnd vpwr scs8hd_diode_2
XPHY_65 vgnd vpwr scs8hd_decap_3
XPHY_54 vgnd vpwr scs8hd_decap_3
XFILLER_25_76 vpwr vgnd scs8hd_fill_2
XFILLER_25_65 vpwr vgnd scs8hd_fill_2
XPHY_43 vgnd vpwr scs8hd_decap_3
XPHY_32 vgnd vpwr scs8hd_decap_3
XPHY_21 vgnd vpwr scs8hd_decap_3
XPHY_76 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_87 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_10 vgnd vpwr scs8hd_decap_3
XPHY_98 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_32_178 vgnd vpwr scs8hd_decap_12
XANTENNA__137__A address[5] vgnd vpwr scs8hd_diode_2
XFILLER_23_123 vgnd vpwr scs8hd_decap_12
XFILLER_35_7 vgnd vpwr scs8hd_decap_12
X_175_ _181_/A _174_/B data_out[38] vgnd vpwr scs8hd_nor2_4
XFILLER_14_178 vgnd vpwr scs8hd_decap_12
XFILLER_28_215 vgnd vpwr scs8hd_decap_12
XFILLER_9_171 vgnd vpwr scs8hd_decap_12
XFILLER_11_159 vgnd vpwr scs8hd_decap_12
XANTENNA__150__A _144_/A vgnd vpwr scs8hd_diode_2
X_158_ _146_/A _155_/X data_out[49] vgnd vpwr scs8hd_nor2_4
XFILLER_26_3 vpwr vgnd scs8hd_fill_2
X_089_ _089_/A _082_/X data_out[25] vgnd vpwr scs8hd_nor2_4
XFILLER_6_141 vgnd vpwr scs8hd_decap_12
XANTENNA__134__B _134_/B vgnd vpwr scs8hd_diode_2
XPHY_202 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_33_98 vgnd vpwr scs8hd_decap_12
XANTENNA__145__A _151_/A vgnd vpwr scs8hd_diode_2
XFILLER_21_232 vgnd vpwr scs8hd_fill_1
XANTENNA__115__D _064_/X vgnd vpwr scs8hd_diode_2
XFILLER_0_125 vgnd vpwr scs8hd_decap_12
XFILLER_29_184 vgnd vpwr scs8hd_decap_12
XFILLER_14_89 vgnd vpwr scs8hd_decap_3
XFILLER_14_56 vpwr vgnd scs8hd_fill_2
XFILLER_14_23 vpwr vgnd scs8hd_fill_2
XFILLER_35_187 vgnd vpwr scs8hd_decap_12
XANTENNA__142__B _142_/B vgnd vpwr scs8hd_diode_2
XPHY_66 vgnd vpwr scs8hd_decap_3
XPHY_55 vgnd vpwr scs8hd_decap_3
XFILLER_26_154 vgnd vpwr scs8hd_decap_12
XPHY_44 vgnd vpwr scs8hd_decap_3
XPHY_33 vgnd vpwr scs8hd_decap_3
XPHY_22 vgnd vpwr scs8hd_decap_3
XPHY_77 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_88 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_11 vgnd vpwr scs8hd_decap_3
XPHY_99 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_17_110 vgnd vpwr scs8hd_decap_12
XFILLER_2_15 vpwr vgnd scs8hd_fill_2
XFILLER_1_220 vgnd vpwr scs8hd_decap_12
XANTENNA__153__A _147_/A vgnd vpwr scs8hd_diode_2
XANTENNA__063__A _063_/A vgnd vpwr scs8hd_diode_2
XFILLER_23_135 vgnd vpwr scs8hd_decap_12
XFILLER_11_13 vpwr vgnd scs8hd_fill_2
X_174_ _144_/A _174_/B data_out[39] vgnd vpwr scs8hd_nor2_4
XFILLER_22_190 vgnd vpwr scs8hd_decap_12
XANTENNA__148__A _148_/A vgnd vpwr scs8hd_diode_2
XFILLER_20_105 vgnd vpwr scs8hd_decap_12
XFILLER_28_227 vgnd vpwr scs8hd_decap_6
XFILLER_22_67 vpwr vgnd scs8hd_fill_2
XFILLER_22_56 vgnd vpwr scs8hd_decap_4
XANTENNA__150__B _149_/X vgnd vpwr scs8hd_diode_2
X_157_ _151_/A _155_/X data_out[50] vgnd vpwr scs8hd_nor2_4
XFILLER_25_208 vgnd vpwr scs8hd_decap_12
XFILLER_19_3 vgnd vpwr scs8hd_fill_1
X_088_ _176_/A _089_/A vgnd vpwr scs8hd_buf_1
XPHY_203 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_17_56 vgnd vpwr scs8hd_decap_3
XFILLER_17_45 vpwr vgnd scs8hd_fill_2
XFILLER_17_34 vpwr vgnd scs8hd_fill_2
XFILLER_17_12 vpwr vgnd scs8hd_fill_2
XFILLER_3_123 vgnd vpwr scs8hd_decap_12
XANTENNA__145__B _147_/B vgnd vpwr scs8hd_diode_2
XANTENNA__161__A _161_/A vgnd vpwr scs8hd_diode_2
XANTENNA__071__A _071_/A vgnd vpwr scs8hd_diode_2
XFILLER_0_137 vgnd vpwr scs8hd_decap_12
XFILLER_8_215 vgnd vpwr scs8hd_decap_12
XANTENNA__156__A _144_/A vgnd vpwr scs8hd_diode_2
XFILLER_30_56 vgnd vpwr scs8hd_decap_12
XANTENNA__066__A address[3] vgnd vpwr scs8hd_diode_2
XFILLER_14_35 vpwr vgnd scs8hd_fill_2
XFILLER_29_196 vgnd vpwr scs8hd_decap_12
XANTENNA__142__C _063_/X vgnd vpwr scs8hd_diode_2
XFILLER_35_199 vgnd vpwr scs8hd_decap_12
XPHY_12 vgnd vpwr scs8hd_decap_3
XPHY_67 vgnd vpwr scs8hd_decap_3
XPHY_56 vgnd vpwr scs8hd_decap_3
XFILLER_26_166 vgnd vpwr scs8hd_decap_12
XFILLER_25_56 vpwr vgnd scs8hd_fill_2
XPHY_45 vgnd vpwr scs8hd_decap_3
XPHY_34 vgnd vpwr scs8hd_decap_3
XPHY_23 vgnd vpwr scs8hd_decap_3
XFILLER_2_27 vpwr vgnd scs8hd_fill_2
XFILLER_1_232 vgnd vpwr scs8hd_fill_1
XPHY_78 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_89 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__153__B _149_/X vgnd vpwr scs8hd_diode_2
XFILLER_23_147 vgnd vpwr scs8hd_decap_12
X_173_ _172_/X _174_/B vgnd vpwr scs8hd_buf_1
XFILLER_11_58 vgnd vpwr scs8hd_decap_3
XANTENNA__148__B _148_/B vgnd vpwr scs8hd_diode_2
XANTENNA__164__A _146_/A vgnd vpwr scs8hd_diode_2
XFILLER_20_117 vgnd vpwr scs8hd_decap_12
XFILLER_9_184 vgnd vpwr scs8hd_decap_12
XFILLER_22_35 vgnd vpwr scs8hd_decap_4
XANTENNA__074__A address[0] vgnd vpwr scs8hd_diode_2
X_156_ _144_/A _155_/X data_out[51] vgnd vpwr scs8hd_nor2_4
X_087_ _086_/X _082_/X data_out[26] vgnd vpwr scs8hd_nor2_4
XFILLER_6_154 vgnd vpwr scs8hd_decap_12
XFILLER_8_26 vpwr vgnd scs8hd_fill_2
XFILLER_33_220 vgnd vpwr scs8hd_decap_12
XANTENNA__159__A _147_/A vgnd vpwr scs8hd_diode_2
XANTENNA__069__A enable vgnd vpwr scs8hd_diode_2
XPHY_204 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_33_34 vpwr vgnd scs8hd_fill_2
XFILLER_33_12 vpwr vgnd scs8hd_fill_2
XFILLER_15_220 vgnd vpwr scs8hd_decap_12
XFILLER_3_135 vgnd vpwr scs8hd_decap_12
XFILLER_31_3 vpwr vgnd scs8hd_fill_2
X_139_ _148_/A _142_/B _063_/X _148_/D _139_/X vgnd vpwr scs8hd_or4_4
XFILLER_2_190 vgnd vpwr scs8hd_decap_12
XFILLER_28_89 vgnd vpwr scs8hd_decap_3
XFILLER_28_56 vpwr vgnd scs8hd_fill_2
XFILLER_28_12 vpwr vgnd scs8hd_fill_2
XANTENNA__071__B address[0] vgnd vpwr scs8hd_diode_2
XFILLER_0_149 vgnd vpwr scs8hd_decap_6
XFILLER_8_227 vgnd vpwr scs8hd_decap_6
XANTENNA__156__B _155_/X vgnd vpwr scs8hd_diode_2
XANTENNA__172__A _148_/A vgnd vpwr scs8hd_diode_2
XFILLER_30_68 vgnd vpwr scs8hd_decap_12
XFILLER_30_46 vgnd vpwr scs8hd_decap_3
XFILLER_30_24 vgnd vpwr scs8hd_decap_4
XANTENNA__082__A _081_/X vgnd vpwr scs8hd_diode_2
XFILLER_14_69 vgnd vpwr scs8hd_decap_12
XFILLER_5_208 vgnd vpwr scs8hd_decap_12
XANTENNA__142__D _148_/D vgnd vpwr scs8hd_diode_2
XFILLER_35_156 vgnd vpwr scs8hd_decap_12
XANTENNA__167__A _167_/A vgnd vpwr scs8hd_diode_2
XPHY_68 vgnd vpwr scs8hd_decap_3
XPHY_57 vgnd vpwr scs8hd_decap_3
XFILLER_26_178 vgnd vpwr scs8hd_decap_12
XFILLER_25_35 vpwr vgnd scs8hd_fill_2
XPHY_46 vgnd vpwr scs8hd_decap_3
XPHY_35 vgnd vpwr scs8hd_decap_3
XANTENNA__077__A _068_/X vgnd vpwr scs8hd_diode_2
XPHY_24 vgnd vpwr scs8hd_decap_3
XPHY_79 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_13 vgnd vpwr scs8hd_decap_3
XFILLER_9_3 vgnd vpwr scs8hd_fill_1
XFILLER_17_123 vgnd vpwr scs8hd_decap_12
XFILLER_23_159 vgnd vpwr scs8hd_decap_12
XFILLER_11_37 vpwr vgnd scs8hd_fill_2
XANTENNA__148__C _063_/A vgnd vpwr scs8hd_diode_2
XANTENNA__164__B _165_/B vgnd vpwr scs8hd_diode_2
X_172_ _148_/A _148_/B address[4] _138_/A _172_/X vgnd vpwr scs8hd_or4_4
XFILLER_20_129 vgnd vpwr scs8hd_decap_12
XFILLER_22_25 vgnd vpwr scs8hd_decap_4
XANTENNA__180__A _180_/A vgnd vpwr scs8hd_diode_2
XFILLER_9_196 vgnd vpwr scs8hd_decap_12
X_155_ _155_/A _155_/X vgnd vpwr scs8hd_buf_1
XANTENNA__090__A _171_/A vgnd vpwr scs8hd_diode_2
X_086_ _181_/A _086_/X vgnd vpwr scs8hd_buf_1
XFILLER_6_166 vgnd vpwr scs8hd_decap_12
XFILLER_8_16 vpwr vgnd scs8hd_fill_2
XFILLER_33_232 vgnd vpwr scs8hd_fill_1
XANTENNA__159__B _155_/X vgnd vpwr scs8hd_diode_2
XANTENNA__175__A _181_/A vgnd vpwr scs8hd_diode_2
XANTENNA__085__A _082_/X vgnd vpwr scs8hd_diode_2
XFILLER_3_147 vgnd vpwr scs8hd_decap_12
XFILLER_30_202 vgnd vpwr scs8hd_decap_12
X_138_ _138_/A _148_/D vgnd vpwr scs8hd_buf_1
XFILLER_24_3 vpwr vgnd scs8hd_fill_2
XFILLER_15_232 vgnd vpwr scs8hd_fill_1
X_069_ enable _071_/A vgnd vpwr scs8hd_inv_8
XFILLER_28_35 vpwr vgnd scs8hd_fill_2
XANTENNA__071__C _071_/C vgnd vpwr scs8hd_diode_2
XFILLER_0_106 vgnd vpwr scs8hd_decap_12
XFILLER_0_94 vgnd vpwr scs8hd_decap_12
XFILLER_0_61 vgnd vpwr scs8hd_fill_1
XFILLER_12_202 vgnd vpwr scs8hd_decap_12
XFILLER_5_17 vpwr vgnd scs8hd_fill_2
XANTENNA__172__B _148_/B vgnd vpwr scs8hd_diode_2
XFILLER_29_121 vgnd vpwr scs8hd_fill_1
XFILLER_35_168 vgnd vpwr scs8hd_decap_12
XANTENNA__183__A _171_/A vgnd vpwr scs8hd_diode_2
XFILLER_6_93 vgnd vpwr scs8hd_decap_12
XPHY_69 vgnd vpwr scs8hd_decap_3
XFILLER_34_190 vgnd vpwr scs8hd_decap_12
XPHY_58 vgnd vpwr scs8hd_decap_3
XFILLER_25_69 vpwr vgnd scs8hd_fill_2
XFILLER_25_14 vpwr vgnd scs8hd_fill_2
XPHY_47 vgnd vpwr scs8hd_decap_3
XPHY_36 vgnd vpwr scs8hd_decap_3
XANTENNA__093__A _063_/X vgnd vpwr scs8hd_diode_2
XANTENNA__077__B _176_/A vgnd vpwr scs8hd_diode_2
XPHY_25 vgnd vpwr scs8hd_decap_3
XPHY_14 vgnd vpwr scs8hd_decap_3
XFILLER_32_105 vgnd vpwr scs8hd_decap_12
XFILLER_17_135 vgnd vpwr scs8hd_decap_12
XFILLER_31_171 vgnd vpwr scs8hd_decap_12
XANTENNA__178__A _154_/A vgnd vpwr scs8hd_diode_2
XFILLER_16_190 vgnd vpwr scs8hd_decap_12
XANTENNA__088__A _176_/A vgnd vpwr scs8hd_diode_2
XANTENNA__148__D _148_/D vgnd vpwr scs8hd_diode_2
X_171_ _171_/A _167_/X data_out[40] vgnd vpwr scs8hd_nor2_4
XFILLER_14_105 vgnd vpwr scs8hd_decap_12
XANTENNA__180__B _179_/X vgnd vpwr scs8hd_diode_2
XFILLER_13_171 vgnd vpwr scs8hd_decap_12
XFILLER_19_208 vgnd vpwr scs8hd_decap_12
XFILLER_10_141 vgnd vpwr scs8hd_decap_12
X_154_ _154_/A _148_/B _063_/A _148_/D _155_/A vgnd vpwr scs8hd_or4_4
XFILLER_26_7 vgnd vpwr scs8hd_decap_3
XANTENNA__175__B _174_/B vgnd vpwr scs8hd_diode_2
X_085_ _082_/X _180_/A data_out[27] vgnd vpwr scs8hd_nor2_4
XFILLER_6_178 vgnd vpwr scs8hd_decap_12
XFILLER_33_47 vgnd vpwr scs8hd_decap_12
XANTENNA__085__B _180_/A vgnd vpwr scs8hd_diode_2
XFILLER_3_159 vgnd vpwr scs8hd_decap_12
X_137_ address[5] _138_/A vgnd vpwr scs8hd_inv_8
X_068_ _067_/X _068_/X vgnd vpwr scs8hd_buf_1
XFILLER_0_118 vgnd vpwr scs8hd_decap_6
XFILLER_9_71 vgnd vpwr scs8hd_decap_12
XFILLER_28_69 vgnd vpwr scs8hd_decap_12
XFILLER_18_80 vgnd vpwr scs8hd_decap_12
XANTENNA__096__A _086_/X vgnd vpwr scs8hd_diode_2
XANTENNA__172__C address[4] vgnd vpwr scs8hd_diode_2
XFILLER_30_15 vpwr vgnd scs8hd_fill_2
XFILLER_14_27 vpwr vgnd scs8hd_fill_2
XFILLER_35_125 vgnd vpwr scs8hd_decap_12
XANTENNA__183__B _179_/X vgnd vpwr scs8hd_diode_2
XPHY_59 vgnd vpwr scs8hd_decap_3
XFILLER_25_48 vpwr vgnd scs8hd_fill_2
XPHY_48 vgnd vpwr scs8hd_decap_3
XPHY_37 vgnd vpwr scs8hd_decap_3
XANTENNA__093__B _064_/X vgnd vpwr scs8hd_diode_2
XPHY_26 vgnd vpwr scs8hd_decap_3
XPHY_15 vgnd vpwr scs8hd_decap_3
XFILLER_32_117 vgnd vpwr scs8hd_decap_12
XFILLER_17_147 vgnd vpwr scs8hd_decap_12
XFILLER_2_19 vpwr vgnd scs8hd_fill_2
XANTENNA__178__B _148_/B vgnd vpwr scs8hd_diode_2
XFILLER_11_17 vpwr vgnd scs8hd_fill_2
X_170_ _146_/A _167_/X data_out[41] vgnd vpwr scs8hd_nor2_4
XFILLER_14_117 vgnd vpwr scs8hd_decap_12
XFILLER_3_40 vpwr vgnd scs8hd_fill_2
XFILLER_3_51 vgnd vpwr scs8hd_decap_8
XFILLER_3_62 vgnd vpwr scs8hd_decap_12
XFILLER_27_220 vgnd vpwr scs8hd_decap_12
XANTENNA__099__A _063_/X vgnd vpwr scs8hd_diode_2
X_153_ _147_/A _149_/X data_out[52] vgnd vpwr scs8hd_nor2_4
XFILLER_19_7 vpwr vgnd scs8hd_fill_2
XFILLER_12_93 vgnd vpwr scs8hd_decap_12
X_084_ _083_/X _180_/A vgnd vpwr scs8hd_buf_1
XFILLER_33_59 vpwr vgnd scs8hd_fill_2
XFILLER_17_16 vgnd vpwr scs8hd_decap_3
XFILLER_30_215 vgnd vpwr scs8hd_decap_12
X_136_ _147_/A _134_/B data_out[0] vgnd vpwr scs8hd_nor2_4
X_067_ _063_/X _064_/X _065_/Y _066_/Y _067_/X vgnd vpwr scs8hd_or4_4
XFILLER_0_63 vgnd vpwr scs8hd_decap_12
XFILLER_0_41 vgnd vpwr scs8hd_decap_12
XFILLER_9_50 vgnd vpwr scs8hd_decap_4
XFILLER_9_83 vgnd vpwr scs8hd_decap_12
XFILLER_28_26 vgnd vpwr scs8hd_decap_3
XFILLER_12_215 vgnd vpwr scs8hd_decap_12
XANTENNA__096__B _096_/B vgnd vpwr scs8hd_diode_2
XANTENNA__172__D _138_/A vgnd vpwr scs8hd_diode_2
X_119_ _089_/A _116_/X data_out[9] vgnd vpwr scs8hd_nor2_4
XFILLER_29_123 vgnd vpwr scs8hd_decap_12
XFILLER_14_39 vpwr vgnd scs8hd_fill_2
XFILLER_35_137 vgnd vpwr scs8hd_decap_12
XFILLER_20_93 vgnd vpwr scs8hd_decap_12
XFILLER_20_60 vpwr vgnd scs8hd_fill_2
XPHY_49 vgnd vpwr scs8hd_decap_3
XPHY_38 vgnd vpwr scs8hd_decap_3
XPHY_27 vgnd vpwr scs8hd_decap_3
XPHY_16 vgnd vpwr scs8hd_decap_3
XFILLER_32_129 vgnd vpwr scs8hd_decap_12
XFILLER_17_159 vgnd vpwr scs8hd_decap_12
XANTENNA__093__C _065_/Y vgnd vpwr scs8hd_diode_2
XFILLER_31_184 vgnd vpwr scs8hd_decap_12
XFILLER_31_81 vgnd vpwr scs8hd_decap_12
XANTENNA__178__C address[4] vgnd vpwr scs8hd_diode_2
XFILLER_14_129 vgnd vpwr scs8hd_decap_12
XFILLER_13_184 vgnd vpwr scs8hd_decap_12
XFILLER_3_74 vgnd vpwr scs8hd_decap_12
XANTENNA__099__B _064_/X vgnd vpwr scs8hd_diode_2
X_152_ _146_/A _149_/X data_out[53] vgnd vpwr scs8hd_nor2_4
XFILLER_27_232 vgnd vpwr scs8hd_fill_1
X_083_ _071_/A _074_/Y _071_/C _083_/X vgnd vpwr scs8hd_or3_4
XFILLER_10_154 vgnd vpwr scs8hd_decap_12
XFILLER_33_16 vpwr vgnd scs8hd_fill_2
XFILLER_24_202 vgnd vpwr scs8hd_decap_12
XFILLER_30_227 vgnd vpwr scs8hd_decap_6
XFILLER_31_7 vpwr vgnd scs8hd_fill_2
XFILLER_23_71 vpwr vgnd scs8hd_fill_2
X_066_ address[3] _066_/Y vgnd vpwr scs8hd_inv_8
X_135_ _171_/A _147_/A vgnd vpwr scs8hd_buf_1
XFILLER_0_75 vgnd vpwr scs8hd_decap_12
XFILLER_0_53 vgnd vpwr scs8hd_decap_8
XFILLER_9_95 vgnd vpwr scs8hd_decap_12
XFILLER_28_16 vpwr vgnd scs8hd_fill_2
XFILLER_12_227 vgnd vpwr scs8hd_decap_6
XFILLER_34_81 vgnd vpwr scs8hd_decap_8
XFILLER_18_93 vgnd vpwr scs8hd_decap_12
X_118_ _086_/X _116_/X data_out[10] vgnd vpwr scs8hd_nor2_4
XFILLER_7_220 vgnd vpwr scs8hd_decap_12
XFILLER_30_28 vgnd vpwr scs8hd_fill_1
XFILLER_22_3 vgnd vpwr scs8hd_decap_4
XFILLER_29_135 vgnd vpwr scs8hd_decap_12
XFILLER_29_81 vgnd vpwr scs8hd_decap_12
XFILLER_35_149 vgnd vpwr scs8hd_decap_6
XFILLER_28_190 vgnd vpwr scs8hd_decap_12
XFILLER_26_105 vgnd vpwr scs8hd_decap_12
XPHY_28 vgnd vpwr scs8hd_decap_3
XFILLER_6_41 vgnd vpwr scs8hd_decap_12
XPHY_17 vgnd vpwr scs8hd_decap_3
XFILLER_25_171 vgnd vpwr scs8hd_decap_12
XPHY_39 vgnd vpwr scs8hd_decap_3
XANTENNA__093__D address[3] vgnd vpwr scs8hd_diode_2
XFILLER_31_93 vgnd vpwr scs8hd_decap_12
XANTENNA__178__D _138_/A vgnd vpwr scs8hd_diode_2
XFILLER_23_119 vgnd vpwr scs8hd_decap_3
XFILLER_31_196 vgnd vpwr scs8hd_decap_12
XFILLER_22_141 vgnd vpwr scs8hd_decap_12
XFILLER_26_93 vgnd vpwr scs8hd_decap_12
XFILLER_13_196 vgnd vpwr scs8hd_decap_12
XFILLER_9_123 vgnd vpwr scs8hd_decap_12
XFILLER_3_86 vgnd vpwr scs8hd_decap_12
X_151_ _151_/A _149_/X data_out[54] vgnd vpwr scs8hd_nor2_4
XANTENNA__099__C address[2] vgnd vpwr scs8hd_diode_2
X_082_ _081_/X _082_/X vgnd vpwr scs8hd_buf_1
XFILLER_12_62 vgnd vpwr scs8hd_decap_12
XFILLER_10_166 vgnd vpwr scs8hd_decap_12
X_065_ address[2] _065_/Y vgnd vpwr scs8hd_inv_8
XFILLER_0_87 vgnd vpwr scs8hd_decap_6
X_134_ _146_/A _134_/B data_out[1] vgnd vpwr scs8hd_nor2_4
XFILLER_28_39 vpwr vgnd scs8hd_fill_2
XFILLER_34_93 vgnd vpwr scs8hd_decap_12
X_117_ _092_/X _116_/X data_out[11] vgnd vpwr scs8hd_nor2_4
XFILLER_7_232 vgnd vpwr scs8hd_fill_1
XFILLER_29_147 vgnd vpwr scs8hd_decap_12
XFILLER_4_202 vgnd vpwr scs8hd_decap_12
XFILLER_35_106 vgnd vpwr scs8hd_decap_12
XFILLER_29_93 vgnd vpwr scs8hd_decap_12
XFILLER_6_53 vgnd vpwr scs8hd_decap_12
XFILLER_26_117 vgnd vpwr scs8hd_decap_12
XFILLER_25_18 vpwr vgnd scs8hd_fill_2
XPHY_29 vgnd vpwr scs8hd_decap_3
XPHY_18 vgnd vpwr scs8hd_decap_3
XFILLER_31_50 vpwr vgnd scs8hd_fill_2
XFILLER_15_73 vpwr vgnd scs8hd_fill_2
XFILLER_15_51 vpwr vgnd scs8hd_fill_2
XANTENNA__102__A _086_/X vgnd vpwr scs8hd_diode_2
XFILLER_9_135 vgnd vpwr scs8hd_decap_12
XFILLER_3_98 vgnd vpwr scs8hd_decap_12
XFILLER_8_190 vgnd vpwr scs8hd_decap_12
X_150_ _144_/A _149_/X data_out[55] vgnd vpwr scs8hd_nor2_4
X_081_ _063_/X _064_/X address[2] _066_/Y _081_/X vgnd vpwr scs8hd_or4_4
XANTENNA__099__D address[3] vgnd vpwr scs8hd_diode_2
XFILLER_12_74 vgnd vpwr scs8hd_decap_12
XFILLER_12_30 vgnd vpwr scs8hd_fill_1
XFILLER_10_178 vgnd vpwr scs8hd_decap_12
XFILLER_6_105 vgnd vpwr scs8hd_decap_12
XFILLER_5_171 vgnd vpwr scs8hd_decap_12
XFILLER_24_215 vgnd vpwr scs8hd_decap_12
XFILLER_23_40 vpwr vgnd scs8hd_fill_2
X_064_ address[5] _064_/X vgnd vpwr scs8hd_buf_1
X_133_ _176_/A _146_/A vgnd vpwr scs8hd_buf_1
XFILLER_2_141 vgnd vpwr scs8hd_decap_12
XANTENNA__110__A _092_/X vgnd vpwr scs8hd_diode_2
XANTENNA__105__A _065_/Y vgnd vpwr scs8hd_diode_2
X_116_ _115_/X _116_/X vgnd vpwr scs8hd_buf_1
XFILLER_30_19 vgnd vpwr scs8hd_decap_3
XFILLER_29_159 vgnd vpwr scs8hd_decap_12
XFILLER_35_118 vgnd vpwr scs8hd_decap_6
XFILLER_6_65 vgnd vpwr scs8hd_decap_12
XFILLER_26_129 vgnd vpwr scs8hd_decap_12
XPHY_19 vgnd vpwr scs8hd_decap_3
XFILLER_25_184 vgnd vpwr scs8hd_decap_12
XANTENNA__102__B _100_/X vgnd vpwr scs8hd_diode_2
XPHY_190 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_31_121 vgnd vpwr scs8hd_fill_1
XFILLER_22_154 vgnd vpwr scs8hd_decap_12
XFILLER_3_22 vgnd vpwr scs8hd_decap_3
XANTENNA__113__A _090_/X vgnd vpwr scs8hd_diode_2
XFILLER_9_147 vgnd vpwr scs8hd_decap_12
X_080_ _068_/X _171_/A data_out[28] vgnd vpwr scs8hd_nor2_4
XFILLER_6_117 vgnd vpwr scs8hd_decap_12
XANTENNA__108__A _148_/A vgnd vpwr scs8hd_diode_2
XFILLER_18_202 vgnd vpwr scs8hd_decap_12
XFILLER_12_86 vgnd vpwr scs8hd_decap_6
XFILLER_12_53 vgnd vpwr scs8hd_decap_6
XFILLER_5_3 vgnd vpwr scs8hd_fill_1
XFILLER_24_227 vgnd vpwr scs8hd_decap_6
X_063_ _063_/A _063_/X vgnd vpwr scs8hd_buf_1
X_132_ _151_/A _134_/B data_out[2] vgnd vpwr scs8hd_nor2_4
XFILLER_21_208 vgnd vpwr scs8hd_decap_12
XFILLER_0_23 vpwr vgnd scs8hd_fill_2
XANTENNA__110__B _112_/B vgnd vpwr scs8hd_diode_2
XFILLER_9_21 vgnd vpwr scs8hd_decap_3
XFILLER_9_43 vpwr vgnd scs8hd_fill_2
XFILLER_18_63 vpwr vgnd scs8hd_fill_2
XFILLER_18_41 vpwr vgnd scs8hd_fill_2
XANTENNA__121__A address[3] vgnd vpwr scs8hd_diode_2
X_115_ _154_/A _142_/B _107_/X _064_/X _115_/X vgnd vpwr scs8hd_or4_4
XFILLER_29_105 vgnd vpwr scs8hd_decap_12
XFILLER_20_64 vpwr vgnd scs8hd_fill_2
XFILLER_20_53 vpwr vgnd scs8hd_fill_2
XANTENNA__116__A _115_/X vgnd vpwr scs8hd_diode_2
XFILLER_4_215 vgnd vpwr scs8hd_decap_12
XFILLER_34_141 vgnd vpwr scs8hd_decap_12
XFILLER_19_171 vgnd vpwr scs8hd_decap_12
XFILLER_6_77 vgnd vpwr scs8hd_decap_12
XFILLER_25_196 vgnd vpwr scs8hd_decap_12
XPHY_191 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_180 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_16_141 vgnd vpwr scs8hd_decap_12
.ends

