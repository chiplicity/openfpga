VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sb_2__0_
  CLASS BLOCK ;
  FOREIGN sb_2__0_ ;
  ORIGIN 0.000 0.000 ;
  SIZE 140.000 BY 140.000 ;
  PIN ccff_head
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 70.080 140.000 70.680 ;
    END
  END ccff_head
  PIN ccff_tail
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 104.970 0.000 105.250 2.400 ;
    END
  END ccff_tail
  PIN chanx_left_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 19.080 2.400 19.680 ;
    END
  END chanx_left_in[0]
  PIN chanx_left_in[10]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 49.680 2.400 50.280 ;
    END
  END chanx_left_in[10]
  PIN chanx_left_in[11]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 53.080 2.400 53.680 ;
    END
  END chanx_left_in[11]
  PIN chanx_left_in[12]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 55.800 2.400 56.400 ;
    END
  END chanx_left_in[12]
  PIN chanx_left_in[13]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 59.200 2.400 59.800 ;
    END
  END chanx_left_in[13]
  PIN chanx_left_in[14]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 61.920 2.400 62.520 ;
    END
  END chanx_left_in[14]
  PIN chanx_left_in[15]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 65.320 2.400 65.920 ;
    END
  END chanx_left_in[15]
  PIN chanx_left_in[16]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 68.040 2.400 68.640 ;
    END
  END chanx_left_in[16]
  PIN chanx_left_in[17]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 71.440 2.400 72.040 ;
    END
  END chanx_left_in[17]
  PIN chanx_left_in[18]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 74.160 2.400 74.760 ;
    END
  END chanx_left_in[18]
  PIN chanx_left_in[19]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 76.880 2.400 77.480 ;
    END
  END chanx_left_in[19]
  PIN chanx_left_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 22.480 2.400 23.080 ;
    END
  END chanx_left_in[1]
  PIN chanx_left_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 25.200 2.400 25.800 ;
    END
  END chanx_left_in[2]
  PIN chanx_left_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 28.600 2.400 29.200 ;
    END
  END chanx_left_in[3]
  PIN chanx_left_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 31.320 2.400 31.920 ;
    END
  END chanx_left_in[4]
  PIN chanx_left_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 34.720 2.400 35.320 ;
    END
  END chanx_left_in[5]
  PIN chanx_left_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 37.440 2.400 38.040 ;
    END
  END chanx_left_in[6]
  PIN chanx_left_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 40.840 2.400 41.440 ;
    END
  END chanx_left_in[7]
  PIN chanx_left_in[8]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 43.560 2.400 44.160 ;
    END
  END chanx_left_in[8]
  PIN chanx_left_in[9]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 46.960 2.400 47.560 ;
    END
  END chanx_left_in[9]
  PIN chanx_left_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 80.280 2.400 80.880 ;
    END
  END chanx_left_out[0]
  PIN chanx_left_out[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 110.880 2.400 111.480 ;
    END
  END chanx_left_out[10]
  PIN chanx_left_out[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 113.600 2.400 114.200 ;
    END
  END chanx_left_out[11]
  PIN chanx_left_out[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 117.000 2.400 117.600 ;
    END
  END chanx_left_out[12]
  PIN chanx_left_out[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 119.720 2.400 120.320 ;
    END
  END chanx_left_out[13]
  PIN chanx_left_out[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 123.120 2.400 123.720 ;
    END
  END chanx_left_out[14]
  PIN chanx_left_out[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 125.840 2.400 126.440 ;
    END
  END chanx_left_out[15]
  PIN chanx_left_out[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 129.240 2.400 129.840 ;
    END
  END chanx_left_out[16]
  PIN chanx_left_out[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 131.960 2.400 132.560 ;
    END
  END chanx_left_out[17]
  PIN chanx_left_out[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 135.360 2.400 135.960 ;
    END
  END chanx_left_out[18]
  PIN chanx_left_out[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 138.080 2.400 138.680 ;
    END
  END chanx_left_out[19]
  PIN chanx_left_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 83.000 2.400 83.600 ;
    END
  END chanx_left_out[1]
  PIN chanx_left_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 86.400 2.400 87.000 ;
    END
  END chanx_left_out[2]
  PIN chanx_left_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 89.120 2.400 89.720 ;
    END
  END chanx_left_out[3]
  PIN chanx_left_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 92.520 2.400 93.120 ;
    END
  END chanx_left_out[4]
  PIN chanx_left_out[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 95.240 2.400 95.840 ;
    END
  END chanx_left_out[5]
  PIN chanx_left_out[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 98.640 2.400 99.240 ;
    END
  END chanx_left_out[6]
  PIN chanx_left_out[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 101.360 2.400 101.960 ;
    END
  END chanx_left_out[7]
  PIN chanx_left_out[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 104.760 2.400 105.360 ;
    END
  END chanx_left_out[8]
  PIN chanx_left_out[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 107.480 2.400 108.080 ;
    END
  END chanx_left_out[9]
  PIN chany_top_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 24.010 137.600 24.290 140.000 ;
    END
  END chany_top_in[0]
  PIN chany_top_in[10]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 52.530 137.600 52.810 140.000 ;
    END
  END chany_top_in[10]
  PIN chany_top_in[11]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 55.290 137.600 55.570 140.000 ;
    END
  END chany_top_in[11]
  PIN chany_top_in[12]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 58.510 137.600 58.790 140.000 ;
    END
  END chany_top_in[12]
  PIN chany_top_in[13]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 61.270 137.600 61.550 140.000 ;
    END
  END chany_top_in[13]
  PIN chany_top_in[14]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 64.030 137.600 64.310 140.000 ;
    END
  END chany_top_in[14]
  PIN chany_top_in[15]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 66.790 137.600 67.070 140.000 ;
    END
  END chany_top_in[15]
  PIN chany_top_in[16]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 69.550 137.600 69.830 140.000 ;
    END
  END chany_top_in[16]
  PIN chany_top_in[17]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 72.770 137.600 73.050 140.000 ;
    END
  END chany_top_in[17]
  PIN chany_top_in[18]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 75.530 137.600 75.810 140.000 ;
    END
  END chany_top_in[18]
  PIN chany_top_in[19]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 78.290 137.600 78.570 140.000 ;
    END
  END chany_top_in[19]
  PIN chany_top_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 26.770 137.600 27.050 140.000 ;
    END
  END chany_top_in[1]
  PIN chany_top_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 29.990 137.600 30.270 140.000 ;
    END
  END chany_top_in[2]
  PIN chany_top_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 32.750 137.600 33.030 140.000 ;
    END
  END chany_top_in[3]
  PIN chany_top_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 35.510 137.600 35.790 140.000 ;
    END
  END chany_top_in[4]
  PIN chany_top_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 38.270 137.600 38.550 140.000 ;
    END
  END chany_top_in[5]
  PIN chany_top_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 41.030 137.600 41.310 140.000 ;
    END
  END chany_top_in[6]
  PIN chany_top_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 44.250 137.600 44.530 140.000 ;
    END
  END chany_top_in[7]
  PIN chany_top_in[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 47.010 137.600 47.290 140.000 ;
    END
  END chany_top_in[8]
  PIN chany_top_in[9]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 49.770 137.600 50.050 140.000 ;
    END
  END chany_top_in[9]
  PIN chany_top_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 81.050 137.600 81.330 140.000 ;
    END
  END chany_top_out[0]
  PIN chany_top_out[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 109.570 137.600 109.850 140.000 ;
    END
  END chany_top_out[10]
  PIN chany_top_out[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 112.330 137.600 112.610 140.000 ;
    END
  END chany_top_out[11]
  PIN chany_top_out[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 115.550 137.600 115.830 140.000 ;
    END
  END chany_top_out[12]
  PIN chany_top_out[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 118.310 137.600 118.590 140.000 ;
    END
  END chany_top_out[13]
  PIN chany_top_out[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 121.070 137.600 121.350 140.000 ;
    END
  END chany_top_out[14]
  PIN chany_top_out[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 123.830 137.600 124.110 140.000 ;
    END
  END chany_top_out[15]
  PIN chany_top_out[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 126.590 137.600 126.870 140.000 ;
    END
  END chany_top_out[16]
  PIN chany_top_out[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 129.810 137.600 130.090 140.000 ;
    END
  END chany_top_out[17]
  PIN chany_top_out[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 132.570 137.600 132.850 140.000 ;
    END
  END chany_top_out[18]
  PIN chany_top_out[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 135.330 137.600 135.610 140.000 ;
    END
  END chany_top_out[19]
  PIN chany_top_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 83.810 137.600 84.090 140.000 ;
    END
  END chany_top_out[1]
  PIN chany_top_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 87.030 137.600 87.310 140.000 ;
    END
  END chany_top_out[2]
  PIN chany_top_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 89.790 137.600 90.070 140.000 ;
    END
  END chany_top_out[3]
  PIN chany_top_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 92.550 137.600 92.830 140.000 ;
    END
  END chany_top_out[4]
  PIN chany_top_out[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 95.310 137.600 95.590 140.000 ;
    END
  END chany_top_out[5]
  PIN chany_top_out[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 98.070 137.600 98.350 140.000 ;
    END
  END chany_top_out[6]
  PIN chany_top_out[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 101.290 137.600 101.570 140.000 ;
    END
  END chany_top_out[7]
  PIN chany_top_out[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 104.050 137.600 104.330 140.000 ;
    END
  END chany_top_out[8]
  PIN chany_top_out[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 106.810 137.600 107.090 140.000 ;
    END
  END chany_top_out[9]
  PIN left_bottom_grid_pin_11_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 16.360 2.400 16.960 ;
    END
  END left_bottom_grid_pin_11_
  PIN left_bottom_grid_pin_1_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 1.400 2.400 2.000 ;
    END
  END left_bottom_grid_pin_1_
  PIN left_bottom_grid_pin_3_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 4.120 2.400 4.720 ;
    END
  END left_bottom_grid_pin_3_
  PIN left_bottom_grid_pin_5_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 6.840 2.400 7.440 ;
    END
  END left_bottom_grid_pin_5_
  PIN left_bottom_grid_pin_7_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 10.240 2.400 10.840 ;
    END
  END left_bottom_grid_pin_7_
  PIN left_bottom_grid_pin_9_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 12.960 2.400 13.560 ;
    END
  END left_bottom_grid_pin_9_
  PIN prog_clk
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 35.050 0.000 35.330 2.400 ;
    END
  END prog_clk
  PIN top_left_grid_pin_42_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1.470 137.600 1.750 140.000 ;
    END
  END top_left_grid_pin_42_
  PIN top_left_grid_pin_43_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 4.230 137.600 4.510 140.000 ;
    END
  END top_left_grid_pin_43_
  PIN top_left_grid_pin_44_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 6.990 137.600 7.270 140.000 ;
    END
  END top_left_grid_pin_44_
  PIN top_left_grid_pin_45_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 9.750 137.600 10.030 140.000 ;
    END
  END top_left_grid_pin_45_
  PIN top_left_grid_pin_46_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 12.510 137.600 12.790 140.000 ;
    END
  END top_left_grid_pin_46_
  PIN top_left_grid_pin_47_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 15.730 137.600 16.010 140.000 ;
    END
  END top_left_grid_pin_47_
  PIN top_left_grid_pin_48_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 18.490 137.600 18.770 140.000 ;
    END
  END top_left_grid_pin_48_
  PIN top_left_grid_pin_49_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 21.250 137.600 21.530 140.000 ;
    END
  END top_left_grid_pin_49_
  PIN top_right_grid_pin_1_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 138.090 137.600 138.370 140.000 ;
    END
  END top_right_grid_pin_1_
  PIN VPWR
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 28.055 10.640 29.655 128.080 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 51.385 10.640 52.985 128.080 ;
    END
  END VGND
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 134.320 127.925 ;
      LAYER met1 ;
        RECT 2.830 10.640 134.320 133.580 ;
      LAYER met2 ;
        RECT 2.030 137.320 3.950 138.565 ;
        RECT 4.790 137.320 6.710 138.565 ;
        RECT 7.550 137.320 9.470 138.565 ;
        RECT 10.310 137.320 12.230 138.565 ;
        RECT 13.070 137.320 15.450 138.565 ;
        RECT 16.290 137.320 18.210 138.565 ;
        RECT 19.050 137.320 20.970 138.565 ;
        RECT 21.810 137.320 23.730 138.565 ;
        RECT 24.570 137.320 26.490 138.565 ;
        RECT 27.330 137.320 29.710 138.565 ;
        RECT 30.550 137.320 32.470 138.565 ;
        RECT 33.310 137.320 35.230 138.565 ;
        RECT 36.070 137.320 37.990 138.565 ;
        RECT 38.830 137.320 40.750 138.565 ;
        RECT 41.590 137.320 43.970 138.565 ;
        RECT 44.810 137.320 46.730 138.565 ;
        RECT 47.570 137.320 49.490 138.565 ;
        RECT 50.330 137.320 52.250 138.565 ;
        RECT 53.090 137.320 55.010 138.565 ;
        RECT 55.850 137.320 58.230 138.565 ;
        RECT 59.070 137.320 60.990 138.565 ;
        RECT 61.830 137.320 63.750 138.565 ;
        RECT 64.590 137.320 66.510 138.565 ;
        RECT 67.350 137.320 69.270 138.565 ;
        RECT 70.110 137.320 72.490 138.565 ;
        RECT 73.330 137.320 75.250 138.565 ;
        RECT 76.090 137.320 78.010 138.565 ;
        RECT 78.850 137.320 80.770 138.565 ;
        RECT 81.610 137.320 83.530 138.565 ;
        RECT 84.370 137.320 86.750 138.565 ;
        RECT 87.590 137.320 89.510 138.565 ;
        RECT 90.350 137.320 92.270 138.565 ;
        RECT 93.110 137.320 95.030 138.565 ;
        RECT 95.870 137.320 97.790 138.565 ;
        RECT 98.630 137.320 101.010 138.565 ;
        RECT 101.850 137.320 103.770 138.565 ;
        RECT 104.610 137.320 106.530 138.565 ;
        RECT 107.370 137.320 109.290 138.565 ;
        RECT 110.130 137.320 112.050 138.565 ;
        RECT 112.890 137.320 115.270 138.565 ;
        RECT 116.110 137.320 118.030 138.565 ;
        RECT 118.870 137.320 120.790 138.565 ;
        RECT 121.630 137.320 123.550 138.565 ;
        RECT 124.390 137.320 126.310 138.565 ;
        RECT 127.150 137.320 129.530 138.565 ;
        RECT 130.370 137.320 132.290 138.565 ;
        RECT 133.130 137.320 135.050 138.565 ;
        RECT 135.890 137.320 137.810 138.565 ;
        RECT 1.470 2.680 138.370 137.320 ;
        RECT 1.470 1.515 34.770 2.680 ;
        RECT 35.610 1.515 104.690 2.680 ;
        RECT 105.530 1.515 138.370 2.680 ;
      LAYER met3 ;
        RECT 2.800 137.680 138.395 138.545 ;
        RECT 1.445 136.360 138.395 137.680 ;
        RECT 2.800 134.960 138.395 136.360 ;
        RECT 1.445 132.960 138.395 134.960 ;
        RECT 2.800 131.560 138.395 132.960 ;
        RECT 1.445 130.240 138.395 131.560 ;
        RECT 2.800 128.840 138.395 130.240 ;
        RECT 1.445 126.840 138.395 128.840 ;
        RECT 2.800 125.440 138.395 126.840 ;
        RECT 1.445 124.120 138.395 125.440 ;
        RECT 2.800 122.720 138.395 124.120 ;
        RECT 1.445 120.720 138.395 122.720 ;
        RECT 2.800 119.320 138.395 120.720 ;
        RECT 1.445 118.000 138.395 119.320 ;
        RECT 2.800 116.600 138.395 118.000 ;
        RECT 1.445 114.600 138.395 116.600 ;
        RECT 2.800 113.200 138.395 114.600 ;
        RECT 1.445 111.880 138.395 113.200 ;
        RECT 2.800 110.480 138.395 111.880 ;
        RECT 1.445 108.480 138.395 110.480 ;
        RECT 2.800 107.080 138.395 108.480 ;
        RECT 1.445 105.760 138.395 107.080 ;
        RECT 2.800 104.360 138.395 105.760 ;
        RECT 1.445 102.360 138.395 104.360 ;
        RECT 2.800 100.960 138.395 102.360 ;
        RECT 1.445 99.640 138.395 100.960 ;
        RECT 2.800 98.240 138.395 99.640 ;
        RECT 1.445 96.240 138.395 98.240 ;
        RECT 2.800 94.840 138.395 96.240 ;
        RECT 1.445 93.520 138.395 94.840 ;
        RECT 2.800 92.120 138.395 93.520 ;
        RECT 1.445 90.120 138.395 92.120 ;
        RECT 2.800 88.720 138.395 90.120 ;
        RECT 1.445 87.400 138.395 88.720 ;
        RECT 2.800 86.000 138.395 87.400 ;
        RECT 1.445 84.000 138.395 86.000 ;
        RECT 2.800 82.600 138.395 84.000 ;
        RECT 1.445 81.280 138.395 82.600 ;
        RECT 2.800 79.880 138.395 81.280 ;
        RECT 1.445 77.880 138.395 79.880 ;
        RECT 2.800 76.480 138.395 77.880 ;
        RECT 1.445 75.160 138.395 76.480 ;
        RECT 2.800 73.760 138.395 75.160 ;
        RECT 1.445 72.440 138.395 73.760 ;
        RECT 2.800 71.080 138.395 72.440 ;
        RECT 2.800 71.040 137.200 71.080 ;
        RECT 1.445 69.680 137.200 71.040 ;
        RECT 1.445 69.040 138.395 69.680 ;
        RECT 2.800 67.640 138.395 69.040 ;
        RECT 1.445 66.320 138.395 67.640 ;
        RECT 2.800 64.920 138.395 66.320 ;
        RECT 1.445 62.920 138.395 64.920 ;
        RECT 2.800 61.520 138.395 62.920 ;
        RECT 1.445 60.200 138.395 61.520 ;
        RECT 2.800 58.800 138.395 60.200 ;
        RECT 1.445 56.800 138.395 58.800 ;
        RECT 2.800 55.400 138.395 56.800 ;
        RECT 1.445 54.080 138.395 55.400 ;
        RECT 2.800 52.680 138.395 54.080 ;
        RECT 1.445 50.680 138.395 52.680 ;
        RECT 2.800 49.280 138.395 50.680 ;
        RECT 1.445 47.960 138.395 49.280 ;
        RECT 2.800 46.560 138.395 47.960 ;
        RECT 1.445 44.560 138.395 46.560 ;
        RECT 2.800 43.160 138.395 44.560 ;
        RECT 1.445 41.840 138.395 43.160 ;
        RECT 2.800 40.440 138.395 41.840 ;
        RECT 1.445 38.440 138.395 40.440 ;
        RECT 2.800 37.040 138.395 38.440 ;
        RECT 1.445 35.720 138.395 37.040 ;
        RECT 2.800 34.320 138.395 35.720 ;
        RECT 1.445 32.320 138.395 34.320 ;
        RECT 2.800 30.920 138.395 32.320 ;
        RECT 1.445 29.600 138.395 30.920 ;
        RECT 2.800 28.200 138.395 29.600 ;
        RECT 1.445 26.200 138.395 28.200 ;
        RECT 2.800 24.800 138.395 26.200 ;
        RECT 1.445 23.480 138.395 24.800 ;
        RECT 2.800 22.080 138.395 23.480 ;
        RECT 1.445 20.080 138.395 22.080 ;
        RECT 2.800 18.680 138.395 20.080 ;
        RECT 1.445 17.360 138.395 18.680 ;
        RECT 2.800 15.960 138.395 17.360 ;
        RECT 1.445 13.960 138.395 15.960 ;
        RECT 2.800 12.560 138.395 13.960 ;
        RECT 1.445 11.240 138.395 12.560 ;
        RECT 2.800 9.840 138.395 11.240 ;
        RECT 1.445 7.840 138.395 9.840 ;
        RECT 2.800 6.440 138.395 7.840 ;
        RECT 1.445 5.120 138.395 6.440 ;
        RECT 2.800 3.720 138.395 5.120 ;
        RECT 1.445 2.400 138.395 3.720 ;
        RECT 2.800 1.535 138.395 2.400 ;
      LAYER met4 ;
        RECT 9.990 10.640 27.655 128.080 ;
        RECT 30.055 10.640 50.985 128.080 ;
        RECT 53.385 10.640 122.985 128.080 ;
      LAYER met5 ;
        RECT 9.780 106.300 49.100 107.900 ;
  END
END sb_2__0_
END LIBRARY

