magic
tech EFS8A
magscale 1 2
timestamp 1602076583
<< locali >>
rect 7699 16609 7734 16643
rect 10735 16609 10770 16643
rect 7843 14569 7849 14603
rect 7843 14501 7877 14569
rect 10091 14433 10126 14467
rect 18199 14025 18337 14059
rect 15847 12393 15853 12427
rect 15847 12325 15881 12393
rect 19199 10081 19234 10115
rect 7199 9367 7233 9435
rect 7199 9333 7205 9367
rect 18647 8993 18682 9027
rect 10051 8041 10057 8075
rect 10051 7973 10085 8041
rect 8493 7905 8654 7939
rect 8493 7735 8527 7905
rect 15243 6817 15370 6851
<< viali >>
rect 8861 20553 8895 20587
rect 19441 20553 19475 20587
rect 21097 20553 21131 20587
rect 8677 20349 8711 20383
rect 19257 20349 19291 20383
rect 19809 20349 19843 20383
rect 20913 20349 20947 20383
rect 21465 20349 21499 20383
rect 9321 20213 9355 20247
rect 7021 17289 7055 17323
rect 6837 17085 6871 17119
rect 7976 17085 8010 17119
rect 8401 17085 8435 17119
rect 7481 16949 7515 16983
rect 8079 16949 8113 16983
rect 8217 16745 8251 16779
rect 7665 16609 7699 16643
rect 10701 16609 10735 16643
rect 7803 16405 7837 16439
rect 10839 16405 10873 16439
rect 7757 16201 7791 16235
rect 8033 16065 8067 16099
rect 11044 15997 11078 16031
rect 11437 15997 11471 16031
rect 7389 15929 7423 15963
rect 8125 15929 8159 15963
rect 8677 15929 8711 15963
rect 10793 15929 10827 15963
rect 11115 15861 11149 15895
rect 5319 15657 5353 15691
rect 10793 15657 10827 15691
rect 8217 15589 8251 15623
rect 9873 15589 9907 15623
rect 11437 15589 11471 15623
rect 5248 15521 5282 15555
rect 12884 15521 12918 15555
rect 15644 15521 15678 15555
rect 8125 15453 8159 15487
rect 8769 15453 8803 15487
rect 9781 15453 9815 15487
rect 10057 15453 10091 15487
rect 11345 15453 11379 15487
rect 11805 15453 11839 15487
rect 15715 15385 15749 15419
rect 16405 15385 16439 15419
rect 12955 15317 12989 15351
rect 16037 15317 16071 15351
rect 7757 15113 7791 15147
rect 8033 15113 8067 15147
rect 10149 15113 10183 15147
rect 11805 15113 11839 15147
rect 12173 15113 12207 15147
rect 14841 15113 14875 15147
rect 15669 15113 15703 15147
rect 21097 15113 21131 15147
rect 21557 15113 21591 15147
rect 5273 14977 5307 15011
rect 9505 14977 9539 15011
rect 10885 14977 10919 15011
rect 11161 14977 11195 15011
rect 12541 14977 12575 15011
rect 16037 14977 16071 15011
rect 6837 14909 6871 14943
rect 14968 14909 15002 14943
rect 20913 14909 20947 14943
rect 7158 14841 7192 14875
rect 8861 14841 8895 14875
rect 8953 14841 8987 14875
rect 10701 14841 10735 14875
rect 10977 14841 11011 14875
rect 12633 14841 12667 14875
rect 13185 14841 13219 14875
rect 16129 14841 16163 14875
rect 16681 14841 16715 14875
rect 5549 14773 5583 14807
rect 6561 14773 6595 14807
rect 8677 14773 8711 14807
rect 9781 14773 9815 14807
rect 13553 14773 13587 14807
rect 15071 14773 15105 14807
rect 7849 14569 7883 14603
rect 8401 14569 8435 14603
rect 12081 14569 12115 14603
rect 12541 14569 12575 14603
rect 5733 14501 5767 14535
rect 6285 14501 6319 14535
rect 8677 14501 8711 14535
rect 11253 14501 11287 14535
rect 11805 14501 11839 14535
rect 16129 14501 16163 14535
rect 16681 14501 16715 14535
rect 10057 14433 10091 14467
rect 5641 14365 5675 14399
rect 7481 14365 7515 14399
rect 10195 14365 10229 14399
rect 11161 14365 11195 14399
rect 16037 14365 16071 14399
rect 9137 14297 9171 14331
rect 6929 14229 6963 14263
rect 10609 14229 10643 14263
rect 1593 14025 1627 14059
rect 5917 14025 5951 14059
rect 6561 14025 6595 14059
rect 9229 14025 9263 14059
rect 11529 14025 11563 14059
rect 12173 14025 12207 14059
rect 15209 14025 15243 14059
rect 18337 14025 18371 14059
rect 6193 13957 6227 13991
rect 11805 13957 11839 13991
rect 2053 13889 2087 13923
rect 10057 13889 10091 13923
rect 10609 13889 10643 13923
rect 16405 13889 16439 13923
rect 16681 13889 16715 13923
rect 18521 13889 18555 13923
rect 1409 13821 1443 13855
rect 4997 13821 5031 13855
rect 8309 13821 8343 13855
rect 15577 13821 15611 13855
rect 16037 13821 16071 13855
rect 18096 13821 18130 13855
rect 4905 13753 4939 13787
rect 5359 13753 5393 13787
rect 7573 13753 7607 13787
rect 8217 13753 8251 13787
rect 8671 13753 8705 13787
rect 10930 13753 10964 13787
rect 7113 13685 7147 13719
rect 10517 13685 10551 13719
rect 5089 13481 5123 13515
rect 5641 13481 5675 13515
rect 11437 13481 11471 13515
rect 16221 13481 16255 13515
rect 10879 13413 10913 13447
rect 15663 13413 15697 13447
rect 17233 13413 17267 13447
rect 5825 13345 5859 13379
rect 6193 13345 6227 13379
rect 6469 13345 6503 13379
rect 6929 13345 6963 13379
rect 10517 13277 10551 13311
rect 15301 13277 15335 13311
rect 17141 13277 17175 13311
rect 17785 13277 17819 13311
rect 7389 13141 7423 13175
rect 8309 13141 8343 13175
rect 10057 13141 10091 13175
rect 13369 13141 13403 13175
rect 13829 13141 13863 13175
rect 5273 12937 5307 12971
rect 16405 12937 16439 12971
rect 17141 12937 17175 12971
rect 17509 12869 17543 12903
rect 11437 12801 11471 12835
rect 12081 12801 12115 12835
rect 14841 12801 14875 12835
rect 15669 12801 15703 12835
rect 18061 12801 18095 12835
rect 5641 12733 5675 12767
rect 6285 12733 6319 12767
rect 7113 12733 7147 12767
rect 7573 12733 7607 12767
rect 7665 12733 7699 12767
rect 8217 12733 8251 12767
rect 10057 12733 10091 12767
rect 10425 12733 10459 12767
rect 10793 12733 10827 12767
rect 11345 12733 11379 12767
rect 13369 12733 13403 12767
rect 13829 12733 13863 12767
rect 14197 12733 14231 12767
rect 14565 12733 14599 12767
rect 16221 12733 16255 12767
rect 16773 12733 16807 12767
rect 9781 12665 9815 12699
rect 12909 12665 12943 12699
rect 4905 12597 4939 12631
rect 6561 12597 6595 12631
rect 7113 12597 7147 12631
rect 9505 12597 9539 12631
rect 11713 12597 11747 12631
rect 13277 12597 13311 12631
rect 15393 12597 15427 12631
rect 7021 12393 7055 12427
rect 10609 12393 10643 12427
rect 12817 12393 12851 12427
rect 15853 12393 15887 12427
rect 16405 12393 16439 12427
rect 7665 12325 7699 12359
rect 8493 12325 8527 12359
rect 9505 12325 9539 12359
rect 17417 12325 17451 12359
rect 5825 12257 5859 12291
rect 6285 12257 6319 12291
rect 6653 12257 6687 12291
rect 7205 12257 7239 12291
rect 10333 12257 10367 12291
rect 10793 12257 10827 12291
rect 11161 12257 11195 12291
rect 11529 12257 11563 12291
rect 13185 12257 13219 12291
rect 13369 12257 13403 12291
rect 13921 12257 13955 12291
rect 14289 12257 14323 12291
rect 18864 12257 18898 12291
rect 5641 12189 5675 12223
rect 14381 12189 14415 12223
rect 15485 12189 15519 12223
rect 17325 12189 17359 12223
rect 17785 12189 17819 12223
rect 8125 12053 8159 12087
rect 10057 12053 10091 12087
rect 12449 12053 12483 12087
rect 18935 12053 18969 12087
rect 1593 11849 1627 11883
rect 5549 11849 5583 11883
rect 10333 11849 10367 11883
rect 12725 11849 12759 11883
rect 14657 11849 14691 11883
rect 16773 11849 16807 11883
rect 17325 11849 17359 11883
rect 18889 11849 18923 11883
rect 1409 11645 1443 11679
rect 1961 11645 1995 11679
rect 6653 11645 6687 11679
rect 7573 11645 7607 11679
rect 8309 11645 8343 11679
rect 8493 11645 8527 11679
rect 8861 11645 8895 11679
rect 9413 11645 9447 11679
rect 10057 11645 10091 11679
rect 11345 11645 11379 11679
rect 11529 11645 11563 11679
rect 13185 11645 13219 11679
rect 13369 11645 13403 11679
rect 13737 11645 13771 11679
rect 14289 11645 14323 11679
rect 14381 11645 14415 11679
rect 15577 11645 15611 11679
rect 15898 11577 15932 11611
rect 5825 11509 5859 11543
rect 6285 11509 6319 11543
rect 7849 11509 7883 11543
rect 8309 11509 8343 11543
rect 11805 11509 11839 11543
rect 12173 11509 12207 11543
rect 15117 11509 15151 11543
rect 15393 11509 15427 11543
rect 16497 11509 16531 11543
rect 17693 11509 17727 11543
rect 5549 11305 5583 11339
rect 10057 11305 10091 11339
rect 15485 11305 15519 11339
rect 16221 11305 16255 11339
rect 8211 11237 8245 11271
rect 17233 11237 17267 11271
rect 17785 11237 17819 11271
rect 18705 11237 18739 11271
rect 18797 11237 18831 11271
rect 5733 11169 5767 11203
rect 6193 11169 6227 11203
rect 6469 11169 6503 11203
rect 6653 11169 6687 11203
rect 9505 11169 9539 11203
rect 10057 11169 10091 11203
rect 10241 11169 10275 11203
rect 10609 11169 10643 11203
rect 10977 11169 11011 11203
rect 15301 11169 15335 11203
rect 7849 11101 7883 11135
rect 13001 11101 13035 11135
rect 17141 11101 17175 11135
rect 18981 11101 19015 11135
rect 12265 11033 12299 11067
rect 12633 11033 12667 11067
rect 7757 10965 7791 10999
rect 8769 10965 8803 10999
rect 13277 10965 13311 10999
rect 13645 10965 13679 10999
rect 15853 10965 15887 10999
rect 18153 10965 18187 10999
rect 1961 10761 1995 10795
rect 5181 10761 5215 10795
rect 12909 10761 12943 10795
rect 15209 10761 15243 10795
rect 17141 10761 17175 10795
rect 17417 10761 17451 10795
rect 19441 10761 19475 10795
rect 5917 10693 5951 10727
rect 6285 10693 6319 10727
rect 9781 10693 9815 10727
rect 21097 10693 21131 10727
rect 10241 10625 10275 10659
rect 11805 10625 11839 10659
rect 14565 10625 14599 10659
rect 15393 10625 15427 10659
rect 18429 10625 18463 10659
rect 1568 10557 1602 10591
rect 5549 10557 5583 10591
rect 7389 10557 7423 10591
rect 8125 10557 8159 10591
rect 8585 10557 8619 10591
rect 8677 10557 8711 10591
rect 9045 10557 9079 10591
rect 12265 10557 12299 10591
rect 13369 10557 13403 10591
rect 13553 10557 13587 10591
rect 13921 10557 13955 10591
rect 14289 10557 14323 10591
rect 16313 10557 16347 10591
rect 17785 10557 17819 10591
rect 20913 10557 20947 10591
rect 21465 10557 21499 10591
rect 7757 10489 7791 10523
rect 10603 10489 10637 10523
rect 14933 10489 14967 10523
rect 15714 10489 15748 10523
rect 18153 10489 18187 10523
rect 18245 10489 18279 10523
rect 1639 10421 1673 10455
rect 4353 10421 4387 10455
rect 7941 10421 7975 10455
rect 11161 10421 11195 10455
rect 11529 10421 11563 10455
rect 19073 10421 19107 10455
rect 7941 10217 7975 10251
rect 9505 10217 9539 10251
rect 14105 10217 14139 10251
rect 19303 10217 19337 10251
rect 4439 10149 4473 10183
rect 10333 10149 10367 10183
rect 13001 10149 13035 10183
rect 16221 10149 16255 10183
rect 17785 10149 17819 10183
rect 18337 10149 18371 10183
rect 4077 10081 4111 10115
rect 6101 10081 6135 10115
rect 6377 10081 6411 10115
rect 6653 10081 6687 10115
rect 7021 10081 7055 10115
rect 8585 10081 8619 10115
rect 12357 10081 12391 10115
rect 13277 10081 13311 10115
rect 19165 10081 19199 10115
rect 10241 10013 10275 10047
rect 10885 10013 10919 10047
rect 16129 10013 16163 10047
rect 16773 10013 16807 10047
rect 17693 10013 17727 10047
rect 7205 9945 7239 9979
rect 4997 9877 5031 9911
rect 8309 9877 8343 9911
rect 9873 9877 9907 9911
rect 11161 9877 11195 9911
rect 13645 9877 13679 9911
rect 15577 9877 15611 9911
rect 3709 9673 3743 9707
rect 4077 9673 4111 9707
rect 4537 9673 4571 9707
rect 5917 9673 5951 9707
rect 9781 9673 9815 9707
rect 10241 9673 10275 9707
rect 10609 9673 10643 9707
rect 12633 9673 12667 9707
rect 19165 9673 19199 9707
rect 18705 9605 18739 9639
rect 4813 9537 4847 9571
rect 5089 9537 5123 9571
rect 6837 9537 6871 9571
rect 8953 9537 8987 9571
rect 14749 9537 14783 9571
rect 15577 9537 15611 9571
rect 19763 9537 19797 9571
rect 13277 9469 13311 9503
rect 13737 9469 13771 9503
rect 14289 9469 14323 9503
rect 14473 9469 14507 9503
rect 16497 9469 16531 9503
rect 17417 9469 17451 9503
rect 17785 9469 17819 9503
rect 19660 9469 19694 9503
rect 20085 9469 20119 9503
rect 4905 9401 4939 9435
rect 8125 9401 8159 9435
rect 8677 9401 8711 9435
rect 8769 9401 8803 9435
rect 10885 9401 10919 9435
rect 10977 9401 11011 9435
rect 11529 9401 11563 9435
rect 15939 9401 15973 9435
rect 18153 9401 18187 9435
rect 18245 9401 18279 9435
rect 6285 9333 6319 9367
rect 6561 9333 6595 9367
rect 7205 9333 7239 9367
rect 7757 9333 7791 9367
rect 8493 9333 8527 9367
rect 13185 9333 13219 9367
rect 15485 9333 15519 9367
rect 16865 9333 16899 9367
rect 4813 9129 4847 9163
rect 5917 9129 5951 9163
rect 6285 9129 6319 9163
rect 6929 9129 6963 9163
rect 10011 9129 10045 9163
rect 16221 9129 16255 9163
rect 18061 9129 18095 9163
rect 21051 9129 21085 9163
rect 1547 9061 1581 9095
rect 7849 9061 7883 9095
rect 10333 9061 10367 9095
rect 11069 9061 11103 9095
rect 15663 9061 15697 9095
rect 17233 9061 17267 9095
rect 17785 9061 17819 9095
rect 1460 8993 1494 9027
rect 9908 8993 9942 9027
rect 13185 8993 13219 9027
rect 13461 8993 13495 9027
rect 13737 8993 13771 9027
rect 14105 8993 14139 9027
rect 18613 8993 18647 9027
rect 19676 8993 19710 9027
rect 20948 8993 20982 9027
rect 7757 8925 7791 8959
rect 8033 8925 8067 8959
rect 10977 8925 11011 8959
rect 11253 8925 11287 8959
rect 14381 8925 14415 8959
rect 15301 8925 15335 8959
rect 17141 8925 17175 8959
rect 18521 8925 18555 8959
rect 19763 8925 19797 8959
rect 10701 8789 10735 8823
rect 16497 8789 16531 8823
rect 18751 8789 18785 8823
rect 1593 8585 1627 8619
rect 7205 8585 7239 8619
rect 9781 8585 9815 8619
rect 11253 8585 11287 8619
rect 12587 8585 12621 8619
rect 13645 8585 13679 8619
rect 14841 8585 14875 8619
rect 15163 8585 15197 8619
rect 16819 8585 16853 8619
rect 17509 8585 17543 8619
rect 20085 8585 20119 8619
rect 21189 8585 21223 8619
rect 8953 8517 8987 8551
rect 18613 8517 18647 8551
rect 20729 8517 20763 8551
rect 7435 8449 7469 8483
rect 9965 8449 9999 8483
rect 1409 8381 1443 8415
rect 7348 8381 7382 8415
rect 12265 8381 12299 8415
rect 12516 8381 12550 8415
rect 15060 8381 15094 8415
rect 15485 8381 15519 8415
rect 16748 8381 16782 8415
rect 19073 8381 19107 8415
rect 20545 8381 20579 8415
rect 7849 8313 7883 8347
rect 8401 8313 8435 8347
rect 8493 8313 8527 8347
rect 10057 8313 10091 8347
rect 10609 8313 10643 8347
rect 13369 8313 13403 8347
rect 21465 8313 21499 8347
rect 2053 8245 2087 8279
rect 8125 8245 8159 8279
rect 9321 8245 9355 8279
rect 10977 8245 11011 8279
rect 12909 8245 12943 8279
rect 14013 8245 14047 8279
rect 15853 8245 15887 8279
rect 17233 8245 17267 8279
rect 19441 8245 19475 8279
rect 1685 8041 1719 8075
rect 7665 8041 7699 8075
rect 10057 8041 10091 8075
rect 10609 8041 10643 8075
rect 17049 8041 17083 8075
rect 7066 7973 7100 8007
rect 7941 7973 7975 8007
rect 11621 7973 11655 8007
rect 15755 7973 15789 8007
rect 17877 7973 17911 8007
rect 19441 7973 19475 8007
rect 8723 7905 8757 7939
rect 6745 7837 6779 7871
rect 9689 7837 9723 7871
rect 11529 7837 11563 7871
rect 11897 7837 11931 7871
rect 15393 7837 15427 7871
rect 17785 7837 17819 7871
rect 19349 7837 19383 7871
rect 20913 7837 20947 7871
rect 9137 7769 9171 7803
rect 18337 7769 18371 7803
rect 19901 7769 19935 7803
rect 8401 7701 8435 7735
rect 8493 7701 8527 7735
rect 10885 7701 10919 7735
rect 13185 7701 13219 7735
rect 13645 7701 13679 7735
rect 16313 7701 16347 7735
rect 18981 7701 19015 7735
rect 10885 7497 10919 7531
rect 11529 7497 11563 7531
rect 11805 7497 11839 7531
rect 18337 7497 18371 7531
rect 18889 7497 18923 7531
rect 19993 7497 20027 7531
rect 10609 7361 10643 7395
rect 14657 7361 14691 7395
rect 19717 7361 19751 7395
rect 6653 7293 6687 7327
rect 7113 7293 7147 7327
rect 7297 7293 7331 7327
rect 7849 7293 7883 7327
rect 8217 7293 8251 7327
rect 9413 7293 9447 7327
rect 9689 7293 9723 7327
rect 9965 7293 9999 7327
rect 10333 7293 10367 7327
rect 13185 7293 13219 7327
rect 13645 7293 13679 7327
rect 14013 7293 14047 7327
rect 14381 7293 14415 7327
rect 15669 7293 15703 7327
rect 5917 7225 5951 7259
rect 15990 7225 16024 7259
rect 19073 7225 19107 7259
rect 19165 7225 19199 7259
rect 6193 7157 6227 7191
rect 6929 7157 6963 7191
rect 8677 7157 8711 7191
rect 8953 7157 8987 7191
rect 12633 7157 12667 7191
rect 13093 7157 13127 7191
rect 15025 7157 15059 7191
rect 15485 7157 15519 7191
rect 16589 7157 16623 7191
rect 17785 7157 17819 7191
rect 7665 6953 7699 6987
rect 8631 6953 8665 6987
rect 9229 6953 9263 6987
rect 9965 6953 9999 6987
rect 11069 6953 11103 6987
rect 16129 6953 16163 6987
rect 19073 6953 19107 6987
rect 14381 6885 14415 6919
rect 17969 6885 18003 6919
rect 7297 6817 7331 6851
rect 8560 6817 8594 6851
rect 10425 6817 10459 6851
rect 12909 6817 12943 6851
rect 13461 6817 13495 6851
rect 13737 6817 13771 6851
rect 14289 6817 14323 6851
rect 15209 6817 15243 6851
rect 16840 6817 16874 6851
rect 10793 6749 10827 6783
rect 17877 6749 17911 6783
rect 18337 6749 18371 6783
rect 19349 6749 19383 6783
rect 12357 6681 12391 6715
rect 6837 6613 6871 6647
rect 10333 6613 10367 6647
rect 10563 6613 10597 6647
rect 10701 6613 10735 6647
rect 12725 6613 12759 6647
rect 15439 6613 15473 6647
rect 15853 6613 15887 6647
rect 16911 6613 16945 6647
rect 11621 6409 11655 6443
rect 15301 6409 15335 6443
rect 16681 6409 16715 6443
rect 17417 6409 17451 6443
rect 17877 6409 17911 6443
rect 12909 6341 12943 6375
rect 13277 6341 13311 6375
rect 9781 6273 9815 6307
rect 10609 6273 10643 6307
rect 18061 6273 18095 6307
rect 9137 6205 9171 6239
rect 9413 6205 9447 6239
rect 11253 6205 11287 6239
rect 13461 6205 13495 6239
rect 13921 6205 13955 6239
rect 14289 6205 14323 6239
rect 14657 6205 14691 6239
rect 14933 6205 14967 6239
rect 15761 6205 15795 6239
rect 18153 6205 18187 6239
rect 9229 6137 9263 6171
rect 10517 6137 10551 6171
rect 16082 6137 16116 6171
rect 17049 6137 17083 6171
rect 8585 6069 8619 6103
rect 10057 6069 10091 6103
rect 12173 6069 12207 6103
rect 16129 5865 16163 5899
rect 18061 5865 18095 5899
rect 11345 5797 11379 5831
rect 12909 5797 12943 5831
rect 16957 5797 16991 5831
rect 9321 5729 9355 5763
rect 10057 5729 10091 5763
rect 10609 5729 10643 5763
rect 12173 5729 12207 5763
rect 18337 5729 18371 5763
rect 10977 5661 11011 5695
rect 12541 5661 12575 5695
rect 16865 5661 16899 5695
rect 10774 5593 10808 5627
rect 12081 5593 12115 5627
rect 12449 5593 12483 5627
rect 13829 5593 13863 5627
rect 17417 5593 17451 5627
rect 18521 5593 18555 5627
rect 10425 5525 10459 5559
rect 10885 5525 10919 5559
rect 12338 5525 12372 5559
rect 13461 5525 13495 5559
rect 14289 5525 14323 5559
rect 15761 5525 15795 5559
rect 9873 5321 9907 5355
rect 10793 5321 10827 5355
rect 11805 5321 11839 5355
rect 17233 5321 17267 5355
rect 18337 5321 18371 5355
rect 12633 5253 12667 5287
rect 7665 5185 7699 5219
rect 13185 5185 13219 5219
rect 15117 5185 15151 5219
rect 7021 5117 7055 5151
rect 10425 5117 10459 5151
rect 13369 5117 13403 5151
rect 13829 5117 13863 5151
rect 14381 5117 14415 5151
rect 14565 5117 14599 5151
rect 14841 5117 14875 5151
rect 15669 5117 15703 5151
rect 10149 5049 10183 5083
rect 15990 5049 16024 5083
rect 16957 5049 16991 5083
rect 6561 4981 6595 5015
rect 11437 4981 11471 5015
rect 12173 4981 12207 5015
rect 15485 4981 15519 5015
rect 16589 4981 16623 5015
rect 9965 4777 9999 4811
rect 10793 4777 10827 4811
rect 11529 4777 11563 4811
rect 13461 4777 13495 4811
rect 13921 4777 13955 4811
rect 15669 4777 15703 4811
rect 17049 4709 17083 4743
rect 18429 4709 18463 4743
rect 9781 4641 9815 4675
rect 11621 4641 11655 4675
rect 12081 4641 12115 4675
rect 12449 4641 12483 4675
rect 13001 4641 13035 4675
rect 18521 4641 18555 4675
rect 14197 4573 14231 4607
rect 16957 4573 16991 4607
rect 17417 4573 17451 4607
rect 13001 4505 13035 4539
rect 9689 4233 9723 4267
rect 10701 4233 10735 4267
rect 11897 4233 11931 4267
rect 12265 4233 12299 4267
rect 18521 4233 18555 4267
rect 17233 4165 17267 4199
rect 11529 4097 11563 4131
rect 12909 4097 12943 4131
rect 13277 4097 13311 4131
rect 16957 4097 16991 4131
rect 10977 4029 11011 4063
rect 13461 4029 13495 4063
rect 13921 4029 13955 4063
rect 14289 4029 14323 4063
rect 14657 4029 14691 4063
rect 15669 4029 15703 4063
rect 15853 4029 15887 4063
rect 18096 4029 18130 4063
rect 18889 4029 18923 4063
rect 14933 3961 14967 3995
rect 16497 3961 16531 3995
rect 18199 3961 18233 3995
rect 12449 3893 12483 3927
rect 12265 3689 12299 3723
rect 12725 3689 12759 3723
rect 14289 3689 14323 3723
rect 16221 3689 16255 3723
rect 17141 3689 17175 3723
rect 11989 3621 12023 3655
rect 13461 3621 13495 3655
rect 15622 3621 15656 3655
rect 11437 3553 11471 3587
rect 11621 3553 11655 3587
rect 13369 3485 13403 3519
rect 15301 3485 15335 3519
rect 13921 3417 13955 3451
rect 10701 3145 10735 3179
rect 14013 3145 14047 3179
rect 16497 3145 16531 3179
rect 16773 3145 16807 3179
rect 10977 3077 11011 3111
rect 16037 3077 16071 3111
rect 12449 3009 12483 3043
rect 15485 3009 15519 3043
rect 17141 3009 17175 3043
rect 11161 2941 11195 2975
rect 14197 2941 14231 2975
rect 14749 2941 14783 2975
rect 12265 2873 12299 2907
rect 12770 2873 12804 2907
rect 15209 2873 15243 2907
rect 15577 2873 15611 2907
rect 11345 2805 11379 2839
rect 11805 2805 11839 2839
rect 13369 2805 13403 2839
rect 13645 2805 13679 2839
rect 14381 2805 14415 2839
rect 12449 2601 12483 2635
rect 15301 2601 15335 2635
rect 17187 2601 17221 2635
rect 7481 2533 7515 2567
rect 13185 2533 13219 2567
rect 13737 2533 13771 2567
rect 14933 2533 14967 2567
rect 15577 2533 15611 2567
rect 15669 2533 15703 2567
rect 6996 2465 7030 2499
rect 9781 2465 9815 2499
rect 10333 2465 10367 2499
rect 10885 2465 10919 2499
rect 11069 2465 11103 2499
rect 17084 2465 17118 2499
rect 18337 2465 18371 2499
rect 18889 2465 18923 2499
rect 21189 2465 21223 2499
rect 21741 2465 21775 2499
rect 11713 2397 11747 2431
rect 12817 2397 12851 2431
rect 13093 2397 13127 2431
rect 15853 2397 15887 2431
rect 17509 2397 17543 2431
rect 18521 2329 18555 2363
rect 21373 2329 21407 2363
rect 7067 2261 7101 2295
rect 9965 2261 9999 2295
<< metal1 >>
rect 13906 23536 13912 23588
rect 13964 23576 13970 23588
rect 14918 23576 14924 23588
rect 13964 23548 14924 23576
rect 13964 23536 13970 23548
rect 14918 23536 14924 23548
rect 14976 23536 14982 23588
rect 1104 21786 22816 21808
rect 1104 21734 4982 21786
rect 5034 21734 5046 21786
rect 5098 21734 5110 21786
rect 5162 21734 5174 21786
rect 5226 21734 12982 21786
rect 13034 21734 13046 21786
rect 13098 21734 13110 21786
rect 13162 21734 13174 21786
rect 13226 21734 20982 21786
rect 21034 21734 21046 21786
rect 21098 21734 21110 21786
rect 21162 21734 21174 21786
rect 21226 21734 22816 21786
rect 1104 21712 22816 21734
rect 1104 21242 22816 21264
rect 1104 21190 8982 21242
rect 9034 21190 9046 21242
rect 9098 21190 9110 21242
rect 9162 21190 9174 21242
rect 9226 21190 16982 21242
rect 17034 21190 17046 21242
rect 17098 21190 17110 21242
rect 17162 21190 17174 21242
rect 17226 21190 22816 21242
rect 1104 21168 22816 21190
rect 1104 20698 22816 20720
rect 1104 20646 4982 20698
rect 5034 20646 5046 20698
rect 5098 20646 5110 20698
rect 5162 20646 5174 20698
rect 5226 20646 12982 20698
rect 13034 20646 13046 20698
rect 13098 20646 13110 20698
rect 13162 20646 13174 20698
rect 13226 20646 20982 20698
rect 21034 20646 21046 20698
rect 21098 20646 21110 20698
rect 21162 20646 21174 20698
rect 21226 20646 22816 20698
rect 1104 20624 22816 20646
rect 8846 20584 8852 20596
rect 8807 20556 8852 20584
rect 8846 20544 8852 20556
rect 8904 20544 8910 20596
rect 19429 20587 19487 20593
rect 19429 20553 19441 20587
rect 19475 20584 19487 20587
rect 20622 20584 20628 20596
rect 19475 20556 20628 20584
rect 19475 20553 19487 20556
rect 19429 20547 19487 20553
rect 20622 20544 20628 20556
rect 20680 20544 20686 20596
rect 21085 20587 21143 20593
rect 21085 20553 21097 20587
rect 21131 20584 21143 20587
rect 22646 20584 22652 20596
rect 21131 20556 22652 20584
rect 21131 20553 21143 20556
rect 21085 20547 21143 20553
rect 22646 20544 22652 20556
rect 22704 20544 22710 20596
rect 8665 20383 8723 20389
rect 8665 20349 8677 20383
rect 8711 20380 8723 20383
rect 8711 20352 9352 20380
rect 8711 20349 8723 20352
rect 8665 20343 8723 20349
rect 9324 20253 9352 20352
rect 15838 20340 15844 20392
rect 15896 20380 15902 20392
rect 19245 20383 19303 20389
rect 19245 20380 19257 20383
rect 15896 20352 19257 20380
rect 15896 20340 15902 20352
rect 19245 20349 19257 20352
rect 19291 20380 19303 20383
rect 19797 20383 19855 20389
rect 19797 20380 19809 20383
rect 19291 20352 19809 20380
rect 19291 20349 19303 20352
rect 19245 20343 19303 20349
rect 19797 20349 19809 20352
rect 19843 20349 19855 20383
rect 19797 20343 19855 20349
rect 20806 20340 20812 20392
rect 20864 20380 20870 20392
rect 20901 20383 20959 20389
rect 20901 20380 20913 20383
rect 20864 20352 20913 20380
rect 20864 20340 20870 20352
rect 20901 20349 20913 20352
rect 20947 20380 20959 20383
rect 21453 20383 21511 20389
rect 21453 20380 21465 20383
rect 20947 20352 21465 20380
rect 20947 20349 20959 20352
rect 20901 20343 20959 20349
rect 21453 20349 21465 20352
rect 21499 20349 21511 20383
rect 21453 20343 21511 20349
rect 9309 20247 9367 20253
rect 9309 20213 9321 20247
rect 9355 20244 9367 20247
rect 10778 20244 10784 20256
rect 9355 20216 10784 20244
rect 9355 20213 9367 20216
rect 9309 20207 9367 20213
rect 10778 20204 10784 20216
rect 10836 20204 10842 20256
rect 1104 20154 22816 20176
rect 1104 20102 8982 20154
rect 9034 20102 9046 20154
rect 9098 20102 9110 20154
rect 9162 20102 9174 20154
rect 9226 20102 16982 20154
rect 17034 20102 17046 20154
rect 17098 20102 17110 20154
rect 17162 20102 17174 20154
rect 17226 20102 22816 20154
rect 1104 20080 22816 20102
rect 1104 19610 22816 19632
rect 1104 19558 4982 19610
rect 5034 19558 5046 19610
rect 5098 19558 5110 19610
rect 5162 19558 5174 19610
rect 5226 19558 12982 19610
rect 13034 19558 13046 19610
rect 13098 19558 13110 19610
rect 13162 19558 13174 19610
rect 13226 19558 20982 19610
rect 21034 19558 21046 19610
rect 21098 19558 21110 19610
rect 21162 19558 21174 19610
rect 21226 19558 22816 19610
rect 1104 19536 22816 19558
rect 1104 19066 22816 19088
rect 1104 19014 8982 19066
rect 9034 19014 9046 19066
rect 9098 19014 9110 19066
rect 9162 19014 9174 19066
rect 9226 19014 16982 19066
rect 17034 19014 17046 19066
rect 17098 19014 17110 19066
rect 17162 19014 17174 19066
rect 17226 19014 22816 19066
rect 1104 18992 22816 19014
rect 1104 18522 22816 18544
rect 1104 18470 4982 18522
rect 5034 18470 5046 18522
rect 5098 18470 5110 18522
rect 5162 18470 5174 18522
rect 5226 18470 12982 18522
rect 13034 18470 13046 18522
rect 13098 18470 13110 18522
rect 13162 18470 13174 18522
rect 13226 18470 20982 18522
rect 21034 18470 21046 18522
rect 21098 18470 21110 18522
rect 21162 18470 21174 18522
rect 21226 18470 22816 18522
rect 1104 18448 22816 18470
rect 1104 17978 22816 18000
rect 1104 17926 8982 17978
rect 9034 17926 9046 17978
rect 9098 17926 9110 17978
rect 9162 17926 9174 17978
rect 9226 17926 16982 17978
rect 17034 17926 17046 17978
rect 17098 17926 17110 17978
rect 17162 17926 17174 17978
rect 17226 17926 22816 17978
rect 1104 17904 22816 17926
rect 11146 17620 11152 17672
rect 11204 17660 11210 17672
rect 14182 17660 14188 17672
rect 11204 17632 14188 17660
rect 11204 17620 11210 17632
rect 14182 17620 14188 17632
rect 14240 17620 14246 17672
rect 1104 17434 22816 17456
rect 1104 17382 4982 17434
rect 5034 17382 5046 17434
rect 5098 17382 5110 17434
rect 5162 17382 5174 17434
rect 5226 17382 12982 17434
rect 13034 17382 13046 17434
rect 13098 17382 13110 17434
rect 13162 17382 13174 17434
rect 13226 17382 20982 17434
rect 21034 17382 21046 17434
rect 21098 17382 21110 17434
rect 21162 17382 21174 17434
rect 21226 17382 22816 17434
rect 1104 17360 22816 17382
rect 7006 17320 7012 17332
rect 6967 17292 7012 17320
rect 7006 17280 7012 17292
rect 7064 17280 7070 17332
rect 5350 17144 5356 17196
rect 5408 17184 5414 17196
rect 5408 17156 7189 17184
rect 5408 17144 5414 17156
rect 6825 17119 6883 17125
rect 6825 17085 6837 17119
rect 6871 17085 6883 17119
rect 7161 17116 7189 17156
rect 7964 17119 8022 17125
rect 7964 17116 7976 17119
rect 7161 17088 7976 17116
rect 6825 17079 6883 17085
rect 7964 17085 7976 17088
rect 8010 17116 8022 17119
rect 8386 17116 8392 17128
rect 8010 17088 8392 17116
rect 8010 17085 8022 17088
rect 7964 17079 8022 17085
rect 6840 16980 6868 17079
rect 8386 17076 8392 17088
rect 8444 17076 8450 17128
rect 7469 16983 7527 16989
rect 7469 16980 7481 16983
rect 6840 16952 7481 16980
rect 7469 16949 7481 16952
rect 7515 16980 7527 16983
rect 7742 16980 7748 16992
rect 7515 16952 7748 16980
rect 7515 16949 7527 16952
rect 7469 16943 7527 16949
rect 7742 16940 7748 16952
rect 7800 16940 7806 16992
rect 8067 16983 8125 16989
rect 8067 16949 8079 16983
rect 8113 16980 8125 16983
rect 8202 16980 8208 16992
rect 8113 16952 8208 16980
rect 8113 16949 8125 16952
rect 8067 16943 8125 16949
rect 8202 16940 8208 16952
rect 8260 16940 8266 16992
rect 1104 16890 22816 16912
rect 1104 16838 8982 16890
rect 9034 16838 9046 16890
rect 9098 16838 9110 16890
rect 9162 16838 9174 16890
rect 9226 16838 16982 16890
rect 17034 16838 17046 16890
rect 17098 16838 17110 16890
rect 17162 16838 17174 16890
rect 17226 16838 22816 16890
rect 1104 16816 22816 16838
rect 8202 16776 8208 16788
rect 8163 16748 8208 16776
rect 8202 16736 8208 16748
rect 8260 16736 8266 16788
rect 7653 16643 7711 16649
rect 7653 16609 7665 16643
rect 7699 16640 7711 16643
rect 7742 16640 7748 16652
rect 7699 16612 7748 16640
rect 7699 16609 7711 16612
rect 7653 16603 7711 16609
rect 7742 16600 7748 16612
rect 7800 16600 7806 16652
rect 10689 16643 10747 16649
rect 10689 16609 10701 16643
rect 10735 16640 10747 16643
rect 10778 16640 10784 16652
rect 10735 16612 10784 16640
rect 10735 16609 10747 16612
rect 10689 16603 10747 16609
rect 10778 16600 10784 16612
rect 10836 16600 10842 16652
rect 7791 16439 7849 16445
rect 7791 16405 7803 16439
rect 7837 16436 7849 16439
rect 8110 16436 8116 16448
rect 7837 16408 8116 16436
rect 7837 16405 7849 16408
rect 7791 16399 7849 16405
rect 8110 16396 8116 16408
rect 8168 16396 8174 16448
rect 10686 16396 10692 16448
rect 10744 16436 10750 16448
rect 10827 16439 10885 16445
rect 10827 16436 10839 16439
rect 10744 16408 10839 16436
rect 10744 16396 10750 16408
rect 10827 16405 10839 16408
rect 10873 16405 10885 16439
rect 10827 16399 10885 16405
rect 1104 16346 22816 16368
rect 1104 16294 4982 16346
rect 5034 16294 5046 16346
rect 5098 16294 5110 16346
rect 5162 16294 5174 16346
rect 5226 16294 12982 16346
rect 13034 16294 13046 16346
rect 13098 16294 13110 16346
rect 13162 16294 13174 16346
rect 13226 16294 20982 16346
rect 21034 16294 21046 16346
rect 21098 16294 21110 16346
rect 21162 16294 21174 16346
rect 21226 16294 22816 16346
rect 1104 16272 22816 16294
rect 7742 16232 7748 16244
rect 7703 16204 7748 16232
rect 7742 16192 7748 16204
rect 7800 16192 7806 16244
rect 8021 16099 8079 16105
rect 8021 16065 8033 16099
rect 8067 16096 8079 16099
rect 8202 16096 8208 16108
rect 8067 16068 8208 16096
rect 8067 16065 8079 16068
rect 8021 16059 8079 16065
rect 8202 16056 8208 16068
rect 8260 16056 8266 16108
rect 11032 16031 11090 16037
rect 11032 15997 11044 16031
rect 11078 16028 11090 16031
rect 11422 16028 11428 16040
rect 11078 16000 11428 16028
rect 11078 15997 11090 16000
rect 11032 15991 11090 15997
rect 11422 15988 11428 16000
rect 11480 15988 11486 16040
rect 7377 15963 7435 15969
rect 7377 15929 7389 15963
rect 7423 15960 7435 15963
rect 8113 15963 8171 15969
rect 8113 15960 8125 15963
rect 7423 15932 8125 15960
rect 7423 15929 7435 15932
rect 7377 15923 7435 15929
rect 8113 15929 8125 15932
rect 8159 15960 8171 15963
rect 8202 15960 8208 15972
rect 8159 15932 8208 15960
rect 8159 15929 8171 15932
rect 8113 15923 8171 15929
rect 8202 15920 8208 15932
rect 8260 15920 8266 15972
rect 8665 15963 8723 15969
rect 8665 15929 8677 15963
rect 8711 15960 8723 15963
rect 9582 15960 9588 15972
rect 8711 15932 9588 15960
rect 8711 15929 8723 15932
rect 8665 15923 8723 15929
rect 9582 15920 9588 15932
rect 9640 15920 9646 15972
rect 10778 15960 10784 15972
rect 10691 15932 10784 15960
rect 10778 15920 10784 15932
rect 10836 15960 10842 15972
rect 14826 15960 14832 15972
rect 10836 15932 14832 15960
rect 10836 15920 10842 15932
rect 14826 15920 14832 15932
rect 14884 15960 14890 15972
rect 16758 15960 16764 15972
rect 14884 15932 16764 15960
rect 14884 15920 14890 15932
rect 16758 15920 16764 15932
rect 16816 15920 16822 15972
rect 11103 15895 11161 15901
rect 11103 15861 11115 15895
rect 11149 15892 11161 15895
rect 11330 15892 11336 15904
rect 11149 15864 11336 15892
rect 11149 15861 11161 15864
rect 11103 15855 11161 15861
rect 11330 15852 11336 15864
rect 11388 15852 11394 15904
rect 11422 15852 11428 15904
rect 11480 15892 11486 15904
rect 15838 15892 15844 15904
rect 11480 15864 15844 15892
rect 11480 15852 11486 15864
rect 15838 15852 15844 15864
rect 15896 15852 15902 15904
rect 1104 15802 22816 15824
rect 1104 15750 8982 15802
rect 9034 15750 9046 15802
rect 9098 15750 9110 15802
rect 9162 15750 9174 15802
rect 9226 15750 16982 15802
rect 17034 15750 17046 15802
rect 17098 15750 17110 15802
rect 17162 15750 17174 15802
rect 17226 15750 22816 15802
rect 1104 15728 22816 15750
rect 106 15648 112 15700
rect 164 15688 170 15700
rect 5307 15691 5365 15697
rect 5307 15688 5319 15691
rect 164 15660 5319 15688
rect 164 15648 170 15660
rect 5307 15657 5319 15660
rect 5353 15657 5365 15691
rect 5307 15651 5365 15657
rect 10686 15648 10692 15700
rect 10744 15688 10750 15700
rect 10781 15691 10839 15697
rect 10781 15688 10793 15691
rect 10744 15660 10793 15688
rect 10744 15648 10750 15660
rect 10781 15657 10793 15660
rect 10827 15657 10839 15691
rect 10781 15651 10839 15657
rect 8202 15620 8208 15632
rect 8163 15592 8208 15620
rect 8202 15580 8208 15592
rect 8260 15580 8266 15632
rect 9766 15580 9772 15632
rect 9824 15620 9830 15632
rect 9861 15623 9919 15629
rect 9861 15620 9873 15623
rect 9824 15592 9873 15620
rect 9824 15580 9830 15592
rect 9861 15589 9873 15592
rect 9907 15589 9919 15623
rect 11422 15620 11428 15632
rect 11383 15592 11428 15620
rect 9861 15583 9919 15589
rect 11422 15580 11428 15592
rect 11480 15580 11486 15632
rect 5236 15555 5294 15561
rect 5236 15521 5248 15555
rect 5282 15552 5294 15555
rect 5350 15552 5356 15564
rect 5282 15524 5356 15552
rect 5282 15521 5294 15524
rect 5236 15515 5294 15521
rect 5350 15512 5356 15524
rect 5408 15512 5414 15564
rect 12872 15555 12930 15561
rect 12872 15521 12884 15555
rect 12918 15552 12930 15555
rect 13538 15552 13544 15564
rect 12918 15524 13544 15552
rect 12918 15521 12930 15524
rect 12872 15515 12930 15521
rect 13538 15512 13544 15524
rect 13596 15512 13602 15564
rect 15632 15555 15690 15561
rect 15632 15521 15644 15555
rect 15678 15552 15690 15555
rect 15838 15552 15844 15564
rect 15678 15524 15844 15552
rect 15678 15521 15690 15524
rect 15632 15515 15690 15521
rect 15838 15512 15844 15524
rect 15896 15512 15902 15564
rect 8110 15484 8116 15496
rect 8071 15456 8116 15484
rect 8110 15444 8116 15456
rect 8168 15444 8174 15496
rect 8757 15487 8815 15493
rect 8757 15453 8769 15487
rect 8803 15484 8815 15487
rect 8846 15484 8852 15496
rect 8803 15456 8852 15484
rect 8803 15453 8815 15456
rect 8757 15447 8815 15453
rect 8846 15444 8852 15456
rect 8904 15444 8910 15496
rect 9582 15444 9588 15496
rect 9640 15484 9646 15496
rect 9769 15487 9827 15493
rect 9769 15484 9781 15487
rect 9640 15456 9781 15484
rect 9640 15444 9646 15456
rect 9769 15453 9781 15456
rect 9815 15453 9827 15487
rect 10042 15484 10048 15496
rect 10003 15456 10048 15484
rect 9769 15447 9827 15453
rect 10042 15444 10048 15456
rect 10100 15444 10106 15496
rect 11330 15484 11336 15496
rect 11291 15456 11336 15484
rect 11330 15444 11336 15456
rect 11388 15444 11394 15496
rect 11790 15484 11796 15496
rect 11751 15456 11796 15484
rect 11790 15444 11796 15456
rect 11848 15444 11854 15496
rect 15703 15419 15761 15425
rect 15703 15385 15715 15419
rect 15749 15416 15761 15419
rect 16114 15416 16120 15428
rect 15749 15388 16120 15416
rect 15749 15385 15761 15388
rect 15703 15379 15761 15385
rect 16114 15376 16120 15388
rect 16172 15416 16178 15428
rect 16393 15419 16451 15425
rect 16393 15416 16405 15419
rect 16172 15388 16405 15416
rect 16172 15376 16178 15388
rect 16393 15385 16405 15388
rect 16439 15385 16451 15419
rect 16393 15379 16451 15385
rect 12526 15308 12532 15360
rect 12584 15348 12590 15360
rect 12943 15351 13001 15357
rect 12943 15348 12955 15351
rect 12584 15320 12955 15348
rect 12584 15308 12590 15320
rect 12943 15317 12955 15320
rect 12989 15317 13001 15351
rect 16022 15348 16028 15360
rect 15983 15320 16028 15348
rect 12943 15311 13001 15317
rect 16022 15308 16028 15320
rect 16080 15308 16086 15360
rect 1104 15258 22816 15280
rect 1104 15206 4982 15258
rect 5034 15206 5046 15258
rect 5098 15206 5110 15258
rect 5162 15206 5174 15258
rect 5226 15206 12982 15258
rect 13034 15206 13046 15258
rect 13098 15206 13110 15258
rect 13162 15206 13174 15258
rect 13226 15206 20982 15258
rect 21034 15206 21046 15258
rect 21098 15206 21110 15258
rect 21162 15206 21174 15258
rect 21226 15206 22816 15258
rect 1104 15184 22816 15206
rect 7745 15147 7803 15153
rect 7745 15113 7757 15147
rect 7791 15144 7803 15147
rect 8021 15147 8079 15153
rect 8021 15144 8033 15147
rect 7791 15116 8033 15144
rect 7791 15113 7803 15116
rect 7745 15107 7803 15113
rect 8021 15113 8033 15116
rect 8067 15144 8079 15147
rect 8202 15144 8208 15156
rect 8067 15116 8208 15144
rect 8067 15113 8079 15116
rect 8021 15107 8079 15113
rect 8202 15104 8208 15116
rect 8260 15104 8266 15156
rect 9582 15104 9588 15156
rect 9640 15144 9646 15156
rect 10137 15147 10195 15153
rect 10137 15144 10149 15147
rect 9640 15116 10149 15144
rect 9640 15104 9646 15116
rect 10137 15113 10149 15116
rect 10183 15113 10195 15147
rect 10137 15107 10195 15113
rect 10152 15076 10180 15107
rect 11422 15104 11428 15156
rect 11480 15144 11486 15156
rect 11793 15147 11851 15153
rect 11793 15144 11805 15147
rect 11480 15116 11805 15144
rect 11480 15104 11486 15116
rect 11793 15113 11805 15116
rect 11839 15144 11851 15147
rect 12161 15147 12219 15153
rect 12161 15144 12173 15147
rect 11839 15116 12173 15144
rect 11839 15113 11851 15116
rect 11793 15107 11851 15113
rect 12161 15113 12173 15116
rect 12207 15113 12219 15147
rect 14826 15144 14832 15156
rect 14787 15116 14832 15144
rect 12161 15107 12219 15113
rect 10152 15048 11192 15076
rect 5261 15011 5319 15017
rect 5261 14977 5273 15011
rect 5307 15008 5319 15011
rect 5350 15008 5356 15020
rect 5307 14980 5356 15008
rect 5307 14977 5319 14980
rect 5261 14971 5319 14977
rect 5350 14968 5356 14980
rect 5408 15008 5414 15020
rect 6270 15008 6276 15020
rect 5408 14980 6276 15008
rect 5408 14968 5414 14980
rect 6270 14968 6276 14980
rect 6328 15008 6334 15020
rect 9493 15011 9551 15017
rect 9493 15008 9505 15011
rect 6328 14980 9505 15008
rect 6328 14968 6334 14980
rect 9493 14977 9505 14980
rect 9539 15008 9551 15011
rect 10042 15008 10048 15020
rect 9539 14980 10048 15008
rect 9539 14977 9551 14980
rect 9493 14971 9551 14977
rect 10042 14968 10048 14980
rect 10100 14968 10106 15020
rect 10686 14968 10692 15020
rect 10744 15008 10750 15020
rect 11164 15017 11192 15048
rect 10873 15011 10931 15017
rect 10873 15008 10885 15011
rect 10744 14980 10885 15008
rect 10744 14968 10750 14980
rect 10873 14977 10885 14980
rect 10919 14977 10931 15011
rect 10873 14971 10931 14977
rect 11149 15011 11207 15017
rect 11149 14977 11161 15011
rect 11195 15008 11207 15011
rect 11195 14980 12112 15008
rect 11195 14977 11207 14980
rect 11149 14971 11207 14977
rect 6825 14943 6883 14949
rect 6825 14909 6837 14943
rect 6871 14940 6883 14943
rect 7006 14940 7012 14952
rect 6871 14912 7012 14940
rect 6871 14909 6883 14912
rect 6825 14903 6883 14909
rect 7006 14900 7012 14912
rect 7064 14900 7070 14952
rect 7146 14875 7204 14881
rect 7146 14872 7158 14875
rect 6564 14844 7158 14872
rect 6564 14816 6592 14844
rect 7146 14841 7158 14844
rect 7192 14841 7204 14875
rect 8846 14872 8852 14884
rect 8807 14844 8852 14872
rect 7146 14835 7204 14841
rect 8846 14832 8852 14844
rect 8904 14832 8910 14884
rect 8941 14875 8999 14881
rect 8941 14841 8953 14875
rect 8987 14841 8999 14875
rect 8941 14835 8999 14841
rect 10689 14875 10747 14881
rect 10689 14841 10701 14875
rect 10735 14872 10747 14875
rect 10965 14875 11023 14881
rect 10965 14872 10977 14875
rect 10735 14844 10977 14872
rect 10735 14841 10747 14844
rect 10689 14835 10747 14841
rect 10965 14841 10977 14844
rect 11011 14872 11023 14875
rect 11238 14872 11244 14884
rect 11011 14844 11244 14872
rect 11011 14841 11023 14844
rect 10965 14835 11023 14841
rect 5537 14807 5595 14813
rect 5537 14773 5549 14807
rect 5583 14804 5595 14807
rect 5626 14804 5632 14816
rect 5583 14776 5632 14804
rect 5583 14773 5595 14776
rect 5537 14767 5595 14773
rect 5626 14764 5632 14776
rect 5684 14764 5690 14816
rect 6546 14804 6552 14816
rect 6507 14776 6552 14804
rect 6546 14764 6552 14776
rect 6604 14764 6610 14816
rect 8665 14807 8723 14813
rect 8665 14773 8677 14807
rect 8711 14804 8723 14807
rect 8754 14804 8760 14816
rect 8711 14776 8760 14804
rect 8711 14773 8723 14776
rect 8665 14767 8723 14773
rect 8754 14764 8760 14776
rect 8812 14804 8818 14816
rect 8956 14804 8984 14835
rect 11238 14832 11244 14844
rect 11296 14832 11302 14884
rect 9766 14804 9772 14816
rect 8812 14776 8984 14804
rect 9727 14776 9772 14804
rect 8812 14764 8818 14776
rect 9766 14764 9772 14776
rect 9824 14764 9830 14816
rect 12084 14804 12112 14980
rect 12176 14872 12204 15107
rect 14826 15104 14832 15116
rect 14884 15104 14890 15156
rect 15657 15147 15715 15153
rect 15657 15113 15669 15147
rect 15703 15144 15715 15147
rect 15838 15144 15844 15156
rect 15703 15116 15844 15144
rect 15703 15113 15715 15116
rect 15657 15107 15715 15113
rect 15838 15104 15844 15116
rect 15896 15104 15902 15156
rect 21085 15147 21143 15153
rect 21085 15113 21097 15147
rect 21131 15144 21143 15147
rect 21266 15144 21272 15156
rect 21131 15116 21272 15144
rect 21131 15113 21143 15116
rect 21085 15107 21143 15113
rect 21266 15104 21272 15116
rect 21324 15104 21330 15156
rect 21542 15144 21548 15156
rect 21503 15116 21548 15144
rect 21542 15104 21548 15116
rect 21600 15104 21606 15156
rect 13538 15036 13544 15088
rect 13596 15076 13602 15088
rect 18598 15076 18604 15088
rect 13596 15048 18604 15076
rect 13596 15036 13602 15048
rect 18598 15036 18604 15048
rect 18656 15036 18662 15088
rect 12526 15008 12532 15020
rect 12487 14980 12532 15008
rect 12526 14968 12532 14980
rect 12584 14968 12590 15020
rect 16025 15011 16083 15017
rect 16025 14977 16037 15011
rect 16071 15008 16083 15011
rect 16114 15008 16120 15020
rect 16071 14980 16120 15008
rect 16071 14977 16083 14980
rect 16025 14971 16083 14977
rect 16114 14968 16120 14980
rect 16172 14968 16178 15020
rect 14826 14900 14832 14952
rect 14884 14940 14890 14952
rect 14956 14943 15014 14949
rect 14956 14940 14968 14943
rect 14884 14912 14968 14940
rect 14884 14900 14890 14912
rect 14956 14909 14968 14912
rect 15002 14909 15014 14943
rect 14956 14903 15014 14909
rect 20806 14900 20812 14952
rect 20864 14940 20870 14952
rect 20901 14943 20959 14949
rect 20901 14940 20913 14943
rect 20864 14912 20913 14940
rect 20864 14900 20870 14912
rect 20901 14909 20913 14912
rect 20947 14940 20959 14943
rect 21542 14940 21548 14952
rect 20947 14912 21548 14940
rect 20947 14909 20959 14912
rect 20901 14903 20959 14909
rect 21542 14900 21548 14912
rect 21600 14900 21606 14952
rect 12621 14875 12679 14881
rect 12621 14872 12633 14875
rect 12176 14844 12633 14872
rect 12621 14841 12633 14844
rect 12667 14841 12679 14875
rect 12621 14835 12679 14841
rect 13173 14875 13231 14881
rect 13173 14841 13185 14875
rect 13219 14841 13231 14875
rect 13173 14835 13231 14841
rect 13188 14804 13216 14835
rect 16022 14832 16028 14884
rect 16080 14872 16086 14884
rect 16117 14875 16175 14881
rect 16117 14872 16129 14875
rect 16080 14844 16129 14872
rect 16080 14832 16086 14844
rect 16117 14841 16129 14844
rect 16163 14841 16175 14875
rect 16666 14872 16672 14884
rect 16627 14844 16672 14872
rect 16117 14835 16175 14841
rect 16666 14832 16672 14844
rect 16724 14832 16730 14884
rect 13538 14804 13544 14816
rect 12084 14776 13216 14804
rect 13499 14776 13544 14804
rect 13538 14764 13544 14776
rect 13596 14764 13602 14816
rect 15059 14807 15117 14813
rect 15059 14773 15071 14807
rect 15105 14804 15117 14807
rect 15194 14804 15200 14816
rect 15105 14776 15200 14804
rect 15105 14773 15117 14776
rect 15059 14767 15117 14773
rect 15194 14764 15200 14776
rect 15252 14764 15258 14816
rect 1104 14714 22816 14736
rect 1104 14662 8982 14714
rect 9034 14662 9046 14714
rect 9098 14662 9110 14714
rect 9162 14662 9174 14714
rect 9226 14662 16982 14714
rect 17034 14662 17046 14714
rect 17098 14662 17110 14714
rect 17162 14662 17174 14714
rect 17226 14662 22816 14714
rect 1104 14640 22816 14662
rect 7834 14600 7840 14612
rect 7795 14572 7840 14600
rect 7834 14560 7840 14572
rect 7892 14560 7898 14612
rect 8389 14603 8447 14609
rect 8389 14569 8401 14603
rect 8435 14600 8447 14603
rect 9766 14600 9772 14612
rect 8435 14572 9772 14600
rect 8435 14569 8447 14572
rect 8389 14563 8447 14569
rect 9766 14560 9772 14572
rect 9824 14560 9830 14612
rect 11330 14560 11336 14612
rect 11388 14600 11394 14612
rect 12069 14603 12127 14609
rect 12069 14600 12081 14603
rect 11388 14572 12081 14600
rect 11388 14560 11394 14572
rect 12069 14569 12081 14572
rect 12115 14569 12127 14603
rect 12526 14600 12532 14612
rect 12487 14572 12532 14600
rect 12069 14563 12127 14569
rect 12526 14560 12532 14572
rect 12584 14560 12590 14612
rect 5718 14532 5724 14544
rect 5679 14504 5724 14532
rect 5718 14492 5724 14504
rect 5776 14492 5782 14544
rect 6270 14532 6276 14544
rect 6231 14504 6276 14532
rect 6270 14492 6276 14504
rect 6328 14492 6334 14544
rect 8110 14492 8116 14544
rect 8168 14532 8174 14544
rect 8665 14535 8723 14541
rect 8665 14532 8677 14535
rect 8168 14504 8677 14532
rect 8168 14492 8174 14504
rect 8665 14501 8677 14504
rect 8711 14501 8723 14535
rect 11238 14532 11244 14544
rect 11199 14504 11244 14532
rect 8665 14495 8723 14501
rect 11238 14492 11244 14504
rect 11296 14492 11302 14544
rect 11790 14532 11796 14544
rect 11751 14504 11796 14532
rect 11790 14492 11796 14504
rect 11848 14492 11854 14544
rect 16114 14532 16120 14544
rect 16075 14504 16120 14532
rect 16114 14492 16120 14504
rect 16172 14492 16178 14544
rect 16666 14532 16672 14544
rect 16627 14504 16672 14532
rect 16666 14492 16672 14504
rect 16724 14492 16730 14544
rect 10042 14464 10048 14476
rect 10003 14436 10048 14464
rect 10042 14424 10048 14436
rect 10100 14424 10106 14476
rect 5626 14396 5632 14408
rect 5587 14368 5632 14396
rect 5626 14356 5632 14368
rect 5684 14356 5690 14408
rect 7098 14356 7104 14408
rect 7156 14396 7162 14408
rect 7469 14399 7527 14405
rect 7469 14396 7481 14399
rect 7156 14368 7481 14396
rect 7156 14356 7162 14368
rect 7469 14365 7481 14368
rect 7515 14365 7527 14399
rect 7469 14359 7527 14365
rect 10183 14399 10241 14405
rect 10183 14365 10195 14399
rect 10229 14396 10241 14399
rect 11149 14399 11207 14405
rect 11149 14396 11161 14399
rect 10229 14368 11161 14396
rect 10229 14365 10241 14368
rect 10183 14359 10241 14365
rect 11149 14365 11161 14368
rect 11195 14396 11207 14399
rect 12158 14396 12164 14408
rect 11195 14368 12164 14396
rect 11195 14365 11207 14368
rect 11149 14359 11207 14365
rect 12158 14356 12164 14368
rect 12216 14356 12222 14408
rect 15194 14356 15200 14408
rect 15252 14396 15258 14408
rect 16025 14399 16083 14405
rect 16025 14396 16037 14399
rect 15252 14368 16037 14396
rect 15252 14356 15258 14368
rect 16025 14365 16037 14368
rect 16071 14365 16083 14399
rect 16025 14359 16083 14365
rect 8846 14288 8852 14340
rect 8904 14328 8910 14340
rect 9125 14331 9183 14337
rect 9125 14328 9137 14331
rect 8904 14300 9137 14328
rect 8904 14288 8910 14300
rect 9125 14297 9137 14300
rect 9171 14328 9183 14331
rect 11790 14328 11796 14340
rect 9171 14300 11796 14328
rect 9171 14297 9183 14300
rect 9125 14291 9183 14297
rect 11790 14288 11796 14300
rect 11848 14288 11854 14340
rect 6917 14263 6975 14269
rect 6917 14229 6929 14263
rect 6963 14260 6975 14263
rect 7006 14260 7012 14272
rect 6963 14232 7012 14260
rect 6963 14229 6975 14232
rect 6917 14223 6975 14229
rect 7006 14220 7012 14232
rect 7064 14220 7070 14272
rect 10594 14260 10600 14272
rect 10555 14232 10600 14260
rect 10594 14220 10600 14232
rect 10652 14220 10658 14272
rect 1104 14170 22816 14192
rect 1104 14118 4982 14170
rect 5034 14118 5046 14170
rect 5098 14118 5110 14170
rect 5162 14118 5174 14170
rect 5226 14118 12982 14170
rect 13034 14118 13046 14170
rect 13098 14118 13110 14170
rect 13162 14118 13174 14170
rect 13226 14118 20982 14170
rect 21034 14118 21046 14170
rect 21098 14118 21110 14170
rect 21162 14118 21174 14170
rect 21226 14118 22816 14170
rect 1104 14096 22816 14118
rect 1486 14016 1492 14068
rect 1544 14056 1550 14068
rect 1581 14059 1639 14065
rect 1581 14056 1593 14059
rect 1544 14028 1593 14056
rect 1544 14016 1550 14028
rect 1581 14025 1593 14028
rect 1627 14025 1639 14059
rect 1581 14019 1639 14025
rect 5718 14016 5724 14068
rect 5776 14056 5782 14068
rect 5905 14059 5963 14065
rect 5905 14056 5917 14059
rect 5776 14028 5917 14056
rect 5776 14016 5782 14028
rect 5905 14025 5917 14028
rect 5951 14056 5963 14059
rect 6549 14059 6607 14065
rect 6549 14056 6561 14059
rect 5951 14028 6561 14056
rect 5951 14025 5963 14028
rect 5905 14019 5963 14025
rect 6549 14025 6561 14028
rect 6595 14025 6607 14059
rect 6549 14019 6607 14025
rect 8754 14016 8760 14068
rect 8812 14056 8818 14068
rect 9217 14059 9275 14065
rect 9217 14056 9229 14059
rect 8812 14028 9229 14056
rect 8812 14016 8818 14028
rect 9217 14025 9229 14028
rect 9263 14025 9275 14059
rect 9217 14019 9275 14025
rect 11422 14016 11428 14068
rect 11480 14056 11486 14068
rect 11517 14059 11575 14065
rect 11517 14056 11529 14059
rect 11480 14028 11529 14056
rect 11480 14016 11486 14028
rect 11517 14025 11529 14028
rect 11563 14025 11575 14059
rect 12158 14056 12164 14068
rect 12119 14028 12164 14056
rect 11517 14019 11575 14025
rect 12158 14016 12164 14028
rect 12216 14016 12222 14068
rect 15194 14056 15200 14068
rect 15155 14028 15200 14056
rect 15194 14016 15200 14028
rect 15252 14016 15258 14068
rect 18322 14056 18328 14068
rect 18283 14028 18328 14056
rect 18322 14016 18328 14028
rect 18380 14016 18386 14068
rect 5626 13948 5632 14000
rect 5684 13988 5690 14000
rect 6181 13991 6239 13997
rect 6181 13988 6193 13991
rect 5684 13960 6193 13988
rect 5684 13948 5690 13960
rect 6181 13957 6193 13960
rect 6227 13957 6239 13991
rect 6181 13951 6239 13957
rect 11238 13948 11244 14000
rect 11296 13988 11302 14000
rect 11793 13991 11851 13997
rect 11793 13988 11805 13991
rect 11296 13960 11805 13988
rect 11296 13948 11302 13960
rect 11793 13957 11805 13960
rect 11839 13957 11851 13991
rect 11793 13951 11851 13957
rect 2041 13923 2099 13929
rect 2041 13920 2053 13923
rect 1412 13892 2053 13920
rect 1412 13861 1440 13892
rect 2041 13889 2053 13892
rect 2087 13920 2099 13923
rect 9398 13920 9404 13932
rect 2087 13892 9404 13920
rect 2087 13889 2099 13892
rect 2041 13883 2099 13889
rect 9398 13880 9404 13892
rect 9456 13920 9462 13932
rect 10042 13920 10048 13932
rect 9456 13892 10048 13920
rect 9456 13880 9462 13892
rect 10042 13880 10048 13892
rect 10100 13880 10106 13932
rect 10594 13920 10600 13932
rect 10555 13892 10600 13920
rect 10594 13880 10600 13892
rect 10652 13880 10658 13932
rect 16114 13880 16120 13932
rect 16172 13920 16178 13932
rect 16393 13923 16451 13929
rect 16393 13920 16405 13923
rect 16172 13892 16405 13920
rect 16172 13880 16178 13892
rect 16393 13889 16405 13892
rect 16439 13920 16451 13923
rect 16669 13923 16727 13929
rect 16669 13920 16681 13923
rect 16439 13892 16681 13920
rect 16439 13889 16451 13892
rect 16393 13883 16451 13889
rect 16669 13889 16681 13892
rect 16715 13889 16727 13923
rect 18509 13923 18567 13929
rect 18509 13920 18521 13923
rect 16669 13883 16727 13889
rect 18099 13892 18521 13920
rect 1397 13855 1455 13861
rect 1397 13821 1409 13855
rect 1443 13821 1455 13855
rect 4982 13852 4988 13864
rect 4943 13824 4988 13852
rect 1397 13815 1455 13821
rect 4982 13812 4988 13824
rect 5040 13812 5046 13864
rect 8294 13852 8300 13864
rect 8255 13824 8300 13852
rect 8294 13812 8300 13824
rect 8352 13812 8358 13864
rect 15565 13855 15623 13861
rect 15565 13821 15577 13855
rect 15611 13852 15623 13855
rect 16022 13852 16028 13864
rect 15611 13824 16028 13852
rect 15611 13821 15623 13824
rect 15565 13815 15623 13821
rect 16022 13812 16028 13824
rect 16080 13812 16086 13864
rect 17770 13812 17776 13864
rect 17828 13852 17834 13864
rect 18099 13861 18127 13892
rect 18509 13889 18521 13892
rect 18555 13889 18567 13923
rect 18509 13883 18567 13889
rect 18084 13855 18142 13861
rect 18084 13852 18096 13855
rect 17828 13824 18096 13852
rect 17828 13812 17834 13824
rect 18084 13821 18096 13824
rect 18130 13821 18142 13855
rect 18084 13815 18142 13821
rect 4893 13787 4951 13793
rect 4893 13753 4905 13787
rect 4939 13784 4951 13787
rect 5347 13787 5405 13793
rect 5347 13784 5359 13787
rect 4939 13756 5359 13784
rect 4939 13753 4951 13756
rect 4893 13747 4951 13753
rect 5347 13753 5359 13756
rect 5393 13784 5405 13787
rect 6638 13784 6644 13796
rect 5393 13756 6644 13784
rect 5393 13753 5405 13756
rect 5347 13747 5405 13753
rect 6638 13744 6644 13756
rect 6696 13784 6702 13796
rect 7561 13787 7619 13793
rect 7561 13784 7573 13787
rect 6696 13756 7573 13784
rect 6696 13744 6702 13756
rect 7561 13753 7573 13756
rect 7607 13784 7619 13787
rect 7834 13784 7840 13796
rect 7607 13756 7840 13784
rect 7607 13753 7619 13756
rect 7561 13747 7619 13753
rect 7834 13744 7840 13756
rect 7892 13784 7898 13796
rect 8205 13787 8263 13793
rect 8205 13784 8217 13787
rect 7892 13756 8217 13784
rect 7892 13744 7898 13756
rect 8205 13753 8217 13756
rect 8251 13784 8263 13787
rect 8659 13787 8717 13793
rect 8659 13784 8671 13787
rect 8251 13756 8671 13784
rect 8251 13753 8263 13756
rect 8205 13747 8263 13753
rect 8659 13753 8671 13756
rect 8705 13753 8717 13787
rect 8659 13747 8717 13753
rect 10918 13787 10976 13793
rect 10918 13753 10930 13787
rect 10964 13753 10976 13787
rect 10918 13747 10976 13753
rect 7098 13716 7104 13728
rect 7059 13688 7104 13716
rect 7098 13676 7104 13688
rect 7156 13676 7162 13728
rect 8680 13716 8708 13747
rect 10502 13716 10508 13728
rect 8680 13688 10508 13716
rect 10502 13676 10508 13688
rect 10560 13716 10566 13728
rect 10933 13716 10961 13747
rect 10560 13688 10961 13716
rect 10560 13676 10566 13688
rect 1104 13626 22816 13648
rect 1104 13574 8982 13626
rect 9034 13574 9046 13626
rect 9098 13574 9110 13626
rect 9162 13574 9174 13626
rect 9226 13574 16982 13626
rect 17034 13574 17046 13626
rect 17098 13574 17110 13626
rect 17162 13574 17174 13626
rect 17226 13574 22816 13626
rect 1104 13552 22816 13574
rect 4982 13472 4988 13524
rect 5040 13512 5046 13524
rect 5077 13515 5135 13521
rect 5077 13512 5089 13515
rect 5040 13484 5089 13512
rect 5040 13472 5046 13484
rect 5077 13481 5089 13484
rect 5123 13512 5135 13515
rect 5629 13515 5687 13521
rect 5629 13512 5641 13515
rect 5123 13484 5641 13512
rect 5123 13481 5135 13484
rect 5077 13475 5135 13481
rect 5629 13481 5641 13484
rect 5675 13481 5687 13515
rect 5629 13475 5687 13481
rect 11238 13472 11244 13524
rect 11296 13512 11302 13524
rect 11425 13515 11483 13521
rect 11425 13512 11437 13515
rect 11296 13484 11437 13512
rect 11296 13472 11302 13484
rect 11425 13481 11437 13484
rect 11471 13481 11483 13515
rect 11425 13475 11483 13481
rect 16209 13515 16267 13521
rect 16209 13481 16221 13515
rect 16255 13512 16267 13515
rect 16255 13484 17264 13512
rect 16255 13481 16267 13484
rect 16209 13475 16267 13481
rect 10502 13404 10508 13456
rect 10560 13444 10566 13456
rect 10867 13447 10925 13453
rect 10867 13444 10879 13447
rect 10560 13416 10879 13444
rect 10560 13404 10566 13416
rect 10867 13413 10879 13416
rect 10913 13444 10925 13447
rect 11698 13444 11704 13456
rect 10913 13416 11704 13444
rect 10913 13413 10925 13416
rect 10867 13407 10925 13413
rect 11698 13404 11704 13416
rect 11756 13404 11762 13456
rect 15651 13447 15709 13453
rect 15651 13413 15663 13447
rect 15697 13444 15709 13447
rect 15838 13444 15844 13456
rect 15697 13416 15844 13444
rect 15697 13413 15709 13416
rect 15651 13407 15709 13413
rect 15838 13404 15844 13416
rect 15896 13404 15902 13456
rect 17236 13453 17264 13484
rect 17221 13447 17279 13453
rect 17221 13413 17233 13447
rect 17267 13444 17279 13447
rect 17494 13444 17500 13456
rect 17267 13416 17500 13444
rect 17267 13413 17279 13416
rect 17221 13407 17279 13413
rect 17494 13404 17500 13416
rect 17552 13404 17558 13456
rect 5810 13376 5816 13388
rect 5771 13348 5816 13376
rect 5810 13336 5816 13348
rect 5868 13336 5874 13388
rect 6181 13379 6239 13385
rect 6181 13345 6193 13379
rect 6227 13345 6239 13379
rect 6454 13376 6460 13388
rect 6415 13348 6460 13376
rect 6181 13339 6239 13345
rect 6196 13184 6224 13339
rect 6454 13336 6460 13348
rect 6512 13336 6518 13388
rect 6914 13376 6920 13388
rect 6875 13348 6920 13376
rect 6914 13336 6920 13348
rect 6972 13336 6978 13388
rect 10502 13308 10508 13320
rect 10463 13280 10508 13308
rect 10502 13268 10508 13280
rect 10560 13268 10566 13320
rect 15286 13308 15292 13320
rect 15247 13280 15292 13308
rect 15286 13268 15292 13280
rect 15344 13268 15350 13320
rect 17126 13308 17132 13320
rect 17087 13280 17132 13308
rect 17126 13268 17132 13280
rect 17184 13268 17190 13320
rect 17770 13308 17776 13320
rect 17731 13280 17776 13308
rect 17770 13268 17776 13280
rect 17828 13268 17834 13320
rect 6178 13172 6184 13184
rect 6091 13144 6184 13172
rect 6178 13132 6184 13144
rect 6236 13172 6242 13184
rect 7374 13172 7380 13184
rect 6236 13144 7380 13172
rect 6236 13132 6242 13144
rect 7374 13132 7380 13144
rect 7432 13132 7438 13184
rect 8294 13172 8300 13184
rect 8255 13144 8300 13172
rect 8294 13132 8300 13144
rect 8352 13132 8358 13184
rect 10045 13175 10103 13181
rect 10045 13141 10057 13175
rect 10091 13172 10103 13175
rect 10134 13172 10140 13184
rect 10091 13144 10140 13172
rect 10091 13141 10103 13144
rect 10045 13135 10103 13141
rect 10134 13132 10140 13144
rect 10192 13132 10198 13184
rect 13354 13172 13360 13184
rect 13315 13144 13360 13172
rect 13354 13132 13360 13144
rect 13412 13132 13418 13184
rect 13817 13175 13875 13181
rect 13817 13141 13829 13175
rect 13863 13172 13875 13175
rect 14550 13172 14556 13184
rect 13863 13144 14556 13172
rect 13863 13141 13875 13144
rect 13817 13135 13875 13141
rect 14550 13132 14556 13144
rect 14608 13132 14614 13184
rect 1104 13082 22816 13104
rect 1104 13030 4982 13082
rect 5034 13030 5046 13082
rect 5098 13030 5110 13082
rect 5162 13030 5174 13082
rect 5226 13030 12982 13082
rect 13034 13030 13046 13082
rect 13098 13030 13110 13082
rect 13162 13030 13174 13082
rect 13226 13030 20982 13082
rect 21034 13030 21046 13082
rect 21098 13030 21110 13082
rect 21162 13030 21174 13082
rect 21226 13030 22816 13082
rect 1104 13008 22816 13030
rect 5261 12971 5319 12977
rect 5261 12937 5273 12971
rect 5307 12968 5319 12971
rect 6178 12968 6184 12980
rect 5307 12940 6184 12968
rect 5307 12937 5319 12940
rect 5261 12931 5319 12937
rect 6178 12928 6184 12940
rect 6236 12928 6242 12980
rect 10042 12968 10048 12980
rect 7852 12940 10048 12968
rect 7852 12900 7880 12940
rect 10042 12928 10048 12940
rect 10100 12928 10106 12980
rect 16390 12968 16396 12980
rect 16351 12940 16396 12968
rect 16390 12928 16396 12940
rect 16448 12928 16454 12980
rect 17126 12968 17132 12980
rect 17087 12940 17132 12968
rect 17126 12928 17132 12940
rect 17184 12968 17190 12980
rect 17184 12940 18092 12968
rect 17184 12928 17190 12940
rect 13354 12900 13360 12912
rect 7300 12872 7880 12900
rect 9646 12872 13360 12900
rect 5629 12767 5687 12773
rect 5629 12733 5641 12767
rect 5675 12764 5687 12767
rect 5810 12764 5816 12776
rect 5675 12736 5816 12764
rect 5675 12733 5687 12736
rect 5629 12727 5687 12733
rect 5810 12724 5816 12736
rect 5868 12764 5874 12776
rect 6273 12767 6331 12773
rect 6273 12764 6285 12767
rect 5868 12736 6285 12764
rect 5868 12724 5874 12736
rect 6273 12733 6285 12736
rect 6319 12764 6331 12767
rect 7101 12767 7159 12773
rect 7101 12764 7113 12767
rect 6319 12736 7113 12764
rect 6319 12733 6331 12736
rect 6273 12727 6331 12733
rect 7101 12733 7113 12736
rect 7147 12764 7159 12767
rect 7300 12764 7328 12872
rect 7374 12792 7380 12844
rect 7432 12832 7438 12844
rect 9646 12832 9674 12872
rect 13354 12860 13360 12872
rect 13412 12860 13418 12912
rect 17494 12900 17500 12912
rect 17455 12872 17500 12900
rect 17494 12860 17500 12872
rect 17552 12860 17558 12912
rect 7432 12804 9674 12832
rect 7432 12792 7438 12804
rect 7576 12773 7604 12804
rect 10502 12792 10508 12844
rect 10560 12832 10566 12844
rect 11425 12835 11483 12841
rect 11425 12832 11437 12835
rect 10560 12804 11437 12832
rect 10560 12792 10566 12804
rect 11425 12801 11437 12804
rect 11471 12832 11483 12835
rect 12069 12835 12127 12841
rect 12069 12832 12081 12835
rect 11471 12804 12081 12832
rect 11471 12801 11483 12804
rect 11425 12795 11483 12801
rect 12069 12801 12081 12804
rect 12115 12801 12127 12835
rect 12069 12795 12127 12801
rect 14829 12835 14887 12841
rect 14829 12801 14841 12835
rect 14875 12832 14887 12835
rect 15286 12832 15292 12844
rect 14875 12804 15292 12832
rect 14875 12801 14887 12804
rect 14829 12795 14887 12801
rect 15286 12792 15292 12804
rect 15344 12832 15350 12844
rect 18064 12841 18092 12940
rect 15657 12835 15715 12841
rect 15657 12832 15669 12835
rect 15344 12804 15669 12832
rect 15344 12792 15350 12804
rect 15657 12801 15669 12804
rect 15703 12801 15715 12835
rect 15657 12795 15715 12801
rect 18049 12835 18107 12841
rect 18049 12801 18061 12835
rect 18095 12801 18107 12835
rect 18049 12795 18107 12801
rect 7147 12736 7328 12764
rect 7561 12767 7619 12773
rect 7147 12733 7159 12736
rect 7101 12727 7159 12733
rect 7561 12733 7573 12767
rect 7607 12733 7619 12767
rect 7561 12727 7619 12733
rect 7653 12767 7711 12773
rect 7653 12733 7665 12767
rect 7699 12733 7711 12767
rect 8202 12764 8208 12776
rect 8163 12736 8208 12764
rect 7653 12727 7711 12733
rect 7668 12696 7696 12727
rect 8202 12724 8208 12736
rect 8260 12724 8266 12776
rect 10042 12764 10048 12776
rect 10003 12736 10048 12764
rect 10042 12724 10048 12736
rect 10100 12724 10106 12776
rect 10134 12724 10140 12776
rect 10192 12764 10198 12776
rect 10413 12767 10471 12773
rect 10413 12764 10425 12767
rect 10192 12736 10425 12764
rect 10192 12724 10198 12736
rect 10413 12733 10425 12736
rect 10459 12733 10471 12767
rect 10413 12727 10471 12733
rect 10781 12767 10839 12773
rect 10781 12733 10793 12767
rect 10827 12733 10839 12767
rect 11330 12764 11336 12776
rect 11291 12736 11336 12764
rect 10781 12727 10839 12733
rect 9766 12696 9772 12708
rect 6564 12668 9772 12696
rect 6564 12640 6592 12668
rect 9766 12656 9772 12668
rect 9824 12696 9830 12708
rect 10796 12696 10824 12727
rect 11330 12724 11336 12736
rect 11388 12724 11394 12776
rect 13262 12724 13268 12776
rect 13320 12764 13326 12776
rect 13357 12767 13415 12773
rect 13357 12764 13369 12767
rect 13320 12736 13369 12764
rect 13320 12724 13326 12736
rect 13357 12733 13369 12736
rect 13403 12733 13415 12767
rect 13357 12727 13415 12733
rect 13446 12724 13452 12776
rect 13504 12764 13510 12776
rect 13817 12767 13875 12773
rect 13817 12764 13829 12767
rect 13504 12736 13829 12764
rect 13504 12724 13510 12736
rect 13817 12733 13829 12736
rect 13863 12733 13875 12767
rect 14185 12767 14243 12773
rect 14185 12764 14197 12767
rect 13817 12727 13875 12733
rect 13924 12736 14197 12764
rect 9824 12668 10824 12696
rect 9824 12656 9830 12668
rect 12802 12656 12808 12708
rect 12860 12696 12866 12708
rect 12897 12699 12955 12705
rect 12897 12696 12909 12699
rect 12860 12668 12909 12696
rect 12860 12656 12866 12668
rect 12897 12665 12909 12668
rect 12943 12696 12955 12699
rect 13630 12696 13636 12708
rect 12943 12668 13636 12696
rect 12943 12665 12955 12668
rect 12897 12659 12955 12665
rect 13630 12656 13636 12668
rect 13688 12696 13694 12708
rect 13924 12696 13952 12736
rect 14185 12733 14197 12736
rect 14231 12733 14243 12767
rect 14550 12764 14556 12776
rect 14511 12736 14556 12764
rect 14185 12727 14243 12733
rect 14550 12724 14556 12736
rect 14608 12724 14614 12776
rect 15930 12724 15936 12776
rect 15988 12764 15994 12776
rect 16209 12767 16267 12773
rect 16209 12764 16221 12767
rect 15988 12736 16221 12764
rect 15988 12724 15994 12736
rect 16209 12733 16221 12736
rect 16255 12764 16267 12767
rect 16761 12767 16819 12773
rect 16761 12764 16773 12767
rect 16255 12736 16773 12764
rect 16255 12733 16267 12736
rect 16209 12727 16267 12733
rect 16761 12733 16773 12736
rect 16807 12733 16819 12767
rect 16761 12727 16819 12733
rect 13688 12668 13952 12696
rect 13688 12656 13694 12668
rect 4893 12631 4951 12637
rect 4893 12597 4905 12631
rect 4939 12628 4951 12631
rect 5350 12628 5356 12640
rect 4939 12600 5356 12628
rect 4939 12597 4951 12600
rect 4893 12591 4951 12597
rect 5350 12588 5356 12600
rect 5408 12588 5414 12640
rect 6546 12628 6552 12640
rect 6507 12600 6552 12628
rect 6546 12588 6552 12600
rect 6604 12588 6610 12640
rect 7098 12628 7104 12640
rect 7059 12600 7104 12628
rect 7098 12588 7104 12600
rect 7156 12588 7162 12640
rect 9490 12628 9496 12640
rect 9451 12600 9496 12628
rect 9490 12588 9496 12600
rect 9548 12588 9554 12640
rect 11698 12628 11704 12640
rect 11659 12600 11704 12628
rect 11698 12588 11704 12600
rect 11756 12588 11762 12640
rect 13262 12628 13268 12640
rect 13223 12600 13268 12628
rect 13262 12588 13268 12600
rect 13320 12588 13326 12640
rect 15381 12631 15439 12637
rect 15381 12597 15393 12631
rect 15427 12628 15439 12631
rect 15838 12628 15844 12640
rect 15427 12600 15844 12628
rect 15427 12597 15439 12600
rect 15381 12591 15439 12597
rect 15838 12588 15844 12600
rect 15896 12588 15902 12640
rect 1104 12538 22816 12560
rect 1104 12486 8982 12538
rect 9034 12486 9046 12538
rect 9098 12486 9110 12538
rect 9162 12486 9174 12538
rect 9226 12486 16982 12538
rect 17034 12486 17046 12538
rect 17098 12486 17110 12538
rect 17162 12486 17174 12538
rect 17226 12486 22816 12538
rect 1104 12464 22816 12486
rect 7006 12424 7012 12436
rect 6967 12396 7012 12424
rect 7006 12384 7012 12396
rect 7064 12384 7070 12436
rect 10594 12424 10600 12436
rect 10555 12396 10600 12424
rect 10594 12384 10600 12396
rect 10652 12384 10658 12436
rect 12802 12424 12808 12436
rect 12763 12396 12808 12424
rect 12802 12384 12808 12396
rect 12860 12384 12866 12436
rect 15838 12424 15844 12436
rect 15799 12396 15844 12424
rect 15838 12384 15844 12396
rect 15896 12384 15902 12436
rect 16393 12427 16451 12433
rect 16393 12393 16405 12427
rect 16439 12424 16451 12427
rect 17310 12424 17316 12436
rect 16439 12396 17316 12424
rect 16439 12393 16451 12396
rect 16393 12387 16451 12393
rect 17310 12384 17316 12396
rect 17368 12424 17374 12436
rect 17368 12396 17448 12424
rect 17368 12384 17374 12396
rect 6914 12316 6920 12368
rect 6972 12356 6978 12368
rect 7653 12359 7711 12365
rect 7653 12356 7665 12359
rect 6972 12328 7665 12356
rect 6972 12316 6978 12328
rect 5718 12248 5724 12300
rect 5776 12288 5782 12300
rect 5813 12291 5871 12297
rect 5813 12288 5825 12291
rect 5776 12260 5825 12288
rect 5776 12248 5782 12260
rect 5813 12257 5825 12260
rect 5859 12257 5871 12291
rect 6270 12288 6276 12300
rect 6231 12260 6276 12288
rect 5813 12251 5871 12257
rect 6270 12248 6276 12260
rect 6328 12248 6334 12300
rect 6454 12248 6460 12300
rect 6512 12288 6518 12300
rect 7208 12297 7236 12328
rect 7653 12325 7665 12328
rect 7699 12356 7711 12359
rect 8202 12356 8208 12368
rect 7699 12328 8208 12356
rect 7699 12325 7711 12328
rect 7653 12319 7711 12325
rect 8202 12316 8208 12328
rect 8260 12356 8266 12368
rect 8481 12359 8539 12365
rect 8481 12356 8493 12359
rect 8260 12328 8493 12356
rect 8260 12316 8266 12328
rect 8481 12325 8493 12328
rect 8527 12356 8539 12359
rect 9490 12356 9496 12368
rect 8527 12328 9496 12356
rect 8527 12325 8539 12328
rect 8481 12319 8539 12325
rect 9490 12316 9496 12328
rect 9548 12356 9554 12368
rect 17420 12365 17448 12396
rect 17405 12359 17463 12365
rect 9548 12328 11376 12356
rect 9548 12316 9554 12328
rect 11348 12300 11376 12328
rect 17405 12325 17417 12359
rect 17451 12325 17463 12359
rect 17405 12319 17463 12325
rect 6641 12291 6699 12297
rect 6641 12288 6653 12291
rect 6512 12260 6653 12288
rect 6512 12248 6518 12260
rect 6641 12257 6653 12260
rect 6687 12257 6699 12291
rect 6641 12251 6699 12257
rect 7193 12291 7251 12297
rect 7193 12257 7205 12291
rect 7239 12257 7251 12291
rect 10318 12288 10324 12300
rect 10279 12260 10324 12288
rect 7193 12251 7251 12257
rect 10318 12248 10324 12260
rect 10376 12248 10382 12300
rect 10781 12291 10839 12297
rect 10781 12288 10793 12291
rect 10520 12260 10793 12288
rect 5629 12223 5687 12229
rect 5629 12189 5641 12223
rect 5675 12220 5687 12223
rect 6472 12220 6500 12248
rect 5675 12192 6500 12220
rect 5675 12189 5687 12192
rect 5629 12183 5687 12189
rect 10134 12180 10140 12232
rect 10192 12220 10198 12232
rect 10520 12220 10548 12260
rect 10781 12257 10793 12260
rect 10827 12257 10839 12291
rect 10781 12251 10839 12257
rect 11149 12291 11207 12297
rect 11149 12257 11161 12291
rect 11195 12257 11207 12291
rect 11149 12251 11207 12257
rect 10192 12192 10548 12220
rect 10192 12180 10198 12192
rect 10594 12180 10600 12232
rect 10652 12220 10658 12232
rect 11164 12220 11192 12251
rect 11330 12248 11336 12300
rect 11388 12288 11394 12300
rect 11517 12291 11575 12297
rect 11517 12288 11529 12291
rect 11388 12260 11529 12288
rect 11388 12248 11394 12260
rect 11517 12257 11529 12260
rect 11563 12257 11575 12291
rect 11517 12251 11575 12257
rect 13173 12291 13231 12297
rect 13173 12257 13185 12291
rect 13219 12257 13231 12291
rect 13354 12288 13360 12300
rect 13315 12260 13360 12288
rect 13173 12251 13231 12257
rect 10652 12192 11192 12220
rect 13188 12220 13216 12251
rect 13354 12248 13360 12260
rect 13412 12248 13418 12300
rect 13906 12288 13912 12300
rect 13867 12260 13912 12288
rect 13906 12248 13912 12260
rect 13964 12248 13970 12300
rect 14274 12288 14280 12300
rect 14187 12260 14280 12288
rect 14274 12248 14280 12260
rect 14332 12288 14338 12300
rect 14550 12288 14556 12300
rect 14332 12260 14556 12288
rect 14332 12248 14338 12260
rect 14550 12248 14556 12260
rect 14608 12248 14614 12300
rect 18874 12297 18880 12300
rect 18852 12291 18880 12297
rect 18852 12288 18864 12291
rect 18787 12260 18864 12288
rect 18852 12257 18864 12260
rect 18932 12288 18938 12300
rect 20806 12288 20812 12300
rect 18932 12260 20812 12288
rect 18852 12251 18880 12257
rect 18874 12248 18880 12251
rect 18932 12248 18938 12260
rect 20806 12248 20812 12260
rect 20864 12248 20870 12300
rect 13262 12220 13268 12232
rect 13188 12192 13268 12220
rect 10652 12180 10658 12192
rect 13262 12180 13268 12192
rect 13320 12180 13326 12232
rect 14369 12223 14427 12229
rect 14369 12189 14381 12223
rect 14415 12220 14427 12223
rect 15473 12223 15531 12229
rect 15473 12220 15485 12223
rect 14415 12192 15485 12220
rect 14415 12189 14427 12192
rect 14369 12183 14427 12189
rect 15473 12189 15485 12192
rect 15519 12220 15531 12223
rect 16758 12220 16764 12232
rect 15519 12192 16764 12220
rect 15519 12189 15531 12192
rect 15473 12183 15531 12189
rect 16758 12180 16764 12192
rect 16816 12180 16822 12232
rect 17313 12223 17371 12229
rect 17313 12189 17325 12223
rect 17359 12220 17371 12223
rect 17402 12220 17408 12232
rect 17359 12192 17408 12220
rect 17359 12189 17371 12192
rect 17313 12183 17371 12189
rect 17402 12180 17408 12192
rect 17460 12180 17466 12232
rect 17770 12220 17776 12232
rect 17731 12192 17776 12220
rect 17770 12180 17776 12192
rect 17828 12180 17834 12232
rect 8110 12084 8116 12096
rect 8071 12056 8116 12084
rect 8110 12044 8116 12056
rect 8168 12044 8174 12096
rect 10042 12084 10048 12096
rect 10003 12056 10048 12084
rect 10042 12044 10048 12056
rect 10100 12044 10106 12096
rect 12434 12084 12440 12096
rect 12395 12056 12440 12084
rect 12434 12044 12440 12056
rect 12492 12044 12498 12096
rect 18690 12044 18696 12096
rect 18748 12084 18754 12096
rect 18923 12087 18981 12093
rect 18923 12084 18935 12087
rect 18748 12056 18935 12084
rect 18748 12044 18754 12056
rect 18923 12053 18935 12056
rect 18969 12053 18981 12087
rect 18923 12047 18981 12053
rect 1104 11994 22816 12016
rect 1104 11942 4982 11994
rect 5034 11942 5046 11994
rect 5098 11942 5110 11994
rect 5162 11942 5174 11994
rect 5226 11942 12982 11994
rect 13034 11942 13046 11994
rect 13098 11942 13110 11994
rect 13162 11942 13174 11994
rect 13226 11942 20982 11994
rect 21034 11942 21046 11994
rect 21098 11942 21110 11994
rect 21162 11942 21174 11994
rect 21226 11942 22816 11994
rect 1104 11920 22816 11942
rect 1486 11840 1492 11892
rect 1544 11880 1550 11892
rect 1581 11883 1639 11889
rect 1581 11880 1593 11883
rect 1544 11852 1593 11880
rect 1544 11840 1550 11852
rect 1581 11849 1593 11852
rect 1627 11849 1639 11883
rect 1581 11843 1639 11849
rect 5350 11840 5356 11892
rect 5408 11880 5414 11892
rect 5537 11883 5595 11889
rect 5537 11880 5549 11883
rect 5408 11852 5549 11880
rect 5408 11840 5414 11852
rect 5537 11849 5549 11852
rect 5583 11880 5595 11883
rect 6914 11880 6920 11892
rect 5583 11852 6920 11880
rect 5583 11849 5595 11852
rect 5537 11843 5595 11849
rect 6914 11840 6920 11852
rect 6972 11840 6978 11892
rect 9766 11840 9772 11892
rect 9824 11880 9830 11892
rect 10321 11883 10379 11889
rect 10321 11880 10333 11883
rect 9824 11852 10333 11880
rect 9824 11840 9830 11852
rect 10321 11849 10333 11852
rect 10367 11880 10379 11883
rect 10594 11880 10600 11892
rect 10367 11852 10600 11880
rect 10367 11849 10379 11852
rect 10321 11843 10379 11849
rect 10594 11840 10600 11852
rect 10652 11880 10658 11892
rect 12713 11883 12771 11889
rect 12713 11880 12725 11883
rect 10652 11852 12725 11880
rect 10652 11840 10658 11852
rect 12713 11849 12725 11852
rect 12759 11880 12771 11883
rect 12802 11880 12808 11892
rect 12759 11852 12808 11880
rect 12759 11849 12771 11852
rect 12713 11843 12771 11849
rect 12802 11840 12808 11852
rect 12860 11840 12866 11892
rect 13354 11840 13360 11892
rect 13412 11880 13418 11892
rect 14645 11883 14703 11889
rect 14645 11880 14657 11883
rect 13412 11852 14657 11880
rect 13412 11840 13418 11852
rect 14645 11849 14657 11852
rect 14691 11849 14703 11883
rect 16758 11880 16764 11892
rect 16719 11852 16764 11880
rect 14645 11843 14703 11849
rect 16758 11840 16764 11852
rect 16816 11840 16822 11892
rect 17310 11880 17316 11892
rect 17271 11852 17316 11880
rect 17310 11840 17316 11852
rect 17368 11840 17374 11892
rect 18874 11880 18880 11892
rect 18835 11852 18880 11880
rect 18874 11840 18880 11852
rect 18932 11840 18938 11892
rect 8202 11772 8208 11824
rect 8260 11812 8266 11824
rect 8260 11784 8661 11812
rect 8260 11772 8266 11784
rect 7834 11704 7840 11756
rect 7892 11744 7898 11756
rect 7892 11716 8524 11744
rect 7892 11704 7898 11716
rect 106 11636 112 11688
rect 164 11676 170 11688
rect 1397 11679 1455 11685
rect 1397 11676 1409 11679
rect 164 11648 1409 11676
rect 164 11636 170 11648
rect 1397 11645 1409 11648
rect 1443 11676 1455 11679
rect 1946 11676 1952 11688
rect 1443 11648 1952 11676
rect 1443 11645 1455 11648
rect 1397 11639 1455 11645
rect 1946 11636 1952 11648
rect 2004 11636 2010 11688
rect 6454 11636 6460 11688
rect 6512 11676 6518 11688
rect 6641 11679 6699 11685
rect 6641 11676 6653 11679
rect 6512 11648 6653 11676
rect 6512 11636 6518 11648
rect 6641 11645 6653 11648
rect 6687 11676 6699 11679
rect 7561 11679 7619 11685
rect 7561 11676 7573 11679
rect 6687 11648 7573 11676
rect 6687 11645 6699 11648
rect 6641 11639 6699 11645
rect 7561 11645 7573 11648
rect 7607 11676 7619 11679
rect 8202 11676 8208 11688
rect 7607 11648 8208 11676
rect 7607 11645 7619 11648
rect 7561 11639 7619 11645
rect 8202 11636 8208 11648
rect 8260 11636 8266 11688
rect 8496 11685 8524 11716
rect 8297 11679 8355 11685
rect 8297 11645 8309 11679
rect 8343 11645 8355 11679
rect 8297 11639 8355 11645
rect 8481 11679 8539 11685
rect 8481 11645 8493 11679
rect 8527 11645 8539 11679
rect 8633 11676 8661 11784
rect 9490 11744 9496 11756
rect 9416 11716 9496 11744
rect 9416 11685 9444 11716
rect 9490 11704 9496 11716
rect 9548 11704 9554 11756
rect 8849 11679 8907 11685
rect 8849 11676 8861 11679
rect 8633 11648 8861 11676
rect 8481 11639 8539 11645
rect 8849 11645 8861 11648
rect 8895 11645 8907 11679
rect 8849 11639 8907 11645
rect 9401 11679 9459 11685
rect 9401 11645 9413 11679
rect 9447 11645 9459 11679
rect 9401 11639 9459 11645
rect 8110 11568 8116 11620
rect 8168 11608 8174 11620
rect 8312 11608 8340 11639
rect 9582 11636 9588 11688
rect 9640 11676 9646 11688
rect 10042 11676 10048 11688
rect 9640 11648 10048 11676
rect 9640 11636 9646 11648
rect 10042 11636 10048 11648
rect 10100 11676 10106 11688
rect 11333 11679 11391 11685
rect 11333 11676 11345 11679
rect 10100 11648 11345 11676
rect 10100 11636 10106 11648
rect 11333 11645 11345 11648
rect 11379 11645 11391 11679
rect 11514 11676 11520 11688
rect 11427 11648 11520 11676
rect 11333 11639 11391 11645
rect 9490 11608 9496 11620
rect 8168 11580 9496 11608
rect 8168 11568 8174 11580
rect 9490 11568 9496 11580
rect 9548 11568 9554 11620
rect 11348 11608 11376 11639
rect 11514 11636 11520 11648
rect 11572 11676 11578 11688
rect 13173 11679 13231 11685
rect 13173 11676 13185 11679
rect 11572 11648 13185 11676
rect 11572 11636 11578 11648
rect 13173 11645 13185 11648
rect 13219 11676 13231 11679
rect 13262 11676 13268 11688
rect 13219 11648 13268 11676
rect 13219 11645 13231 11648
rect 13173 11639 13231 11645
rect 13262 11636 13268 11648
rect 13320 11636 13326 11688
rect 13357 11679 13415 11685
rect 13357 11645 13369 11679
rect 13403 11645 13415 11679
rect 13357 11639 13415 11645
rect 13078 11608 13084 11620
rect 11348 11580 13084 11608
rect 13078 11568 13084 11580
rect 13136 11568 13142 11620
rect 5718 11500 5724 11552
rect 5776 11540 5782 11552
rect 5813 11543 5871 11549
rect 5813 11540 5825 11543
rect 5776 11512 5825 11540
rect 5776 11500 5782 11512
rect 5813 11509 5825 11512
rect 5859 11509 5871 11543
rect 6270 11540 6276 11552
rect 6231 11512 6276 11540
rect 5813 11503 5871 11509
rect 6270 11500 6276 11512
rect 6328 11500 6334 11552
rect 7834 11540 7840 11552
rect 7795 11512 7840 11540
rect 7834 11500 7840 11512
rect 7892 11500 7898 11552
rect 8294 11540 8300 11552
rect 8255 11512 8300 11540
rect 8294 11500 8300 11512
rect 8352 11500 8358 11552
rect 10134 11500 10140 11552
rect 10192 11540 10198 11552
rect 11793 11543 11851 11549
rect 11793 11540 11805 11543
rect 10192 11512 11805 11540
rect 10192 11500 10198 11512
rect 11793 11509 11805 11512
rect 11839 11540 11851 11543
rect 12161 11543 12219 11549
rect 12161 11540 12173 11543
rect 11839 11512 12173 11540
rect 11839 11509 11851 11512
rect 11793 11503 11851 11509
rect 12161 11509 12173 11512
rect 12207 11540 12219 11543
rect 12342 11540 12348 11552
rect 12207 11512 12348 11540
rect 12207 11509 12219 11512
rect 12161 11503 12219 11509
rect 12342 11500 12348 11512
rect 12400 11540 12406 11552
rect 13372 11540 13400 11639
rect 13630 11636 13636 11688
rect 13688 11676 13694 11688
rect 13725 11679 13783 11685
rect 13725 11676 13737 11679
rect 13688 11648 13737 11676
rect 13688 11636 13694 11648
rect 13725 11645 13737 11648
rect 13771 11645 13783 11679
rect 14274 11676 14280 11688
rect 14235 11648 14280 11676
rect 13725 11639 13783 11645
rect 14274 11636 14280 11648
rect 14332 11636 14338 11688
rect 14369 11679 14427 11685
rect 14369 11645 14381 11679
rect 14415 11676 14427 11679
rect 15562 11676 15568 11688
rect 14415 11648 15568 11676
rect 14415 11645 14427 11648
rect 14369 11639 14427 11645
rect 15562 11636 15568 11648
rect 15620 11636 15626 11688
rect 14292 11608 14320 11636
rect 15838 11608 15844 11620
rect 13740 11580 14320 11608
rect 15396 11580 15844 11608
rect 13740 11552 13768 11580
rect 12400 11512 13400 11540
rect 12400 11500 12406 11512
rect 13722 11500 13728 11552
rect 13780 11500 13786 11552
rect 15102 11540 15108 11552
rect 15063 11512 15108 11540
rect 15102 11500 15108 11512
rect 15160 11540 15166 11552
rect 15396 11549 15424 11580
rect 15838 11568 15844 11580
rect 15896 11617 15902 11620
rect 15896 11611 15944 11617
rect 15896 11577 15898 11611
rect 15932 11577 15944 11611
rect 15896 11571 15944 11577
rect 15896 11568 15902 11571
rect 15381 11543 15439 11549
rect 15381 11540 15393 11543
rect 15160 11512 15393 11540
rect 15160 11500 15166 11512
rect 15381 11509 15393 11512
rect 15427 11509 15439 11543
rect 16482 11540 16488 11552
rect 16443 11512 16488 11540
rect 15381 11503 15439 11509
rect 16482 11500 16488 11512
rect 16540 11500 16546 11552
rect 17402 11500 17408 11552
rect 17460 11540 17466 11552
rect 17681 11543 17739 11549
rect 17681 11540 17693 11543
rect 17460 11512 17693 11540
rect 17460 11500 17466 11512
rect 17681 11509 17693 11512
rect 17727 11540 17739 11543
rect 18966 11540 18972 11552
rect 17727 11512 18972 11540
rect 17727 11509 17739 11512
rect 17681 11503 17739 11509
rect 18966 11500 18972 11512
rect 19024 11500 19030 11552
rect 1104 11450 22816 11472
rect 1104 11398 8982 11450
rect 9034 11398 9046 11450
rect 9098 11398 9110 11450
rect 9162 11398 9174 11450
rect 9226 11398 16982 11450
rect 17034 11398 17046 11450
rect 17098 11398 17110 11450
rect 17162 11398 17174 11450
rect 17226 11398 22816 11450
rect 1104 11376 22816 11398
rect 5534 11336 5540 11348
rect 5495 11308 5540 11336
rect 5534 11296 5540 11308
rect 5592 11296 5598 11348
rect 10042 11336 10048 11348
rect 10003 11308 10048 11336
rect 10042 11296 10048 11308
rect 10100 11296 10106 11348
rect 15470 11336 15476 11348
rect 15431 11308 15476 11336
rect 15470 11296 15476 11308
rect 15528 11296 15534 11348
rect 15562 11296 15568 11348
rect 15620 11336 15626 11348
rect 16209 11339 16267 11345
rect 16209 11336 16221 11339
rect 15620 11308 16221 11336
rect 15620 11296 15626 11308
rect 16209 11305 16221 11308
rect 16255 11305 16267 11339
rect 16209 11299 16267 11305
rect 8018 11228 8024 11280
rect 8076 11268 8082 11280
rect 8199 11271 8257 11277
rect 8199 11268 8211 11271
rect 8076 11240 8211 11268
rect 8076 11228 8082 11240
rect 8199 11237 8211 11240
rect 8245 11268 8257 11271
rect 9950 11268 9956 11280
rect 8245 11240 9956 11268
rect 8245 11237 8257 11240
rect 8199 11231 8257 11237
rect 9950 11228 9956 11240
rect 10008 11228 10014 11280
rect 10318 11268 10324 11280
rect 10060 11240 10324 11268
rect 5718 11200 5724 11212
rect 5679 11172 5724 11200
rect 5718 11160 5724 11172
rect 5776 11160 5782 11212
rect 6178 11200 6184 11212
rect 6139 11172 6184 11200
rect 6178 11160 6184 11172
rect 6236 11160 6242 11212
rect 6454 11200 6460 11212
rect 6415 11172 6460 11200
rect 6454 11160 6460 11172
rect 6512 11160 6518 11212
rect 6638 11200 6644 11212
rect 6599 11172 6644 11200
rect 6638 11160 6644 11172
rect 6696 11160 6702 11212
rect 9490 11200 9496 11212
rect 9403 11172 9496 11200
rect 9490 11160 9496 11172
rect 9548 11200 9554 11212
rect 10060 11209 10088 11240
rect 10318 11228 10324 11240
rect 10376 11268 10382 11280
rect 11514 11268 11520 11280
rect 10376 11240 11520 11268
rect 10376 11228 10382 11240
rect 11514 11228 11520 11240
rect 11572 11228 11578 11280
rect 16482 11228 16488 11280
rect 16540 11268 16546 11280
rect 17126 11268 17132 11280
rect 16540 11240 17132 11268
rect 16540 11228 16546 11240
rect 17126 11228 17132 11240
rect 17184 11268 17190 11280
rect 17221 11271 17279 11277
rect 17221 11268 17233 11271
rect 17184 11240 17233 11268
rect 17184 11228 17190 11240
rect 17221 11237 17233 11240
rect 17267 11237 17279 11271
rect 17770 11268 17776 11280
rect 17731 11240 17776 11268
rect 17221 11231 17279 11237
rect 17770 11228 17776 11240
rect 17828 11228 17834 11280
rect 18690 11268 18696 11280
rect 18651 11240 18696 11268
rect 18690 11228 18696 11240
rect 18748 11228 18754 11280
rect 18785 11271 18843 11277
rect 18785 11237 18797 11271
rect 18831 11268 18843 11271
rect 18874 11268 18880 11280
rect 18831 11240 18880 11268
rect 18831 11237 18843 11240
rect 18785 11231 18843 11237
rect 18874 11228 18880 11240
rect 18932 11228 18938 11280
rect 10045 11203 10103 11209
rect 10045 11200 10057 11203
rect 9548 11172 10057 11200
rect 9548 11160 9554 11172
rect 10045 11169 10057 11172
rect 10091 11169 10103 11203
rect 10045 11163 10103 11169
rect 10134 11160 10140 11212
rect 10192 11200 10198 11212
rect 10229 11203 10287 11209
rect 10229 11200 10241 11203
rect 10192 11172 10241 11200
rect 10192 11160 10198 11172
rect 10229 11169 10241 11172
rect 10275 11169 10287 11203
rect 10594 11200 10600 11212
rect 10555 11172 10600 11200
rect 10229 11163 10287 11169
rect 10594 11160 10600 11172
rect 10652 11160 10658 11212
rect 10965 11203 11023 11209
rect 10965 11169 10977 11203
rect 11011 11169 11023 11203
rect 10965 11163 11023 11169
rect 7837 11135 7895 11141
rect 7837 11101 7849 11135
rect 7883 11101 7895 11135
rect 7837 11095 7895 11101
rect 7745 10999 7803 11005
rect 7745 10965 7757 10999
rect 7791 10996 7803 10999
rect 7852 10996 7880 11095
rect 8846 11092 8852 11144
rect 8904 11132 8910 11144
rect 10980 11132 11008 11163
rect 13998 11160 14004 11212
rect 14056 11200 14062 11212
rect 15194 11200 15200 11212
rect 14056 11172 15200 11200
rect 14056 11160 14062 11172
rect 15194 11160 15200 11172
rect 15252 11200 15258 11212
rect 15289 11203 15347 11209
rect 15289 11200 15301 11203
rect 15252 11172 15301 11200
rect 15252 11160 15258 11172
rect 15289 11169 15301 11172
rect 15335 11169 15347 11203
rect 15289 11163 15347 11169
rect 8904 11104 11008 11132
rect 12989 11135 13047 11141
rect 8904 11092 8910 11104
rect 12989 11101 13001 11135
rect 13035 11132 13047 11135
rect 13262 11132 13268 11144
rect 13035 11104 13268 11132
rect 13035 11101 13047 11104
rect 12989 11095 13047 11101
rect 13262 11092 13268 11104
rect 13320 11092 13326 11144
rect 17129 11135 17187 11141
rect 17129 11101 17141 11135
rect 17175 11132 17187 11135
rect 17402 11132 17408 11144
rect 17175 11104 17408 11132
rect 17175 11101 17187 11104
rect 17129 11095 17187 11101
rect 17402 11092 17408 11104
rect 17460 11092 17466 11144
rect 18966 11132 18972 11144
rect 18927 11104 18972 11132
rect 18966 11092 18972 11104
rect 19024 11092 19030 11144
rect 12253 11067 12311 11073
rect 12253 11033 12265 11067
rect 12299 11064 12311 11067
rect 12434 11064 12440 11076
rect 12299 11036 12440 11064
rect 12299 11033 12311 11036
rect 12253 11027 12311 11033
rect 12434 11024 12440 11036
rect 12492 11064 12498 11076
rect 12621 11067 12679 11073
rect 12621 11064 12633 11067
rect 12492 11036 12633 11064
rect 12492 11024 12498 11036
rect 12621 11033 12633 11036
rect 12667 11064 12679 11067
rect 13722 11064 13728 11076
rect 12667 11036 13728 11064
rect 12667 11033 12679 11036
rect 12621 11027 12679 11033
rect 13722 11024 13728 11036
rect 13780 11024 13786 11076
rect 7926 10996 7932 11008
rect 7791 10968 7932 10996
rect 7791 10965 7803 10968
rect 7745 10959 7803 10965
rect 7926 10956 7932 10968
rect 7984 10956 7990 11008
rect 8754 10996 8760 11008
rect 8715 10968 8760 10996
rect 8754 10956 8760 10968
rect 8812 10956 8818 11008
rect 12342 10956 12348 11008
rect 12400 10996 12406 11008
rect 13265 10999 13323 11005
rect 13265 10996 13277 10999
rect 12400 10968 13277 10996
rect 12400 10956 12406 10968
rect 13265 10965 13277 10968
rect 13311 10965 13323 10999
rect 13265 10959 13323 10965
rect 13354 10956 13360 11008
rect 13412 10996 13418 11008
rect 13633 10999 13691 11005
rect 13633 10996 13645 10999
rect 13412 10968 13645 10996
rect 13412 10956 13418 10968
rect 13633 10965 13645 10968
rect 13679 10965 13691 10999
rect 15838 10996 15844 11008
rect 15799 10968 15844 10996
rect 13633 10959 13691 10965
rect 15838 10956 15844 10968
rect 15896 10956 15902 11008
rect 18138 10996 18144 11008
rect 18099 10968 18144 10996
rect 18138 10956 18144 10968
rect 18196 10956 18202 11008
rect 1104 10906 22816 10928
rect 1104 10854 4982 10906
rect 5034 10854 5046 10906
rect 5098 10854 5110 10906
rect 5162 10854 5174 10906
rect 5226 10854 12982 10906
rect 13034 10854 13046 10906
rect 13098 10854 13110 10906
rect 13162 10854 13174 10906
rect 13226 10854 20982 10906
rect 21034 10854 21046 10906
rect 21098 10854 21110 10906
rect 21162 10854 21174 10906
rect 21226 10854 22816 10906
rect 1104 10832 22816 10854
rect 1946 10792 1952 10804
rect 1907 10764 1952 10792
rect 1946 10752 1952 10764
rect 2004 10752 2010 10804
rect 5169 10795 5227 10801
rect 5169 10761 5181 10795
rect 5215 10792 5227 10795
rect 6638 10792 6644 10804
rect 5215 10764 6644 10792
rect 5215 10761 5227 10764
rect 5169 10755 5227 10761
rect 6638 10752 6644 10764
rect 6696 10752 6702 10804
rect 12802 10752 12808 10804
rect 12860 10792 12866 10804
rect 12897 10795 12955 10801
rect 12897 10792 12909 10795
rect 12860 10764 12909 10792
rect 12860 10752 12866 10764
rect 12897 10761 12909 10764
rect 12943 10761 12955 10795
rect 15194 10792 15200 10804
rect 15155 10764 15200 10792
rect 12897 10755 12955 10761
rect 5905 10727 5963 10733
rect 5905 10693 5917 10727
rect 5951 10724 5963 10727
rect 6178 10724 6184 10736
rect 5951 10696 6184 10724
rect 5951 10693 5963 10696
rect 5905 10687 5963 10693
rect 6178 10684 6184 10696
rect 6236 10684 6242 10736
rect 6273 10727 6331 10733
rect 6273 10693 6285 10727
rect 6319 10724 6331 10727
rect 6454 10724 6460 10736
rect 6319 10696 6460 10724
rect 6319 10693 6331 10696
rect 6273 10687 6331 10693
rect 6454 10684 6460 10696
rect 6512 10684 6518 10736
rect 6546 10684 6552 10736
rect 6604 10724 6610 10736
rect 9769 10727 9827 10733
rect 9769 10724 9781 10727
rect 6604 10696 9781 10724
rect 6604 10684 6610 10696
rect 9769 10693 9781 10696
rect 9815 10693 9827 10727
rect 9769 10687 9827 10693
rect 8294 10616 8300 10668
rect 8352 10656 8358 10668
rect 8352 10628 8708 10656
rect 8352 10616 8358 10628
rect 1556 10591 1614 10597
rect 1556 10557 1568 10591
rect 1602 10588 1614 10591
rect 1946 10588 1952 10600
rect 1602 10560 1952 10588
rect 1602 10557 1614 10560
rect 1556 10551 1614 10557
rect 1946 10548 1952 10560
rect 2004 10548 2010 10600
rect 5537 10591 5595 10597
rect 5537 10557 5549 10591
rect 5583 10588 5595 10591
rect 5718 10588 5724 10600
rect 5583 10560 5724 10588
rect 5583 10557 5595 10560
rect 5537 10551 5595 10557
rect 5718 10548 5724 10560
rect 5776 10548 5782 10600
rect 7377 10591 7435 10597
rect 7377 10557 7389 10591
rect 7423 10588 7435 10591
rect 8110 10588 8116 10600
rect 7423 10560 8116 10588
rect 7423 10557 7435 10560
rect 7377 10551 7435 10557
rect 8110 10548 8116 10560
rect 8168 10548 8174 10600
rect 8680 10597 8708 10628
rect 10042 10616 10048 10668
rect 10100 10656 10106 10668
rect 10229 10659 10287 10665
rect 10229 10656 10241 10659
rect 10100 10628 10241 10656
rect 10100 10616 10106 10628
rect 10229 10625 10241 10628
rect 10275 10656 10287 10659
rect 11793 10659 11851 10665
rect 11793 10656 11805 10659
rect 10275 10628 11805 10656
rect 10275 10625 10287 10628
rect 10229 10619 10287 10625
rect 11793 10625 11805 10628
rect 11839 10625 11851 10659
rect 12912 10656 12940 10755
rect 15194 10752 15200 10764
rect 15252 10752 15258 10804
rect 17126 10792 17132 10804
rect 17087 10764 17132 10792
rect 17126 10752 17132 10764
rect 17184 10752 17190 10804
rect 17402 10792 17408 10804
rect 17363 10764 17408 10792
rect 17402 10752 17408 10764
rect 17460 10752 17466 10804
rect 18690 10752 18696 10804
rect 18748 10792 18754 10804
rect 19429 10795 19487 10801
rect 19429 10792 19441 10795
rect 18748 10764 19441 10792
rect 18748 10752 18754 10764
rect 19429 10761 19441 10764
rect 19475 10761 19487 10795
rect 19429 10755 19487 10761
rect 13170 10684 13176 10736
rect 13228 10724 13234 10736
rect 15102 10724 15108 10736
rect 13228 10696 15108 10724
rect 13228 10684 13234 10696
rect 15102 10684 15108 10696
rect 15160 10684 15166 10736
rect 14553 10659 14611 10665
rect 12912 10628 13814 10656
rect 11793 10619 11851 10625
rect 8573 10591 8631 10597
rect 8573 10557 8585 10591
rect 8619 10557 8631 10591
rect 8573 10551 8631 10557
rect 8665 10591 8723 10597
rect 8665 10557 8677 10591
rect 8711 10557 8723 10591
rect 8665 10551 8723 10557
rect 6270 10480 6276 10532
rect 6328 10520 6334 10532
rect 7745 10523 7803 10529
rect 7745 10520 7757 10523
rect 6328 10492 7757 10520
rect 6328 10480 6334 10492
rect 7745 10489 7757 10492
rect 7791 10520 7803 10523
rect 7834 10520 7840 10532
rect 7791 10492 7840 10520
rect 7791 10489 7803 10492
rect 7745 10483 7803 10489
rect 7834 10480 7840 10492
rect 7892 10520 7898 10532
rect 8588 10520 8616 10551
rect 8846 10548 8852 10600
rect 8904 10588 8910 10600
rect 9033 10591 9091 10597
rect 9033 10588 9045 10591
rect 8904 10560 9045 10588
rect 8904 10548 8910 10560
rect 9033 10557 9045 10560
rect 9079 10557 9091 10591
rect 10134 10588 10140 10600
rect 9033 10551 9091 10557
rect 9692 10560 10140 10588
rect 9692 10532 9720 10560
rect 10134 10548 10140 10560
rect 10192 10548 10198 10600
rect 12253 10591 12311 10597
rect 12253 10557 12265 10591
rect 12299 10588 12311 10591
rect 13354 10588 13360 10600
rect 12299 10560 13360 10588
rect 12299 10557 12311 10560
rect 12253 10551 12311 10557
rect 13354 10548 13360 10560
rect 13412 10548 13418 10600
rect 13541 10591 13599 10597
rect 13541 10557 13553 10591
rect 13587 10557 13599 10591
rect 13786 10588 13814 10628
rect 14553 10625 14565 10659
rect 14599 10656 14611 10659
rect 15381 10659 15439 10665
rect 15381 10656 15393 10659
rect 14599 10628 15393 10656
rect 14599 10625 14611 10628
rect 14553 10619 14611 10625
rect 15381 10625 15393 10628
rect 15427 10656 15439 10659
rect 15838 10656 15844 10668
rect 15427 10628 15844 10656
rect 15427 10625 15439 10628
rect 15381 10619 15439 10625
rect 15838 10616 15844 10628
rect 15896 10616 15902 10668
rect 17420 10656 17448 10752
rect 21085 10727 21143 10733
rect 21085 10693 21097 10727
rect 21131 10724 21143 10727
rect 21358 10724 21364 10736
rect 21131 10696 21364 10724
rect 21131 10693 21143 10696
rect 21085 10687 21143 10693
rect 21358 10684 21364 10696
rect 21416 10684 21422 10736
rect 18322 10656 18328 10668
rect 17420 10628 18328 10656
rect 18322 10616 18328 10628
rect 18380 10656 18386 10668
rect 18417 10659 18475 10665
rect 18417 10656 18429 10659
rect 18380 10628 18429 10656
rect 18380 10616 18386 10628
rect 18417 10625 18429 10628
rect 18463 10625 18475 10659
rect 18417 10619 18475 10625
rect 13906 10588 13912 10600
rect 13786 10560 13912 10588
rect 13541 10551 13599 10557
rect 9674 10520 9680 10532
rect 7892 10492 9680 10520
rect 7892 10480 7898 10492
rect 9674 10480 9680 10492
rect 9732 10480 9738 10532
rect 10042 10480 10048 10532
rect 10100 10520 10106 10532
rect 10591 10523 10649 10529
rect 10591 10520 10603 10523
rect 10100 10492 10603 10520
rect 10100 10480 10106 10492
rect 10591 10489 10603 10492
rect 10637 10520 10649 10523
rect 10637 10492 11560 10520
rect 10637 10489 10649 10492
rect 10591 10483 10649 10489
rect 1627 10455 1685 10461
rect 1627 10421 1639 10455
rect 1673 10452 1685 10455
rect 3326 10452 3332 10464
rect 1673 10424 3332 10452
rect 1673 10421 1685 10424
rect 1627 10415 1685 10421
rect 3326 10412 3332 10424
rect 3384 10412 3390 10464
rect 4338 10452 4344 10464
rect 4299 10424 4344 10452
rect 4338 10412 4344 10424
rect 4396 10412 4402 10464
rect 7926 10452 7932 10464
rect 7887 10424 7932 10452
rect 7926 10412 7932 10424
rect 7984 10412 7990 10464
rect 11146 10452 11152 10464
rect 11107 10424 11152 10452
rect 11146 10412 11152 10424
rect 11204 10412 11210 10464
rect 11532 10461 11560 10492
rect 12342 10480 12348 10532
rect 12400 10520 12406 10532
rect 13556 10520 13584 10551
rect 13906 10548 13912 10560
rect 13964 10548 13970 10600
rect 14274 10588 14280 10600
rect 14235 10560 14280 10588
rect 14274 10548 14280 10560
rect 14332 10548 14338 10600
rect 16301 10591 16359 10597
rect 16301 10557 16313 10591
rect 16347 10588 16359 10591
rect 17773 10591 17831 10597
rect 17773 10588 17785 10591
rect 16347 10560 17785 10588
rect 16347 10557 16359 10560
rect 16301 10551 16359 10557
rect 17773 10557 17785 10560
rect 17819 10557 17831 10591
rect 17773 10551 17831 10557
rect 12400 10492 13584 10520
rect 14921 10523 14979 10529
rect 12400 10480 12406 10492
rect 14921 10489 14933 10523
rect 14967 10520 14979 10523
rect 15102 10520 15108 10532
rect 14967 10492 15108 10520
rect 14967 10489 14979 10492
rect 14921 10483 14979 10489
rect 15102 10480 15108 10492
rect 15160 10520 15166 10532
rect 15470 10520 15476 10532
rect 15160 10492 15476 10520
rect 15160 10480 15166 10492
rect 15470 10480 15476 10492
rect 15528 10520 15534 10532
rect 15702 10523 15760 10529
rect 15702 10520 15714 10523
rect 15528 10492 15714 10520
rect 15528 10480 15534 10492
rect 15702 10489 15714 10492
rect 15748 10489 15760 10523
rect 15702 10483 15760 10489
rect 11517 10455 11575 10461
rect 11517 10421 11529 10455
rect 11563 10452 11575 10455
rect 11698 10452 11704 10464
rect 11563 10424 11704 10452
rect 11563 10421 11575 10424
rect 11517 10415 11575 10421
rect 11698 10412 11704 10424
rect 11756 10452 11762 10464
rect 13170 10452 13176 10464
rect 11756 10424 13176 10452
rect 11756 10412 11762 10424
rect 13170 10412 13176 10424
rect 13228 10412 13234 10464
rect 17788 10452 17816 10551
rect 20070 10548 20076 10600
rect 20128 10588 20134 10600
rect 20901 10591 20959 10597
rect 20901 10588 20913 10591
rect 20128 10560 20913 10588
rect 20128 10548 20134 10560
rect 20901 10557 20913 10560
rect 20947 10588 20959 10591
rect 21453 10591 21511 10597
rect 21453 10588 21465 10591
rect 20947 10560 21465 10588
rect 20947 10557 20959 10560
rect 20901 10551 20959 10557
rect 21453 10557 21465 10560
rect 21499 10557 21511 10591
rect 21453 10551 21511 10557
rect 18138 10520 18144 10532
rect 18099 10492 18144 10520
rect 18138 10480 18144 10492
rect 18196 10480 18202 10532
rect 18233 10523 18291 10529
rect 18233 10489 18245 10523
rect 18279 10489 18291 10523
rect 18233 10483 18291 10489
rect 18248 10452 18276 10483
rect 18874 10452 18880 10464
rect 17788 10424 18880 10452
rect 18874 10412 18880 10424
rect 18932 10452 18938 10464
rect 19061 10455 19119 10461
rect 19061 10452 19073 10455
rect 18932 10424 19073 10452
rect 18932 10412 18938 10424
rect 19061 10421 19073 10424
rect 19107 10421 19119 10455
rect 19061 10415 19119 10421
rect 1104 10362 22816 10384
rect 1104 10310 8982 10362
rect 9034 10310 9046 10362
rect 9098 10310 9110 10362
rect 9162 10310 9174 10362
rect 9226 10310 16982 10362
rect 17034 10310 17046 10362
rect 17098 10310 17110 10362
rect 17162 10310 17174 10362
rect 17226 10310 22816 10362
rect 1104 10288 22816 10310
rect 7929 10251 7987 10257
rect 7929 10217 7941 10251
rect 7975 10248 7987 10251
rect 8018 10248 8024 10260
rect 7975 10220 8024 10248
rect 7975 10217 7987 10220
rect 7929 10211 7987 10217
rect 8018 10208 8024 10220
rect 8076 10208 8082 10260
rect 9490 10248 9496 10260
rect 9451 10220 9496 10248
rect 9490 10208 9496 10220
rect 9548 10208 9554 10260
rect 13722 10208 13728 10260
rect 13780 10248 13786 10260
rect 14093 10251 14151 10257
rect 14093 10248 14105 10251
rect 13780 10220 14105 10248
rect 13780 10208 13786 10220
rect 14093 10217 14105 10220
rect 14139 10248 14151 10251
rect 14274 10248 14280 10260
rect 14139 10220 14280 10248
rect 14139 10217 14151 10220
rect 14093 10211 14151 10217
rect 14274 10208 14280 10220
rect 14332 10208 14338 10260
rect 18138 10208 18144 10260
rect 18196 10248 18202 10260
rect 19291 10251 19349 10257
rect 19291 10248 19303 10251
rect 18196 10220 19303 10248
rect 18196 10208 18202 10220
rect 19291 10217 19303 10220
rect 19337 10217 19349 10251
rect 19291 10211 19349 10217
rect 3786 10140 3792 10192
rect 3844 10180 3850 10192
rect 4427 10183 4485 10189
rect 4427 10180 4439 10183
rect 3844 10152 4439 10180
rect 3844 10140 3850 10152
rect 4427 10149 4439 10152
rect 4473 10180 4485 10183
rect 5442 10180 5448 10192
rect 4473 10152 5448 10180
rect 4473 10149 4485 10152
rect 4427 10143 4485 10149
rect 5442 10140 5448 10152
rect 5500 10140 5506 10192
rect 5902 10140 5908 10192
rect 5960 10180 5966 10192
rect 6178 10180 6184 10192
rect 5960 10152 6184 10180
rect 5960 10140 5966 10152
rect 6178 10140 6184 10152
rect 6236 10180 6242 10192
rect 10321 10183 10379 10189
rect 6236 10152 6408 10180
rect 6236 10140 6242 10152
rect 3694 10072 3700 10124
rect 3752 10112 3758 10124
rect 4065 10115 4123 10121
rect 4065 10112 4077 10115
rect 3752 10084 4077 10112
rect 3752 10072 3758 10084
rect 4065 10081 4077 10084
rect 4111 10112 4123 10115
rect 5534 10112 5540 10124
rect 4111 10084 5540 10112
rect 4111 10081 4123 10084
rect 4065 10075 4123 10081
rect 5534 10072 5540 10084
rect 5592 10072 5598 10124
rect 5718 10072 5724 10124
rect 5776 10112 5782 10124
rect 6089 10115 6147 10121
rect 6089 10112 6101 10115
rect 5776 10084 6101 10112
rect 5776 10072 5782 10084
rect 6089 10081 6101 10084
rect 6135 10112 6147 10115
rect 6270 10112 6276 10124
rect 6135 10084 6276 10112
rect 6135 10081 6147 10084
rect 6089 10075 6147 10081
rect 6270 10072 6276 10084
rect 6328 10072 6334 10124
rect 6380 10121 6408 10152
rect 10321 10149 10333 10183
rect 10367 10180 10379 10183
rect 10594 10180 10600 10192
rect 10367 10152 10600 10180
rect 10367 10149 10379 10152
rect 10321 10143 10379 10149
rect 10594 10140 10600 10152
rect 10652 10180 10658 10192
rect 11146 10180 11152 10192
rect 10652 10152 11152 10180
rect 10652 10140 10658 10152
rect 11146 10140 11152 10152
rect 11204 10140 11210 10192
rect 12989 10183 13047 10189
rect 12989 10149 13001 10183
rect 13035 10180 13047 10183
rect 13446 10180 13452 10192
rect 13035 10152 13452 10180
rect 13035 10149 13047 10152
rect 12989 10143 13047 10149
rect 13446 10140 13452 10152
rect 13504 10140 13510 10192
rect 16206 10180 16212 10192
rect 16167 10152 16212 10180
rect 16206 10140 16212 10152
rect 16264 10140 16270 10192
rect 17770 10180 17776 10192
rect 17731 10152 17776 10180
rect 17770 10140 17776 10152
rect 17828 10140 17834 10192
rect 18322 10180 18328 10192
rect 18283 10152 18328 10180
rect 18322 10140 18328 10152
rect 18380 10140 18386 10192
rect 6365 10115 6423 10121
rect 6365 10081 6377 10115
rect 6411 10081 6423 10115
rect 6365 10075 6423 10081
rect 6546 10072 6552 10124
rect 6604 10112 6610 10124
rect 6641 10115 6699 10121
rect 6641 10112 6653 10115
rect 6604 10084 6653 10112
rect 6604 10072 6610 10084
rect 6641 10081 6653 10084
rect 6687 10081 6699 10115
rect 6641 10075 6699 10081
rect 6730 10072 6736 10124
rect 6788 10112 6794 10124
rect 7009 10115 7067 10121
rect 7009 10112 7021 10115
rect 6788 10084 7021 10112
rect 6788 10072 6794 10084
rect 7009 10081 7021 10084
rect 7055 10112 7067 10115
rect 8573 10115 8631 10121
rect 8573 10112 8585 10115
rect 7055 10084 8585 10112
rect 7055 10081 7067 10084
rect 7009 10075 7067 10081
rect 8573 10081 8585 10084
rect 8619 10112 8631 10115
rect 8846 10112 8852 10124
rect 8619 10084 8852 10112
rect 8619 10081 8631 10084
rect 8573 10075 8631 10081
rect 8846 10072 8852 10084
rect 8904 10072 8910 10124
rect 12342 10112 12348 10124
rect 12303 10084 12348 10112
rect 12342 10072 12348 10084
rect 12400 10112 12406 10124
rect 13265 10115 13323 10121
rect 13265 10112 13277 10115
rect 12400 10084 13277 10112
rect 12400 10072 12406 10084
rect 13265 10081 13277 10084
rect 13311 10112 13323 10115
rect 19150 10112 19156 10124
rect 13311 10084 13492 10112
rect 19111 10084 19156 10112
rect 13311 10081 13323 10084
rect 13265 10075 13323 10081
rect 13464 10056 13492 10084
rect 19150 10072 19156 10084
rect 19208 10072 19214 10124
rect 10226 10044 10232 10056
rect 4126 10016 10232 10044
rect 3326 9936 3332 9988
rect 3384 9976 3390 9988
rect 4126 9976 4154 10016
rect 10226 10004 10232 10016
rect 10284 10004 10290 10056
rect 10873 10047 10931 10053
rect 10873 10013 10885 10047
rect 10919 10044 10931 10047
rect 11882 10044 11888 10056
rect 10919 10016 11888 10044
rect 10919 10013 10931 10016
rect 10873 10007 10931 10013
rect 11882 10004 11888 10016
rect 11940 10004 11946 10056
rect 13446 10004 13452 10056
rect 13504 10004 13510 10056
rect 16117 10047 16175 10053
rect 16117 10013 16129 10047
rect 16163 10044 16175 10047
rect 16482 10044 16488 10056
rect 16163 10016 16488 10044
rect 16163 10013 16175 10016
rect 16117 10007 16175 10013
rect 16482 10004 16488 10016
rect 16540 10004 16546 10056
rect 16758 10044 16764 10056
rect 16719 10016 16764 10044
rect 16758 10004 16764 10016
rect 16816 10004 16822 10056
rect 17678 10044 17684 10056
rect 17639 10016 17684 10044
rect 17678 10004 17684 10016
rect 17736 10004 17742 10056
rect 7190 9976 7196 9988
rect 3384 9948 4154 9976
rect 7151 9948 7196 9976
rect 3384 9936 3390 9948
rect 7190 9936 7196 9948
rect 7248 9936 7254 9988
rect 3970 9868 3976 9920
rect 4028 9908 4034 9920
rect 4985 9911 5043 9917
rect 4985 9908 4997 9911
rect 4028 9880 4997 9908
rect 4028 9868 4034 9880
rect 4985 9877 4997 9880
rect 5031 9877 5043 9911
rect 8294 9908 8300 9920
rect 8255 9880 8300 9908
rect 4985 9871 5043 9877
rect 8294 9868 8300 9880
rect 8352 9868 8358 9920
rect 9674 9868 9680 9920
rect 9732 9908 9738 9920
rect 9861 9911 9919 9917
rect 9861 9908 9873 9911
rect 9732 9880 9873 9908
rect 9732 9868 9738 9880
rect 9861 9877 9873 9880
rect 9907 9877 9919 9911
rect 11146 9908 11152 9920
rect 11107 9880 11152 9908
rect 9861 9871 9919 9877
rect 11146 9868 11152 9880
rect 11204 9868 11210 9920
rect 13630 9908 13636 9920
rect 13591 9880 13636 9908
rect 13630 9868 13636 9880
rect 13688 9868 13694 9920
rect 15562 9908 15568 9920
rect 15523 9880 15568 9908
rect 15562 9868 15568 9880
rect 15620 9868 15626 9920
rect 1104 9818 22816 9840
rect 1104 9766 4982 9818
rect 5034 9766 5046 9818
rect 5098 9766 5110 9818
rect 5162 9766 5174 9818
rect 5226 9766 12982 9818
rect 13034 9766 13046 9818
rect 13098 9766 13110 9818
rect 13162 9766 13174 9818
rect 13226 9766 20982 9818
rect 21034 9766 21046 9818
rect 21098 9766 21110 9818
rect 21162 9766 21174 9818
rect 21226 9766 22816 9818
rect 1104 9744 22816 9766
rect 3694 9704 3700 9716
rect 3655 9676 3700 9704
rect 3694 9664 3700 9676
rect 3752 9664 3758 9716
rect 3786 9664 3792 9716
rect 3844 9704 3850 9716
rect 4065 9707 4123 9713
rect 4065 9704 4077 9707
rect 3844 9676 4077 9704
rect 3844 9664 3850 9676
rect 4065 9673 4077 9676
rect 4111 9673 4123 9707
rect 4065 9667 4123 9673
rect 4338 9664 4344 9716
rect 4396 9704 4402 9716
rect 4525 9707 4583 9713
rect 4525 9704 4537 9707
rect 4396 9676 4537 9704
rect 4396 9664 4402 9676
rect 4525 9673 4537 9676
rect 4571 9673 4583 9707
rect 4525 9667 4583 9673
rect 5905 9707 5963 9713
rect 5905 9673 5917 9707
rect 5951 9704 5963 9707
rect 6546 9704 6552 9716
rect 5951 9676 6552 9704
rect 5951 9673 5963 9676
rect 5905 9667 5963 9673
rect 6546 9664 6552 9676
rect 6604 9664 6610 9716
rect 8846 9664 8852 9716
rect 8904 9704 8910 9716
rect 9766 9704 9772 9716
rect 8904 9676 9772 9704
rect 8904 9664 8910 9676
rect 9766 9664 9772 9676
rect 9824 9664 9830 9716
rect 10229 9707 10287 9713
rect 10229 9673 10241 9707
rect 10275 9704 10287 9707
rect 10594 9704 10600 9716
rect 10275 9676 10600 9704
rect 10275 9673 10287 9676
rect 10229 9667 10287 9673
rect 10594 9664 10600 9676
rect 10652 9664 10658 9716
rect 12342 9664 12348 9716
rect 12400 9704 12406 9716
rect 12621 9707 12679 9713
rect 12621 9704 12633 9707
rect 12400 9676 12633 9704
rect 12400 9664 12406 9676
rect 12621 9673 12633 9676
rect 12667 9673 12679 9707
rect 12621 9667 12679 9673
rect 17954 9664 17960 9716
rect 18012 9704 18018 9716
rect 19150 9704 19156 9716
rect 18012 9676 19156 9704
rect 18012 9664 18018 9676
rect 19150 9664 19156 9676
rect 19208 9664 19214 9716
rect 2314 9596 2320 9648
rect 2372 9636 2378 9648
rect 8018 9636 8024 9648
rect 2372 9608 8024 9636
rect 2372 9596 2378 9608
rect 4062 9528 4068 9580
rect 4120 9568 4126 9580
rect 5092 9577 5120 9608
rect 8018 9596 8024 9608
rect 8076 9636 8082 9648
rect 8076 9608 8984 9636
rect 8076 9596 8082 9608
rect 4801 9571 4859 9577
rect 4801 9568 4813 9571
rect 4120 9540 4813 9568
rect 4120 9528 4126 9540
rect 4801 9537 4813 9540
rect 4847 9537 4859 9571
rect 4801 9531 4859 9537
rect 5077 9571 5135 9577
rect 5077 9537 5089 9571
rect 5123 9537 5135 9571
rect 5077 9531 5135 9537
rect 6825 9571 6883 9577
rect 6825 9537 6837 9571
rect 6871 9568 6883 9571
rect 7190 9568 7196 9580
rect 6871 9540 7196 9568
rect 6871 9537 6883 9540
rect 6825 9531 6883 9537
rect 7190 9528 7196 9540
rect 7248 9528 7254 9580
rect 8956 9577 8984 9608
rect 10134 9596 10140 9648
rect 10192 9636 10198 9648
rect 16666 9636 16672 9648
rect 10192 9608 16672 9636
rect 10192 9596 10198 9608
rect 16666 9596 16672 9608
rect 16724 9596 16730 9648
rect 16758 9596 16764 9648
rect 16816 9636 16822 9648
rect 18693 9639 18751 9645
rect 18693 9636 18705 9639
rect 16816 9608 18705 9636
rect 16816 9596 16822 9608
rect 18693 9605 18705 9608
rect 18739 9636 18751 9639
rect 18966 9636 18972 9648
rect 18739 9608 18972 9636
rect 18739 9605 18751 9608
rect 18693 9599 18751 9605
rect 18966 9596 18972 9608
rect 19024 9596 19030 9648
rect 8941 9571 8999 9577
rect 8941 9537 8953 9571
rect 8987 9537 8999 9571
rect 8941 9531 8999 9537
rect 13630 9528 13636 9580
rect 13688 9568 13694 9580
rect 14737 9571 14795 9577
rect 13688 9540 14320 9568
rect 13688 9528 13694 9540
rect 14292 9512 14320 9540
rect 14737 9537 14749 9571
rect 14783 9568 14795 9571
rect 15562 9568 15568 9580
rect 14783 9540 15568 9568
rect 14783 9537 14795 9540
rect 14737 9531 14795 9537
rect 15562 9528 15568 9540
rect 15620 9528 15626 9580
rect 17678 9528 17684 9580
rect 17736 9568 17742 9580
rect 19751 9571 19809 9577
rect 19751 9568 19763 9571
rect 17736 9540 19763 9568
rect 17736 9528 17742 9540
rect 19751 9537 19763 9540
rect 19797 9537 19809 9571
rect 19751 9531 19809 9537
rect 13265 9503 13323 9509
rect 13265 9469 13277 9503
rect 13311 9469 13323 9503
rect 13265 9463 13323 9469
rect 3970 9392 3976 9444
rect 4028 9432 4034 9444
rect 4798 9432 4804 9444
rect 4028 9404 4804 9432
rect 4028 9392 4034 9404
rect 4798 9392 4804 9404
rect 4856 9432 4862 9444
rect 4893 9435 4951 9441
rect 4893 9432 4905 9435
rect 4856 9404 4905 9432
rect 4856 9392 4862 9404
rect 4893 9401 4905 9404
rect 4939 9401 4951 9435
rect 4893 9395 4951 9401
rect 5442 9392 5448 9444
rect 5500 9432 5506 9444
rect 7926 9432 7932 9444
rect 5500 9404 6592 9432
rect 5500 9392 5506 9404
rect 6564 9376 6592 9404
rect 7208 9404 7932 9432
rect 6270 9364 6276 9376
rect 6231 9336 6276 9364
rect 6270 9324 6276 9336
rect 6328 9324 6334 9376
rect 6546 9364 6552 9376
rect 6507 9336 6552 9364
rect 6546 9324 6552 9336
rect 6604 9364 6610 9376
rect 7208 9373 7236 9404
rect 7926 9392 7932 9404
rect 7984 9392 7990 9444
rect 8113 9435 8171 9441
rect 8113 9401 8125 9435
rect 8159 9432 8171 9435
rect 8662 9432 8668 9444
rect 8159 9404 8668 9432
rect 8159 9401 8171 9404
rect 8113 9395 8171 9401
rect 8662 9392 8668 9404
rect 8720 9392 8726 9444
rect 8754 9392 8760 9444
rect 8812 9432 8818 9444
rect 10870 9432 10876 9444
rect 8812 9404 8857 9432
rect 10831 9404 10876 9432
rect 8812 9392 8818 9404
rect 10870 9392 10876 9404
rect 10928 9392 10934 9444
rect 10965 9435 11023 9441
rect 10965 9401 10977 9435
rect 11011 9401 11023 9435
rect 10965 9395 11023 9401
rect 7193 9367 7251 9373
rect 7193 9364 7205 9367
rect 6604 9336 7205 9364
rect 6604 9324 6610 9336
rect 7193 9333 7205 9336
rect 7239 9333 7251 9367
rect 7193 9327 7251 9333
rect 7745 9367 7803 9373
rect 7745 9333 7757 9367
rect 7791 9364 7803 9367
rect 7834 9364 7840 9376
rect 7791 9336 7840 9364
rect 7791 9333 7803 9336
rect 7745 9327 7803 9333
rect 7834 9324 7840 9336
rect 7892 9324 7898 9376
rect 8481 9367 8539 9373
rect 8481 9333 8493 9367
rect 8527 9364 8539 9367
rect 8772 9364 8800 9392
rect 8527 9336 8800 9364
rect 8527 9333 8539 9336
rect 8481 9327 8539 9333
rect 10594 9324 10600 9376
rect 10652 9364 10658 9376
rect 10980 9364 11008 9395
rect 11238 9392 11244 9444
rect 11296 9432 11302 9444
rect 11517 9435 11575 9441
rect 11517 9432 11529 9435
rect 11296 9404 11529 9432
rect 11296 9392 11302 9404
rect 11517 9401 11529 9404
rect 11563 9401 11575 9435
rect 11517 9395 11575 9401
rect 13280 9376 13308 9463
rect 13446 9460 13452 9512
rect 13504 9500 13510 9512
rect 13725 9503 13783 9509
rect 13725 9500 13737 9503
rect 13504 9472 13737 9500
rect 13504 9460 13510 9472
rect 13725 9469 13737 9472
rect 13771 9469 13783 9503
rect 14274 9500 14280 9512
rect 14235 9472 14280 9500
rect 13725 9463 13783 9469
rect 14274 9460 14280 9472
rect 14332 9460 14338 9512
rect 14461 9503 14519 9509
rect 14461 9469 14473 9503
rect 14507 9469 14519 9503
rect 16485 9503 16543 9509
rect 14461 9463 14519 9469
rect 15488 9472 15976 9500
rect 13998 9392 14004 9444
rect 14056 9432 14062 9444
rect 14476 9432 14504 9463
rect 14056 9404 14504 9432
rect 14056 9392 14062 9404
rect 15488 9376 15516 9472
rect 15948 9441 15976 9472
rect 16485 9469 16497 9503
rect 16531 9500 16543 9503
rect 17405 9503 17463 9509
rect 17405 9500 17417 9503
rect 16531 9472 17417 9500
rect 16531 9469 16543 9472
rect 16485 9463 16543 9469
rect 17405 9469 17417 9472
rect 17451 9500 17463 9503
rect 17770 9500 17776 9512
rect 17451 9472 17776 9500
rect 17451 9469 17463 9472
rect 17405 9463 17463 9469
rect 17770 9460 17776 9472
rect 17828 9460 17834 9512
rect 19648 9503 19706 9509
rect 19648 9500 19660 9503
rect 19444 9472 19660 9500
rect 15927 9435 15985 9441
rect 15927 9401 15939 9435
rect 15973 9401 15985 9435
rect 15927 9395 15985 9401
rect 10652 9336 11008 9364
rect 13173 9367 13231 9373
rect 10652 9324 10658 9336
rect 13173 9333 13185 9367
rect 13219 9364 13231 9367
rect 13262 9364 13268 9376
rect 13219 9336 13268 9364
rect 13219 9333 13231 9336
rect 13173 9327 13231 9333
rect 13262 9324 13268 9336
rect 13320 9324 13326 9376
rect 15470 9364 15476 9376
rect 15431 9336 15476 9364
rect 15470 9324 15476 9336
rect 15528 9324 15534 9376
rect 16853 9367 16911 9373
rect 16853 9333 16865 9367
rect 16899 9364 16911 9367
rect 17494 9364 17500 9376
rect 16899 9336 17500 9364
rect 16899 9333 16911 9336
rect 16853 9327 16911 9333
rect 17494 9324 17500 9336
rect 17552 9324 17558 9376
rect 17788 9364 17816 9460
rect 18138 9432 18144 9444
rect 18099 9404 18144 9432
rect 18138 9392 18144 9404
rect 18196 9392 18202 9444
rect 18233 9435 18291 9441
rect 18233 9401 18245 9435
rect 18279 9401 18291 9435
rect 18233 9395 18291 9401
rect 18248 9364 18276 9395
rect 18598 9392 18604 9444
rect 18656 9432 18662 9444
rect 19444 9432 19472 9472
rect 19648 9469 19660 9472
rect 19694 9500 19706 9503
rect 20070 9500 20076 9512
rect 19694 9472 20076 9500
rect 19694 9469 19706 9472
rect 19648 9463 19706 9469
rect 20070 9460 20076 9472
rect 20128 9460 20134 9512
rect 18656 9404 19472 9432
rect 18656 9392 18662 9404
rect 17788 9336 18276 9364
rect 1104 9274 22816 9296
rect 1104 9222 8982 9274
rect 9034 9222 9046 9274
rect 9098 9222 9110 9274
rect 9162 9222 9174 9274
rect 9226 9222 16982 9274
rect 17034 9222 17046 9274
rect 17098 9222 17110 9274
rect 17162 9222 17174 9274
rect 17226 9222 22816 9274
rect 1104 9200 22816 9222
rect 4798 9160 4804 9172
rect 4759 9132 4804 9160
rect 4798 9120 4804 9132
rect 4856 9120 4862 9172
rect 5902 9160 5908 9172
rect 5863 9132 5908 9160
rect 5902 9120 5908 9132
rect 5960 9120 5966 9172
rect 6273 9163 6331 9169
rect 6273 9129 6285 9163
rect 6319 9160 6331 9163
rect 6638 9160 6644 9172
rect 6319 9132 6644 9160
rect 6319 9129 6331 9132
rect 6273 9123 6331 9129
rect 6638 9120 6644 9132
rect 6696 9120 6702 9172
rect 6917 9163 6975 9169
rect 6917 9129 6929 9163
rect 6963 9160 6975 9163
rect 7190 9160 7196 9172
rect 6963 9132 7196 9160
rect 6963 9129 6975 9132
rect 6917 9123 6975 9129
rect 7190 9120 7196 9132
rect 7248 9120 7254 9172
rect 9999 9163 10057 9169
rect 9999 9129 10011 9163
rect 10045 9160 10057 9163
rect 10870 9160 10876 9172
rect 10045 9132 10876 9160
rect 10045 9129 10057 9132
rect 9999 9123 10057 9129
rect 10870 9120 10876 9132
rect 10928 9120 10934 9172
rect 13722 9120 13728 9172
rect 13780 9160 13786 9172
rect 16206 9160 16212 9172
rect 13780 9132 14044 9160
rect 16119 9132 16212 9160
rect 13780 9120 13786 9132
rect 106 9052 112 9104
rect 164 9092 170 9104
rect 1535 9095 1593 9101
rect 1535 9092 1547 9095
rect 164 9064 1547 9092
rect 164 9052 170 9064
rect 1535 9061 1547 9064
rect 1581 9061 1593 9095
rect 7834 9092 7840 9104
rect 7795 9064 7840 9092
rect 1535 9055 1593 9061
rect 7834 9052 7840 9064
rect 7892 9052 7898 9104
rect 10134 9092 10140 9104
rect 9911 9064 10140 9092
rect 1448 9027 1506 9033
rect 1448 8993 1460 9027
rect 1494 9024 1506 9027
rect 1670 9024 1676 9036
rect 1494 8996 1676 9024
rect 1494 8993 1506 8996
rect 1448 8987 1506 8993
rect 1670 8984 1676 8996
rect 1728 9024 1734 9036
rect 2314 9024 2320 9036
rect 1728 8996 2320 9024
rect 1728 8984 1734 8996
rect 2314 8984 2320 8996
rect 2372 8984 2378 9036
rect 9911 9033 9939 9064
rect 10134 9052 10140 9064
rect 10192 9052 10198 9104
rect 10226 9052 10232 9104
rect 10284 9092 10290 9104
rect 10321 9095 10379 9101
rect 10321 9092 10333 9095
rect 10284 9064 10333 9092
rect 10284 9052 10290 9064
rect 10321 9061 10333 9064
rect 10367 9061 10379 9095
rect 11054 9092 11060 9104
rect 11015 9064 11060 9092
rect 10321 9055 10379 9061
rect 11054 9052 11060 9064
rect 11112 9052 11118 9104
rect 14016 9036 14044 9132
rect 16206 9120 16212 9132
rect 16264 9120 16270 9172
rect 17678 9120 17684 9172
rect 17736 9160 17742 9172
rect 18049 9163 18107 9169
rect 18049 9160 18061 9163
rect 17736 9132 18061 9160
rect 17736 9120 17742 9132
rect 18049 9129 18061 9132
rect 18095 9129 18107 9163
rect 18049 9123 18107 9129
rect 21039 9163 21097 9169
rect 21039 9129 21051 9163
rect 21085 9160 21097 9163
rect 21266 9160 21272 9172
rect 21085 9132 21272 9160
rect 21085 9129 21097 9132
rect 21039 9123 21097 9129
rect 21266 9120 21272 9132
rect 21324 9120 21330 9172
rect 15470 9052 15476 9104
rect 15528 9092 15534 9104
rect 15651 9095 15709 9101
rect 15651 9092 15663 9095
rect 15528 9064 15663 9092
rect 15528 9052 15534 9064
rect 15651 9061 15663 9064
rect 15697 9092 15709 9095
rect 15838 9092 15844 9104
rect 15697 9064 15844 9092
rect 15697 9061 15709 9064
rect 15651 9055 15709 9061
rect 15838 9052 15844 9064
rect 15896 9052 15902 9104
rect 16224 9092 16252 9120
rect 17221 9095 17279 9101
rect 17221 9092 17233 9095
rect 16224 9064 17233 9092
rect 17221 9061 17233 9064
rect 17267 9092 17279 9095
rect 17494 9092 17500 9104
rect 17267 9064 17500 9092
rect 17267 9061 17279 9064
rect 17221 9055 17279 9061
rect 17494 9052 17500 9064
rect 17552 9052 17558 9104
rect 17773 9095 17831 9101
rect 17773 9061 17785 9095
rect 17819 9092 17831 9095
rect 18322 9092 18328 9104
rect 17819 9064 18328 9092
rect 17819 9061 17831 9064
rect 17773 9055 17831 9061
rect 18322 9052 18328 9064
rect 18380 9052 18386 9104
rect 9896 9027 9954 9033
rect 9896 8993 9908 9027
rect 9942 8993 9954 9027
rect 9896 8987 9954 8993
rect 13173 9027 13231 9033
rect 13173 8993 13185 9027
rect 13219 9024 13231 9027
rect 13262 9024 13268 9036
rect 13219 8996 13268 9024
rect 13219 8993 13231 8996
rect 13173 8987 13231 8993
rect 13262 8984 13268 8996
rect 13320 8984 13326 9036
rect 13446 9024 13452 9036
rect 13407 8996 13452 9024
rect 13446 8984 13452 8996
rect 13504 8984 13510 9036
rect 13725 9027 13783 9033
rect 13725 8993 13737 9027
rect 13771 9024 13783 9027
rect 13906 9024 13912 9036
rect 13771 8996 13912 9024
rect 13771 8993 13783 8996
rect 13725 8987 13783 8993
rect 7742 8956 7748 8968
rect 7703 8928 7748 8956
rect 7742 8916 7748 8928
rect 7800 8916 7806 8968
rect 8018 8956 8024 8968
rect 7979 8928 8024 8956
rect 8018 8916 8024 8928
rect 8076 8916 8082 8968
rect 10962 8956 10968 8968
rect 10923 8928 10968 8956
rect 10962 8916 10968 8928
rect 11020 8916 11026 8968
rect 11238 8956 11244 8968
rect 11151 8928 11244 8956
rect 11238 8916 11244 8928
rect 11296 8916 11302 8968
rect 12802 8916 12808 8968
rect 12860 8956 12866 8968
rect 13740 8956 13768 8987
rect 13906 8984 13912 8996
rect 13964 8984 13970 9036
rect 13998 8984 14004 9036
rect 14056 9024 14062 9036
rect 14093 9027 14151 9033
rect 14093 9024 14105 9027
rect 14056 8996 14105 9024
rect 14056 8984 14062 8996
rect 14093 8993 14105 8996
rect 14139 8993 14151 9027
rect 18598 9024 18604 9036
rect 18559 8996 18604 9024
rect 14093 8987 14151 8993
rect 18598 8984 18604 8996
rect 18656 8984 18662 9036
rect 19664 9027 19722 9033
rect 19664 8993 19676 9027
rect 19710 9024 19722 9027
rect 20070 9024 20076 9036
rect 19710 8996 20076 9024
rect 19710 8993 19722 8996
rect 19664 8987 19722 8993
rect 20070 8984 20076 8996
rect 20128 8984 20134 9036
rect 20806 8984 20812 9036
rect 20864 9024 20870 9036
rect 20936 9027 20994 9033
rect 20936 9024 20948 9027
rect 20864 8996 20948 9024
rect 20864 8984 20870 8996
rect 20936 8993 20948 8996
rect 20982 8993 20994 9027
rect 20936 8987 20994 8993
rect 12860 8928 13768 8956
rect 14369 8959 14427 8965
rect 12860 8916 12866 8928
rect 14369 8925 14381 8959
rect 14415 8956 14427 8959
rect 14826 8956 14832 8968
rect 14415 8928 14832 8956
rect 14415 8925 14427 8928
rect 14369 8919 14427 8925
rect 14826 8916 14832 8928
rect 14884 8956 14890 8968
rect 15289 8959 15347 8965
rect 15289 8956 15301 8959
rect 14884 8928 15301 8956
rect 14884 8916 14890 8928
rect 15289 8925 15301 8928
rect 15335 8925 15347 8959
rect 17126 8956 17132 8968
rect 17087 8928 17132 8956
rect 15289 8919 15347 8925
rect 17126 8916 17132 8928
rect 17184 8916 17190 8968
rect 18138 8916 18144 8968
rect 18196 8956 18202 8968
rect 18509 8959 18567 8965
rect 18509 8956 18521 8959
rect 18196 8928 18521 8956
rect 18196 8916 18202 8928
rect 18509 8925 18521 8928
rect 18555 8956 18567 8959
rect 19751 8959 19809 8965
rect 19751 8956 19763 8959
rect 18555 8928 19763 8956
rect 18555 8925 18567 8928
rect 18509 8919 18567 8925
rect 19751 8925 19763 8928
rect 19797 8925 19809 8959
rect 19751 8919 19809 8925
rect 10410 8848 10416 8900
rect 10468 8888 10474 8900
rect 11256 8888 11284 8916
rect 10468 8860 11284 8888
rect 10468 8848 10474 8860
rect 10686 8820 10692 8832
rect 10647 8792 10692 8820
rect 10686 8780 10692 8792
rect 10744 8780 10750 8832
rect 16482 8820 16488 8832
rect 16443 8792 16488 8820
rect 16482 8780 16488 8792
rect 16540 8780 16546 8832
rect 18506 8780 18512 8832
rect 18564 8820 18570 8832
rect 18739 8823 18797 8829
rect 18739 8820 18751 8823
rect 18564 8792 18751 8820
rect 18564 8780 18570 8792
rect 18739 8789 18751 8792
rect 18785 8789 18797 8823
rect 18739 8783 18797 8789
rect 1104 8730 22816 8752
rect 1104 8678 4982 8730
rect 5034 8678 5046 8730
rect 5098 8678 5110 8730
rect 5162 8678 5174 8730
rect 5226 8678 12982 8730
rect 13034 8678 13046 8730
rect 13098 8678 13110 8730
rect 13162 8678 13174 8730
rect 13226 8678 20982 8730
rect 21034 8678 21046 8730
rect 21098 8678 21110 8730
rect 21162 8678 21174 8730
rect 21226 8678 22816 8730
rect 1104 8656 22816 8678
rect 1581 8619 1639 8625
rect 1581 8585 1593 8619
rect 1627 8616 1639 8619
rect 1762 8616 1768 8628
rect 1627 8588 1768 8616
rect 1627 8585 1639 8588
rect 1581 8579 1639 8585
rect 1762 8576 1768 8588
rect 1820 8576 1826 8628
rect 7193 8619 7251 8625
rect 7193 8585 7205 8619
rect 7239 8616 7251 8619
rect 7834 8616 7840 8628
rect 7239 8588 7840 8616
rect 7239 8585 7251 8588
rect 7193 8579 7251 8585
rect 7834 8576 7840 8588
rect 7892 8576 7898 8628
rect 9769 8619 9827 8625
rect 9769 8585 9781 8619
rect 9815 8616 9827 8619
rect 10134 8616 10140 8628
rect 9815 8588 10140 8616
rect 9815 8585 9827 8588
rect 9769 8579 9827 8585
rect 10134 8576 10140 8588
rect 10192 8576 10198 8628
rect 10962 8576 10968 8628
rect 11020 8616 11026 8628
rect 11241 8619 11299 8625
rect 11241 8616 11253 8619
rect 11020 8588 11253 8616
rect 11020 8576 11026 8588
rect 11241 8585 11253 8588
rect 11287 8616 11299 8619
rect 12575 8619 12633 8625
rect 12575 8616 12587 8619
rect 11287 8588 12587 8616
rect 11287 8585 11299 8588
rect 11241 8579 11299 8585
rect 12575 8585 12587 8588
rect 12621 8585 12633 8619
rect 12575 8579 12633 8585
rect 13446 8576 13452 8628
rect 13504 8616 13510 8628
rect 13633 8619 13691 8625
rect 13633 8616 13645 8619
rect 13504 8588 13645 8616
rect 13504 8576 13510 8588
rect 13633 8585 13645 8588
rect 13679 8585 13691 8619
rect 14826 8616 14832 8628
rect 14787 8588 14832 8616
rect 13633 8579 13691 8585
rect 14826 8576 14832 8588
rect 14884 8576 14890 8628
rect 15151 8619 15209 8625
rect 15151 8585 15163 8619
rect 15197 8616 15209 8619
rect 16482 8616 16488 8628
rect 15197 8588 16488 8616
rect 15197 8585 15209 8588
rect 15151 8579 15209 8585
rect 16482 8576 16488 8588
rect 16540 8576 16546 8628
rect 16850 8625 16856 8628
rect 16807 8619 16856 8625
rect 16807 8616 16819 8619
rect 16763 8588 16819 8616
rect 16807 8585 16819 8588
rect 16853 8585 16856 8619
rect 16807 8579 16856 8585
rect 16850 8576 16856 8579
rect 16908 8616 16914 8628
rect 17126 8616 17132 8628
rect 16908 8588 17132 8616
rect 16908 8576 16914 8588
rect 17126 8576 17132 8588
rect 17184 8576 17190 8628
rect 17494 8616 17500 8628
rect 17455 8588 17500 8616
rect 17494 8576 17500 8588
rect 17552 8576 17558 8628
rect 20070 8616 20076 8628
rect 19983 8588 20076 8616
rect 20070 8576 20076 8588
rect 20128 8616 20134 8628
rect 21177 8619 21235 8625
rect 21177 8616 21189 8619
rect 20128 8588 21189 8616
rect 20128 8576 20134 8588
rect 8662 8508 8668 8560
rect 8720 8548 8726 8560
rect 8941 8551 8999 8557
rect 8941 8548 8953 8551
rect 8720 8520 8953 8548
rect 8720 8508 8726 8520
rect 8941 8517 8953 8520
rect 8987 8548 8999 8551
rect 11882 8548 11888 8560
rect 8987 8520 11888 8548
rect 8987 8517 8999 8520
rect 8941 8511 8999 8517
rect 11882 8508 11888 8520
rect 11940 8508 11946 8560
rect 14182 8508 14188 8560
rect 14240 8548 14246 8560
rect 18598 8548 18604 8560
rect 14240 8520 18604 8548
rect 14240 8508 14246 8520
rect 18598 8508 18604 8520
rect 18656 8508 18662 8560
rect 7423 8483 7481 8489
rect 7423 8449 7435 8483
rect 7469 8480 7481 8483
rect 9953 8483 10011 8489
rect 9953 8480 9965 8483
rect 7469 8452 9965 8480
rect 7469 8449 7481 8452
rect 7423 8443 7481 8449
rect 9953 8449 9965 8452
rect 9999 8480 10011 8483
rect 10686 8480 10692 8492
rect 9999 8452 10692 8480
rect 9999 8449 10011 8452
rect 9953 8443 10011 8449
rect 10686 8440 10692 8452
rect 10744 8440 10750 8492
rect 12618 8440 12624 8492
rect 12676 8480 12682 8492
rect 12676 8452 14872 8480
rect 12676 8440 12682 8452
rect 1397 8415 1455 8421
rect 1397 8381 1409 8415
rect 1443 8412 1455 8415
rect 1443 8384 2084 8412
rect 1443 8381 1455 8384
rect 1397 8375 1455 8381
rect 2056 8288 2084 8384
rect 2774 8372 2780 8424
rect 2832 8412 2838 8424
rect 7336 8415 7394 8421
rect 7336 8412 7348 8415
rect 2832 8384 7348 8412
rect 2832 8372 2838 8384
rect 7336 8381 7348 8384
rect 7382 8412 7394 8415
rect 12253 8415 12311 8421
rect 7382 8384 7880 8412
rect 7382 8381 7394 8384
rect 7336 8375 7394 8381
rect 7852 8353 7880 8384
rect 12253 8381 12265 8415
rect 12299 8412 12311 8415
rect 12504 8415 12562 8421
rect 12504 8412 12516 8415
rect 12299 8384 12516 8412
rect 12299 8381 12311 8384
rect 12253 8375 12311 8381
rect 12504 8381 12516 8384
rect 12550 8412 12562 8415
rect 14090 8412 14096 8424
rect 12550 8384 14096 8412
rect 12550 8381 12562 8384
rect 12504 8375 12562 8381
rect 14090 8372 14096 8384
rect 14148 8372 14154 8424
rect 14844 8412 14872 8452
rect 15048 8415 15106 8421
rect 15048 8412 15060 8415
rect 14844 8384 15060 8412
rect 15048 8381 15060 8384
rect 15094 8412 15106 8415
rect 15473 8415 15531 8421
rect 15473 8412 15485 8415
rect 15094 8384 15485 8412
rect 15094 8381 15106 8384
rect 15048 8375 15106 8381
rect 15473 8381 15485 8384
rect 15519 8381 15531 8415
rect 15473 8375 15531 8381
rect 16736 8415 16794 8421
rect 16736 8381 16748 8415
rect 16782 8412 16794 8415
rect 19058 8412 19064 8424
rect 16782 8384 17264 8412
rect 19019 8384 19064 8412
rect 16782 8381 16794 8384
rect 16736 8375 16794 8381
rect 7837 8347 7895 8353
rect 7837 8313 7849 8347
rect 7883 8344 7895 8347
rect 8018 8344 8024 8356
rect 7883 8316 8024 8344
rect 7883 8313 7895 8316
rect 7837 8307 7895 8313
rect 8018 8304 8024 8316
rect 8076 8304 8082 8356
rect 8386 8344 8392 8356
rect 8347 8316 8392 8344
rect 8386 8304 8392 8316
rect 8444 8304 8450 8356
rect 8481 8347 8539 8353
rect 8481 8313 8493 8347
rect 8527 8313 8539 8347
rect 10045 8347 10103 8353
rect 10045 8344 10057 8347
rect 8481 8307 8539 8313
rect 9324 8316 10057 8344
rect 2038 8276 2044 8288
rect 1999 8248 2044 8276
rect 2038 8236 2044 8248
rect 2096 8236 2102 8288
rect 8110 8276 8116 8288
rect 8071 8248 8116 8276
rect 8110 8236 8116 8248
rect 8168 8276 8174 8288
rect 8496 8276 8524 8307
rect 9324 8285 9352 8316
rect 10045 8313 10057 8316
rect 10091 8313 10103 8347
rect 10045 8307 10103 8313
rect 10410 8304 10416 8356
rect 10468 8344 10474 8356
rect 10597 8347 10655 8353
rect 10597 8344 10609 8347
rect 10468 8316 10609 8344
rect 10468 8304 10474 8316
rect 10597 8313 10609 8316
rect 10643 8313 10655 8347
rect 10597 8307 10655 8313
rect 13262 8304 13268 8356
rect 13320 8344 13326 8356
rect 13357 8347 13415 8353
rect 13357 8344 13369 8347
rect 13320 8316 13369 8344
rect 13320 8304 13326 8316
rect 13357 8313 13369 8316
rect 13403 8344 13415 8347
rect 13814 8344 13820 8356
rect 13403 8316 13820 8344
rect 13403 8313 13415 8316
rect 13357 8307 13415 8313
rect 13814 8304 13820 8316
rect 13872 8304 13878 8356
rect 9309 8279 9367 8285
rect 9309 8276 9321 8279
rect 8168 8248 9321 8276
rect 8168 8236 8174 8248
rect 9309 8245 9321 8248
rect 9355 8245 9367 8279
rect 9309 8239 9367 8245
rect 10965 8279 11023 8285
rect 10965 8245 10977 8279
rect 11011 8276 11023 8279
rect 11054 8276 11060 8288
rect 11011 8248 11060 8276
rect 11011 8245 11023 8248
rect 10965 8239 11023 8245
rect 11054 8236 11060 8248
rect 11112 8276 11118 8288
rect 11514 8276 11520 8288
rect 11112 8248 11520 8276
rect 11112 8236 11118 8248
rect 11514 8236 11520 8248
rect 11572 8236 11578 8288
rect 12802 8236 12808 8288
rect 12860 8276 12866 8288
rect 12897 8279 12955 8285
rect 12897 8276 12909 8279
rect 12860 8248 12909 8276
rect 12860 8236 12866 8248
rect 12897 8245 12909 8248
rect 12943 8245 12955 8279
rect 13998 8276 14004 8288
rect 13959 8248 14004 8276
rect 12897 8239 12955 8245
rect 13998 8236 14004 8248
rect 14056 8236 14062 8288
rect 15838 8276 15844 8288
rect 15799 8248 15844 8276
rect 15838 8236 15844 8248
rect 15896 8236 15902 8288
rect 17236 8285 17264 8384
rect 19058 8372 19064 8384
rect 19116 8372 19122 8424
rect 20548 8421 20576 8588
rect 21177 8585 21189 8588
rect 21223 8616 21235 8619
rect 21358 8616 21364 8628
rect 21223 8588 21364 8616
rect 21223 8585 21235 8588
rect 21177 8579 21235 8585
rect 21358 8576 21364 8588
rect 21416 8576 21422 8628
rect 20717 8551 20775 8557
rect 20717 8517 20729 8551
rect 20763 8548 20775 8551
rect 21266 8548 21272 8560
rect 20763 8520 21272 8548
rect 20763 8517 20775 8520
rect 20717 8511 20775 8517
rect 21266 8508 21272 8520
rect 21324 8508 21330 8560
rect 20533 8415 20591 8421
rect 20533 8381 20545 8415
rect 20579 8381 20591 8415
rect 20533 8375 20591 8381
rect 19702 8304 19708 8356
rect 19760 8344 19766 8356
rect 20806 8344 20812 8356
rect 19760 8316 20812 8344
rect 19760 8304 19766 8316
rect 20806 8304 20812 8316
rect 20864 8344 20870 8356
rect 21453 8347 21511 8353
rect 21453 8344 21465 8347
rect 20864 8316 21465 8344
rect 20864 8304 20870 8316
rect 21453 8313 21465 8316
rect 21499 8313 21511 8347
rect 21453 8307 21511 8313
rect 17221 8279 17279 8285
rect 17221 8245 17233 8279
rect 17267 8276 17279 8279
rect 17310 8276 17316 8288
rect 17267 8248 17316 8276
rect 17267 8245 17279 8248
rect 17221 8239 17279 8245
rect 17310 8236 17316 8248
rect 17368 8236 17374 8288
rect 19426 8276 19432 8288
rect 19387 8248 19432 8276
rect 19426 8236 19432 8248
rect 19484 8236 19490 8288
rect 1104 8186 22816 8208
rect 1104 8134 8982 8186
rect 9034 8134 9046 8186
rect 9098 8134 9110 8186
rect 9162 8134 9174 8186
rect 9226 8134 16982 8186
rect 17034 8134 17046 8186
rect 17098 8134 17110 8186
rect 17162 8134 17174 8186
rect 17226 8134 22816 8186
rect 1104 8112 22816 8134
rect 1670 8072 1676 8084
rect 1631 8044 1676 8072
rect 1670 8032 1676 8044
rect 1728 8032 1734 8084
rect 7653 8075 7711 8081
rect 7653 8041 7665 8075
rect 7699 8072 7711 8075
rect 8110 8072 8116 8084
rect 7699 8044 8116 8072
rect 7699 8041 7711 8044
rect 7653 8035 7711 8041
rect 8110 8032 8116 8044
rect 8168 8032 8174 8084
rect 10042 8072 10048 8084
rect 10003 8044 10048 8072
rect 10042 8032 10048 8044
rect 10100 8032 10106 8084
rect 10597 8075 10655 8081
rect 10597 8041 10609 8075
rect 10643 8041 10655 8075
rect 10597 8035 10655 8041
rect 6638 7964 6644 8016
rect 6696 8004 6702 8016
rect 7054 8007 7112 8013
rect 7054 8004 7066 8007
rect 6696 7976 7066 8004
rect 6696 7964 6702 7976
rect 7054 7973 7066 7976
rect 7100 7973 7112 8007
rect 7054 7967 7112 7973
rect 7742 7964 7748 8016
rect 7800 8004 7806 8016
rect 7929 8007 7987 8013
rect 7929 8004 7941 8007
rect 7800 7976 7941 8004
rect 7800 7964 7806 7976
rect 7929 7973 7941 7976
rect 7975 8004 7987 8007
rect 10410 8004 10416 8016
rect 7975 7976 10416 8004
rect 7975 7973 7987 7976
rect 7929 7967 7987 7973
rect 10410 7964 10416 7976
rect 10468 7964 10474 8016
rect 10612 8004 10640 8035
rect 16850 8032 16856 8084
rect 16908 8072 16914 8084
rect 17037 8075 17095 8081
rect 17037 8072 17049 8075
rect 16908 8044 17049 8072
rect 16908 8032 16914 8044
rect 17037 8041 17049 8044
rect 17083 8041 17095 8075
rect 17037 8035 17095 8041
rect 11514 8004 11520 8016
rect 10612 7976 11520 8004
rect 11514 7964 11520 7976
rect 11572 8004 11578 8016
rect 11609 8007 11667 8013
rect 11609 8004 11621 8007
rect 11572 7976 11621 8004
rect 11572 7964 11578 7976
rect 11609 7973 11621 7976
rect 11655 7973 11667 8007
rect 11609 7967 11667 7973
rect 15743 8007 15801 8013
rect 15743 7973 15755 8007
rect 15789 8004 15801 8007
rect 15838 8004 15844 8016
rect 15789 7976 15844 8004
rect 15789 7973 15801 7976
rect 15743 7967 15801 7973
rect 15838 7964 15844 7976
rect 15896 7964 15902 8016
rect 17865 8007 17923 8013
rect 17865 7973 17877 8007
rect 17911 8004 17923 8007
rect 18046 8004 18052 8016
rect 17911 7976 18052 8004
rect 17911 7973 17923 7976
rect 17865 7967 17923 7973
rect 18046 7964 18052 7976
rect 18104 7964 18110 8016
rect 19426 8004 19432 8016
rect 19387 7976 19432 8004
rect 19426 7964 19432 7976
rect 19484 7964 19490 8016
rect 8711 7939 8769 7945
rect 8711 7905 8723 7939
rect 8757 7936 8769 7939
rect 8757 7908 11100 7936
rect 8757 7905 8769 7908
rect 8711 7899 8769 7905
rect 6730 7868 6736 7880
rect 6691 7840 6736 7868
rect 6730 7828 6736 7840
rect 6788 7828 6794 7880
rect 9677 7871 9735 7877
rect 9677 7837 9689 7871
rect 9723 7868 9735 7871
rect 11072 7868 11100 7908
rect 11517 7871 11575 7877
rect 11517 7868 11529 7871
rect 9723 7840 10916 7868
rect 11072 7840 11529 7868
rect 9723 7837 9735 7840
rect 9677 7831 9735 7837
rect 7282 7760 7288 7812
rect 7340 7800 7346 7812
rect 9125 7803 9183 7809
rect 9125 7800 9137 7803
rect 7340 7772 9137 7800
rect 7340 7760 7346 7772
rect 9125 7769 9137 7772
rect 9171 7769 9183 7803
rect 9125 7763 9183 7769
rect 8386 7732 8392 7744
rect 8347 7704 8392 7732
rect 8386 7692 8392 7704
rect 8444 7692 8450 7744
rect 8481 7735 8539 7741
rect 8481 7701 8493 7735
rect 8527 7732 8539 7735
rect 8662 7732 8668 7744
rect 8527 7704 8668 7732
rect 8527 7701 8539 7704
rect 8481 7695 8539 7701
rect 8662 7692 8668 7704
rect 8720 7692 8726 7744
rect 9140 7732 9168 7763
rect 10888 7744 10916 7840
rect 11517 7837 11529 7840
rect 11563 7868 11575 7871
rect 11790 7868 11796 7880
rect 11563 7840 11796 7868
rect 11563 7837 11575 7840
rect 11517 7831 11575 7837
rect 11790 7828 11796 7840
rect 11848 7828 11854 7880
rect 11882 7828 11888 7880
rect 11940 7868 11946 7880
rect 15378 7868 15384 7880
rect 11940 7840 11985 7868
rect 15339 7840 15384 7868
rect 11940 7828 11946 7840
rect 15378 7828 15384 7840
rect 15436 7828 15442 7880
rect 17773 7871 17831 7877
rect 17773 7837 17785 7871
rect 17819 7868 17831 7871
rect 18506 7868 18512 7880
rect 17819 7840 18512 7868
rect 17819 7837 17831 7840
rect 17773 7831 17831 7837
rect 18506 7828 18512 7840
rect 18564 7828 18570 7880
rect 18874 7828 18880 7880
rect 18932 7868 18938 7880
rect 19337 7871 19395 7877
rect 19337 7868 19349 7871
rect 18932 7840 19349 7868
rect 18932 7828 18938 7840
rect 19337 7837 19349 7840
rect 19383 7868 19395 7871
rect 20901 7871 20959 7877
rect 20901 7868 20913 7871
rect 19383 7840 20913 7868
rect 19383 7837 19395 7840
rect 19337 7831 19395 7837
rect 20901 7837 20913 7840
rect 20947 7837 20959 7871
rect 20901 7831 20959 7837
rect 18322 7800 18328 7812
rect 18283 7772 18328 7800
rect 18322 7760 18328 7772
rect 18380 7760 18386 7812
rect 19702 7760 19708 7812
rect 19760 7800 19766 7812
rect 19889 7803 19947 7809
rect 19889 7800 19901 7803
rect 19760 7772 19901 7800
rect 19760 7760 19766 7772
rect 19889 7769 19901 7772
rect 19935 7769 19947 7803
rect 19889 7763 19947 7769
rect 9674 7732 9680 7744
rect 9140 7704 9680 7732
rect 9674 7692 9680 7704
rect 9732 7692 9738 7744
rect 10870 7732 10876 7744
rect 10831 7704 10876 7732
rect 10870 7692 10876 7704
rect 10928 7692 10934 7744
rect 12710 7692 12716 7744
rect 12768 7732 12774 7744
rect 13173 7735 13231 7741
rect 13173 7732 13185 7735
rect 12768 7704 13185 7732
rect 12768 7692 12774 7704
rect 13173 7701 13185 7704
rect 13219 7701 13231 7735
rect 13173 7695 13231 7701
rect 13633 7735 13691 7741
rect 13633 7701 13645 7735
rect 13679 7732 13691 7735
rect 13722 7732 13728 7744
rect 13679 7704 13728 7732
rect 13679 7701 13691 7704
rect 13633 7695 13691 7701
rect 13722 7692 13728 7704
rect 13780 7692 13786 7744
rect 16301 7735 16359 7741
rect 16301 7701 16313 7735
rect 16347 7732 16359 7735
rect 18969 7735 19027 7741
rect 18969 7732 18981 7735
rect 16347 7704 18981 7732
rect 16347 7701 16359 7704
rect 16301 7695 16359 7701
rect 18969 7701 18981 7704
rect 19015 7732 19027 7735
rect 19058 7732 19064 7744
rect 19015 7704 19064 7732
rect 19015 7701 19027 7704
rect 18969 7695 19027 7701
rect 19058 7692 19064 7704
rect 19116 7692 19122 7744
rect 1104 7642 22816 7664
rect 1104 7590 4982 7642
rect 5034 7590 5046 7642
rect 5098 7590 5110 7642
rect 5162 7590 5174 7642
rect 5226 7590 12982 7642
rect 13034 7590 13046 7642
rect 13098 7590 13110 7642
rect 13162 7590 13174 7642
rect 13226 7590 20982 7642
rect 21034 7590 21046 7642
rect 21098 7590 21110 7642
rect 21162 7590 21174 7642
rect 21226 7590 22816 7642
rect 1104 7568 22816 7590
rect 9766 7488 9772 7540
rect 9824 7528 9830 7540
rect 10873 7531 10931 7537
rect 10873 7528 10885 7531
rect 9824 7500 10885 7528
rect 9824 7488 9830 7500
rect 8294 7460 8300 7472
rect 7852 7432 8300 7460
rect 6270 7284 6276 7336
rect 6328 7324 6334 7336
rect 6641 7327 6699 7333
rect 6641 7324 6653 7327
rect 6328 7296 6653 7324
rect 6328 7284 6334 7296
rect 6641 7293 6653 7296
rect 6687 7324 6699 7327
rect 7101 7327 7159 7333
rect 7101 7324 7113 7327
rect 6687 7296 7113 7324
rect 6687 7293 6699 7296
rect 6641 7287 6699 7293
rect 7101 7293 7113 7296
rect 7147 7293 7159 7327
rect 7282 7324 7288 7336
rect 7243 7296 7288 7324
rect 7101 7287 7159 7293
rect 5905 7259 5963 7265
rect 5905 7225 5917 7259
rect 5951 7256 5963 7259
rect 7116 7256 7144 7287
rect 7282 7284 7288 7296
rect 7340 7284 7346 7336
rect 7650 7284 7656 7336
rect 7708 7324 7714 7336
rect 7852 7333 7880 7432
rect 8294 7420 8300 7432
rect 8352 7460 8358 7472
rect 9306 7460 9312 7472
rect 8352 7432 9312 7460
rect 8352 7420 8358 7432
rect 9306 7420 9312 7432
rect 9364 7420 9370 7472
rect 9784 7392 9812 7488
rect 8220 7364 9812 7392
rect 8220 7336 8248 7364
rect 7837 7327 7895 7333
rect 7837 7324 7849 7327
rect 7708 7296 7849 7324
rect 7708 7284 7714 7296
rect 7837 7293 7849 7296
rect 7883 7293 7895 7327
rect 8202 7324 8208 7336
rect 8115 7296 8208 7324
rect 7837 7287 7895 7293
rect 8202 7284 8208 7296
rect 8260 7284 8266 7336
rect 9401 7327 9459 7333
rect 9401 7324 9413 7327
rect 8312 7296 9413 7324
rect 8312 7256 8340 7296
rect 9401 7293 9413 7296
rect 9447 7324 9459 7327
rect 9490 7324 9496 7336
rect 9447 7296 9496 7324
rect 9447 7293 9459 7296
rect 9401 7287 9459 7293
rect 9490 7284 9496 7296
rect 9548 7284 9554 7336
rect 9674 7324 9680 7336
rect 9635 7296 9680 7324
rect 9674 7284 9680 7296
rect 9732 7284 9738 7336
rect 10336 7333 10364 7500
rect 10873 7497 10885 7500
rect 10919 7528 10931 7531
rect 11054 7528 11060 7540
rect 10919 7500 11060 7528
rect 10919 7497 10931 7500
rect 10873 7491 10931 7497
rect 11054 7488 11060 7500
rect 11112 7488 11118 7540
rect 11514 7528 11520 7540
rect 11475 7500 11520 7528
rect 11514 7488 11520 7500
rect 11572 7488 11578 7540
rect 11790 7528 11796 7540
rect 11751 7500 11796 7528
rect 11790 7488 11796 7500
rect 11848 7488 11854 7540
rect 18325 7531 18383 7537
rect 18325 7497 18337 7531
rect 18371 7528 18383 7531
rect 18506 7528 18512 7540
rect 18371 7500 18512 7528
rect 18371 7497 18383 7500
rect 18325 7491 18383 7497
rect 18506 7488 18512 7500
rect 18564 7488 18570 7540
rect 18874 7528 18880 7540
rect 18835 7500 18880 7528
rect 18874 7488 18880 7500
rect 18932 7488 18938 7540
rect 19426 7488 19432 7540
rect 19484 7528 19490 7540
rect 19981 7531 20039 7537
rect 19981 7528 19993 7531
rect 19484 7500 19993 7528
rect 19484 7488 19490 7500
rect 19981 7497 19993 7500
rect 20027 7497 20039 7531
rect 19981 7491 20039 7497
rect 10597 7395 10655 7401
rect 10597 7361 10609 7395
rect 10643 7392 10655 7395
rect 10870 7392 10876 7404
rect 10643 7364 10876 7392
rect 10643 7361 10655 7364
rect 10597 7355 10655 7361
rect 10870 7352 10876 7364
rect 10928 7352 10934 7404
rect 14645 7395 14703 7401
rect 14645 7361 14657 7395
rect 14691 7392 14703 7395
rect 15378 7392 15384 7404
rect 14691 7364 15384 7392
rect 14691 7361 14703 7364
rect 14645 7355 14703 7361
rect 15378 7352 15384 7364
rect 15436 7352 15442 7404
rect 19702 7392 19708 7404
rect 19663 7364 19708 7392
rect 19702 7352 19708 7364
rect 19760 7352 19766 7404
rect 9953 7327 10011 7333
rect 9953 7293 9965 7327
rect 9999 7293 10011 7327
rect 9953 7287 10011 7293
rect 10321 7327 10379 7333
rect 10321 7293 10333 7327
rect 10367 7293 10379 7327
rect 10321 7287 10379 7293
rect 9968 7256 9996 7287
rect 12710 7284 12716 7336
rect 12768 7324 12774 7336
rect 13173 7327 13231 7333
rect 13173 7324 13185 7327
rect 12768 7296 13185 7324
rect 12768 7284 12774 7296
rect 13173 7293 13185 7296
rect 13219 7293 13231 7327
rect 13633 7327 13691 7333
rect 13633 7324 13645 7327
rect 13173 7287 13231 7293
rect 13464 7296 13645 7324
rect 5951 7228 6776 7256
rect 7116 7228 8340 7256
rect 8956 7228 9996 7256
rect 5951 7225 5963 7228
rect 5905 7219 5963 7225
rect 6748 7200 6776 7228
rect 3050 7148 3056 7200
rect 3108 7188 3114 7200
rect 6181 7191 6239 7197
rect 6181 7188 6193 7191
rect 3108 7160 6193 7188
rect 3108 7148 3114 7160
rect 6181 7157 6193 7160
rect 6227 7188 6239 7191
rect 6638 7188 6644 7200
rect 6227 7160 6644 7188
rect 6227 7157 6239 7160
rect 6181 7151 6239 7157
rect 6638 7148 6644 7160
rect 6696 7148 6702 7200
rect 6730 7148 6736 7200
rect 6788 7188 6794 7200
rect 6917 7191 6975 7197
rect 6917 7188 6929 7191
rect 6788 7160 6929 7188
rect 6788 7148 6794 7160
rect 6917 7157 6929 7160
rect 6963 7157 6975 7191
rect 8662 7188 8668 7200
rect 8623 7160 8668 7188
rect 6917 7151 6975 7157
rect 8662 7148 8668 7160
rect 8720 7148 8726 7200
rect 8846 7148 8852 7200
rect 8904 7188 8910 7200
rect 8956 7197 8984 7228
rect 13464 7200 13492 7296
rect 13633 7293 13645 7296
rect 13679 7293 13691 7327
rect 13633 7287 13691 7293
rect 13722 7284 13728 7336
rect 13780 7324 13786 7336
rect 14001 7327 14059 7333
rect 14001 7324 14013 7327
rect 13780 7296 14013 7324
rect 13780 7284 13786 7296
rect 14001 7293 14013 7296
rect 14047 7293 14059 7327
rect 14001 7287 14059 7293
rect 14274 7284 14280 7336
rect 14332 7324 14338 7336
rect 14369 7327 14427 7333
rect 14369 7324 14381 7327
rect 14332 7296 14381 7324
rect 14332 7284 14338 7296
rect 14369 7293 14381 7296
rect 14415 7293 14427 7327
rect 15657 7327 15715 7333
rect 15657 7324 15669 7327
rect 14369 7287 14427 7293
rect 15028 7296 15669 7324
rect 8941 7191 8999 7197
rect 8941 7188 8953 7191
rect 8904 7160 8953 7188
rect 8904 7148 8910 7160
rect 8941 7157 8953 7160
rect 8987 7157 8999 7191
rect 8941 7151 8999 7157
rect 9306 7148 9312 7200
rect 9364 7188 9370 7200
rect 12526 7188 12532 7200
rect 9364 7160 12532 7188
rect 9364 7148 9370 7160
rect 12526 7148 12532 7160
rect 12584 7188 12590 7200
rect 12621 7191 12679 7197
rect 12621 7188 12633 7191
rect 12584 7160 12633 7188
rect 12584 7148 12590 7160
rect 12621 7157 12633 7160
rect 12667 7157 12679 7191
rect 12621 7151 12679 7157
rect 13081 7191 13139 7197
rect 13081 7157 13093 7191
rect 13127 7188 13139 7191
rect 13446 7188 13452 7200
rect 13127 7160 13452 7188
rect 13127 7157 13139 7160
rect 13081 7151 13139 7157
rect 13446 7148 13452 7160
rect 13504 7148 13510 7200
rect 13630 7148 13636 7200
rect 13688 7188 13694 7200
rect 14384 7188 14412 7287
rect 15028 7200 15056 7296
rect 15657 7293 15669 7296
rect 15703 7293 15715 7327
rect 15657 7287 15715 7293
rect 15978 7259 16036 7265
rect 15978 7225 15990 7259
rect 16024 7225 16036 7259
rect 15978 7219 16036 7225
rect 15010 7188 15016 7200
rect 13688 7160 14412 7188
rect 14971 7160 15016 7188
rect 13688 7148 13694 7160
rect 15010 7148 15016 7160
rect 15068 7148 15074 7200
rect 15473 7191 15531 7197
rect 15473 7157 15485 7191
rect 15519 7188 15531 7191
rect 15838 7188 15844 7200
rect 15519 7160 15844 7188
rect 15519 7157 15531 7160
rect 15473 7151 15531 7157
rect 15838 7148 15844 7160
rect 15896 7188 15902 7200
rect 15993 7188 16021 7219
rect 18322 7216 18328 7268
rect 18380 7256 18386 7268
rect 19061 7259 19119 7265
rect 19061 7256 19073 7259
rect 18380 7228 19073 7256
rect 18380 7216 18386 7228
rect 19061 7225 19073 7228
rect 19107 7225 19119 7259
rect 19061 7219 19119 7225
rect 19150 7216 19156 7268
rect 19208 7256 19214 7268
rect 19208 7228 19253 7256
rect 19208 7216 19214 7228
rect 16574 7188 16580 7200
rect 15896 7160 16021 7188
rect 16535 7160 16580 7188
rect 15896 7148 15902 7160
rect 16574 7148 16580 7160
rect 16632 7148 16638 7200
rect 17773 7191 17831 7197
rect 17773 7157 17785 7191
rect 17819 7188 17831 7191
rect 18046 7188 18052 7200
rect 17819 7160 18052 7188
rect 17819 7157 17831 7160
rect 17773 7151 17831 7157
rect 18046 7148 18052 7160
rect 18104 7148 18110 7200
rect 1104 7098 22816 7120
rect 1104 7046 8982 7098
rect 9034 7046 9046 7098
rect 9098 7046 9110 7098
rect 9162 7046 9174 7098
rect 9226 7046 16982 7098
rect 17034 7046 17046 7098
rect 17098 7046 17110 7098
rect 17162 7046 17174 7098
rect 17226 7046 22816 7098
rect 1104 7024 22816 7046
rect 7653 6987 7711 6993
rect 7653 6953 7665 6987
rect 7699 6984 7711 6987
rect 8202 6984 8208 6996
rect 7699 6956 8208 6984
rect 7699 6953 7711 6956
rect 7653 6947 7711 6953
rect 8202 6944 8208 6956
rect 8260 6944 8266 6996
rect 8386 6944 8392 6996
rect 8444 6984 8450 6996
rect 8619 6987 8677 6993
rect 8619 6984 8631 6987
rect 8444 6956 8631 6984
rect 8444 6944 8450 6956
rect 8619 6953 8631 6956
rect 8665 6953 8677 6987
rect 8619 6947 8677 6953
rect 9217 6987 9275 6993
rect 9217 6953 9229 6987
rect 9263 6984 9275 6987
rect 9490 6984 9496 6996
rect 9263 6956 9496 6984
rect 9263 6953 9275 6956
rect 9217 6947 9275 6953
rect 9490 6944 9496 6956
rect 9548 6944 9554 6996
rect 9953 6987 10011 6993
rect 9953 6953 9965 6987
rect 9999 6984 10011 6987
rect 10042 6984 10048 6996
rect 9999 6956 10048 6984
rect 9999 6953 10011 6956
rect 9953 6947 10011 6953
rect 10042 6944 10048 6956
rect 10100 6944 10106 6996
rect 11054 6984 11060 6996
rect 11015 6956 11060 6984
rect 11054 6944 11060 6956
rect 11112 6944 11118 6996
rect 12526 6944 12532 6996
rect 12584 6984 12590 6996
rect 13630 6984 13636 6996
rect 12584 6956 13636 6984
rect 12584 6944 12590 6956
rect 13630 6944 13636 6956
rect 13688 6944 13694 6996
rect 15378 6944 15384 6996
rect 15436 6984 15442 6996
rect 16117 6987 16175 6993
rect 16117 6984 16129 6987
rect 15436 6956 16129 6984
rect 15436 6944 15442 6956
rect 16117 6953 16129 6956
rect 16163 6953 16175 6987
rect 19058 6984 19064 6996
rect 19019 6956 19064 6984
rect 16117 6947 16175 6953
rect 19058 6944 19064 6956
rect 19116 6944 19122 6996
rect 9582 6876 9588 6928
rect 9640 6916 9646 6928
rect 12618 6916 12624 6928
rect 9640 6888 12624 6916
rect 9640 6876 9646 6888
rect 12618 6876 12624 6888
rect 12676 6876 12682 6928
rect 14369 6919 14427 6925
rect 14369 6885 14381 6919
rect 14415 6916 14427 6919
rect 15010 6916 15016 6928
rect 14415 6888 15016 6916
rect 14415 6885 14427 6888
rect 14369 6879 14427 6885
rect 15010 6876 15016 6888
rect 15068 6876 15074 6928
rect 16574 6876 16580 6928
rect 16632 6916 16638 6928
rect 17862 6916 17868 6928
rect 16632 6888 17868 6916
rect 16632 6876 16638 6888
rect 17862 6876 17868 6888
rect 17920 6916 17926 6928
rect 17957 6919 18015 6925
rect 17957 6916 17969 6919
rect 17920 6888 17969 6916
rect 17920 6876 17926 6888
rect 17957 6885 17969 6888
rect 18003 6885 18015 6919
rect 17957 6879 18015 6885
rect 7285 6851 7343 6857
rect 7285 6817 7297 6851
rect 7331 6848 7343 6851
rect 7650 6848 7656 6860
rect 7331 6820 7656 6848
rect 7331 6817 7343 6820
rect 7285 6811 7343 6817
rect 7650 6808 7656 6820
rect 7708 6808 7714 6860
rect 8548 6851 8606 6857
rect 8548 6817 8560 6851
rect 8594 6848 8606 6851
rect 9600 6848 9628 6876
rect 10410 6848 10416 6860
rect 8594 6820 9628 6848
rect 10371 6820 10416 6848
rect 8594 6817 8606 6820
rect 8548 6811 8606 6817
rect 10410 6808 10416 6820
rect 10468 6808 10474 6860
rect 12710 6808 12716 6860
rect 12768 6848 12774 6860
rect 12897 6851 12955 6857
rect 12897 6848 12909 6851
rect 12768 6820 12909 6848
rect 12768 6808 12774 6820
rect 12897 6817 12909 6820
rect 12943 6817 12955 6851
rect 13446 6848 13452 6860
rect 13407 6820 13452 6848
rect 12897 6811 12955 6817
rect 13446 6808 13452 6820
rect 13504 6808 13510 6860
rect 13722 6848 13728 6860
rect 13635 6820 13728 6848
rect 13722 6808 13728 6820
rect 13780 6808 13786 6860
rect 14277 6851 14335 6857
rect 14277 6817 14289 6851
rect 14323 6848 14335 6851
rect 14642 6848 14648 6860
rect 14323 6820 14648 6848
rect 14323 6817 14335 6820
rect 14277 6811 14335 6817
rect 14642 6808 14648 6820
rect 14700 6808 14706 6860
rect 15197 6851 15255 6857
rect 15197 6817 15209 6851
rect 15243 6848 15255 6851
rect 15286 6848 15292 6860
rect 15243 6820 15292 6848
rect 15243 6817 15255 6820
rect 15197 6811 15255 6817
rect 15286 6808 15292 6820
rect 15344 6808 15350 6860
rect 16828 6851 16886 6857
rect 16828 6817 16840 6851
rect 16874 6848 16886 6851
rect 17034 6848 17040 6860
rect 16874 6820 17040 6848
rect 16874 6817 16886 6820
rect 16828 6811 16886 6817
rect 17034 6808 17040 6820
rect 17092 6848 17098 6860
rect 17310 6848 17316 6860
rect 17092 6820 17316 6848
rect 17092 6808 17098 6820
rect 17310 6808 17316 6820
rect 17368 6808 17374 6860
rect 10042 6740 10048 6792
rect 10100 6780 10106 6792
rect 10781 6783 10839 6789
rect 10781 6780 10793 6783
rect 10100 6752 10793 6780
rect 10100 6740 10106 6752
rect 10781 6749 10793 6752
rect 10827 6749 10839 6783
rect 13740 6780 13768 6808
rect 17865 6783 17923 6789
rect 17865 6780 17877 6783
rect 10781 6743 10839 6749
rect 12360 6752 13768 6780
rect 17420 6752 17877 6780
rect 7282 6712 7288 6724
rect 6840 6684 7288 6712
rect 4798 6604 4804 6656
rect 4856 6644 4862 6656
rect 6840 6653 6868 6684
rect 7282 6672 7288 6684
rect 7340 6672 7346 6724
rect 9766 6672 9772 6724
rect 9824 6712 9830 6724
rect 11514 6712 11520 6724
rect 9824 6684 11520 6712
rect 9824 6672 9830 6684
rect 11514 6672 11520 6684
rect 11572 6712 11578 6724
rect 12360 6721 12388 6752
rect 12345 6715 12403 6721
rect 12345 6712 12357 6715
rect 11572 6684 12357 6712
rect 11572 6672 11578 6684
rect 12345 6681 12357 6684
rect 12391 6681 12403 6715
rect 12345 6675 12403 6681
rect 17420 6656 17448 6752
rect 17865 6749 17877 6752
rect 17911 6749 17923 6783
rect 18322 6780 18328 6792
rect 18283 6752 18328 6780
rect 17865 6743 17923 6749
rect 18322 6740 18328 6752
rect 18380 6780 18386 6792
rect 19337 6783 19395 6789
rect 19337 6780 19349 6783
rect 18380 6752 19349 6780
rect 18380 6740 18386 6752
rect 19337 6749 19349 6752
rect 19383 6749 19395 6783
rect 19337 6743 19395 6749
rect 10594 6653 10600 6656
rect 6825 6647 6883 6653
rect 6825 6644 6837 6647
rect 4856 6616 6837 6644
rect 4856 6604 4862 6616
rect 6825 6613 6837 6616
rect 6871 6613 6883 6647
rect 6825 6607 6883 6613
rect 10321 6647 10379 6653
rect 10321 6613 10333 6647
rect 10367 6644 10379 6647
rect 10551 6647 10600 6653
rect 10551 6644 10563 6647
rect 10367 6616 10563 6644
rect 10367 6613 10379 6616
rect 10321 6607 10379 6613
rect 10551 6613 10563 6616
rect 10597 6613 10600 6647
rect 10551 6607 10600 6613
rect 10594 6604 10600 6607
rect 10652 6604 10658 6656
rect 10686 6604 10692 6656
rect 10744 6644 10750 6656
rect 12710 6644 12716 6656
rect 10744 6616 10789 6644
rect 12671 6616 12716 6644
rect 10744 6604 10750 6616
rect 12710 6604 12716 6616
rect 12768 6604 12774 6656
rect 15427 6647 15485 6653
rect 15427 6613 15439 6647
rect 15473 6644 15485 6647
rect 15562 6644 15568 6656
rect 15473 6616 15568 6644
rect 15473 6613 15485 6616
rect 15427 6607 15485 6613
rect 15562 6604 15568 6616
rect 15620 6604 15626 6656
rect 15838 6644 15844 6656
rect 15799 6616 15844 6644
rect 15838 6604 15844 6616
rect 15896 6604 15902 6656
rect 16899 6647 16957 6653
rect 16899 6613 16911 6647
rect 16945 6644 16957 6647
rect 17402 6644 17408 6656
rect 16945 6616 17408 6644
rect 16945 6613 16957 6616
rect 16899 6607 16957 6613
rect 17402 6604 17408 6616
rect 17460 6604 17466 6656
rect 1104 6554 22816 6576
rect 1104 6502 4982 6554
rect 5034 6502 5046 6554
rect 5098 6502 5110 6554
rect 5162 6502 5174 6554
rect 5226 6502 12982 6554
rect 13034 6502 13046 6554
rect 13098 6502 13110 6554
rect 13162 6502 13174 6554
rect 13226 6502 20982 6554
rect 21034 6502 21046 6554
rect 21098 6502 21110 6554
rect 21162 6502 21174 6554
rect 21226 6502 22816 6554
rect 1104 6480 22816 6502
rect 10686 6400 10692 6452
rect 10744 6440 10750 6452
rect 11609 6443 11667 6449
rect 11609 6440 11621 6443
rect 10744 6412 11621 6440
rect 10744 6400 10750 6412
rect 11609 6409 11621 6412
rect 11655 6409 11667 6443
rect 15286 6440 15292 6452
rect 15247 6412 15292 6440
rect 11609 6403 11667 6409
rect 15286 6400 15292 6412
rect 15344 6400 15350 6452
rect 16022 6400 16028 6452
rect 16080 6440 16086 6452
rect 16669 6443 16727 6449
rect 16669 6440 16681 6443
rect 16080 6412 16681 6440
rect 16080 6400 16086 6412
rect 16669 6409 16681 6412
rect 16715 6409 16727 6443
rect 17402 6440 17408 6452
rect 17363 6412 17408 6440
rect 16669 6403 16727 6409
rect 17402 6400 17408 6412
rect 17460 6400 17466 6452
rect 17862 6440 17868 6452
rect 17823 6412 17868 6440
rect 17862 6400 17868 6412
rect 17920 6400 17926 6452
rect 8846 6332 8852 6384
rect 8904 6372 8910 6384
rect 12802 6372 12808 6384
rect 8904 6344 12808 6372
rect 8904 6332 8910 6344
rect 12802 6332 12808 6344
rect 12860 6372 12866 6384
rect 12897 6375 12955 6381
rect 12897 6372 12909 6375
rect 12860 6344 12909 6372
rect 12860 6332 12866 6344
rect 12897 6341 12909 6344
rect 12943 6372 12955 6375
rect 13262 6372 13268 6384
rect 12943 6344 13268 6372
rect 12943 6341 12955 6344
rect 12897 6335 12955 6341
rect 13262 6332 13268 6344
rect 13320 6372 13326 6384
rect 13630 6372 13636 6384
rect 13320 6344 13636 6372
rect 13320 6332 13326 6344
rect 13630 6332 13636 6344
rect 13688 6332 13694 6384
rect 9766 6304 9772 6316
rect 9727 6276 9772 6304
rect 9766 6264 9772 6276
rect 9824 6264 9830 6316
rect 10594 6304 10600 6316
rect 10555 6276 10600 6304
rect 10594 6264 10600 6276
rect 10652 6264 10658 6316
rect 18046 6304 18052 6316
rect 18007 6276 18052 6304
rect 18046 6264 18052 6276
rect 18104 6264 18110 6316
rect 9125 6239 9183 6245
rect 9125 6205 9137 6239
rect 9171 6236 9183 6239
rect 9401 6239 9459 6245
rect 9401 6236 9413 6239
rect 9171 6208 9413 6236
rect 9171 6205 9183 6208
rect 9125 6199 9183 6205
rect 9401 6205 9413 6208
rect 9447 6236 9459 6239
rect 10612 6236 10640 6264
rect 11238 6236 11244 6248
rect 9447 6208 10640 6236
rect 11199 6208 11244 6236
rect 9447 6205 9459 6208
rect 9401 6199 9459 6205
rect 11238 6196 11244 6208
rect 11296 6196 11302 6248
rect 13354 6196 13360 6248
rect 13412 6236 13418 6248
rect 13449 6239 13507 6245
rect 13449 6236 13461 6239
rect 13412 6208 13461 6236
rect 13412 6196 13418 6208
rect 13449 6205 13461 6208
rect 13495 6205 13507 6239
rect 13909 6239 13967 6245
rect 13909 6236 13921 6239
rect 13449 6199 13507 6205
rect 13556 6208 13921 6236
rect 9217 6171 9275 6177
rect 9217 6137 9229 6171
rect 9263 6168 9275 6171
rect 9306 6168 9312 6180
rect 9263 6140 9312 6168
rect 9263 6137 9275 6140
rect 9217 6131 9275 6137
rect 9306 6128 9312 6140
rect 9364 6128 9370 6180
rect 10505 6171 10563 6177
rect 10505 6137 10517 6171
rect 10551 6168 10563 6171
rect 11256 6168 11284 6196
rect 10551 6140 11284 6168
rect 10551 6137 10563 6140
rect 10505 6131 10563 6137
rect 8573 6103 8631 6109
rect 8573 6069 8585 6103
rect 8619 6100 8631 6103
rect 9582 6100 9588 6112
rect 8619 6072 9588 6100
rect 8619 6069 8631 6072
rect 8573 6063 8631 6069
rect 9582 6060 9588 6072
rect 9640 6060 9646 6112
rect 10042 6100 10048 6112
rect 10003 6072 10048 6100
rect 10042 6060 10048 6072
rect 10100 6060 10106 6112
rect 12066 6060 12072 6112
rect 12124 6100 12130 6112
rect 12161 6103 12219 6109
rect 12161 6100 12173 6103
rect 12124 6072 12173 6100
rect 12124 6060 12130 6072
rect 12161 6069 12173 6072
rect 12207 6069 12219 6103
rect 12161 6063 12219 6069
rect 13446 6060 13452 6112
rect 13504 6100 13510 6112
rect 13556 6100 13584 6208
rect 13909 6205 13921 6208
rect 13955 6205 13967 6239
rect 14274 6236 14280 6248
rect 14235 6208 14280 6236
rect 13909 6199 13967 6205
rect 14274 6196 14280 6208
rect 14332 6196 14338 6248
rect 14642 6236 14648 6248
rect 14603 6208 14648 6236
rect 14642 6196 14648 6208
rect 14700 6196 14706 6248
rect 14921 6239 14979 6245
rect 14921 6205 14933 6239
rect 14967 6236 14979 6239
rect 15746 6236 15752 6248
rect 14967 6208 15752 6236
rect 14967 6205 14979 6208
rect 14921 6199 14979 6205
rect 15746 6196 15752 6208
rect 15804 6196 15810 6248
rect 17862 6196 17868 6248
rect 17920 6236 17926 6248
rect 18141 6239 18199 6245
rect 18141 6236 18153 6239
rect 17920 6208 18153 6236
rect 17920 6196 17926 6208
rect 18141 6205 18153 6208
rect 18187 6205 18199 6239
rect 18141 6199 18199 6205
rect 13504 6072 13584 6100
rect 13504 6060 13510 6072
rect 13630 6060 13636 6112
rect 13688 6100 13694 6112
rect 14660 6100 14688 6196
rect 15838 6128 15844 6180
rect 15896 6168 15902 6180
rect 16070 6171 16128 6177
rect 16070 6168 16082 6171
rect 15896 6140 16082 6168
rect 15896 6128 15902 6140
rect 16070 6137 16082 6140
rect 16116 6137 16128 6171
rect 17034 6168 17040 6180
rect 16947 6140 17040 6168
rect 16070 6131 16128 6137
rect 17034 6128 17040 6140
rect 17092 6168 17098 6180
rect 18322 6168 18328 6180
rect 17092 6140 18328 6168
rect 17092 6128 17098 6140
rect 18322 6128 18328 6140
rect 18380 6128 18386 6180
rect 13688 6072 14688 6100
rect 13688 6060 13694 6072
rect 1104 6010 22816 6032
rect 1104 5958 8982 6010
rect 9034 5958 9046 6010
rect 9098 5958 9110 6010
rect 9162 5958 9174 6010
rect 9226 5958 16982 6010
rect 17034 5958 17046 6010
rect 17098 5958 17110 6010
rect 17162 5958 17174 6010
rect 17226 5958 22816 6010
rect 1104 5936 22816 5958
rect 15746 5856 15752 5908
rect 15804 5896 15810 5908
rect 16117 5899 16175 5905
rect 16117 5896 16129 5899
rect 15804 5868 16129 5896
rect 15804 5856 15810 5868
rect 16117 5865 16129 5868
rect 16163 5865 16175 5899
rect 16117 5859 16175 5865
rect 17862 5856 17868 5908
rect 17920 5896 17926 5908
rect 18049 5899 18107 5905
rect 18049 5896 18061 5899
rect 17920 5868 18061 5896
rect 17920 5856 17926 5868
rect 18049 5865 18061 5868
rect 18095 5865 18107 5899
rect 18049 5859 18107 5865
rect 11330 5828 11336 5840
rect 11291 5800 11336 5828
rect 11330 5788 11336 5800
rect 11388 5788 11394 5840
rect 12897 5831 12955 5837
rect 12897 5797 12909 5831
rect 12943 5828 12955 5831
rect 13998 5828 14004 5840
rect 12943 5800 14004 5828
rect 12943 5797 12955 5800
rect 12897 5791 12955 5797
rect 13998 5788 14004 5800
rect 14056 5788 14062 5840
rect 16942 5828 16948 5840
rect 16903 5800 16948 5828
rect 16942 5788 16948 5800
rect 17000 5788 17006 5840
rect 9306 5760 9312 5772
rect 9219 5732 9312 5760
rect 9306 5720 9312 5732
rect 9364 5760 9370 5772
rect 9858 5760 9864 5772
rect 9364 5732 9864 5760
rect 9364 5720 9370 5732
rect 9858 5720 9864 5732
rect 9916 5760 9922 5772
rect 10045 5763 10103 5769
rect 10045 5760 10057 5763
rect 9916 5732 10057 5760
rect 9916 5720 9922 5732
rect 10045 5729 10057 5732
rect 10091 5760 10103 5763
rect 10410 5760 10416 5772
rect 10091 5732 10416 5760
rect 10091 5729 10103 5732
rect 10045 5723 10103 5729
rect 10410 5720 10416 5732
rect 10468 5760 10474 5772
rect 10597 5763 10655 5769
rect 10597 5760 10609 5763
rect 10468 5732 10609 5760
rect 10468 5720 10474 5732
rect 10597 5729 10609 5732
rect 10643 5760 10655 5763
rect 11882 5760 11888 5772
rect 10643 5732 11888 5760
rect 10643 5729 10655 5732
rect 10597 5723 10655 5729
rect 11882 5720 11888 5732
rect 11940 5720 11946 5772
rect 12158 5760 12164 5772
rect 12119 5732 12164 5760
rect 12158 5720 12164 5732
rect 12216 5720 12222 5772
rect 18322 5760 18328 5772
rect 18283 5732 18328 5760
rect 18322 5720 18328 5732
rect 18380 5720 18386 5772
rect 10134 5652 10140 5704
rect 10192 5692 10198 5704
rect 10870 5692 10876 5704
rect 10192 5664 10876 5692
rect 10192 5652 10198 5664
rect 10870 5652 10876 5664
rect 10928 5692 10934 5704
rect 10965 5695 11023 5701
rect 10965 5692 10977 5695
rect 10928 5664 10977 5692
rect 10928 5652 10934 5664
rect 10965 5661 10977 5664
rect 11011 5661 11023 5695
rect 10965 5655 11023 5661
rect 11790 5652 11796 5704
rect 11848 5692 11854 5704
rect 12529 5695 12587 5701
rect 12529 5692 12541 5695
rect 11848 5664 12541 5692
rect 11848 5652 11854 5664
rect 12529 5661 12541 5664
rect 12575 5661 12587 5695
rect 12529 5655 12587 5661
rect 16853 5695 16911 5701
rect 16853 5661 16865 5695
rect 16899 5661 16911 5695
rect 16853 5655 16911 5661
rect 10762 5627 10820 5633
rect 10762 5593 10774 5627
rect 10808 5624 10820 5627
rect 11238 5624 11244 5636
rect 10808 5596 11244 5624
rect 10808 5593 10820 5596
rect 10762 5587 10820 5593
rect 11238 5584 11244 5596
rect 11296 5624 11302 5636
rect 11808 5624 11836 5652
rect 11296 5596 11836 5624
rect 11296 5584 11302 5596
rect 11882 5584 11888 5636
rect 11940 5624 11946 5636
rect 12069 5627 12127 5633
rect 12069 5624 12081 5627
rect 11940 5596 12081 5624
rect 11940 5584 11946 5596
rect 12069 5593 12081 5596
rect 12115 5624 12127 5627
rect 12437 5627 12495 5633
rect 12437 5624 12449 5627
rect 12115 5596 12449 5624
rect 12115 5593 12127 5596
rect 12069 5587 12127 5593
rect 12437 5593 12449 5596
rect 12483 5593 12495 5627
rect 12437 5587 12495 5593
rect 13354 5584 13360 5636
rect 13412 5624 13418 5636
rect 13817 5627 13875 5633
rect 13817 5624 13829 5627
rect 13412 5596 13829 5624
rect 13412 5584 13418 5596
rect 13817 5593 13829 5596
rect 13863 5593 13875 5627
rect 13817 5587 13875 5593
rect 16758 5584 16764 5636
rect 16816 5624 16822 5636
rect 16868 5624 16896 5655
rect 17402 5624 17408 5636
rect 16816 5596 16896 5624
rect 17363 5596 17408 5624
rect 16816 5584 16822 5596
rect 17402 5584 17408 5596
rect 17460 5584 17466 5636
rect 17770 5584 17776 5636
rect 17828 5624 17834 5636
rect 18509 5627 18567 5633
rect 18509 5624 18521 5627
rect 17828 5596 18521 5624
rect 17828 5584 17834 5596
rect 18509 5593 18521 5596
rect 18555 5593 18567 5627
rect 18509 5587 18567 5593
rect 10410 5556 10416 5568
rect 10371 5528 10416 5556
rect 10410 5516 10416 5528
rect 10468 5556 10474 5568
rect 10873 5559 10931 5565
rect 10873 5556 10885 5559
rect 10468 5528 10885 5556
rect 10468 5516 10474 5528
rect 10873 5525 10885 5528
rect 10919 5525 10931 5559
rect 10873 5519 10931 5525
rect 12326 5559 12384 5565
rect 12326 5525 12338 5559
rect 12372 5556 12384 5559
rect 12710 5556 12716 5568
rect 12372 5528 12716 5556
rect 12372 5525 12384 5528
rect 12326 5519 12384 5525
rect 12710 5516 12716 5528
rect 12768 5516 12774 5568
rect 13446 5556 13452 5568
rect 13407 5528 13452 5556
rect 13446 5516 13452 5528
rect 13504 5516 13510 5568
rect 14274 5556 14280 5568
rect 14235 5528 14280 5556
rect 14274 5516 14280 5528
rect 14332 5516 14338 5568
rect 15746 5556 15752 5568
rect 15707 5528 15752 5556
rect 15746 5516 15752 5528
rect 15804 5516 15810 5568
rect 1104 5466 22816 5488
rect 1104 5414 4982 5466
rect 5034 5414 5046 5466
rect 5098 5414 5110 5466
rect 5162 5414 5174 5466
rect 5226 5414 12982 5466
rect 13034 5414 13046 5466
rect 13098 5414 13110 5466
rect 13162 5414 13174 5466
rect 13226 5414 20982 5466
rect 21034 5414 21046 5466
rect 21098 5414 21110 5466
rect 21162 5414 21174 5466
rect 21226 5414 22816 5466
rect 1104 5392 22816 5414
rect 9858 5352 9864 5364
rect 9819 5324 9864 5352
rect 9858 5312 9864 5324
rect 9916 5312 9922 5364
rect 10686 5312 10692 5364
rect 10744 5352 10750 5364
rect 10781 5355 10839 5361
rect 10781 5352 10793 5355
rect 10744 5324 10793 5352
rect 10744 5312 10750 5324
rect 10781 5321 10793 5324
rect 10827 5352 10839 5355
rect 11793 5355 11851 5361
rect 11793 5352 11805 5355
rect 10827 5324 11805 5352
rect 10827 5321 10839 5324
rect 10781 5315 10839 5321
rect 11793 5321 11805 5324
rect 11839 5352 11851 5355
rect 12158 5352 12164 5364
rect 11839 5324 12164 5352
rect 11839 5321 11851 5324
rect 11793 5315 11851 5321
rect 12158 5312 12164 5324
rect 12216 5312 12222 5364
rect 16758 5312 16764 5364
rect 16816 5352 16822 5364
rect 17221 5355 17279 5361
rect 17221 5352 17233 5355
rect 16816 5324 17233 5352
rect 16816 5312 16822 5324
rect 17221 5321 17233 5324
rect 17267 5321 17279 5355
rect 18322 5352 18328 5364
rect 18283 5324 18328 5352
rect 17221 5315 17279 5321
rect 18322 5312 18328 5324
rect 18380 5312 18386 5364
rect 10870 5244 10876 5296
rect 10928 5284 10934 5296
rect 12621 5287 12679 5293
rect 12621 5284 12633 5287
rect 10928 5256 12633 5284
rect 10928 5244 10934 5256
rect 12621 5253 12633 5256
rect 12667 5284 12679 5287
rect 12710 5284 12716 5296
rect 12667 5256 12716 5284
rect 12667 5253 12679 5256
rect 12621 5247 12679 5253
rect 12710 5244 12716 5256
rect 12768 5244 12774 5296
rect 7650 5216 7656 5228
rect 7611 5188 7656 5216
rect 7650 5176 7656 5188
rect 7708 5176 7714 5228
rect 12066 5176 12072 5228
rect 12124 5216 12130 5228
rect 13173 5219 13231 5225
rect 13173 5216 13185 5219
rect 12124 5188 13185 5216
rect 12124 5176 12130 5188
rect 13173 5185 13185 5188
rect 13219 5216 13231 5219
rect 13446 5216 13452 5228
rect 13219 5188 13452 5216
rect 13219 5185 13231 5188
rect 13173 5179 13231 5185
rect 13446 5176 13452 5188
rect 13504 5216 13510 5228
rect 13504 5188 13860 5216
rect 13504 5176 13510 5188
rect 6546 5108 6552 5160
rect 6604 5148 6610 5160
rect 7009 5151 7067 5157
rect 7009 5148 7021 5151
rect 6604 5120 7021 5148
rect 6604 5108 6610 5120
rect 7009 5117 7021 5120
rect 7055 5148 7067 5151
rect 8846 5148 8852 5160
rect 7055 5120 8852 5148
rect 7055 5117 7067 5120
rect 7009 5111 7067 5117
rect 8846 5108 8852 5120
rect 8904 5108 8910 5160
rect 10410 5148 10416 5160
rect 10323 5120 10416 5148
rect 10410 5108 10416 5120
rect 10468 5108 10474 5160
rect 13354 5148 13360 5160
rect 13315 5120 13360 5148
rect 13354 5108 13360 5120
rect 13412 5108 13418 5160
rect 13832 5157 13860 5188
rect 14274 5176 14280 5228
rect 14332 5216 14338 5228
rect 15105 5219 15163 5225
rect 15105 5216 15117 5219
rect 14332 5188 15117 5216
rect 14332 5176 14338 5188
rect 14384 5157 14412 5188
rect 15105 5185 15117 5188
rect 15151 5185 15163 5219
rect 15105 5179 15163 5185
rect 13817 5151 13875 5157
rect 13817 5117 13829 5151
rect 13863 5117 13875 5151
rect 13817 5111 13875 5117
rect 14369 5151 14427 5157
rect 14369 5117 14381 5151
rect 14415 5117 14427 5151
rect 14550 5148 14556 5160
rect 14511 5120 14556 5148
rect 14369 5111 14427 5117
rect 106 5040 112 5092
rect 164 5080 170 5092
rect 10137 5083 10195 5089
rect 10137 5080 10149 5083
rect 164 5052 10149 5080
rect 164 5040 170 5052
rect 10137 5049 10149 5052
rect 10183 5080 10195 5083
rect 10428 5080 10456 5108
rect 10183 5052 10456 5080
rect 10183 5049 10195 5052
rect 10137 5043 10195 5049
rect 11974 5040 11980 5092
rect 12032 5080 12038 5092
rect 14384 5080 14412 5111
rect 14550 5108 14556 5120
rect 14608 5108 14614 5160
rect 14829 5151 14887 5157
rect 14829 5117 14841 5151
rect 14875 5148 14887 5151
rect 15654 5148 15660 5160
rect 14875 5120 15660 5148
rect 14875 5117 14887 5120
rect 14829 5111 14887 5117
rect 15654 5108 15660 5120
rect 15712 5108 15718 5160
rect 12032 5052 14412 5080
rect 15978 5083 16036 5089
rect 12032 5040 12038 5052
rect 15978 5049 15990 5083
rect 16024 5049 16036 5083
rect 16942 5080 16948 5092
rect 15978 5043 16036 5049
rect 16592 5052 16948 5080
rect 6546 5012 6552 5024
rect 6507 4984 6552 5012
rect 6546 4972 6552 4984
rect 6604 4972 6610 5024
rect 11425 5015 11483 5021
rect 11425 4981 11437 5015
rect 11471 5012 11483 5015
rect 11790 5012 11796 5024
rect 11471 4984 11796 5012
rect 11471 4981 11483 4984
rect 11425 4975 11483 4981
rect 11790 4972 11796 4984
rect 11848 5012 11854 5024
rect 12161 5015 12219 5021
rect 12161 5012 12173 5015
rect 11848 4984 12173 5012
rect 11848 4972 11854 4984
rect 12161 4981 12173 4984
rect 12207 4981 12219 5015
rect 12161 4975 12219 4981
rect 15194 4972 15200 5024
rect 15252 5012 15258 5024
rect 15473 5015 15531 5021
rect 15473 5012 15485 5015
rect 15252 4984 15485 5012
rect 15252 4972 15258 4984
rect 15473 4981 15485 4984
rect 15519 5012 15531 5015
rect 15746 5012 15752 5024
rect 15519 4984 15752 5012
rect 15519 4981 15531 4984
rect 15473 4975 15531 4981
rect 15746 4972 15752 4984
rect 15804 5012 15810 5024
rect 15993 5012 16021 5043
rect 16592 5021 16620 5052
rect 16942 5040 16948 5052
rect 17000 5080 17006 5092
rect 18506 5080 18512 5092
rect 17000 5052 18512 5080
rect 17000 5040 17006 5052
rect 18506 5040 18512 5052
rect 18564 5040 18570 5092
rect 15804 4984 16021 5012
rect 16577 5015 16635 5021
rect 15804 4972 15810 4984
rect 16577 4981 16589 5015
rect 16623 4981 16635 5015
rect 16577 4975 16635 4981
rect 1104 4922 22816 4944
rect 1104 4870 8982 4922
rect 9034 4870 9046 4922
rect 9098 4870 9110 4922
rect 9162 4870 9174 4922
rect 9226 4870 16982 4922
rect 17034 4870 17046 4922
rect 17098 4870 17110 4922
rect 17162 4870 17174 4922
rect 17226 4870 22816 4922
rect 1104 4848 22816 4870
rect 9858 4768 9864 4820
rect 9916 4808 9922 4820
rect 9953 4811 10011 4817
rect 9953 4808 9965 4811
rect 9916 4780 9965 4808
rect 9916 4768 9922 4780
rect 9953 4777 9965 4780
rect 9999 4808 10011 4811
rect 10686 4808 10692 4820
rect 9999 4780 10692 4808
rect 9999 4777 10011 4780
rect 9953 4771 10011 4777
rect 10686 4768 10692 4780
rect 10744 4768 10750 4820
rect 10781 4811 10839 4817
rect 10781 4777 10793 4811
rect 10827 4808 10839 4811
rect 10870 4808 10876 4820
rect 10827 4780 10876 4808
rect 10827 4777 10839 4780
rect 10781 4771 10839 4777
rect 10870 4768 10876 4780
rect 10928 4768 10934 4820
rect 11514 4808 11520 4820
rect 11475 4780 11520 4808
rect 11514 4768 11520 4780
rect 11572 4768 11578 4820
rect 13446 4808 13452 4820
rect 13407 4780 13452 4808
rect 13446 4768 13452 4780
rect 13504 4808 13510 4820
rect 13630 4808 13636 4820
rect 13504 4780 13636 4808
rect 13504 4768 13510 4780
rect 13630 4768 13636 4780
rect 13688 4768 13694 4820
rect 13909 4811 13967 4817
rect 13909 4808 13921 4811
rect 13786 4780 13921 4808
rect 11532 4740 11560 4768
rect 11532 4712 12480 4740
rect 1210 4632 1216 4684
rect 1268 4672 1274 4684
rect 9674 4672 9680 4684
rect 1268 4644 9680 4672
rect 1268 4632 1274 4644
rect 9674 4632 9680 4644
rect 9732 4672 9738 4684
rect 9769 4675 9827 4681
rect 9769 4672 9781 4675
rect 9732 4644 9781 4672
rect 9732 4632 9738 4644
rect 9769 4641 9781 4644
rect 9815 4641 9827 4675
rect 11606 4672 11612 4684
rect 11567 4644 11612 4672
rect 9769 4635 9827 4641
rect 11606 4632 11612 4644
rect 11664 4632 11670 4684
rect 12066 4672 12072 4684
rect 11979 4644 12072 4672
rect 12066 4632 12072 4644
rect 12124 4632 12130 4684
rect 12452 4681 12480 4712
rect 12437 4675 12495 4681
rect 12437 4641 12449 4675
rect 12483 4641 12495 4675
rect 12437 4635 12495 4641
rect 10410 4564 10416 4616
rect 10468 4604 10474 4616
rect 11882 4604 11888 4616
rect 10468 4576 11888 4604
rect 10468 4564 10474 4576
rect 11882 4564 11888 4576
rect 11940 4604 11946 4616
rect 12084 4604 12112 4632
rect 11940 4576 12112 4604
rect 12452 4604 12480 4635
rect 12526 4632 12532 4684
rect 12584 4672 12590 4684
rect 12989 4675 13047 4681
rect 12989 4672 13001 4675
rect 12584 4644 13001 4672
rect 12584 4632 12590 4644
rect 12989 4641 13001 4644
rect 13035 4672 13047 4675
rect 13786 4672 13814 4780
rect 13909 4777 13921 4780
rect 13955 4808 13967 4811
rect 14550 4808 14556 4820
rect 13955 4780 14556 4808
rect 13955 4777 13967 4780
rect 13909 4771 13967 4777
rect 14550 4768 14556 4780
rect 14608 4768 14614 4820
rect 15654 4808 15660 4820
rect 15615 4780 15660 4808
rect 15654 4768 15660 4780
rect 15712 4768 15718 4820
rect 17034 4740 17040 4752
rect 16947 4712 17040 4740
rect 17034 4700 17040 4712
rect 17092 4740 17098 4752
rect 18417 4743 18475 4749
rect 18417 4740 18429 4743
rect 17092 4712 18429 4740
rect 17092 4700 17098 4712
rect 18417 4709 18429 4712
rect 18463 4709 18475 4743
rect 18417 4703 18475 4709
rect 18506 4672 18512 4684
rect 13035 4644 13814 4672
rect 18467 4644 18512 4672
rect 13035 4641 13047 4644
rect 12989 4635 13047 4641
rect 18506 4632 18512 4644
rect 18564 4632 18570 4684
rect 12452 4576 13124 4604
rect 11940 4564 11946 4576
rect 12710 4496 12716 4548
rect 12768 4536 12774 4548
rect 12989 4539 13047 4545
rect 12989 4536 13001 4539
rect 12768 4508 13001 4536
rect 12768 4496 12774 4508
rect 12989 4505 13001 4508
rect 13035 4505 13047 4539
rect 13096 4536 13124 4576
rect 13354 4564 13360 4616
rect 13412 4604 13418 4616
rect 14185 4607 14243 4613
rect 14185 4604 14197 4607
rect 13412 4576 14197 4604
rect 13412 4564 13418 4576
rect 14185 4573 14197 4576
rect 14231 4573 14243 4607
rect 14185 4567 14243 4573
rect 16945 4607 17003 4613
rect 16945 4573 16957 4607
rect 16991 4573 17003 4607
rect 17402 4604 17408 4616
rect 17363 4576 17408 4604
rect 16945 4567 17003 4573
rect 14274 4536 14280 4548
rect 13096 4508 14280 4536
rect 12989 4499 13047 4505
rect 14274 4496 14280 4508
rect 14332 4496 14338 4548
rect 16850 4496 16856 4548
rect 16908 4536 16914 4548
rect 16960 4536 16988 4567
rect 17402 4564 17408 4576
rect 17460 4564 17466 4616
rect 16908 4508 16988 4536
rect 16908 4496 16914 4508
rect 1104 4378 22816 4400
rect 1104 4326 4982 4378
rect 5034 4326 5046 4378
rect 5098 4326 5110 4378
rect 5162 4326 5174 4378
rect 5226 4326 12982 4378
rect 13034 4326 13046 4378
rect 13098 4326 13110 4378
rect 13162 4326 13174 4378
rect 13226 4326 20982 4378
rect 21034 4326 21046 4378
rect 21098 4326 21110 4378
rect 21162 4326 21174 4378
rect 21226 4326 22816 4378
rect 1104 4304 22816 4326
rect 9674 4264 9680 4276
rect 9635 4236 9680 4264
rect 9674 4224 9680 4236
rect 9732 4224 9738 4276
rect 10689 4267 10747 4273
rect 10689 4233 10701 4267
rect 10735 4264 10747 4267
rect 10870 4264 10876 4276
rect 10735 4236 10876 4264
rect 10735 4233 10747 4236
rect 10689 4227 10747 4233
rect 10870 4224 10876 4236
rect 10928 4224 10934 4276
rect 11882 4264 11888 4276
rect 11843 4236 11888 4264
rect 11882 4224 11888 4236
rect 11940 4224 11946 4276
rect 12253 4267 12311 4273
rect 12253 4233 12265 4267
rect 12299 4264 12311 4267
rect 12526 4264 12532 4276
rect 12299 4236 12532 4264
rect 12299 4233 12311 4236
rect 12253 4227 12311 4233
rect 12526 4224 12532 4236
rect 12584 4224 12590 4276
rect 18506 4264 18512 4276
rect 18467 4236 18512 4264
rect 18506 4224 18512 4236
rect 18564 4224 18570 4276
rect 9582 4156 9588 4208
rect 9640 4196 9646 4208
rect 9766 4196 9772 4208
rect 9640 4168 9772 4196
rect 9640 4156 9646 4168
rect 9766 4156 9772 4168
rect 9824 4156 9830 4208
rect 16850 4156 16856 4208
rect 16908 4196 16914 4208
rect 17221 4199 17279 4205
rect 17221 4196 17233 4199
rect 16908 4168 17233 4196
rect 16908 4156 16914 4168
rect 17221 4165 17233 4168
rect 17267 4165 17279 4199
rect 17221 4159 17279 4165
rect 11514 4128 11520 4140
rect 11475 4100 11520 4128
rect 11514 4088 11520 4100
rect 11572 4128 11578 4140
rect 12897 4131 12955 4137
rect 12897 4128 12909 4131
rect 11572 4100 12909 4128
rect 11572 4088 11578 4100
rect 12897 4097 12909 4100
rect 12943 4097 12955 4131
rect 13262 4128 13268 4140
rect 13223 4100 13268 4128
rect 12897 4091 12955 4097
rect 10962 4060 10968 4072
rect 10923 4032 10968 4060
rect 10962 4020 10968 4032
rect 11020 4020 11026 4072
rect 12912 4060 12940 4091
rect 13262 4088 13268 4100
rect 13320 4088 13326 4140
rect 16945 4131 17003 4137
rect 16945 4097 16957 4131
rect 16991 4128 17003 4131
rect 17034 4128 17040 4140
rect 16991 4100 17040 4128
rect 16991 4097 17003 4100
rect 16945 4091 17003 4097
rect 17034 4088 17040 4100
rect 17092 4088 17098 4140
rect 13354 4060 13360 4072
rect 12912 4032 13360 4060
rect 13354 4020 13360 4032
rect 13412 4060 13418 4072
rect 13449 4063 13507 4069
rect 13449 4060 13461 4063
rect 13412 4032 13461 4060
rect 13412 4020 13418 4032
rect 13449 4029 13461 4032
rect 13495 4029 13507 4063
rect 13449 4023 13507 4029
rect 13630 4020 13636 4072
rect 13688 4060 13694 4072
rect 13909 4063 13967 4069
rect 13909 4060 13921 4063
rect 13688 4032 13921 4060
rect 13688 4020 13694 4032
rect 13909 4029 13921 4032
rect 13955 4029 13967 4063
rect 14274 4060 14280 4072
rect 14235 4032 14280 4060
rect 13909 4023 13967 4029
rect 14274 4020 14280 4032
rect 14332 4020 14338 4072
rect 14645 4063 14703 4069
rect 14645 4060 14657 4063
rect 14384 4032 14657 4060
rect 12434 3924 12440 3936
rect 12395 3896 12440 3924
rect 12434 3884 12440 3896
rect 12492 3884 12498 3936
rect 13262 3884 13268 3936
rect 13320 3924 13326 3936
rect 14384 3924 14412 4032
rect 14645 4029 14657 4032
rect 14691 4029 14703 4063
rect 14645 4023 14703 4029
rect 15657 4063 15715 4069
rect 15657 4029 15669 4063
rect 15703 4060 15715 4063
rect 15841 4063 15899 4069
rect 15841 4060 15853 4063
rect 15703 4032 15853 4060
rect 15703 4029 15715 4032
rect 15657 4023 15715 4029
rect 15841 4029 15853 4032
rect 15887 4060 15899 4063
rect 16206 4060 16212 4072
rect 15887 4032 16212 4060
rect 15887 4029 15899 4032
rect 15841 4023 15899 4029
rect 16206 4020 16212 4032
rect 16264 4020 16270 4072
rect 17402 4020 17408 4072
rect 17460 4060 17466 4072
rect 18084 4063 18142 4069
rect 18084 4060 18096 4063
rect 17460 4032 18096 4060
rect 17460 4020 17466 4032
rect 18084 4029 18096 4032
rect 18130 4060 18142 4063
rect 18877 4063 18935 4069
rect 18877 4060 18889 4063
rect 18130 4032 18889 4060
rect 18130 4029 18142 4032
rect 18084 4023 18142 4029
rect 18877 4029 18889 4032
rect 18923 4029 18935 4063
rect 18877 4023 18935 4029
rect 14918 3992 14924 4004
rect 14879 3964 14924 3992
rect 14918 3952 14924 3964
rect 14976 3952 14982 4004
rect 16482 3992 16488 4004
rect 16443 3964 16488 3992
rect 16482 3952 16488 3964
rect 16540 3952 16546 4004
rect 18187 3995 18245 4001
rect 18187 3961 18199 3995
rect 18233 3992 18245 3995
rect 23566 3992 23572 4004
rect 18233 3964 23572 3992
rect 18233 3961 18245 3964
rect 18187 3955 18245 3961
rect 23566 3952 23572 3964
rect 23624 3952 23630 4004
rect 13320 3896 14412 3924
rect 13320 3884 13326 3896
rect 1104 3834 22816 3856
rect 1104 3782 8982 3834
rect 9034 3782 9046 3834
rect 9098 3782 9110 3834
rect 9162 3782 9174 3834
rect 9226 3782 16982 3834
rect 17034 3782 17046 3834
rect 17098 3782 17110 3834
rect 17162 3782 17174 3834
rect 17226 3782 22816 3834
rect 1104 3760 22816 3782
rect 11514 3680 11520 3732
rect 11572 3720 11578 3732
rect 12253 3723 12311 3729
rect 12253 3720 12265 3723
rect 11572 3692 12265 3720
rect 11572 3680 11578 3692
rect 12253 3689 12265 3692
rect 12299 3689 12311 3723
rect 12710 3720 12716 3732
rect 12671 3692 12716 3720
rect 12253 3683 12311 3689
rect 12710 3680 12716 3692
rect 12768 3680 12774 3732
rect 14274 3720 14280 3732
rect 14235 3692 14280 3720
rect 14274 3680 14280 3692
rect 14332 3680 14338 3732
rect 16206 3720 16212 3732
rect 16167 3692 16212 3720
rect 16206 3680 16212 3692
rect 16264 3680 16270 3732
rect 16850 3680 16856 3732
rect 16908 3720 16914 3732
rect 17129 3723 17187 3729
rect 17129 3720 17141 3723
rect 16908 3692 17141 3720
rect 16908 3680 16914 3692
rect 17129 3689 17141 3692
rect 17175 3689 17187 3723
rect 17129 3683 17187 3689
rect 11974 3652 11980 3664
rect 11935 3624 11980 3652
rect 11974 3612 11980 3624
rect 12032 3612 12038 3664
rect 13446 3652 13452 3664
rect 13407 3624 13452 3652
rect 13446 3612 13452 3624
rect 13504 3612 13510 3664
rect 15194 3612 15200 3664
rect 15252 3652 15258 3664
rect 15610 3655 15668 3661
rect 15610 3652 15622 3655
rect 15252 3624 15622 3652
rect 15252 3612 15258 3624
rect 15610 3621 15622 3624
rect 15656 3621 15668 3655
rect 15610 3615 15668 3621
rect 10686 3544 10692 3596
rect 10744 3584 10750 3596
rect 11425 3587 11483 3593
rect 11425 3584 11437 3587
rect 10744 3556 11437 3584
rect 10744 3544 10750 3556
rect 11425 3553 11437 3556
rect 11471 3553 11483 3587
rect 11425 3547 11483 3553
rect 11609 3587 11667 3593
rect 11609 3553 11621 3587
rect 11655 3584 11667 3587
rect 11790 3584 11796 3596
rect 11655 3556 11796 3584
rect 11655 3553 11667 3556
rect 11609 3547 11667 3553
rect 11790 3544 11796 3556
rect 11848 3544 11854 3596
rect 13357 3519 13415 3525
rect 13357 3485 13369 3519
rect 13403 3516 13415 3519
rect 13998 3516 14004 3528
rect 13403 3488 14004 3516
rect 13403 3485 13415 3488
rect 13357 3479 13415 3485
rect 13998 3476 14004 3488
rect 14056 3476 14062 3528
rect 14918 3476 14924 3528
rect 14976 3516 14982 3528
rect 15289 3519 15347 3525
rect 15289 3516 15301 3519
rect 14976 3488 15301 3516
rect 14976 3476 14982 3488
rect 15289 3485 15301 3488
rect 15335 3516 15347 3519
rect 16758 3516 16764 3528
rect 15335 3488 16764 3516
rect 15335 3485 15347 3488
rect 15289 3479 15347 3485
rect 16758 3476 16764 3488
rect 16816 3476 16822 3528
rect 13722 3408 13728 3460
rect 13780 3448 13786 3460
rect 13909 3451 13967 3457
rect 13909 3448 13921 3451
rect 13780 3420 13921 3448
rect 13780 3408 13786 3420
rect 13909 3417 13921 3420
rect 13955 3417 13967 3451
rect 13909 3411 13967 3417
rect 1104 3290 22816 3312
rect 1104 3238 4982 3290
rect 5034 3238 5046 3290
rect 5098 3238 5110 3290
rect 5162 3238 5174 3290
rect 5226 3238 12982 3290
rect 13034 3238 13046 3290
rect 13098 3238 13110 3290
rect 13162 3238 13174 3290
rect 13226 3238 20982 3290
rect 21034 3238 21046 3290
rect 21098 3238 21110 3290
rect 21162 3238 21174 3290
rect 21226 3238 22816 3290
rect 1104 3216 22816 3238
rect 10686 3176 10692 3188
rect 10647 3148 10692 3176
rect 10686 3136 10692 3148
rect 10744 3136 10750 3188
rect 13998 3176 14004 3188
rect 13959 3148 14004 3176
rect 13998 3136 14004 3148
rect 14056 3136 14062 3188
rect 16482 3176 16488 3188
rect 16443 3148 16488 3176
rect 16482 3136 16488 3148
rect 16540 3136 16546 3188
rect 16758 3176 16764 3188
rect 16719 3148 16764 3176
rect 16758 3136 16764 3148
rect 16816 3136 16822 3188
rect 10134 3068 10140 3120
rect 10192 3108 10198 3120
rect 10965 3111 11023 3117
rect 10965 3108 10977 3111
rect 10192 3080 10977 3108
rect 10192 3068 10198 3080
rect 10965 3077 10977 3080
rect 11011 3077 11023 3111
rect 14016 3108 14044 3136
rect 15838 3108 15844 3120
rect 14016 3080 15844 3108
rect 10965 3071 11023 3077
rect 10980 2972 11008 3071
rect 15838 3068 15844 3080
rect 15896 3108 15902 3120
rect 16025 3111 16083 3117
rect 16025 3108 16037 3111
rect 15896 3080 16037 3108
rect 15896 3068 15902 3080
rect 16025 3077 16037 3080
rect 16071 3077 16083 3111
rect 16025 3071 16083 3077
rect 12437 3043 12495 3049
rect 12437 3009 12449 3043
rect 12483 3040 12495 3043
rect 12710 3040 12716 3052
rect 12483 3012 12716 3040
rect 12483 3009 12495 3012
rect 12437 3003 12495 3009
rect 12710 3000 12716 3012
rect 12768 3000 12774 3052
rect 15473 3043 15531 3049
rect 15473 3009 15485 3043
rect 15519 3040 15531 3043
rect 16850 3040 16856 3052
rect 15519 3012 16856 3040
rect 15519 3009 15531 3012
rect 15473 3003 15531 3009
rect 16850 3000 16856 3012
rect 16908 3040 16914 3052
rect 17129 3043 17187 3049
rect 17129 3040 17141 3043
rect 16908 3012 17141 3040
rect 16908 3000 16914 3012
rect 17129 3009 17141 3012
rect 17175 3009 17187 3043
rect 17129 3003 17187 3009
rect 11149 2975 11207 2981
rect 11149 2972 11161 2975
rect 10980 2944 11161 2972
rect 11149 2941 11161 2944
rect 11195 2941 11207 2975
rect 11149 2935 11207 2941
rect 13538 2932 13544 2984
rect 13596 2972 13602 2984
rect 14185 2975 14243 2981
rect 14185 2972 14197 2975
rect 13596 2944 14197 2972
rect 13596 2932 13602 2944
rect 14185 2941 14197 2944
rect 14231 2972 14243 2975
rect 14737 2975 14795 2981
rect 14737 2972 14749 2975
rect 14231 2944 14749 2972
rect 14231 2941 14243 2944
rect 14185 2935 14243 2941
rect 14737 2941 14749 2944
rect 14783 2941 14795 2975
rect 14737 2935 14795 2941
rect 12253 2907 12311 2913
rect 12253 2873 12265 2907
rect 12299 2904 12311 2907
rect 12758 2907 12816 2913
rect 12758 2904 12770 2907
rect 12299 2876 12770 2904
rect 12299 2873 12311 2876
rect 12253 2867 12311 2873
rect 12758 2873 12770 2876
rect 12804 2904 12816 2907
rect 15194 2904 15200 2916
rect 12804 2876 15200 2904
rect 12804 2873 12816 2876
rect 12758 2867 12816 2873
rect 15194 2864 15200 2876
rect 15252 2864 15258 2916
rect 15565 2907 15623 2913
rect 15565 2873 15577 2907
rect 15611 2873 15623 2907
rect 15565 2867 15623 2873
rect 11333 2839 11391 2845
rect 11333 2805 11345 2839
rect 11379 2836 11391 2839
rect 11606 2836 11612 2848
rect 11379 2808 11612 2836
rect 11379 2805 11391 2808
rect 11333 2799 11391 2805
rect 11606 2796 11612 2808
rect 11664 2796 11670 2848
rect 11790 2836 11796 2848
rect 11751 2808 11796 2836
rect 11790 2796 11796 2808
rect 11848 2796 11854 2848
rect 12526 2796 12532 2848
rect 12584 2836 12590 2848
rect 13357 2839 13415 2845
rect 13357 2836 13369 2839
rect 12584 2808 13369 2836
rect 12584 2796 12590 2808
rect 13357 2805 13369 2808
rect 13403 2836 13415 2839
rect 13446 2836 13452 2848
rect 13403 2808 13452 2836
rect 13403 2805 13415 2808
rect 13357 2799 13415 2805
rect 13446 2796 13452 2808
rect 13504 2836 13510 2848
rect 13633 2839 13691 2845
rect 13633 2836 13645 2839
rect 13504 2808 13645 2836
rect 13504 2796 13510 2808
rect 13633 2805 13645 2808
rect 13679 2805 13691 2839
rect 13633 2799 13691 2805
rect 14090 2796 14096 2848
rect 14148 2836 14154 2848
rect 14369 2839 14427 2845
rect 14369 2836 14381 2839
rect 14148 2808 14381 2836
rect 14148 2796 14154 2808
rect 14369 2805 14381 2808
rect 14415 2805 14427 2839
rect 15580 2836 15608 2867
rect 16482 2836 16488 2848
rect 15580 2808 16488 2836
rect 14369 2799 14427 2805
rect 16482 2796 16488 2808
rect 16540 2796 16546 2848
rect 1104 2746 22816 2768
rect 1104 2694 8982 2746
rect 9034 2694 9046 2746
rect 9098 2694 9110 2746
rect 9162 2694 9174 2746
rect 9226 2694 16982 2746
rect 17034 2694 17046 2746
rect 17098 2694 17110 2746
rect 17162 2694 17174 2746
rect 17226 2694 22816 2746
rect 1104 2672 22816 2694
rect 12434 2632 12440 2644
rect 12395 2604 12440 2632
rect 12434 2592 12440 2604
rect 12492 2592 12498 2644
rect 15289 2635 15347 2641
rect 12544 2604 13768 2632
rect 7469 2567 7527 2573
rect 7469 2564 7481 2567
rect 6999 2536 7481 2564
rect 6999 2505 7027 2536
rect 7469 2533 7481 2536
rect 7515 2564 7527 2567
rect 12544 2564 12572 2604
rect 13740 2576 13768 2604
rect 15289 2601 15301 2635
rect 15335 2632 15347 2635
rect 15335 2604 15700 2632
rect 15335 2601 15347 2604
rect 15289 2595 15347 2601
rect 13173 2567 13231 2573
rect 13173 2564 13185 2567
rect 7515 2536 12572 2564
rect 12820 2536 13185 2564
rect 7515 2533 7527 2536
rect 7469 2527 7527 2533
rect 6984 2499 7042 2505
rect 6984 2465 6996 2499
rect 7030 2465 7042 2499
rect 9766 2496 9772 2508
rect 9727 2468 9772 2496
rect 6984 2459 7042 2465
rect 9766 2456 9772 2468
rect 9824 2496 9830 2508
rect 10321 2499 10379 2505
rect 10321 2496 10333 2499
rect 9824 2468 10333 2496
rect 9824 2456 9830 2468
rect 10321 2465 10333 2468
rect 10367 2465 10379 2499
rect 10321 2459 10379 2465
rect 10873 2499 10931 2505
rect 10873 2465 10885 2499
rect 10919 2496 10931 2499
rect 11057 2499 11115 2505
rect 11057 2496 11069 2499
rect 10919 2468 11069 2496
rect 10919 2465 10931 2468
rect 10873 2459 10931 2465
rect 11057 2465 11069 2468
rect 11103 2496 11115 2499
rect 12526 2496 12532 2508
rect 11103 2468 12532 2496
rect 11103 2465 11115 2468
rect 11057 2459 11115 2465
rect 12526 2456 12532 2468
rect 12584 2456 12590 2508
rect 12820 2437 12848 2536
rect 13173 2533 13185 2536
rect 13219 2533 13231 2567
rect 13722 2564 13728 2576
rect 13683 2536 13728 2564
rect 13173 2527 13231 2533
rect 13722 2524 13728 2536
rect 13780 2524 13786 2576
rect 14921 2567 14979 2573
rect 14921 2533 14933 2567
rect 14967 2564 14979 2567
rect 15562 2564 15568 2576
rect 14967 2536 15568 2564
rect 14967 2533 14979 2536
rect 14921 2527 14979 2533
rect 15562 2524 15568 2536
rect 15620 2524 15626 2576
rect 15672 2573 15700 2604
rect 16850 2592 16856 2644
rect 16908 2632 16914 2644
rect 17175 2635 17233 2641
rect 17175 2632 17187 2635
rect 16908 2604 17187 2632
rect 16908 2592 16914 2604
rect 17175 2601 17187 2604
rect 17221 2601 17233 2635
rect 17175 2595 17233 2601
rect 15657 2567 15715 2573
rect 15657 2533 15669 2567
rect 15703 2564 15715 2567
rect 16206 2564 16212 2576
rect 15703 2536 16212 2564
rect 15703 2533 15715 2536
rect 15657 2527 15715 2533
rect 16206 2524 16212 2536
rect 16264 2524 16270 2576
rect 17072 2499 17130 2505
rect 17072 2465 17084 2499
rect 17118 2465 17130 2499
rect 17072 2459 17130 2465
rect 11701 2431 11759 2437
rect 11701 2397 11713 2431
rect 11747 2428 11759 2431
rect 12805 2431 12863 2437
rect 12805 2428 12817 2431
rect 11747 2400 12817 2428
rect 11747 2397 11759 2400
rect 11701 2391 11759 2397
rect 12805 2397 12817 2400
rect 12851 2397 12863 2431
rect 12805 2391 12863 2397
rect 13081 2431 13139 2437
rect 13081 2397 13093 2431
rect 13127 2397 13139 2431
rect 15838 2428 15844 2440
rect 15799 2400 15844 2428
rect 13081 2391 13139 2397
rect 12434 2320 12440 2372
rect 12492 2360 12498 2372
rect 13096 2360 13124 2391
rect 15838 2388 15844 2400
rect 15896 2388 15902 2440
rect 15930 2388 15936 2440
rect 15988 2428 15994 2440
rect 17087 2428 17115 2459
rect 17954 2456 17960 2508
rect 18012 2496 18018 2508
rect 18325 2499 18383 2505
rect 18325 2496 18337 2499
rect 18012 2468 18337 2496
rect 18012 2456 18018 2468
rect 18325 2465 18337 2468
rect 18371 2496 18383 2499
rect 18877 2499 18935 2505
rect 18877 2496 18889 2499
rect 18371 2468 18889 2496
rect 18371 2465 18383 2468
rect 18325 2459 18383 2465
rect 18877 2465 18889 2468
rect 18923 2465 18935 2499
rect 18877 2459 18935 2465
rect 19886 2456 19892 2508
rect 19944 2496 19950 2508
rect 21177 2499 21235 2505
rect 21177 2496 21189 2499
rect 19944 2468 21189 2496
rect 19944 2456 19950 2468
rect 21177 2465 21189 2468
rect 21223 2496 21235 2499
rect 21729 2499 21787 2505
rect 21729 2496 21741 2499
rect 21223 2468 21741 2496
rect 21223 2465 21235 2468
rect 21177 2459 21235 2465
rect 21729 2465 21741 2468
rect 21775 2465 21787 2499
rect 21729 2459 21787 2465
rect 17497 2431 17555 2437
rect 17497 2428 17509 2431
rect 15988 2400 17509 2428
rect 15988 2388 15994 2400
rect 17497 2397 17509 2400
rect 17543 2397 17555 2431
rect 17497 2391 17555 2397
rect 12492 2332 13124 2360
rect 18509 2363 18567 2369
rect 12492 2320 12498 2332
rect 18509 2329 18521 2363
rect 18555 2360 18567 2363
rect 19426 2360 19432 2372
rect 18555 2332 19432 2360
rect 18555 2329 18567 2332
rect 18509 2323 18567 2329
rect 19426 2320 19432 2332
rect 19484 2320 19490 2372
rect 21361 2363 21419 2369
rect 21361 2329 21373 2363
rect 21407 2360 21419 2363
rect 23106 2360 23112 2372
rect 21407 2332 23112 2360
rect 21407 2329 21419 2332
rect 21361 2323 21419 2329
rect 23106 2320 23112 2332
rect 23164 2320 23170 2372
rect 6730 2252 6736 2304
rect 6788 2292 6794 2304
rect 7055 2295 7113 2301
rect 7055 2292 7067 2295
rect 6788 2264 7067 2292
rect 6788 2252 6794 2264
rect 7055 2261 7067 2264
rect 7101 2261 7113 2295
rect 7055 2255 7113 2261
rect 9953 2295 10011 2301
rect 9953 2261 9965 2295
rect 9999 2292 10011 2295
rect 10226 2292 10232 2304
rect 9999 2264 10232 2292
rect 9999 2261 10011 2264
rect 9953 2255 10011 2261
rect 10226 2252 10232 2264
rect 10284 2252 10290 2304
rect 1104 2202 22816 2224
rect 1104 2150 4982 2202
rect 5034 2150 5046 2202
rect 5098 2150 5110 2202
rect 5162 2150 5174 2202
rect 5226 2150 12982 2202
rect 13034 2150 13046 2202
rect 13098 2150 13110 2202
rect 13162 2150 13174 2202
rect 13226 2150 20982 2202
rect 21034 2150 21046 2202
rect 21098 2150 21110 2202
rect 21162 2150 21174 2202
rect 21226 2150 22816 2202
rect 1104 2128 22816 2150
<< via1 >>
rect 13912 23536 13964 23588
rect 14924 23536 14976 23588
rect 4982 21734 5034 21786
rect 5046 21734 5098 21786
rect 5110 21734 5162 21786
rect 5174 21734 5226 21786
rect 12982 21734 13034 21786
rect 13046 21734 13098 21786
rect 13110 21734 13162 21786
rect 13174 21734 13226 21786
rect 20982 21734 21034 21786
rect 21046 21734 21098 21786
rect 21110 21734 21162 21786
rect 21174 21734 21226 21786
rect 8982 21190 9034 21242
rect 9046 21190 9098 21242
rect 9110 21190 9162 21242
rect 9174 21190 9226 21242
rect 16982 21190 17034 21242
rect 17046 21190 17098 21242
rect 17110 21190 17162 21242
rect 17174 21190 17226 21242
rect 4982 20646 5034 20698
rect 5046 20646 5098 20698
rect 5110 20646 5162 20698
rect 5174 20646 5226 20698
rect 12982 20646 13034 20698
rect 13046 20646 13098 20698
rect 13110 20646 13162 20698
rect 13174 20646 13226 20698
rect 20982 20646 21034 20698
rect 21046 20646 21098 20698
rect 21110 20646 21162 20698
rect 21174 20646 21226 20698
rect 8852 20587 8904 20596
rect 8852 20553 8861 20587
rect 8861 20553 8895 20587
rect 8895 20553 8904 20587
rect 8852 20544 8904 20553
rect 20628 20544 20680 20596
rect 22652 20544 22704 20596
rect 15844 20340 15896 20392
rect 20812 20340 20864 20392
rect 10784 20204 10836 20256
rect 8982 20102 9034 20154
rect 9046 20102 9098 20154
rect 9110 20102 9162 20154
rect 9174 20102 9226 20154
rect 16982 20102 17034 20154
rect 17046 20102 17098 20154
rect 17110 20102 17162 20154
rect 17174 20102 17226 20154
rect 4982 19558 5034 19610
rect 5046 19558 5098 19610
rect 5110 19558 5162 19610
rect 5174 19558 5226 19610
rect 12982 19558 13034 19610
rect 13046 19558 13098 19610
rect 13110 19558 13162 19610
rect 13174 19558 13226 19610
rect 20982 19558 21034 19610
rect 21046 19558 21098 19610
rect 21110 19558 21162 19610
rect 21174 19558 21226 19610
rect 8982 19014 9034 19066
rect 9046 19014 9098 19066
rect 9110 19014 9162 19066
rect 9174 19014 9226 19066
rect 16982 19014 17034 19066
rect 17046 19014 17098 19066
rect 17110 19014 17162 19066
rect 17174 19014 17226 19066
rect 4982 18470 5034 18522
rect 5046 18470 5098 18522
rect 5110 18470 5162 18522
rect 5174 18470 5226 18522
rect 12982 18470 13034 18522
rect 13046 18470 13098 18522
rect 13110 18470 13162 18522
rect 13174 18470 13226 18522
rect 20982 18470 21034 18522
rect 21046 18470 21098 18522
rect 21110 18470 21162 18522
rect 21174 18470 21226 18522
rect 8982 17926 9034 17978
rect 9046 17926 9098 17978
rect 9110 17926 9162 17978
rect 9174 17926 9226 17978
rect 16982 17926 17034 17978
rect 17046 17926 17098 17978
rect 17110 17926 17162 17978
rect 17174 17926 17226 17978
rect 11152 17620 11204 17672
rect 14188 17620 14240 17672
rect 4982 17382 5034 17434
rect 5046 17382 5098 17434
rect 5110 17382 5162 17434
rect 5174 17382 5226 17434
rect 12982 17382 13034 17434
rect 13046 17382 13098 17434
rect 13110 17382 13162 17434
rect 13174 17382 13226 17434
rect 20982 17382 21034 17434
rect 21046 17382 21098 17434
rect 21110 17382 21162 17434
rect 21174 17382 21226 17434
rect 7012 17323 7064 17332
rect 7012 17289 7021 17323
rect 7021 17289 7055 17323
rect 7055 17289 7064 17323
rect 7012 17280 7064 17289
rect 5356 17144 5408 17196
rect 8392 17119 8444 17128
rect 8392 17085 8401 17119
rect 8401 17085 8435 17119
rect 8435 17085 8444 17119
rect 8392 17076 8444 17085
rect 7748 16940 7800 16992
rect 8208 16940 8260 16992
rect 8982 16838 9034 16890
rect 9046 16838 9098 16890
rect 9110 16838 9162 16890
rect 9174 16838 9226 16890
rect 16982 16838 17034 16890
rect 17046 16838 17098 16890
rect 17110 16838 17162 16890
rect 17174 16838 17226 16890
rect 8208 16779 8260 16788
rect 8208 16745 8217 16779
rect 8217 16745 8251 16779
rect 8251 16745 8260 16779
rect 8208 16736 8260 16745
rect 7748 16600 7800 16652
rect 10784 16600 10836 16652
rect 8116 16396 8168 16448
rect 10692 16396 10744 16448
rect 4982 16294 5034 16346
rect 5046 16294 5098 16346
rect 5110 16294 5162 16346
rect 5174 16294 5226 16346
rect 12982 16294 13034 16346
rect 13046 16294 13098 16346
rect 13110 16294 13162 16346
rect 13174 16294 13226 16346
rect 20982 16294 21034 16346
rect 21046 16294 21098 16346
rect 21110 16294 21162 16346
rect 21174 16294 21226 16346
rect 7748 16235 7800 16244
rect 7748 16201 7757 16235
rect 7757 16201 7791 16235
rect 7791 16201 7800 16235
rect 7748 16192 7800 16201
rect 8208 16056 8260 16108
rect 11428 16031 11480 16040
rect 11428 15997 11437 16031
rect 11437 15997 11471 16031
rect 11471 15997 11480 16031
rect 11428 15988 11480 15997
rect 8208 15920 8260 15972
rect 9588 15920 9640 15972
rect 10784 15963 10836 15972
rect 10784 15929 10793 15963
rect 10793 15929 10827 15963
rect 10827 15929 10836 15963
rect 10784 15920 10836 15929
rect 14832 15920 14884 15972
rect 16764 15920 16816 15972
rect 11336 15852 11388 15904
rect 11428 15852 11480 15904
rect 15844 15852 15896 15904
rect 8982 15750 9034 15802
rect 9046 15750 9098 15802
rect 9110 15750 9162 15802
rect 9174 15750 9226 15802
rect 16982 15750 17034 15802
rect 17046 15750 17098 15802
rect 17110 15750 17162 15802
rect 17174 15750 17226 15802
rect 112 15648 164 15700
rect 10692 15648 10744 15700
rect 8208 15623 8260 15632
rect 8208 15589 8217 15623
rect 8217 15589 8251 15623
rect 8251 15589 8260 15623
rect 8208 15580 8260 15589
rect 9772 15580 9824 15632
rect 11428 15623 11480 15632
rect 11428 15589 11437 15623
rect 11437 15589 11471 15623
rect 11471 15589 11480 15623
rect 11428 15580 11480 15589
rect 5356 15512 5408 15564
rect 13544 15512 13596 15564
rect 15844 15512 15896 15564
rect 8116 15487 8168 15496
rect 8116 15453 8125 15487
rect 8125 15453 8159 15487
rect 8159 15453 8168 15487
rect 8116 15444 8168 15453
rect 8852 15444 8904 15496
rect 9588 15444 9640 15496
rect 10048 15487 10100 15496
rect 10048 15453 10057 15487
rect 10057 15453 10091 15487
rect 10091 15453 10100 15487
rect 10048 15444 10100 15453
rect 11336 15487 11388 15496
rect 11336 15453 11345 15487
rect 11345 15453 11379 15487
rect 11379 15453 11388 15487
rect 11336 15444 11388 15453
rect 11796 15487 11848 15496
rect 11796 15453 11805 15487
rect 11805 15453 11839 15487
rect 11839 15453 11848 15487
rect 11796 15444 11848 15453
rect 16120 15376 16172 15428
rect 12532 15308 12584 15360
rect 16028 15351 16080 15360
rect 16028 15317 16037 15351
rect 16037 15317 16071 15351
rect 16071 15317 16080 15351
rect 16028 15308 16080 15317
rect 4982 15206 5034 15258
rect 5046 15206 5098 15258
rect 5110 15206 5162 15258
rect 5174 15206 5226 15258
rect 12982 15206 13034 15258
rect 13046 15206 13098 15258
rect 13110 15206 13162 15258
rect 13174 15206 13226 15258
rect 20982 15206 21034 15258
rect 21046 15206 21098 15258
rect 21110 15206 21162 15258
rect 21174 15206 21226 15258
rect 8208 15104 8260 15156
rect 9588 15104 9640 15156
rect 11428 15104 11480 15156
rect 14832 15147 14884 15156
rect 5356 14968 5408 15020
rect 6276 14968 6328 15020
rect 10048 14968 10100 15020
rect 10692 14968 10744 15020
rect 7012 14900 7064 14952
rect 8852 14875 8904 14884
rect 8852 14841 8861 14875
rect 8861 14841 8895 14875
rect 8895 14841 8904 14875
rect 8852 14832 8904 14841
rect 5632 14764 5684 14816
rect 6552 14807 6604 14816
rect 6552 14773 6561 14807
rect 6561 14773 6595 14807
rect 6595 14773 6604 14807
rect 6552 14764 6604 14773
rect 8760 14764 8812 14816
rect 11244 14832 11296 14884
rect 9772 14807 9824 14816
rect 9772 14773 9781 14807
rect 9781 14773 9815 14807
rect 9815 14773 9824 14807
rect 9772 14764 9824 14773
rect 14832 15113 14841 15147
rect 14841 15113 14875 15147
rect 14875 15113 14884 15147
rect 14832 15104 14884 15113
rect 15844 15104 15896 15156
rect 21272 15104 21324 15156
rect 21548 15147 21600 15156
rect 21548 15113 21557 15147
rect 21557 15113 21591 15147
rect 21591 15113 21600 15147
rect 21548 15104 21600 15113
rect 13544 15036 13596 15088
rect 18604 15036 18656 15088
rect 12532 15011 12584 15020
rect 12532 14977 12541 15011
rect 12541 14977 12575 15011
rect 12575 14977 12584 15011
rect 12532 14968 12584 14977
rect 16120 14968 16172 15020
rect 14832 14900 14884 14952
rect 20812 14900 20864 14952
rect 21548 14900 21600 14952
rect 16028 14832 16080 14884
rect 16672 14875 16724 14884
rect 16672 14841 16681 14875
rect 16681 14841 16715 14875
rect 16715 14841 16724 14875
rect 16672 14832 16724 14841
rect 13544 14807 13596 14816
rect 13544 14773 13553 14807
rect 13553 14773 13587 14807
rect 13587 14773 13596 14807
rect 13544 14764 13596 14773
rect 15200 14764 15252 14816
rect 8982 14662 9034 14714
rect 9046 14662 9098 14714
rect 9110 14662 9162 14714
rect 9174 14662 9226 14714
rect 16982 14662 17034 14714
rect 17046 14662 17098 14714
rect 17110 14662 17162 14714
rect 17174 14662 17226 14714
rect 7840 14603 7892 14612
rect 7840 14569 7849 14603
rect 7849 14569 7883 14603
rect 7883 14569 7892 14603
rect 7840 14560 7892 14569
rect 9772 14560 9824 14612
rect 11336 14560 11388 14612
rect 12532 14603 12584 14612
rect 12532 14569 12541 14603
rect 12541 14569 12575 14603
rect 12575 14569 12584 14603
rect 12532 14560 12584 14569
rect 5724 14535 5776 14544
rect 5724 14501 5733 14535
rect 5733 14501 5767 14535
rect 5767 14501 5776 14535
rect 5724 14492 5776 14501
rect 6276 14535 6328 14544
rect 6276 14501 6285 14535
rect 6285 14501 6319 14535
rect 6319 14501 6328 14535
rect 6276 14492 6328 14501
rect 8116 14492 8168 14544
rect 11244 14535 11296 14544
rect 11244 14501 11253 14535
rect 11253 14501 11287 14535
rect 11287 14501 11296 14535
rect 11244 14492 11296 14501
rect 11796 14535 11848 14544
rect 11796 14501 11805 14535
rect 11805 14501 11839 14535
rect 11839 14501 11848 14535
rect 11796 14492 11848 14501
rect 16120 14535 16172 14544
rect 16120 14501 16129 14535
rect 16129 14501 16163 14535
rect 16163 14501 16172 14535
rect 16120 14492 16172 14501
rect 16672 14535 16724 14544
rect 16672 14501 16681 14535
rect 16681 14501 16715 14535
rect 16715 14501 16724 14535
rect 16672 14492 16724 14501
rect 10048 14467 10100 14476
rect 10048 14433 10057 14467
rect 10057 14433 10091 14467
rect 10091 14433 10100 14467
rect 10048 14424 10100 14433
rect 5632 14399 5684 14408
rect 5632 14365 5641 14399
rect 5641 14365 5675 14399
rect 5675 14365 5684 14399
rect 5632 14356 5684 14365
rect 7104 14356 7156 14408
rect 12164 14356 12216 14408
rect 15200 14356 15252 14408
rect 8852 14288 8904 14340
rect 11796 14288 11848 14340
rect 7012 14220 7064 14272
rect 10600 14263 10652 14272
rect 10600 14229 10609 14263
rect 10609 14229 10643 14263
rect 10643 14229 10652 14263
rect 10600 14220 10652 14229
rect 4982 14118 5034 14170
rect 5046 14118 5098 14170
rect 5110 14118 5162 14170
rect 5174 14118 5226 14170
rect 12982 14118 13034 14170
rect 13046 14118 13098 14170
rect 13110 14118 13162 14170
rect 13174 14118 13226 14170
rect 20982 14118 21034 14170
rect 21046 14118 21098 14170
rect 21110 14118 21162 14170
rect 21174 14118 21226 14170
rect 1492 14016 1544 14068
rect 5724 14016 5776 14068
rect 8760 14016 8812 14068
rect 11428 14016 11480 14068
rect 12164 14059 12216 14068
rect 12164 14025 12173 14059
rect 12173 14025 12207 14059
rect 12207 14025 12216 14059
rect 12164 14016 12216 14025
rect 15200 14059 15252 14068
rect 15200 14025 15209 14059
rect 15209 14025 15243 14059
rect 15243 14025 15252 14059
rect 15200 14016 15252 14025
rect 18328 14059 18380 14068
rect 18328 14025 18337 14059
rect 18337 14025 18371 14059
rect 18371 14025 18380 14059
rect 18328 14016 18380 14025
rect 5632 13948 5684 14000
rect 11244 13948 11296 14000
rect 9404 13880 9456 13932
rect 10048 13923 10100 13932
rect 10048 13889 10057 13923
rect 10057 13889 10091 13923
rect 10091 13889 10100 13923
rect 10048 13880 10100 13889
rect 10600 13923 10652 13932
rect 10600 13889 10609 13923
rect 10609 13889 10643 13923
rect 10643 13889 10652 13923
rect 10600 13880 10652 13889
rect 16120 13880 16172 13932
rect 4988 13855 5040 13864
rect 4988 13821 4997 13855
rect 4997 13821 5031 13855
rect 5031 13821 5040 13855
rect 4988 13812 5040 13821
rect 8300 13855 8352 13864
rect 8300 13821 8309 13855
rect 8309 13821 8343 13855
rect 8343 13821 8352 13855
rect 8300 13812 8352 13821
rect 16028 13855 16080 13864
rect 16028 13821 16037 13855
rect 16037 13821 16071 13855
rect 16071 13821 16080 13855
rect 16028 13812 16080 13821
rect 17776 13812 17828 13864
rect 6644 13744 6696 13796
rect 7840 13744 7892 13796
rect 7104 13719 7156 13728
rect 7104 13685 7113 13719
rect 7113 13685 7147 13719
rect 7147 13685 7156 13719
rect 7104 13676 7156 13685
rect 10508 13719 10560 13728
rect 10508 13685 10517 13719
rect 10517 13685 10551 13719
rect 10551 13685 10560 13719
rect 10508 13676 10560 13685
rect 8982 13574 9034 13626
rect 9046 13574 9098 13626
rect 9110 13574 9162 13626
rect 9174 13574 9226 13626
rect 16982 13574 17034 13626
rect 17046 13574 17098 13626
rect 17110 13574 17162 13626
rect 17174 13574 17226 13626
rect 4988 13472 5040 13524
rect 11244 13472 11296 13524
rect 10508 13404 10560 13456
rect 11704 13404 11756 13456
rect 15844 13404 15896 13456
rect 17500 13404 17552 13456
rect 5816 13379 5868 13388
rect 5816 13345 5825 13379
rect 5825 13345 5859 13379
rect 5859 13345 5868 13379
rect 5816 13336 5868 13345
rect 6460 13379 6512 13388
rect 6460 13345 6469 13379
rect 6469 13345 6503 13379
rect 6503 13345 6512 13379
rect 6460 13336 6512 13345
rect 6920 13379 6972 13388
rect 6920 13345 6929 13379
rect 6929 13345 6963 13379
rect 6963 13345 6972 13379
rect 6920 13336 6972 13345
rect 10508 13311 10560 13320
rect 10508 13277 10517 13311
rect 10517 13277 10551 13311
rect 10551 13277 10560 13311
rect 10508 13268 10560 13277
rect 15292 13311 15344 13320
rect 15292 13277 15301 13311
rect 15301 13277 15335 13311
rect 15335 13277 15344 13311
rect 15292 13268 15344 13277
rect 17132 13311 17184 13320
rect 17132 13277 17141 13311
rect 17141 13277 17175 13311
rect 17175 13277 17184 13311
rect 17132 13268 17184 13277
rect 17776 13311 17828 13320
rect 17776 13277 17785 13311
rect 17785 13277 17819 13311
rect 17819 13277 17828 13311
rect 17776 13268 17828 13277
rect 6184 13132 6236 13184
rect 7380 13175 7432 13184
rect 7380 13141 7389 13175
rect 7389 13141 7423 13175
rect 7423 13141 7432 13175
rect 7380 13132 7432 13141
rect 8300 13175 8352 13184
rect 8300 13141 8309 13175
rect 8309 13141 8343 13175
rect 8343 13141 8352 13175
rect 8300 13132 8352 13141
rect 10140 13132 10192 13184
rect 13360 13175 13412 13184
rect 13360 13141 13369 13175
rect 13369 13141 13403 13175
rect 13403 13141 13412 13175
rect 13360 13132 13412 13141
rect 14556 13132 14608 13184
rect 4982 13030 5034 13082
rect 5046 13030 5098 13082
rect 5110 13030 5162 13082
rect 5174 13030 5226 13082
rect 12982 13030 13034 13082
rect 13046 13030 13098 13082
rect 13110 13030 13162 13082
rect 13174 13030 13226 13082
rect 20982 13030 21034 13082
rect 21046 13030 21098 13082
rect 21110 13030 21162 13082
rect 21174 13030 21226 13082
rect 6184 12928 6236 12980
rect 10048 12928 10100 12980
rect 16396 12971 16448 12980
rect 16396 12937 16405 12971
rect 16405 12937 16439 12971
rect 16439 12937 16448 12971
rect 16396 12928 16448 12937
rect 17132 12971 17184 12980
rect 17132 12937 17141 12971
rect 17141 12937 17175 12971
rect 17175 12937 17184 12971
rect 17132 12928 17184 12937
rect 5816 12724 5868 12776
rect 7380 12792 7432 12844
rect 13360 12860 13412 12912
rect 17500 12903 17552 12912
rect 17500 12869 17509 12903
rect 17509 12869 17543 12903
rect 17543 12869 17552 12903
rect 17500 12860 17552 12869
rect 10508 12792 10560 12844
rect 15292 12792 15344 12844
rect 8208 12767 8260 12776
rect 8208 12733 8217 12767
rect 8217 12733 8251 12767
rect 8251 12733 8260 12767
rect 8208 12724 8260 12733
rect 10048 12767 10100 12776
rect 10048 12733 10057 12767
rect 10057 12733 10091 12767
rect 10091 12733 10100 12767
rect 10048 12724 10100 12733
rect 10140 12724 10192 12776
rect 11336 12767 11388 12776
rect 9772 12699 9824 12708
rect 9772 12665 9781 12699
rect 9781 12665 9815 12699
rect 9815 12665 9824 12699
rect 11336 12733 11345 12767
rect 11345 12733 11379 12767
rect 11379 12733 11388 12767
rect 11336 12724 11388 12733
rect 13268 12724 13320 12776
rect 13452 12724 13504 12776
rect 9772 12656 9824 12665
rect 12808 12656 12860 12708
rect 13636 12656 13688 12708
rect 14556 12767 14608 12776
rect 14556 12733 14565 12767
rect 14565 12733 14599 12767
rect 14599 12733 14608 12767
rect 14556 12724 14608 12733
rect 15936 12724 15988 12776
rect 5356 12588 5408 12640
rect 6552 12631 6604 12640
rect 6552 12597 6561 12631
rect 6561 12597 6595 12631
rect 6595 12597 6604 12631
rect 6552 12588 6604 12597
rect 7104 12631 7156 12640
rect 7104 12597 7113 12631
rect 7113 12597 7147 12631
rect 7147 12597 7156 12631
rect 7104 12588 7156 12597
rect 9496 12631 9548 12640
rect 9496 12597 9505 12631
rect 9505 12597 9539 12631
rect 9539 12597 9548 12631
rect 9496 12588 9548 12597
rect 11704 12631 11756 12640
rect 11704 12597 11713 12631
rect 11713 12597 11747 12631
rect 11747 12597 11756 12631
rect 11704 12588 11756 12597
rect 13268 12631 13320 12640
rect 13268 12597 13277 12631
rect 13277 12597 13311 12631
rect 13311 12597 13320 12631
rect 13268 12588 13320 12597
rect 15844 12588 15896 12640
rect 8982 12486 9034 12538
rect 9046 12486 9098 12538
rect 9110 12486 9162 12538
rect 9174 12486 9226 12538
rect 16982 12486 17034 12538
rect 17046 12486 17098 12538
rect 17110 12486 17162 12538
rect 17174 12486 17226 12538
rect 7012 12427 7064 12436
rect 7012 12393 7021 12427
rect 7021 12393 7055 12427
rect 7055 12393 7064 12427
rect 7012 12384 7064 12393
rect 10600 12427 10652 12436
rect 10600 12393 10609 12427
rect 10609 12393 10643 12427
rect 10643 12393 10652 12427
rect 10600 12384 10652 12393
rect 12808 12427 12860 12436
rect 12808 12393 12817 12427
rect 12817 12393 12851 12427
rect 12851 12393 12860 12427
rect 12808 12384 12860 12393
rect 15844 12427 15896 12436
rect 15844 12393 15853 12427
rect 15853 12393 15887 12427
rect 15887 12393 15896 12427
rect 15844 12384 15896 12393
rect 17316 12384 17368 12436
rect 6920 12316 6972 12368
rect 5724 12248 5776 12300
rect 6276 12291 6328 12300
rect 6276 12257 6285 12291
rect 6285 12257 6319 12291
rect 6319 12257 6328 12291
rect 6276 12248 6328 12257
rect 6460 12248 6512 12300
rect 8208 12316 8260 12368
rect 9496 12359 9548 12368
rect 9496 12325 9505 12359
rect 9505 12325 9539 12359
rect 9539 12325 9548 12359
rect 9496 12316 9548 12325
rect 10324 12291 10376 12300
rect 10324 12257 10333 12291
rect 10333 12257 10367 12291
rect 10367 12257 10376 12291
rect 10324 12248 10376 12257
rect 10140 12180 10192 12232
rect 10600 12180 10652 12232
rect 11336 12248 11388 12300
rect 13360 12291 13412 12300
rect 13360 12257 13369 12291
rect 13369 12257 13403 12291
rect 13403 12257 13412 12291
rect 13360 12248 13412 12257
rect 13912 12291 13964 12300
rect 13912 12257 13921 12291
rect 13921 12257 13955 12291
rect 13955 12257 13964 12291
rect 13912 12248 13964 12257
rect 14280 12291 14332 12300
rect 14280 12257 14289 12291
rect 14289 12257 14323 12291
rect 14323 12257 14332 12291
rect 14280 12248 14332 12257
rect 14556 12248 14608 12300
rect 18880 12291 18932 12300
rect 18880 12257 18898 12291
rect 18898 12257 18932 12291
rect 18880 12248 18932 12257
rect 20812 12248 20864 12300
rect 13268 12180 13320 12232
rect 16764 12180 16816 12232
rect 17408 12180 17460 12232
rect 17776 12223 17828 12232
rect 17776 12189 17785 12223
rect 17785 12189 17819 12223
rect 17819 12189 17828 12223
rect 17776 12180 17828 12189
rect 8116 12087 8168 12096
rect 8116 12053 8125 12087
rect 8125 12053 8159 12087
rect 8159 12053 8168 12087
rect 8116 12044 8168 12053
rect 10048 12087 10100 12096
rect 10048 12053 10057 12087
rect 10057 12053 10091 12087
rect 10091 12053 10100 12087
rect 10048 12044 10100 12053
rect 12440 12087 12492 12096
rect 12440 12053 12449 12087
rect 12449 12053 12483 12087
rect 12483 12053 12492 12087
rect 12440 12044 12492 12053
rect 18696 12044 18748 12096
rect 4982 11942 5034 11994
rect 5046 11942 5098 11994
rect 5110 11942 5162 11994
rect 5174 11942 5226 11994
rect 12982 11942 13034 11994
rect 13046 11942 13098 11994
rect 13110 11942 13162 11994
rect 13174 11942 13226 11994
rect 20982 11942 21034 11994
rect 21046 11942 21098 11994
rect 21110 11942 21162 11994
rect 21174 11942 21226 11994
rect 1492 11840 1544 11892
rect 5356 11840 5408 11892
rect 6920 11840 6972 11892
rect 9772 11840 9824 11892
rect 10600 11840 10652 11892
rect 12808 11840 12860 11892
rect 13360 11840 13412 11892
rect 16764 11883 16816 11892
rect 16764 11849 16773 11883
rect 16773 11849 16807 11883
rect 16807 11849 16816 11883
rect 16764 11840 16816 11849
rect 17316 11883 17368 11892
rect 17316 11849 17325 11883
rect 17325 11849 17359 11883
rect 17359 11849 17368 11883
rect 17316 11840 17368 11849
rect 18880 11883 18932 11892
rect 18880 11849 18889 11883
rect 18889 11849 18923 11883
rect 18923 11849 18932 11883
rect 18880 11840 18932 11849
rect 8208 11772 8260 11824
rect 7840 11704 7892 11756
rect 112 11636 164 11688
rect 1952 11679 2004 11688
rect 1952 11645 1961 11679
rect 1961 11645 1995 11679
rect 1995 11645 2004 11679
rect 1952 11636 2004 11645
rect 6460 11636 6512 11688
rect 8208 11636 8260 11688
rect 9496 11704 9548 11756
rect 8116 11568 8168 11620
rect 9588 11636 9640 11688
rect 10048 11679 10100 11688
rect 10048 11645 10057 11679
rect 10057 11645 10091 11679
rect 10091 11645 10100 11679
rect 10048 11636 10100 11645
rect 11520 11679 11572 11688
rect 9496 11568 9548 11620
rect 11520 11645 11529 11679
rect 11529 11645 11563 11679
rect 11563 11645 11572 11679
rect 11520 11636 11572 11645
rect 13268 11636 13320 11688
rect 13084 11568 13136 11620
rect 5724 11500 5776 11552
rect 6276 11543 6328 11552
rect 6276 11509 6285 11543
rect 6285 11509 6319 11543
rect 6319 11509 6328 11543
rect 6276 11500 6328 11509
rect 7840 11543 7892 11552
rect 7840 11509 7849 11543
rect 7849 11509 7883 11543
rect 7883 11509 7892 11543
rect 7840 11500 7892 11509
rect 8300 11543 8352 11552
rect 8300 11509 8309 11543
rect 8309 11509 8343 11543
rect 8343 11509 8352 11543
rect 8300 11500 8352 11509
rect 10140 11500 10192 11552
rect 12348 11500 12400 11552
rect 13636 11636 13688 11688
rect 14280 11679 14332 11688
rect 14280 11645 14289 11679
rect 14289 11645 14323 11679
rect 14323 11645 14332 11679
rect 14280 11636 14332 11645
rect 15568 11679 15620 11688
rect 15568 11645 15577 11679
rect 15577 11645 15611 11679
rect 15611 11645 15620 11679
rect 15568 11636 15620 11645
rect 13728 11500 13780 11552
rect 15108 11543 15160 11552
rect 15108 11509 15117 11543
rect 15117 11509 15151 11543
rect 15151 11509 15160 11543
rect 15844 11568 15896 11620
rect 15108 11500 15160 11509
rect 16488 11543 16540 11552
rect 16488 11509 16497 11543
rect 16497 11509 16531 11543
rect 16531 11509 16540 11543
rect 16488 11500 16540 11509
rect 17408 11500 17460 11552
rect 18972 11500 19024 11552
rect 8982 11398 9034 11450
rect 9046 11398 9098 11450
rect 9110 11398 9162 11450
rect 9174 11398 9226 11450
rect 16982 11398 17034 11450
rect 17046 11398 17098 11450
rect 17110 11398 17162 11450
rect 17174 11398 17226 11450
rect 5540 11339 5592 11348
rect 5540 11305 5549 11339
rect 5549 11305 5583 11339
rect 5583 11305 5592 11339
rect 5540 11296 5592 11305
rect 10048 11339 10100 11348
rect 10048 11305 10057 11339
rect 10057 11305 10091 11339
rect 10091 11305 10100 11339
rect 10048 11296 10100 11305
rect 15476 11339 15528 11348
rect 15476 11305 15485 11339
rect 15485 11305 15519 11339
rect 15519 11305 15528 11339
rect 15476 11296 15528 11305
rect 15568 11296 15620 11348
rect 8024 11228 8076 11280
rect 9956 11228 10008 11280
rect 5724 11203 5776 11212
rect 5724 11169 5733 11203
rect 5733 11169 5767 11203
rect 5767 11169 5776 11203
rect 5724 11160 5776 11169
rect 6184 11203 6236 11212
rect 6184 11169 6193 11203
rect 6193 11169 6227 11203
rect 6227 11169 6236 11203
rect 6184 11160 6236 11169
rect 6460 11203 6512 11212
rect 6460 11169 6469 11203
rect 6469 11169 6503 11203
rect 6503 11169 6512 11203
rect 6460 11160 6512 11169
rect 6644 11203 6696 11212
rect 6644 11169 6653 11203
rect 6653 11169 6687 11203
rect 6687 11169 6696 11203
rect 6644 11160 6696 11169
rect 9496 11203 9548 11212
rect 9496 11169 9505 11203
rect 9505 11169 9539 11203
rect 9539 11169 9548 11203
rect 10324 11228 10376 11280
rect 11520 11228 11572 11280
rect 16488 11228 16540 11280
rect 17132 11228 17184 11280
rect 17776 11271 17828 11280
rect 17776 11237 17785 11271
rect 17785 11237 17819 11271
rect 17819 11237 17828 11271
rect 17776 11228 17828 11237
rect 18696 11271 18748 11280
rect 18696 11237 18705 11271
rect 18705 11237 18739 11271
rect 18739 11237 18748 11271
rect 18696 11228 18748 11237
rect 18880 11228 18932 11280
rect 9496 11160 9548 11169
rect 10140 11160 10192 11212
rect 10600 11203 10652 11212
rect 10600 11169 10609 11203
rect 10609 11169 10643 11203
rect 10643 11169 10652 11203
rect 10600 11160 10652 11169
rect 8852 11092 8904 11144
rect 14004 11160 14056 11212
rect 15200 11160 15252 11212
rect 13268 11092 13320 11144
rect 17408 11092 17460 11144
rect 18972 11135 19024 11144
rect 18972 11101 18981 11135
rect 18981 11101 19015 11135
rect 19015 11101 19024 11135
rect 18972 11092 19024 11101
rect 12440 11024 12492 11076
rect 13728 11024 13780 11076
rect 7932 10956 7984 11008
rect 8760 10999 8812 11008
rect 8760 10965 8769 10999
rect 8769 10965 8803 10999
rect 8803 10965 8812 10999
rect 8760 10956 8812 10965
rect 12348 10956 12400 11008
rect 13360 10956 13412 11008
rect 15844 10999 15896 11008
rect 15844 10965 15853 10999
rect 15853 10965 15887 10999
rect 15887 10965 15896 10999
rect 15844 10956 15896 10965
rect 18144 10999 18196 11008
rect 18144 10965 18153 10999
rect 18153 10965 18187 10999
rect 18187 10965 18196 10999
rect 18144 10956 18196 10965
rect 4982 10854 5034 10906
rect 5046 10854 5098 10906
rect 5110 10854 5162 10906
rect 5174 10854 5226 10906
rect 12982 10854 13034 10906
rect 13046 10854 13098 10906
rect 13110 10854 13162 10906
rect 13174 10854 13226 10906
rect 20982 10854 21034 10906
rect 21046 10854 21098 10906
rect 21110 10854 21162 10906
rect 21174 10854 21226 10906
rect 1952 10795 2004 10804
rect 1952 10761 1961 10795
rect 1961 10761 1995 10795
rect 1995 10761 2004 10795
rect 1952 10752 2004 10761
rect 6644 10752 6696 10804
rect 12808 10752 12860 10804
rect 15200 10795 15252 10804
rect 6184 10684 6236 10736
rect 6460 10684 6512 10736
rect 6552 10684 6604 10736
rect 8300 10616 8352 10668
rect 1952 10548 2004 10600
rect 5724 10548 5776 10600
rect 8116 10591 8168 10600
rect 8116 10557 8125 10591
rect 8125 10557 8159 10591
rect 8159 10557 8168 10591
rect 8116 10548 8168 10557
rect 10048 10616 10100 10668
rect 15200 10761 15209 10795
rect 15209 10761 15243 10795
rect 15243 10761 15252 10795
rect 15200 10752 15252 10761
rect 17132 10795 17184 10804
rect 17132 10761 17141 10795
rect 17141 10761 17175 10795
rect 17175 10761 17184 10795
rect 17132 10752 17184 10761
rect 17408 10795 17460 10804
rect 17408 10761 17417 10795
rect 17417 10761 17451 10795
rect 17451 10761 17460 10795
rect 17408 10752 17460 10761
rect 18696 10752 18748 10804
rect 13176 10684 13228 10736
rect 15108 10684 15160 10736
rect 6276 10480 6328 10532
rect 7840 10480 7892 10532
rect 8852 10548 8904 10600
rect 10140 10548 10192 10600
rect 13360 10591 13412 10600
rect 13360 10557 13369 10591
rect 13369 10557 13403 10591
rect 13403 10557 13412 10591
rect 13360 10548 13412 10557
rect 15844 10616 15896 10668
rect 21364 10684 21416 10736
rect 18328 10616 18380 10668
rect 13912 10591 13964 10600
rect 9680 10480 9732 10532
rect 10048 10480 10100 10532
rect 3332 10412 3384 10464
rect 4344 10455 4396 10464
rect 4344 10421 4353 10455
rect 4353 10421 4387 10455
rect 4387 10421 4396 10455
rect 4344 10412 4396 10421
rect 7932 10455 7984 10464
rect 7932 10421 7941 10455
rect 7941 10421 7975 10455
rect 7975 10421 7984 10455
rect 7932 10412 7984 10421
rect 11152 10455 11204 10464
rect 11152 10421 11161 10455
rect 11161 10421 11195 10455
rect 11195 10421 11204 10455
rect 11152 10412 11204 10421
rect 12348 10480 12400 10532
rect 13912 10557 13921 10591
rect 13921 10557 13955 10591
rect 13955 10557 13964 10591
rect 13912 10548 13964 10557
rect 14280 10591 14332 10600
rect 14280 10557 14289 10591
rect 14289 10557 14323 10591
rect 14323 10557 14332 10591
rect 14280 10548 14332 10557
rect 15108 10480 15160 10532
rect 15476 10480 15528 10532
rect 11704 10412 11756 10464
rect 13176 10412 13228 10464
rect 20076 10548 20128 10600
rect 18144 10523 18196 10532
rect 18144 10489 18153 10523
rect 18153 10489 18187 10523
rect 18187 10489 18196 10523
rect 18144 10480 18196 10489
rect 18880 10412 18932 10464
rect 8982 10310 9034 10362
rect 9046 10310 9098 10362
rect 9110 10310 9162 10362
rect 9174 10310 9226 10362
rect 16982 10310 17034 10362
rect 17046 10310 17098 10362
rect 17110 10310 17162 10362
rect 17174 10310 17226 10362
rect 8024 10208 8076 10260
rect 9496 10251 9548 10260
rect 9496 10217 9505 10251
rect 9505 10217 9539 10251
rect 9539 10217 9548 10251
rect 9496 10208 9548 10217
rect 13728 10208 13780 10260
rect 14280 10208 14332 10260
rect 18144 10208 18196 10260
rect 3792 10140 3844 10192
rect 5448 10140 5500 10192
rect 5908 10140 5960 10192
rect 6184 10140 6236 10192
rect 3700 10072 3752 10124
rect 5540 10072 5592 10124
rect 5724 10072 5776 10124
rect 6276 10072 6328 10124
rect 10600 10140 10652 10192
rect 11152 10140 11204 10192
rect 13452 10140 13504 10192
rect 16212 10183 16264 10192
rect 16212 10149 16221 10183
rect 16221 10149 16255 10183
rect 16255 10149 16264 10183
rect 16212 10140 16264 10149
rect 17776 10183 17828 10192
rect 17776 10149 17785 10183
rect 17785 10149 17819 10183
rect 17819 10149 17828 10183
rect 17776 10140 17828 10149
rect 18328 10183 18380 10192
rect 18328 10149 18337 10183
rect 18337 10149 18371 10183
rect 18371 10149 18380 10183
rect 18328 10140 18380 10149
rect 6552 10072 6604 10124
rect 6736 10072 6788 10124
rect 8852 10072 8904 10124
rect 12348 10115 12400 10124
rect 12348 10081 12357 10115
rect 12357 10081 12391 10115
rect 12391 10081 12400 10115
rect 12348 10072 12400 10081
rect 19156 10115 19208 10124
rect 19156 10081 19165 10115
rect 19165 10081 19199 10115
rect 19199 10081 19208 10115
rect 19156 10072 19208 10081
rect 10232 10047 10284 10056
rect 3332 9936 3384 9988
rect 10232 10013 10241 10047
rect 10241 10013 10275 10047
rect 10275 10013 10284 10047
rect 10232 10004 10284 10013
rect 11888 10004 11940 10056
rect 13452 10004 13504 10056
rect 16488 10004 16540 10056
rect 16764 10047 16816 10056
rect 16764 10013 16773 10047
rect 16773 10013 16807 10047
rect 16807 10013 16816 10047
rect 16764 10004 16816 10013
rect 17684 10047 17736 10056
rect 17684 10013 17693 10047
rect 17693 10013 17727 10047
rect 17727 10013 17736 10047
rect 17684 10004 17736 10013
rect 7196 9979 7248 9988
rect 7196 9945 7205 9979
rect 7205 9945 7239 9979
rect 7239 9945 7248 9979
rect 7196 9936 7248 9945
rect 3976 9868 4028 9920
rect 8300 9911 8352 9920
rect 8300 9877 8309 9911
rect 8309 9877 8343 9911
rect 8343 9877 8352 9911
rect 8300 9868 8352 9877
rect 9680 9868 9732 9920
rect 11152 9911 11204 9920
rect 11152 9877 11161 9911
rect 11161 9877 11195 9911
rect 11195 9877 11204 9911
rect 11152 9868 11204 9877
rect 13636 9911 13688 9920
rect 13636 9877 13645 9911
rect 13645 9877 13679 9911
rect 13679 9877 13688 9911
rect 13636 9868 13688 9877
rect 15568 9911 15620 9920
rect 15568 9877 15577 9911
rect 15577 9877 15611 9911
rect 15611 9877 15620 9911
rect 15568 9868 15620 9877
rect 4982 9766 5034 9818
rect 5046 9766 5098 9818
rect 5110 9766 5162 9818
rect 5174 9766 5226 9818
rect 12982 9766 13034 9818
rect 13046 9766 13098 9818
rect 13110 9766 13162 9818
rect 13174 9766 13226 9818
rect 20982 9766 21034 9818
rect 21046 9766 21098 9818
rect 21110 9766 21162 9818
rect 21174 9766 21226 9818
rect 3700 9707 3752 9716
rect 3700 9673 3709 9707
rect 3709 9673 3743 9707
rect 3743 9673 3752 9707
rect 3700 9664 3752 9673
rect 3792 9664 3844 9716
rect 4344 9664 4396 9716
rect 6552 9664 6604 9716
rect 8852 9664 8904 9716
rect 9772 9707 9824 9716
rect 9772 9673 9781 9707
rect 9781 9673 9815 9707
rect 9815 9673 9824 9707
rect 9772 9664 9824 9673
rect 10600 9707 10652 9716
rect 10600 9673 10609 9707
rect 10609 9673 10643 9707
rect 10643 9673 10652 9707
rect 10600 9664 10652 9673
rect 12348 9664 12400 9716
rect 17960 9664 18012 9716
rect 19156 9707 19208 9716
rect 19156 9673 19165 9707
rect 19165 9673 19199 9707
rect 19199 9673 19208 9707
rect 19156 9664 19208 9673
rect 2320 9596 2372 9648
rect 4068 9528 4120 9580
rect 8024 9596 8076 9648
rect 7196 9528 7248 9580
rect 10140 9596 10192 9648
rect 16672 9596 16724 9648
rect 16764 9596 16816 9648
rect 18972 9596 19024 9648
rect 13636 9528 13688 9580
rect 15568 9571 15620 9580
rect 15568 9537 15577 9571
rect 15577 9537 15611 9571
rect 15611 9537 15620 9571
rect 15568 9528 15620 9537
rect 17684 9528 17736 9580
rect 3976 9392 4028 9444
rect 4804 9392 4856 9444
rect 5448 9392 5500 9444
rect 6276 9367 6328 9376
rect 6276 9333 6285 9367
rect 6285 9333 6319 9367
rect 6319 9333 6328 9367
rect 6276 9324 6328 9333
rect 6552 9367 6604 9376
rect 6552 9333 6561 9367
rect 6561 9333 6595 9367
rect 6595 9333 6604 9367
rect 7932 9392 7984 9444
rect 8668 9435 8720 9444
rect 8668 9401 8677 9435
rect 8677 9401 8711 9435
rect 8711 9401 8720 9435
rect 8668 9392 8720 9401
rect 8760 9435 8812 9444
rect 8760 9401 8769 9435
rect 8769 9401 8803 9435
rect 8803 9401 8812 9435
rect 10876 9435 10928 9444
rect 8760 9392 8812 9401
rect 10876 9401 10885 9435
rect 10885 9401 10919 9435
rect 10919 9401 10928 9435
rect 10876 9392 10928 9401
rect 6552 9324 6604 9333
rect 7840 9324 7892 9376
rect 10600 9324 10652 9376
rect 11244 9392 11296 9444
rect 13452 9460 13504 9512
rect 14280 9503 14332 9512
rect 14280 9469 14289 9503
rect 14289 9469 14323 9503
rect 14323 9469 14332 9503
rect 14280 9460 14332 9469
rect 14004 9392 14056 9444
rect 17776 9503 17828 9512
rect 17776 9469 17785 9503
rect 17785 9469 17819 9503
rect 17819 9469 17828 9503
rect 17776 9460 17828 9469
rect 13268 9324 13320 9376
rect 15476 9367 15528 9376
rect 15476 9333 15485 9367
rect 15485 9333 15519 9367
rect 15519 9333 15528 9367
rect 15476 9324 15528 9333
rect 17500 9324 17552 9376
rect 18144 9435 18196 9444
rect 18144 9401 18153 9435
rect 18153 9401 18187 9435
rect 18187 9401 18196 9435
rect 18144 9392 18196 9401
rect 18604 9392 18656 9444
rect 20076 9503 20128 9512
rect 20076 9469 20085 9503
rect 20085 9469 20119 9503
rect 20119 9469 20128 9503
rect 20076 9460 20128 9469
rect 8982 9222 9034 9274
rect 9046 9222 9098 9274
rect 9110 9222 9162 9274
rect 9174 9222 9226 9274
rect 16982 9222 17034 9274
rect 17046 9222 17098 9274
rect 17110 9222 17162 9274
rect 17174 9222 17226 9274
rect 4804 9163 4856 9172
rect 4804 9129 4813 9163
rect 4813 9129 4847 9163
rect 4847 9129 4856 9163
rect 4804 9120 4856 9129
rect 5908 9163 5960 9172
rect 5908 9129 5917 9163
rect 5917 9129 5951 9163
rect 5951 9129 5960 9163
rect 5908 9120 5960 9129
rect 6644 9120 6696 9172
rect 7196 9120 7248 9172
rect 10876 9120 10928 9172
rect 13728 9120 13780 9172
rect 16212 9163 16264 9172
rect 112 9052 164 9104
rect 7840 9095 7892 9104
rect 7840 9061 7849 9095
rect 7849 9061 7883 9095
rect 7883 9061 7892 9095
rect 7840 9052 7892 9061
rect 1676 8984 1728 9036
rect 2320 8984 2372 9036
rect 10140 9052 10192 9104
rect 10232 9052 10284 9104
rect 11060 9095 11112 9104
rect 11060 9061 11069 9095
rect 11069 9061 11103 9095
rect 11103 9061 11112 9095
rect 11060 9052 11112 9061
rect 16212 9129 16221 9163
rect 16221 9129 16255 9163
rect 16255 9129 16264 9163
rect 16212 9120 16264 9129
rect 17684 9120 17736 9172
rect 21272 9120 21324 9172
rect 15476 9052 15528 9104
rect 15844 9052 15896 9104
rect 17500 9052 17552 9104
rect 18328 9052 18380 9104
rect 13268 8984 13320 9036
rect 13452 9027 13504 9036
rect 13452 8993 13461 9027
rect 13461 8993 13495 9027
rect 13495 8993 13504 9027
rect 13452 8984 13504 8993
rect 7748 8959 7800 8968
rect 7748 8925 7757 8959
rect 7757 8925 7791 8959
rect 7791 8925 7800 8959
rect 7748 8916 7800 8925
rect 8024 8959 8076 8968
rect 8024 8925 8033 8959
rect 8033 8925 8067 8959
rect 8067 8925 8076 8959
rect 8024 8916 8076 8925
rect 10968 8959 11020 8968
rect 10968 8925 10977 8959
rect 10977 8925 11011 8959
rect 11011 8925 11020 8959
rect 10968 8916 11020 8925
rect 11244 8959 11296 8968
rect 11244 8925 11253 8959
rect 11253 8925 11287 8959
rect 11287 8925 11296 8959
rect 11244 8916 11296 8925
rect 12808 8916 12860 8968
rect 13912 8984 13964 9036
rect 14004 8984 14056 9036
rect 18604 9027 18656 9036
rect 18604 8993 18613 9027
rect 18613 8993 18647 9027
rect 18647 8993 18656 9027
rect 18604 8984 18656 8993
rect 20076 8984 20128 9036
rect 20812 8984 20864 9036
rect 14832 8916 14884 8968
rect 17132 8959 17184 8968
rect 17132 8925 17141 8959
rect 17141 8925 17175 8959
rect 17175 8925 17184 8959
rect 17132 8916 17184 8925
rect 18144 8916 18196 8968
rect 10416 8848 10468 8900
rect 10692 8823 10744 8832
rect 10692 8789 10701 8823
rect 10701 8789 10735 8823
rect 10735 8789 10744 8823
rect 10692 8780 10744 8789
rect 16488 8823 16540 8832
rect 16488 8789 16497 8823
rect 16497 8789 16531 8823
rect 16531 8789 16540 8823
rect 16488 8780 16540 8789
rect 18512 8780 18564 8832
rect 4982 8678 5034 8730
rect 5046 8678 5098 8730
rect 5110 8678 5162 8730
rect 5174 8678 5226 8730
rect 12982 8678 13034 8730
rect 13046 8678 13098 8730
rect 13110 8678 13162 8730
rect 13174 8678 13226 8730
rect 20982 8678 21034 8730
rect 21046 8678 21098 8730
rect 21110 8678 21162 8730
rect 21174 8678 21226 8730
rect 1768 8576 1820 8628
rect 7840 8576 7892 8628
rect 10140 8576 10192 8628
rect 10968 8576 11020 8628
rect 13452 8576 13504 8628
rect 14832 8619 14884 8628
rect 14832 8585 14841 8619
rect 14841 8585 14875 8619
rect 14875 8585 14884 8619
rect 14832 8576 14884 8585
rect 16488 8576 16540 8628
rect 16856 8576 16908 8628
rect 17132 8576 17184 8628
rect 17500 8619 17552 8628
rect 17500 8585 17509 8619
rect 17509 8585 17543 8619
rect 17543 8585 17552 8619
rect 17500 8576 17552 8585
rect 20076 8619 20128 8628
rect 20076 8585 20085 8619
rect 20085 8585 20119 8619
rect 20119 8585 20128 8619
rect 20076 8576 20128 8585
rect 8668 8508 8720 8560
rect 11888 8508 11940 8560
rect 14188 8508 14240 8560
rect 18604 8551 18656 8560
rect 18604 8517 18613 8551
rect 18613 8517 18647 8551
rect 18647 8517 18656 8551
rect 18604 8508 18656 8517
rect 10692 8440 10744 8492
rect 12624 8440 12676 8492
rect 2780 8372 2832 8424
rect 14096 8372 14148 8424
rect 19064 8415 19116 8424
rect 8024 8304 8076 8356
rect 8392 8347 8444 8356
rect 8392 8313 8401 8347
rect 8401 8313 8435 8347
rect 8435 8313 8444 8347
rect 8392 8304 8444 8313
rect 2044 8279 2096 8288
rect 2044 8245 2053 8279
rect 2053 8245 2087 8279
rect 2087 8245 2096 8279
rect 2044 8236 2096 8245
rect 8116 8279 8168 8288
rect 8116 8245 8125 8279
rect 8125 8245 8159 8279
rect 8159 8245 8168 8279
rect 10416 8304 10468 8356
rect 13268 8304 13320 8356
rect 13820 8304 13872 8356
rect 8116 8236 8168 8245
rect 11060 8236 11112 8288
rect 11520 8236 11572 8288
rect 12808 8236 12860 8288
rect 14004 8279 14056 8288
rect 14004 8245 14013 8279
rect 14013 8245 14047 8279
rect 14047 8245 14056 8279
rect 14004 8236 14056 8245
rect 15844 8279 15896 8288
rect 15844 8245 15853 8279
rect 15853 8245 15887 8279
rect 15887 8245 15896 8279
rect 15844 8236 15896 8245
rect 19064 8381 19073 8415
rect 19073 8381 19107 8415
rect 19107 8381 19116 8415
rect 19064 8372 19116 8381
rect 21364 8576 21416 8628
rect 21272 8508 21324 8560
rect 19708 8304 19760 8356
rect 20812 8304 20864 8356
rect 17316 8236 17368 8288
rect 19432 8279 19484 8288
rect 19432 8245 19441 8279
rect 19441 8245 19475 8279
rect 19475 8245 19484 8279
rect 19432 8236 19484 8245
rect 8982 8134 9034 8186
rect 9046 8134 9098 8186
rect 9110 8134 9162 8186
rect 9174 8134 9226 8186
rect 16982 8134 17034 8186
rect 17046 8134 17098 8186
rect 17110 8134 17162 8186
rect 17174 8134 17226 8186
rect 1676 8075 1728 8084
rect 1676 8041 1685 8075
rect 1685 8041 1719 8075
rect 1719 8041 1728 8075
rect 1676 8032 1728 8041
rect 8116 8032 8168 8084
rect 10048 8075 10100 8084
rect 10048 8041 10057 8075
rect 10057 8041 10091 8075
rect 10091 8041 10100 8075
rect 10048 8032 10100 8041
rect 6644 7964 6696 8016
rect 7748 7964 7800 8016
rect 10416 7964 10468 8016
rect 16856 8032 16908 8084
rect 11520 7964 11572 8016
rect 15844 7964 15896 8016
rect 18052 7964 18104 8016
rect 19432 8007 19484 8016
rect 19432 7973 19441 8007
rect 19441 7973 19475 8007
rect 19475 7973 19484 8007
rect 19432 7964 19484 7973
rect 6736 7871 6788 7880
rect 6736 7837 6745 7871
rect 6745 7837 6779 7871
rect 6779 7837 6788 7871
rect 6736 7828 6788 7837
rect 7288 7760 7340 7812
rect 8392 7735 8444 7744
rect 8392 7701 8401 7735
rect 8401 7701 8435 7735
rect 8435 7701 8444 7735
rect 8392 7692 8444 7701
rect 8668 7692 8720 7744
rect 11796 7828 11848 7880
rect 11888 7871 11940 7880
rect 11888 7837 11897 7871
rect 11897 7837 11931 7871
rect 11931 7837 11940 7871
rect 15384 7871 15436 7880
rect 11888 7828 11940 7837
rect 15384 7837 15393 7871
rect 15393 7837 15427 7871
rect 15427 7837 15436 7871
rect 15384 7828 15436 7837
rect 18512 7828 18564 7880
rect 18880 7828 18932 7880
rect 18328 7803 18380 7812
rect 18328 7769 18337 7803
rect 18337 7769 18371 7803
rect 18371 7769 18380 7803
rect 18328 7760 18380 7769
rect 19708 7760 19760 7812
rect 9680 7692 9732 7744
rect 10876 7735 10928 7744
rect 10876 7701 10885 7735
rect 10885 7701 10919 7735
rect 10919 7701 10928 7735
rect 10876 7692 10928 7701
rect 12716 7692 12768 7744
rect 13728 7692 13780 7744
rect 19064 7692 19116 7744
rect 4982 7590 5034 7642
rect 5046 7590 5098 7642
rect 5110 7590 5162 7642
rect 5174 7590 5226 7642
rect 12982 7590 13034 7642
rect 13046 7590 13098 7642
rect 13110 7590 13162 7642
rect 13174 7590 13226 7642
rect 20982 7590 21034 7642
rect 21046 7590 21098 7642
rect 21110 7590 21162 7642
rect 21174 7590 21226 7642
rect 9772 7488 9824 7540
rect 6276 7284 6328 7336
rect 7288 7327 7340 7336
rect 7288 7293 7297 7327
rect 7297 7293 7331 7327
rect 7331 7293 7340 7327
rect 7288 7284 7340 7293
rect 7656 7284 7708 7336
rect 8300 7420 8352 7472
rect 9312 7420 9364 7472
rect 8208 7327 8260 7336
rect 8208 7293 8217 7327
rect 8217 7293 8251 7327
rect 8251 7293 8260 7327
rect 8208 7284 8260 7293
rect 9496 7284 9548 7336
rect 9680 7327 9732 7336
rect 9680 7293 9689 7327
rect 9689 7293 9723 7327
rect 9723 7293 9732 7327
rect 9680 7284 9732 7293
rect 11060 7488 11112 7540
rect 11520 7531 11572 7540
rect 11520 7497 11529 7531
rect 11529 7497 11563 7531
rect 11563 7497 11572 7531
rect 11520 7488 11572 7497
rect 11796 7531 11848 7540
rect 11796 7497 11805 7531
rect 11805 7497 11839 7531
rect 11839 7497 11848 7531
rect 11796 7488 11848 7497
rect 18512 7488 18564 7540
rect 18880 7531 18932 7540
rect 18880 7497 18889 7531
rect 18889 7497 18923 7531
rect 18923 7497 18932 7531
rect 18880 7488 18932 7497
rect 19432 7488 19484 7540
rect 10876 7352 10928 7404
rect 15384 7352 15436 7404
rect 19708 7395 19760 7404
rect 19708 7361 19717 7395
rect 19717 7361 19751 7395
rect 19751 7361 19760 7395
rect 19708 7352 19760 7361
rect 12716 7284 12768 7336
rect 3056 7148 3108 7200
rect 6644 7148 6696 7200
rect 6736 7148 6788 7200
rect 8668 7191 8720 7200
rect 8668 7157 8677 7191
rect 8677 7157 8711 7191
rect 8711 7157 8720 7191
rect 8668 7148 8720 7157
rect 8852 7148 8904 7200
rect 13728 7284 13780 7336
rect 14280 7284 14332 7336
rect 9312 7148 9364 7200
rect 12532 7148 12584 7200
rect 13452 7148 13504 7200
rect 13636 7148 13688 7200
rect 15016 7191 15068 7200
rect 15016 7157 15025 7191
rect 15025 7157 15059 7191
rect 15059 7157 15068 7191
rect 15016 7148 15068 7157
rect 15844 7148 15896 7200
rect 18328 7216 18380 7268
rect 19156 7259 19208 7268
rect 19156 7225 19165 7259
rect 19165 7225 19199 7259
rect 19199 7225 19208 7259
rect 19156 7216 19208 7225
rect 16580 7191 16632 7200
rect 16580 7157 16589 7191
rect 16589 7157 16623 7191
rect 16623 7157 16632 7191
rect 16580 7148 16632 7157
rect 18052 7148 18104 7200
rect 8982 7046 9034 7098
rect 9046 7046 9098 7098
rect 9110 7046 9162 7098
rect 9174 7046 9226 7098
rect 16982 7046 17034 7098
rect 17046 7046 17098 7098
rect 17110 7046 17162 7098
rect 17174 7046 17226 7098
rect 8208 6944 8260 6996
rect 8392 6944 8444 6996
rect 9496 6944 9548 6996
rect 10048 6944 10100 6996
rect 11060 6987 11112 6996
rect 11060 6953 11069 6987
rect 11069 6953 11103 6987
rect 11103 6953 11112 6987
rect 11060 6944 11112 6953
rect 12532 6944 12584 6996
rect 13636 6944 13688 6996
rect 15384 6944 15436 6996
rect 19064 6987 19116 6996
rect 19064 6953 19073 6987
rect 19073 6953 19107 6987
rect 19107 6953 19116 6987
rect 19064 6944 19116 6953
rect 9588 6876 9640 6928
rect 12624 6876 12676 6928
rect 15016 6876 15068 6928
rect 16580 6876 16632 6928
rect 17868 6876 17920 6928
rect 7656 6808 7708 6860
rect 10416 6851 10468 6860
rect 10416 6817 10425 6851
rect 10425 6817 10459 6851
rect 10459 6817 10468 6851
rect 10416 6808 10468 6817
rect 12716 6808 12768 6860
rect 13452 6851 13504 6860
rect 13452 6817 13461 6851
rect 13461 6817 13495 6851
rect 13495 6817 13504 6851
rect 13452 6808 13504 6817
rect 13728 6851 13780 6860
rect 13728 6817 13737 6851
rect 13737 6817 13771 6851
rect 13771 6817 13780 6851
rect 13728 6808 13780 6817
rect 14648 6808 14700 6860
rect 15292 6808 15344 6860
rect 17040 6808 17092 6860
rect 17316 6808 17368 6860
rect 10048 6740 10100 6792
rect 4804 6604 4856 6656
rect 7288 6672 7340 6724
rect 9772 6672 9824 6724
rect 11520 6672 11572 6724
rect 18328 6783 18380 6792
rect 18328 6749 18337 6783
rect 18337 6749 18371 6783
rect 18371 6749 18380 6783
rect 18328 6740 18380 6749
rect 10600 6604 10652 6656
rect 10692 6647 10744 6656
rect 10692 6613 10701 6647
rect 10701 6613 10735 6647
rect 10735 6613 10744 6647
rect 12716 6647 12768 6656
rect 10692 6604 10744 6613
rect 12716 6613 12725 6647
rect 12725 6613 12759 6647
rect 12759 6613 12768 6647
rect 12716 6604 12768 6613
rect 15568 6604 15620 6656
rect 15844 6647 15896 6656
rect 15844 6613 15853 6647
rect 15853 6613 15887 6647
rect 15887 6613 15896 6647
rect 15844 6604 15896 6613
rect 17408 6604 17460 6656
rect 4982 6502 5034 6554
rect 5046 6502 5098 6554
rect 5110 6502 5162 6554
rect 5174 6502 5226 6554
rect 12982 6502 13034 6554
rect 13046 6502 13098 6554
rect 13110 6502 13162 6554
rect 13174 6502 13226 6554
rect 20982 6502 21034 6554
rect 21046 6502 21098 6554
rect 21110 6502 21162 6554
rect 21174 6502 21226 6554
rect 10692 6400 10744 6452
rect 15292 6443 15344 6452
rect 15292 6409 15301 6443
rect 15301 6409 15335 6443
rect 15335 6409 15344 6443
rect 15292 6400 15344 6409
rect 16028 6400 16080 6452
rect 17408 6443 17460 6452
rect 17408 6409 17417 6443
rect 17417 6409 17451 6443
rect 17451 6409 17460 6443
rect 17408 6400 17460 6409
rect 17868 6443 17920 6452
rect 17868 6409 17877 6443
rect 17877 6409 17911 6443
rect 17911 6409 17920 6443
rect 17868 6400 17920 6409
rect 8852 6332 8904 6384
rect 12808 6332 12860 6384
rect 13268 6375 13320 6384
rect 13268 6341 13277 6375
rect 13277 6341 13311 6375
rect 13311 6341 13320 6375
rect 13268 6332 13320 6341
rect 13636 6332 13688 6384
rect 9772 6307 9824 6316
rect 9772 6273 9781 6307
rect 9781 6273 9815 6307
rect 9815 6273 9824 6307
rect 9772 6264 9824 6273
rect 10600 6307 10652 6316
rect 10600 6273 10609 6307
rect 10609 6273 10643 6307
rect 10643 6273 10652 6307
rect 10600 6264 10652 6273
rect 18052 6307 18104 6316
rect 18052 6273 18061 6307
rect 18061 6273 18095 6307
rect 18095 6273 18104 6307
rect 18052 6264 18104 6273
rect 11244 6239 11296 6248
rect 11244 6205 11253 6239
rect 11253 6205 11287 6239
rect 11287 6205 11296 6239
rect 11244 6196 11296 6205
rect 13360 6196 13412 6248
rect 9312 6128 9364 6180
rect 9588 6060 9640 6112
rect 10048 6103 10100 6112
rect 10048 6069 10057 6103
rect 10057 6069 10091 6103
rect 10091 6069 10100 6103
rect 10048 6060 10100 6069
rect 12072 6060 12124 6112
rect 13452 6060 13504 6112
rect 14280 6239 14332 6248
rect 14280 6205 14289 6239
rect 14289 6205 14323 6239
rect 14323 6205 14332 6239
rect 14280 6196 14332 6205
rect 14648 6239 14700 6248
rect 14648 6205 14657 6239
rect 14657 6205 14691 6239
rect 14691 6205 14700 6239
rect 14648 6196 14700 6205
rect 15752 6239 15804 6248
rect 15752 6205 15761 6239
rect 15761 6205 15795 6239
rect 15795 6205 15804 6239
rect 15752 6196 15804 6205
rect 17868 6196 17920 6248
rect 13636 6060 13688 6112
rect 15844 6128 15896 6180
rect 17040 6171 17092 6180
rect 17040 6137 17049 6171
rect 17049 6137 17083 6171
rect 17083 6137 17092 6171
rect 17040 6128 17092 6137
rect 18328 6128 18380 6180
rect 8982 5958 9034 6010
rect 9046 5958 9098 6010
rect 9110 5958 9162 6010
rect 9174 5958 9226 6010
rect 16982 5958 17034 6010
rect 17046 5958 17098 6010
rect 17110 5958 17162 6010
rect 17174 5958 17226 6010
rect 15752 5856 15804 5908
rect 17868 5856 17920 5908
rect 11336 5831 11388 5840
rect 11336 5797 11345 5831
rect 11345 5797 11379 5831
rect 11379 5797 11388 5831
rect 11336 5788 11388 5797
rect 14004 5788 14056 5840
rect 16948 5831 17000 5840
rect 16948 5797 16957 5831
rect 16957 5797 16991 5831
rect 16991 5797 17000 5831
rect 16948 5788 17000 5797
rect 9312 5763 9364 5772
rect 9312 5729 9321 5763
rect 9321 5729 9355 5763
rect 9355 5729 9364 5763
rect 9312 5720 9364 5729
rect 9864 5720 9916 5772
rect 10416 5720 10468 5772
rect 11888 5720 11940 5772
rect 12164 5763 12216 5772
rect 12164 5729 12173 5763
rect 12173 5729 12207 5763
rect 12207 5729 12216 5763
rect 12164 5720 12216 5729
rect 18328 5763 18380 5772
rect 18328 5729 18337 5763
rect 18337 5729 18371 5763
rect 18371 5729 18380 5763
rect 18328 5720 18380 5729
rect 10140 5652 10192 5704
rect 10876 5652 10928 5704
rect 11796 5652 11848 5704
rect 11244 5584 11296 5636
rect 11888 5584 11940 5636
rect 13360 5584 13412 5636
rect 16764 5584 16816 5636
rect 17408 5627 17460 5636
rect 17408 5593 17417 5627
rect 17417 5593 17451 5627
rect 17451 5593 17460 5627
rect 17408 5584 17460 5593
rect 17776 5584 17828 5636
rect 10416 5559 10468 5568
rect 10416 5525 10425 5559
rect 10425 5525 10459 5559
rect 10459 5525 10468 5559
rect 10416 5516 10468 5525
rect 12716 5516 12768 5568
rect 13452 5559 13504 5568
rect 13452 5525 13461 5559
rect 13461 5525 13495 5559
rect 13495 5525 13504 5559
rect 13452 5516 13504 5525
rect 14280 5559 14332 5568
rect 14280 5525 14289 5559
rect 14289 5525 14323 5559
rect 14323 5525 14332 5559
rect 14280 5516 14332 5525
rect 15752 5559 15804 5568
rect 15752 5525 15761 5559
rect 15761 5525 15795 5559
rect 15795 5525 15804 5559
rect 15752 5516 15804 5525
rect 4982 5414 5034 5466
rect 5046 5414 5098 5466
rect 5110 5414 5162 5466
rect 5174 5414 5226 5466
rect 12982 5414 13034 5466
rect 13046 5414 13098 5466
rect 13110 5414 13162 5466
rect 13174 5414 13226 5466
rect 20982 5414 21034 5466
rect 21046 5414 21098 5466
rect 21110 5414 21162 5466
rect 21174 5414 21226 5466
rect 9864 5355 9916 5364
rect 9864 5321 9873 5355
rect 9873 5321 9907 5355
rect 9907 5321 9916 5355
rect 9864 5312 9916 5321
rect 10692 5312 10744 5364
rect 12164 5312 12216 5364
rect 16764 5312 16816 5364
rect 18328 5355 18380 5364
rect 18328 5321 18337 5355
rect 18337 5321 18371 5355
rect 18371 5321 18380 5355
rect 18328 5312 18380 5321
rect 10876 5244 10928 5296
rect 12716 5244 12768 5296
rect 7656 5219 7708 5228
rect 7656 5185 7665 5219
rect 7665 5185 7699 5219
rect 7699 5185 7708 5219
rect 7656 5176 7708 5185
rect 12072 5176 12124 5228
rect 13452 5176 13504 5228
rect 6552 5108 6604 5160
rect 8852 5108 8904 5160
rect 10416 5151 10468 5160
rect 10416 5117 10425 5151
rect 10425 5117 10459 5151
rect 10459 5117 10468 5151
rect 10416 5108 10468 5117
rect 13360 5151 13412 5160
rect 13360 5117 13369 5151
rect 13369 5117 13403 5151
rect 13403 5117 13412 5151
rect 13360 5108 13412 5117
rect 14280 5176 14332 5228
rect 14556 5151 14608 5160
rect 112 5040 164 5092
rect 11980 5040 12032 5092
rect 14556 5117 14565 5151
rect 14565 5117 14599 5151
rect 14599 5117 14608 5151
rect 14556 5108 14608 5117
rect 15660 5151 15712 5160
rect 15660 5117 15669 5151
rect 15669 5117 15703 5151
rect 15703 5117 15712 5151
rect 15660 5108 15712 5117
rect 16948 5083 17000 5092
rect 6552 5015 6604 5024
rect 6552 4981 6561 5015
rect 6561 4981 6595 5015
rect 6595 4981 6604 5015
rect 6552 4972 6604 4981
rect 11796 4972 11848 5024
rect 15200 4972 15252 5024
rect 15752 4972 15804 5024
rect 16948 5049 16957 5083
rect 16957 5049 16991 5083
rect 16991 5049 17000 5083
rect 16948 5040 17000 5049
rect 18512 5040 18564 5092
rect 8982 4870 9034 4922
rect 9046 4870 9098 4922
rect 9110 4870 9162 4922
rect 9174 4870 9226 4922
rect 16982 4870 17034 4922
rect 17046 4870 17098 4922
rect 17110 4870 17162 4922
rect 17174 4870 17226 4922
rect 9864 4768 9916 4820
rect 10692 4768 10744 4820
rect 10876 4768 10928 4820
rect 11520 4811 11572 4820
rect 11520 4777 11529 4811
rect 11529 4777 11563 4811
rect 11563 4777 11572 4811
rect 11520 4768 11572 4777
rect 13452 4811 13504 4820
rect 13452 4777 13461 4811
rect 13461 4777 13495 4811
rect 13495 4777 13504 4811
rect 13452 4768 13504 4777
rect 13636 4768 13688 4820
rect 1216 4632 1268 4684
rect 9680 4632 9732 4684
rect 11612 4675 11664 4684
rect 11612 4641 11621 4675
rect 11621 4641 11655 4675
rect 11655 4641 11664 4675
rect 11612 4632 11664 4641
rect 12072 4675 12124 4684
rect 12072 4641 12081 4675
rect 12081 4641 12115 4675
rect 12115 4641 12124 4675
rect 12072 4632 12124 4641
rect 10416 4564 10468 4616
rect 11888 4564 11940 4616
rect 12532 4632 12584 4684
rect 14556 4768 14608 4820
rect 15660 4811 15712 4820
rect 15660 4777 15669 4811
rect 15669 4777 15703 4811
rect 15703 4777 15712 4811
rect 15660 4768 15712 4777
rect 17040 4743 17092 4752
rect 17040 4709 17049 4743
rect 17049 4709 17083 4743
rect 17083 4709 17092 4743
rect 17040 4700 17092 4709
rect 18512 4675 18564 4684
rect 18512 4641 18521 4675
rect 18521 4641 18555 4675
rect 18555 4641 18564 4675
rect 18512 4632 18564 4641
rect 12716 4496 12768 4548
rect 13360 4564 13412 4616
rect 17408 4607 17460 4616
rect 14280 4496 14332 4548
rect 16856 4496 16908 4548
rect 17408 4573 17417 4607
rect 17417 4573 17451 4607
rect 17451 4573 17460 4607
rect 17408 4564 17460 4573
rect 4982 4326 5034 4378
rect 5046 4326 5098 4378
rect 5110 4326 5162 4378
rect 5174 4326 5226 4378
rect 12982 4326 13034 4378
rect 13046 4326 13098 4378
rect 13110 4326 13162 4378
rect 13174 4326 13226 4378
rect 20982 4326 21034 4378
rect 21046 4326 21098 4378
rect 21110 4326 21162 4378
rect 21174 4326 21226 4378
rect 9680 4267 9732 4276
rect 9680 4233 9689 4267
rect 9689 4233 9723 4267
rect 9723 4233 9732 4267
rect 9680 4224 9732 4233
rect 10876 4224 10928 4276
rect 11888 4267 11940 4276
rect 11888 4233 11897 4267
rect 11897 4233 11931 4267
rect 11931 4233 11940 4267
rect 11888 4224 11940 4233
rect 12532 4224 12584 4276
rect 18512 4267 18564 4276
rect 18512 4233 18521 4267
rect 18521 4233 18555 4267
rect 18555 4233 18564 4267
rect 18512 4224 18564 4233
rect 9588 4156 9640 4208
rect 9772 4156 9824 4208
rect 16856 4156 16908 4208
rect 11520 4131 11572 4140
rect 11520 4097 11529 4131
rect 11529 4097 11563 4131
rect 11563 4097 11572 4131
rect 11520 4088 11572 4097
rect 13268 4131 13320 4140
rect 10968 4063 11020 4072
rect 10968 4029 10977 4063
rect 10977 4029 11011 4063
rect 11011 4029 11020 4063
rect 10968 4020 11020 4029
rect 13268 4097 13277 4131
rect 13277 4097 13311 4131
rect 13311 4097 13320 4131
rect 13268 4088 13320 4097
rect 17040 4088 17092 4140
rect 13360 4020 13412 4072
rect 13636 4020 13688 4072
rect 14280 4063 14332 4072
rect 14280 4029 14289 4063
rect 14289 4029 14323 4063
rect 14323 4029 14332 4063
rect 14280 4020 14332 4029
rect 12440 3927 12492 3936
rect 12440 3893 12449 3927
rect 12449 3893 12483 3927
rect 12483 3893 12492 3927
rect 12440 3884 12492 3893
rect 13268 3884 13320 3936
rect 16212 4020 16264 4072
rect 17408 4020 17460 4072
rect 14924 3995 14976 4004
rect 14924 3961 14933 3995
rect 14933 3961 14967 3995
rect 14967 3961 14976 3995
rect 14924 3952 14976 3961
rect 16488 3995 16540 4004
rect 16488 3961 16497 3995
rect 16497 3961 16531 3995
rect 16531 3961 16540 3995
rect 16488 3952 16540 3961
rect 23572 3952 23624 4004
rect 8982 3782 9034 3834
rect 9046 3782 9098 3834
rect 9110 3782 9162 3834
rect 9174 3782 9226 3834
rect 16982 3782 17034 3834
rect 17046 3782 17098 3834
rect 17110 3782 17162 3834
rect 17174 3782 17226 3834
rect 11520 3680 11572 3732
rect 12716 3723 12768 3732
rect 12716 3689 12725 3723
rect 12725 3689 12759 3723
rect 12759 3689 12768 3723
rect 12716 3680 12768 3689
rect 14280 3723 14332 3732
rect 14280 3689 14289 3723
rect 14289 3689 14323 3723
rect 14323 3689 14332 3723
rect 14280 3680 14332 3689
rect 16212 3723 16264 3732
rect 16212 3689 16221 3723
rect 16221 3689 16255 3723
rect 16255 3689 16264 3723
rect 16212 3680 16264 3689
rect 16856 3680 16908 3732
rect 11980 3655 12032 3664
rect 11980 3621 11989 3655
rect 11989 3621 12023 3655
rect 12023 3621 12032 3655
rect 11980 3612 12032 3621
rect 13452 3655 13504 3664
rect 13452 3621 13461 3655
rect 13461 3621 13495 3655
rect 13495 3621 13504 3655
rect 13452 3612 13504 3621
rect 15200 3612 15252 3664
rect 10692 3544 10744 3596
rect 11796 3544 11848 3596
rect 14004 3476 14056 3528
rect 14924 3476 14976 3528
rect 16764 3476 16816 3528
rect 13728 3408 13780 3460
rect 4982 3238 5034 3290
rect 5046 3238 5098 3290
rect 5110 3238 5162 3290
rect 5174 3238 5226 3290
rect 12982 3238 13034 3290
rect 13046 3238 13098 3290
rect 13110 3238 13162 3290
rect 13174 3238 13226 3290
rect 20982 3238 21034 3290
rect 21046 3238 21098 3290
rect 21110 3238 21162 3290
rect 21174 3238 21226 3290
rect 10692 3179 10744 3188
rect 10692 3145 10701 3179
rect 10701 3145 10735 3179
rect 10735 3145 10744 3179
rect 10692 3136 10744 3145
rect 14004 3179 14056 3188
rect 14004 3145 14013 3179
rect 14013 3145 14047 3179
rect 14047 3145 14056 3179
rect 14004 3136 14056 3145
rect 16488 3179 16540 3188
rect 16488 3145 16497 3179
rect 16497 3145 16531 3179
rect 16531 3145 16540 3179
rect 16488 3136 16540 3145
rect 16764 3179 16816 3188
rect 16764 3145 16773 3179
rect 16773 3145 16807 3179
rect 16807 3145 16816 3179
rect 16764 3136 16816 3145
rect 10140 3068 10192 3120
rect 15844 3068 15896 3120
rect 12716 3000 12768 3052
rect 16856 3000 16908 3052
rect 13544 2932 13596 2984
rect 15200 2907 15252 2916
rect 15200 2873 15209 2907
rect 15209 2873 15243 2907
rect 15243 2873 15252 2907
rect 15200 2864 15252 2873
rect 11612 2796 11664 2848
rect 11796 2839 11848 2848
rect 11796 2805 11805 2839
rect 11805 2805 11839 2839
rect 11839 2805 11848 2839
rect 11796 2796 11848 2805
rect 12532 2796 12584 2848
rect 13452 2796 13504 2848
rect 14096 2796 14148 2848
rect 16488 2796 16540 2848
rect 8982 2694 9034 2746
rect 9046 2694 9098 2746
rect 9110 2694 9162 2746
rect 9174 2694 9226 2746
rect 16982 2694 17034 2746
rect 17046 2694 17098 2746
rect 17110 2694 17162 2746
rect 17174 2694 17226 2746
rect 12440 2635 12492 2644
rect 12440 2601 12449 2635
rect 12449 2601 12483 2635
rect 12483 2601 12492 2635
rect 12440 2592 12492 2601
rect 9772 2499 9824 2508
rect 9772 2465 9781 2499
rect 9781 2465 9815 2499
rect 9815 2465 9824 2499
rect 9772 2456 9824 2465
rect 12532 2456 12584 2508
rect 13728 2567 13780 2576
rect 13728 2533 13737 2567
rect 13737 2533 13771 2567
rect 13771 2533 13780 2567
rect 13728 2524 13780 2533
rect 15568 2567 15620 2576
rect 15568 2533 15577 2567
rect 15577 2533 15611 2567
rect 15611 2533 15620 2567
rect 15568 2524 15620 2533
rect 16856 2592 16908 2644
rect 16212 2524 16264 2576
rect 15844 2431 15896 2440
rect 12440 2320 12492 2372
rect 15844 2397 15853 2431
rect 15853 2397 15887 2431
rect 15887 2397 15896 2431
rect 15844 2388 15896 2397
rect 15936 2388 15988 2440
rect 17960 2456 18012 2508
rect 19892 2456 19944 2508
rect 19432 2320 19484 2372
rect 23112 2320 23164 2372
rect 6736 2252 6788 2304
rect 10232 2252 10284 2304
rect 4982 2150 5034 2202
rect 5046 2150 5098 2202
rect 5110 2150 5162 2202
rect 5174 2150 5226 2202
rect 12982 2150 13034 2202
rect 13046 2150 13098 2202
rect 13110 2150 13162 2202
rect 13174 2150 13226 2202
rect 20982 2150 21034 2202
rect 21046 2150 21098 2202
rect 21110 2150 21162 2202
rect 21174 2150 21226 2202
<< metal2 >>
rect 938 23610 994 24000
rect 2870 23610 2926 24000
rect 938 23582 1256 23610
rect 938 23520 994 23582
rect 110 22536 166 22545
rect 110 22471 166 22480
rect 124 15706 152 22471
rect 1228 18873 1256 23582
rect 2792 23582 2926 23610
rect 1766 19272 1822 19281
rect 1766 19207 1822 19216
rect 1214 18864 1270 18873
rect 1214 18799 1270 18808
rect 1398 16688 1454 16697
rect 1398 16623 1454 16632
rect 112 15700 164 15706
rect 112 15642 164 15648
rect 1412 13814 1440 16623
rect 1490 14240 1546 14249
rect 1490 14175 1546 14184
rect 1504 14074 1532 14175
rect 1492 14068 1544 14074
rect 1492 14010 1544 14016
rect 1412 13786 1532 13814
rect 110 11928 166 11937
rect 1504 11898 1532 13786
rect 110 11863 166 11872
rect 1492 11892 1544 11898
rect 124 11694 152 11863
rect 1492 11834 1544 11840
rect 112 11688 164 11694
rect 112 11630 164 11636
rect 110 9208 166 9217
rect 110 9143 166 9152
rect 124 9110 152 9143
rect 112 9104 164 9110
rect 112 9046 164 9052
rect 1676 9036 1728 9042
rect 1676 8978 1728 8984
rect 1688 8090 1716 8978
rect 1780 8634 1808 19207
rect 1952 11688 2004 11694
rect 1952 11630 2004 11636
rect 1964 10810 1992 11630
rect 1952 10804 2004 10810
rect 1952 10746 2004 10752
rect 1964 10606 1992 10746
rect 1952 10600 2004 10606
rect 1952 10542 2004 10548
rect 2320 9648 2372 9654
rect 2320 9590 2372 9596
rect 2332 9042 2360 9590
rect 2320 9036 2372 9042
rect 2320 8978 2372 8984
rect 1768 8628 1820 8634
rect 1768 8570 1820 8576
rect 2792 8430 2820 23582
rect 2870 23520 2926 23582
rect 4894 23610 4950 24000
rect 6918 23610 6974 24000
rect 8942 23610 8998 24000
rect 4894 23582 5396 23610
rect 4894 23520 4950 23582
rect 4956 21788 5252 21808
rect 5012 21786 5036 21788
rect 5092 21786 5116 21788
rect 5172 21786 5196 21788
rect 5034 21734 5036 21786
rect 5098 21734 5110 21786
rect 5172 21734 5174 21786
rect 5012 21732 5036 21734
rect 5092 21732 5116 21734
rect 5172 21732 5196 21734
rect 4956 21712 5252 21732
rect 4956 20700 5252 20720
rect 5012 20698 5036 20700
rect 5092 20698 5116 20700
rect 5172 20698 5196 20700
rect 5034 20646 5036 20698
rect 5098 20646 5110 20698
rect 5172 20646 5174 20698
rect 5012 20644 5036 20646
rect 5092 20644 5116 20646
rect 5172 20644 5196 20646
rect 4956 20624 5252 20644
rect 4956 19612 5252 19632
rect 5012 19610 5036 19612
rect 5092 19610 5116 19612
rect 5172 19610 5196 19612
rect 5034 19558 5036 19610
rect 5098 19558 5110 19610
rect 5172 19558 5174 19610
rect 5012 19556 5036 19558
rect 5092 19556 5116 19558
rect 5172 19556 5196 19558
rect 4956 19536 5252 19556
rect 4956 18524 5252 18544
rect 5012 18522 5036 18524
rect 5092 18522 5116 18524
rect 5172 18522 5196 18524
rect 5034 18470 5036 18522
rect 5098 18470 5110 18522
rect 5172 18470 5174 18522
rect 5012 18468 5036 18470
rect 5092 18468 5116 18470
rect 5172 18468 5196 18470
rect 4956 18448 5252 18468
rect 4956 17436 5252 17456
rect 5012 17434 5036 17436
rect 5092 17434 5116 17436
rect 5172 17434 5196 17436
rect 5034 17382 5036 17434
rect 5098 17382 5110 17434
rect 5172 17382 5174 17434
rect 5012 17380 5036 17382
rect 5092 17380 5116 17382
rect 5172 17380 5196 17382
rect 4956 17360 5252 17380
rect 5368 17202 5396 23582
rect 6918 23582 7052 23610
rect 6918 23520 6974 23582
rect 7024 17338 7052 23582
rect 8864 23582 8998 23610
rect 8864 20602 8892 23582
rect 8942 23520 8998 23582
rect 10874 23610 10930 24000
rect 12898 23610 12954 24000
rect 10874 23582 11192 23610
rect 10874 23520 10930 23582
rect 8956 21244 9252 21264
rect 9012 21242 9036 21244
rect 9092 21242 9116 21244
rect 9172 21242 9196 21244
rect 9034 21190 9036 21242
rect 9098 21190 9110 21242
rect 9172 21190 9174 21242
rect 9012 21188 9036 21190
rect 9092 21188 9116 21190
rect 9172 21188 9196 21190
rect 8956 21168 9252 21188
rect 8852 20596 8904 20602
rect 8852 20538 8904 20544
rect 10784 20256 10836 20262
rect 10784 20198 10836 20204
rect 8956 20156 9252 20176
rect 9012 20154 9036 20156
rect 9092 20154 9116 20156
rect 9172 20154 9196 20156
rect 9034 20102 9036 20154
rect 9098 20102 9110 20154
rect 9172 20102 9174 20154
rect 9012 20100 9036 20102
rect 9092 20100 9116 20102
rect 9172 20100 9196 20102
rect 8956 20080 9252 20100
rect 8956 19068 9252 19088
rect 9012 19066 9036 19068
rect 9092 19066 9116 19068
rect 9172 19066 9196 19068
rect 9034 19014 9036 19066
rect 9098 19014 9110 19066
rect 9172 19014 9174 19066
rect 9012 19012 9036 19014
rect 9092 19012 9116 19014
rect 9172 19012 9196 19014
rect 8956 18992 9252 19012
rect 8390 18728 8446 18737
rect 8390 18663 8446 18672
rect 7012 17332 7064 17338
rect 7012 17274 7064 17280
rect 5356 17196 5408 17202
rect 5356 17138 5408 17144
rect 8404 17134 8432 18663
rect 8956 17980 9252 18000
rect 9012 17978 9036 17980
rect 9092 17978 9116 17980
rect 9172 17978 9196 17980
rect 9034 17926 9036 17978
rect 9098 17926 9110 17978
rect 9172 17926 9174 17978
rect 9012 17924 9036 17926
rect 9092 17924 9116 17926
rect 9172 17924 9196 17926
rect 8956 17904 9252 17924
rect 8392 17128 8444 17134
rect 8392 17070 8444 17076
rect 7748 16992 7800 16998
rect 7748 16934 7800 16940
rect 8208 16992 8260 16998
rect 8208 16934 8260 16940
rect 7760 16697 7788 16934
rect 8220 16794 8248 16934
rect 8956 16892 9252 16912
rect 9012 16890 9036 16892
rect 9092 16890 9116 16892
rect 9172 16890 9196 16892
rect 9034 16838 9036 16890
rect 9098 16838 9110 16890
rect 9172 16838 9174 16890
rect 9012 16836 9036 16838
rect 9092 16836 9116 16838
rect 9172 16836 9196 16838
rect 8956 16816 9252 16836
rect 8208 16788 8260 16794
rect 8208 16730 8260 16736
rect 7746 16688 7802 16697
rect 7746 16623 7748 16632
rect 7800 16623 7802 16632
rect 7748 16594 7800 16600
rect 4956 16348 5252 16368
rect 5012 16346 5036 16348
rect 5092 16346 5116 16348
rect 5172 16346 5196 16348
rect 5034 16294 5036 16346
rect 5098 16294 5110 16346
rect 5172 16294 5174 16346
rect 5012 16292 5036 16294
rect 5092 16292 5116 16294
rect 5172 16292 5196 16294
rect 4956 16272 5252 16292
rect 7760 16250 7788 16594
rect 8116 16448 8168 16454
rect 8116 16390 8168 16396
rect 7748 16244 7800 16250
rect 7748 16186 7800 16192
rect 5356 15564 5408 15570
rect 5356 15506 5408 15512
rect 4956 15260 5252 15280
rect 5012 15258 5036 15260
rect 5092 15258 5116 15260
rect 5172 15258 5196 15260
rect 5034 15206 5036 15258
rect 5098 15206 5110 15258
rect 5172 15206 5174 15258
rect 5012 15204 5036 15206
rect 5092 15204 5116 15206
rect 5172 15204 5196 15206
rect 4956 15184 5252 15204
rect 5368 15026 5396 15506
rect 8128 15502 8156 16390
rect 8220 16114 8248 16730
rect 10796 16658 10824 20198
rect 11164 17678 11192 23582
rect 12636 23582 12954 23610
rect 11426 18864 11482 18873
rect 11426 18799 11482 18808
rect 11152 17672 11204 17678
rect 11152 17614 11204 17620
rect 10784 16652 10836 16658
rect 10784 16594 10836 16600
rect 10692 16448 10744 16454
rect 10692 16390 10744 16396
rect 8208 16108 8260 16114
rect 8208 16050 8260 16056
rect 8208 15972 8260 15978
rect 8208 15914 8260 15920
rect 9588 15972 9640 15978
rect 9588 15914 9640 15920
rect 8220 15638 8248 15914
rect 8956 15804 9252 15824
rect 9012 15802 9036 15804
rect 9092 15802 9116 15804
rect 9172 15802 9196 15804
rect 9034 15750 9036 15802
rect 9098 15750 9110 15802
rect 9172 15750 9174 15802
rect 9012 15748 9036 15750
rect 9092 15748 9116 15750
rect 9172 15748 9196 15750
rect 8956 15728 9252 15748
rect 8208 15632 8260 15638
rect 8208 15574 8260 15580
rect 8116 15496 8168 15502
rect 8116 15438 8168 15444
rect 5356 15020 5408 15026
rect 5356 14962 5408 14968
rect 6276 15020 6328 15026
rect 6276 14962 6328 14968
rect 5632 14816 5684 14822
rect 5632 14758 5684 14764
rect 5644 14414 5672 14758
rect 6288 14550 6316 14962
rect 7012 14952 7064 14958
rect 7012 14894 7064 14900
rect 6552 14816 6604 14822
rect 6552 14758 6604 14764
rect 5724 14544 5776 14550
rect 5724 14486 5776 14492
rect 6276 14544 6328 14550
rect 6276 14486 6328 14492
rect 5632 14408 5684 14414
rect 5632 14350 5684 14356
rect 4956 14172 5252 14192
rect 5012 14170 5036 14172
rect 5092 14170 5116 14172
rect 5172 14170 5196 14172
rect 5034 14118 5036 14170
rect 5098 14118 5110 14170
rect 5172 14118 5174 14170
rect 5012 14116 5036 14118
rect 5092 14116 5116 14118
rect 5172 14116 5196 14118
rect 4956 14096 5252 14116
rect 5644 14006 5672 14350
rect 5736 14074 5764 14486
rect 5724 14068 5776 14074
rect 5724 14010 5776 14016
rect 5632 14000 5684 14006
rect 5632 13942 5684 13948
rect 4988 13864 5040 13870
rect 4988 13806 5040 13812
rect 6564 13814 6592 14758
rect 7024 14278 7052 14894
rect 7840 14612 7892 14618
rect 7840 14554 7892 14560
rect 7104 14408 7156 14414
rect 7104 14350 7156 14356
rect 7012 14272 7064 14278
rect 7012 14214 7064 14220
rect 5000 13530 5028 13806
rect 6564 13802 6684 13814
rect 6564 13796 6696 13802
rect 6564 13786 6644 13796
rect 6644 13738 6696 13744
rect 4988 13524 5040 13530
rect 4988 13466 5040 13472
rect 5816 13388 5868 13394
rect 5816 13330 5868 13336
rect 6460 13388 6512 13394
rect 6460 13330 6512 13336
rect 6920 13388 6972 13394
rect 6920 13330 6972 13336
rect 4956 13084 5252 13104
rect 5012 13082 5036 13084
rect 5092 13082 5116 13084
rect 5172 13082 5196 13084
rect 5034 13030 5036 13082
rect 5098 13030 5110 13082
rect 5172 13030 5174 13082
rect 5012 13028 5036 13030
rect 5092 13028 5116 13030
rect 5172 13028 5196 13030
rect 4956 13008 5252 13028
rect 5828 12782 5856 13330
rect 6184 13184 6236 13190
rect 6184 13126 6236 13132
rect 6196 12986 6224 13126
rect 6184 12980 6236 12986
rect 6184 12922 6236 12928
rect 5816 12776 5868 12782
rect 5816 12718 5868 12724
rect 5356 12640 5408 12646
rect 5356 12582 5408 12588
rect 4956 11996 5252 12016
rect 5012 11994 5036 11996
rect 5092 11994 5116 11996
rect 5172 11994 5196 11996
rect 5034 11942 5036 11994
rect 5098 11942 5110 11994
rect 5172 11942 5174 11994
rect 5012 11940 5036 11942
rect 5092 11940 5116 11942
rect 5172 11940 5196 11942
rect 4956 11920 5252 11940
rect 5368 11898 5396 12582
rect 5724 12300 5776 12306
rect 5724 12242 5776 12248
rect 5356 11892 5408 11898
rect 5356 11834 5408 11840
rect 5736 11558 5764 12242
rect 5724 11552 5776 11558
rect 5724 11494 5776 11500
rect 5540 11348 5592 11354
rect 5540 11290 5592 11296
rect 4956 10908 5252 10928
rect 5012 10906 5036 10908
rect 5092 10906 5116 10908
rect 5172 10906 5196 10908
rect 5034 10854 5036 10906
rect 5098 10854 5110 10906
rect 5172 10854 5174 10906
rect 5012 10852 5036 10854
rect 5092 10852 5116 10854
rect 5172 10852 5196 10854
rect 4956 10832 5252 10852
rect 3332 10464 3384 10470
rect 3332 10406 3384 10412
rect 4344 10464 4396 10470
rect 4344 10406 4396 10412
rect 3344 9994 3372 10406
rect 3792 10192 3844 10198
rect 3792 10134 3844 10140
rect 3700 10124 3752 10130
rect 3700 10066 3752 10072
rect 3332 9988 3384 9994
rect 3332 9930 3384 9936
rect 3712 9722 3740 10066
rect 3804 9722 3832 10134
rect 4356 10010 4384 10406
rect 5448 10192 5500 10198
rect 5448 10134 5500 10140
rect 4080 9982 4384 10010
rect 3976 9920 4028 9926
rect 3976 9862 4028 9868
rect 3700 9716 3752 9722
rect 3700 9658 3752 9664
rect 3792 9716 3844 9722
rect 3792 9658 3844 9664
rect 3988 9450 4016 9862
rect 4080 9586 4108 9982
rect 4356 9722 4384 9982
rect 4956 9820 5252 9840
rect 5012 9818 5036 9820
rect 5092 9818 5116 9820
rect 5172 9818 5196 9820
rect 5034 9766 5036 9818
rect 5098 9766 5110 9818
rect 5172 9766 5174 9818
rect 5012 9764 5036 9766
rect 5092 9764 5116 9766
rect 5172 9764 5196 9766
rect 4956 9744 5252 9764
rect 4344 9716 4396 9722
rect 4344 9658 4396 9664
rect 4068 9580 4120 9586
rect 4068 9522 4120 9528
rect 5460 9450 5488 10134
rect 5552 10130 5580 11290
rect 5736 11218 5764 11494
rect 6196 11218 6224 12922
rect 6472 12306 6500 13330
rect 6552 12640 6604 12646
rect 6552 12582 6604 12588
rect 6276 12300 6328 12306
rect 6276 12242 6328 12248
rect 6460 12300 6512 12306
rect 6460 12242 6512 12248
rect 6288 11558 6316 12242
rect 6472 11694 6500 12242
rect 6460 11688 6512 11694
rect 6460 11630 6512 11636
rect 6276 11552 6328 11558
rect 6276 11494 6328 11500
rect 5724 11212 5776 11218
rect 5724 11154 5776 11160
rect 6184 11212 6236 11218
rect 6184 11154 6236 11160
rect 5736 10606 5764 11154
rect 6196 10742 6224 11154
rect 6184 10736 6236 10742
rect 6184 10678 6236 10684
rect 5724 10600 5776 10606
rect 5724 10542 5776 10548
rect 5736 10130 5764 10542
rect 6196 10198 6224 10678
rect 6288 10538 6316 11494
rect 6472 11218 6500 11630
rect 6460 11212 6512 11218
rect 6460 11154 6512 11160
rect 6472 10742 6500 11154
rect 6564 10742 6592 12582
rect 6932 12374 6960 13330
rect 7024 12442 7052 14214
rect 7116 13734 7144 14350
rect 7852 13802 7880 14554
rect 8128 14550 8156 15438
rect 8220 15162 8248 15574
rect 9600 15502 9628 15914
rect 10704 15706 10732 16390
rect 10796 15978 10824 16594
rect 11440 16046 11468 18799
rect 11428 16040 11480 16046
rect 11428 15982 11480 15988
rect 10784 15972 10836 15978
rect 10784 15914 10836 15920
rect 11440 15910 11468 15982
rect 11336 15904 11388 15910
rect 11336 15846 11388 15852
rect 11428 15904 11480 15910
rect 11428 15846 11480 15852
rect 10692 15700 10744 15706
rect 10692 15642 10744 15648
rect 9772 15632 9824 15638
rect 9772 15574 9824 15580
rect 8852 15496 8904 15502
rect 8852 15438 8904 15444
rect 9588 15496 9640 15502
rect 9588 15438 9640 15444
rect 8208 15156 8260 15162
rect 8208 15098 8260 15104
rect 8864 14890 8892 15438
rect 9600 15162 9628 15438
rect 9588 15156 9640 15162
rect 9588 15098 9640 15104
rect 8852 14884 8904 14890
rect 8852 14826 8904 14832
rect 8760 14816 8812 14822
rect 8760 14758 8812 14764
rect 8116 14544 8168 14550
rect 8116 14486 8168 14492
rect 8772 14074 8800 14758
rect 8864 14346 8892 14826
rect 9784 14822 9812 15574
rect 10048 15496 10100 15502
rect 10048 15438 10100 15444
rect 10060 15026 10088 15438
rect 10704 15026 10732 15642
rect 11348 15502 11376 15846
rect 11428 15632 11480 15638
rect 11428 15574 11480 15580
rect 11336 15496 11388 15502
rect 11336 15438 11388 15444
rect 10048 15020 10100 15026
rect 10048 14962 10100 14968
rect 10692 15020 10744 15026
rect 10692 14962 10744 14968
rect 11244 14884 11296 14890
rect 11244 14826 11296 14832
rect 9772 14816 9824 14822
rect 9772 14758 9824 14764
rect 8956 14716 9252 14736
rect 9012 14714 9036 14716
rect 9092 14714 9116 14716
rect 9172 14714 9196 14716
rect 9034 14662 9036 14714
rect 9098 14662 9110 14714
rect 9172 14662 9174 14714
rect 9012 14660 9036 14662
rect 9092 14660 9116 14662
rect 9172 14660 9196 14662
rect 8956 14640 9252 14660
rect 9784 14618 9812 14758
rect 9772 14612 9824 14618
rect 9772 14554 9824 14560
rect 11256 14550 11284 14826
rect 11348 14618 11376 15438
rect 11440 15162 11468 15574
rect 11796 15496 11848 15502
rect 11796 15438 11848 15444
rect 11428 15156 11480 15162
rect 11428 15098 11480 15104
rect 11336 14612 11388 14618
rect 11336 14554 11388 14560
rect 11244 14544 11296 14550
rect 11244 14486 11296 14492
rect 10048 14476 10100 14482
rect 10048 14418 10100 14424
rect 8852 14340 8904 14346
rect 8852 14282 8904 14288
rect 8760 14068 8812 14074
rect 8760 14010 8812 14016
rect 10060 13938 10088 14418
rect 10600 14272 10652 14278
rect 10600 14214 10652 14220
rect 10612 13938 10640 14214
rect 11256 14006 11284 14486
rect 11440 14074 11468 15098
rect 11808 14550 11836 15438
rect 12532 15360 12584 15366
rect 12532 15302 12584 15308
rect 12544 15026 12572 15302
rect 12532 15020 12584 15026
rect 12532 14962 12584 14968
rect 12544 14618 12572 14962
rect 12532 14612 12584 14618
rect 12532 14554 12584 14560
rect 11796 14544 11848 14550
rect 11796 14486 11848 14492
rect 11808 14346 11836 14486
rect 12164 14408 12216 14414
rect 12164 14350 12216 14356
rect 11796 14340 11848 14346
rect 11796 14282 11848 14288
rect 12176 14074 12204 14350
rect 11428 14068 11480 14074
rect 11428 14010 11480 14016
rect 12164 14068 12216 14074
rect 12164 14010 12216 14016
rect 11244 14000 11296 14006
rect 11244 13942 11296 13948
rect 9404 13932 9456 13938
rect 9404 13874 9456 13880
rect 10048 13932 10100 13938
rect 10048 13874 10100 13880
rect 10600 13932 10652 13938
rect 10600 13874 10652 13880
rect 8300 13864 8352 13870
rect 8300 13806 8352 13812
rect 7840 13796 7892 13802
rect 7840 13738 7892 13744
rect 7104 13728 7156 13734
rect 7104 13670 7156 13676
rect 7116 12646 7144 13670
rect 8312 13190 8340 13806
rect 8956 13628 9252 13648
rect 9012 13626 9036 13628
rect 9092 13626 9116 13628
rect 9172 13626 9196 13628
rect 9034 13574 9036 13626
rect 9098 13574 9110 13626
rect 9172 13574 9174 13626
rect 9012 13572 9036 13574
rect 9092 13572 9116 13574
rect 9172 13572 9196 13574
rect 8956 13552 9252 13572
rect 7380 13184 7432 13190
rect 7380 13126 7432 13132
rect 8300 13184 8352 13190
rect 8300 13126 8352 13132
rect 7392 12850 7420 13126
rect 7380 12844 7432 12850
rect 7380 12786 7432 12792
rect 8208 12776 8260 12782
rect 8208 12718 8260 12724
rect 7104 12640 7156 12646
rect 7104 12582 7156 12588
rect 7012 12436 7064 12442
rect 7012 12378 7064 12384
rect 8220 12374 8248 12718
rect 6920 12368 6972 12374
rect 6920 12310 6972 12316
rect 8208 12368 8260 12374
rect 8208 12310 8260 12316
rect 6932 11898 6960 12310
rect 8116 12096 8168 12102
rect 8116 12038 8168 12044
rect 6920 11892 6972 11898
rect 6920 11834 6972 11840
rect 7840 11756 7892 11762
rect 7840 11698 7892 11704
rect 7852 11558 7880 11698
rect 8128 11626 8156 12038
rect 8208 11824 8260 11830
rect 8208 11766 8260 11772
rect 8220 11694 8248 11766
rect 8208 11688 8260 11694
rect 8208 11630 8260 11636
rect 8116 11620 8168 11626
rect 8116 11562 8168 11568
rect 7840 11552 7892 11558
rect 7840 11494 7892 11500
rect 6644 11212 6696 11218
rect 6644 11154 6696 11160
rect 6656 10810 6684 11154
rect 6644 10804 6696 10810
rect 6644 10746 6696 10752
rect 6460 10736 6512 10742
rect 6460 10678 6512 10684
rect 6552 10736 6604 10742
rect 6552 10678 6604 10684
rect 6276 10532 6328 10538
rect 6276 10474 6328 10480
rect 5908 10192 5960 10198
rect 5908 10134 5960 10140
rect 6184 10192 6236 10198
rect 6184 10134 6236 10140
rect 5540 10124 5592 10130
rect 5540 10066 5592 10072
rect 5724 10124 5776 10130
rect 5724 10066 5776 10072
rect 3976 9444 4028 9450
rect 3976 9386 4028 9392
rect 4804 9444 4856 9450
rect 4804 9386 4856 9392
rect 5448 9444 5500 9450
rect 5448 9386 5500 9392
rect 4816 9178 4844 9386
rect 5920 9178 5948 10134
rect 6564 10130 6592 10678
rect 6276 10124 6328 10130
rect 6276 10066 6328 10072
rect 6552 10124 6604 10130
rect 6552 10066 6604 10072
rect 6656 10112 6684 10746
rect 7852 10538 7880 11494
rect 8024 11280 8076 11286
rect 8024 11222 8076 11228
rect 7932 11008 7984 11014
rect 7932 10950 7984 10956
rect 7840 10532 7892 10538
rect 7840 10474 7892 10480
rect 7944 10470 7972 10950
rect 7932 10464 7984 10470
rect 7932 10406 7984 10412
rect 8036 10266 8064 11222
rect 8128 10606 8156 11562
rect 8220 10656 8248 11630
rect 8312 11558 8340 13126
rect 8956 12540 9252 12560
rect 9012 12538 9036 12540
rect 9092 12538 9116 12540
rect 9172 12538 9196 12540
rect 9034 12486 9036 12538
rect 9098 12486 9110 12538
rect 9172 12486 9174 12538
rect 9012 12484 9036 12486
rect 9092 12484 9116 12486
rect 9172 12484 9196 12486
rect 8956 12464 9252 12484
rect 8300 11552 8352 11558
rect 8300 11494 8352 11500
rect 8956 11452 9252 11472
rect 9012 11450 9036 11452
rect 9092 11450 9116 11452
rect 9172 11450 9196 11452
rect 9034 11398 9036 11450
rect 9098 11398 9110 11450
rect 9172 11398 9174 11450
rect 9012 11396 9036 11398
rect 9092 11396 9116 11398
rect 9172 11396 9196 11398
rect 8956 11376 9252 11396
rect 8852 11144 8904 11150
rect 8852 11086 8904 11092
rect 8760 11008 8812 11014
rect 8760 10950 8812 10956
rect 8300 10668 8352 10674
rect 8220 10628 8300 10656
rect 8300 10610 8352 10616
rect 8116 10600 8168 10606
rect 8116 10542 8168 10548
rect 8024 10260 8076 10266
rect 7944 10220 8024 10248
rect 6736 10124 6788 10130
rect 6656 10084 6736 10112
rect 6288 9382 6316 10066
rect 6564 9722 6592 10066
rect 6552 9716 6604 9722
rect 6552 9658 6604 9664
rect 6276 9376 6328 9382
rect 6276 9318 6328 9324
rect 6552 9376 6604 9382
rect 6552 9318 6604 9324
rect 4804 9172 4856 9178
rect 4804 9114 4856 9120
rect 5908 9172 5960 9178
rect 5908 9114 5960 9120
rect 4956 8732 5252 8752
rect 5012 8730 5036 8732
rect 5092 8730 5116 8732
rect 5172 8730 5196 8732
rect 5034 8678 5036 8730
rect 5098 8678 5110 8730
rect 5172 8678 5174 8730
rect 5012 8676 5036 8678
rect 5092 8676 5116 8678
rect 5172 8676 5196 8678
rect 4956 8656 5252 8676
rect 2780 8424 2832 8430
rect 2780 8366 2832 8372
rect 2044 8288 2096 8294
rect 2044 8230 2096 8236
rect 1676 8084 1728 8090
rect 1676 8026 1728 8032
rect 2056 7993 2084 8230
rect 2042 7984 2098 7993
rect 2042 7919 2098 7928
rect 4956 7644 5252 7664
rect 5012 7642 5036 7644
rect 5092 7642 5116 7644
rect 5172 7642 5196 7644
rect 5034 7590 5036 7642
rect 5098 7590 5110 7642
rect 5172 7590 5174 7642
rect 5012 7588 5036 7590
rect 5092 7588 5116 7590
rect 5172 7588 5196 7590
rect 4956 7568 5252 7588
rect 6288 7342 6316 9318
rect 6564 8004 6592 9318
rect 6656 9178 6684 10084
rect 6736 10066 6788 10072
rect 7196 9988 7248 9994
rect 7196 9930 7248 9936
rect 7208 9586 7236 9930
rect 7196 9580 7248 9586
rect 7196 9522 7248 9528
rect 7208 9178 7236 9522
rect 7944 9450 7972 10220
rect 8024 10202 8076 10208
rect 8312 9926 8340 10610
rect 8300 9920 8352 9926
rect 8300 9862 8352 9868
rect 8024 9648 8076 9654
rect 8024 9590 8076 9596
rect 7932 9444 7984 9450
rect 7932 9386 7984 9392
rect 7840 9376 7892 9382
rect 7840 9318 7892 9324
rect 6644 9172 6696 9178
rect 6644 9114 6696 9120
rect 7196 9172 7248 9178
rect 7196 9114 7248 9120
rect 7852 9110 7880 9318
rect 7840 9104 7892 9110
rect 7840 9046 7892 9052
rect 7748 8968 7800 8974
rect 7748 8910 7800 8916
rect 7760 8022 7788 8910
rect 7852 8634 7880 9046
rect 8036 8974 8064 9590
rect 8024 8968 8076 8974
rect 8024 8910 8076 8916
rect 7840 8628 7892 8634
rect 7840 8570 7892 8576
rect 8024 8356 8076 8362
rect 8024 8298 8076 8304
rect 6644 8016 6696 8022
rect 6564 7976 6644 8004
rect 6644 7958 6696 7964
rect 7748 8016 7800 8022
rect 7748 7958 7800 7964
rect 6276 7336 6328 7342
rect 6276 7278 6328 7284
rect 6656 7206 6684 7958
rect 6736 7880 6788 7886
rect 6736 7822 6788 7828
rect 6748 7206 6776 7822
rect 7288 7812 7340 7818
rect 7288 7754 7340 7760
rect 7300 7342 7328 7754
rect 7288 7336 7340 7342
rect 7288 7278 7340 7284
rect 7656 7336 7708 7342
rect 7656 7278 7708 7284
rect 3056 7200 3108 7206
rect 3056 7142 3108 7148
rect 6644 7200 6696 7206
rect 6644 7142 6696 7148
rect 6736 7200 6788 7206
rect 6736 7142 6788 7148
rect 112 5092 164 5098
rect 112 5034 164 5040
rect 124 3913 152 5034
rect 1216 4684 1268 4690
rect 1216 4626 1268 4632
rect 110 3904 166 3913
rect 110 3839 166 3848
rect 938 82 994 480
rect 1228 82 1256 4626
rect 938 54 1256 82
rect 2778 82 2834 480
rect 3068 82 3096 7142
rect 7300 6730 7328 7278
rect 7668 6866 7696 7278
rect 7656 6860 7708 6866
rect 7656 6802 7708 6808
rect 7288 6724 7340 6730
rect 7288 6666 7340 6672
rect 4804 6656 4856 6662
rect 4804 6598 4856 6604
rect 2778 54 3096 82
rect 4618 82 4674 480
rect 4816 82 4844 6598
rect 4956 6556 5252 6576
rect 5012 6554 5036 6556
rect 5092 6554 5116 6556
rect 5172 6554 5196 6556
rect 5034 6502 5036 6554
rect 5098 6502 5110 6554
rect 5172 6502 5174 6554
rect 5012 6500 5036 6502
rect 5092 6500 5116 6502
rect 5172 6500 5196 6502
rect 4956 6480 5252 6500
rect 4956 5468 5252 5488
rect 5012 5466 5036 5468
rect 5092 5466 5116 5468
rect 5172 5466 5196 5468
rect 5034 5414 5036 5466
rect 5098 5414 5110 5466
rect 5172 5414 5174 5466
rect 5012 5412 5036 5414
rect 5092 5412 5116 5414
rect 5172 5412 5196 5414
rect 4956 5392 5252 5412
rect 7668 5234 7696 6802
rect 7656 5228 7708 5234
rect 7656 5170 7708 5176
rect 6552 5160 6604 5166
rect 6552 5102 6604 5108
rect 6564 5030 6592 5102
rect 6552 5024 6604 5030
rect 6552 4966 6604 4972
rect 4956 4380 5252 4400
rect 5012 4378 5036 4380
rect 5092 4378 5116 4380
rect 5172 4378 5196 4380
rect 5034 4326 5036 4378
rect 5098 4326 5110 4378
rect 5172 4326 5174 4378
rect 5012 4324 5036 4326
rect 5092 4324 5116 4326
rect 5172 4324 5196 4326
rect 4956 4304 5252 4324
rect 4956 3292 5252 3312
rect 5012 3290 5036 3292
rect 5092 3290 5116 3292
rect 5172 3290 5196 3292
rect 5034 3238 5036 3290
rect 5098 3238 5110 3290
rect 5172 3238 5174 3290
rect 5012 3236 5036 3238
rect 5092 3236 5116 3238
rect 5172 3236 5196 3238
rect 4956 3216 5252 3236
rect 4956 2204 5252 2224
rect 5012 2202 5036 2204
rect 5092 2202 5116 2204
rect 5172 2202 5196 2204
rect 5034 2150 5036 2202
rect 5098 2150 5110 2202
rect 5172 2150 5174 2202
rect 5012 2148 5036 2150
rect 5092 2148 5116 2150
rect 5172 2148 5196 2150
rect 4956 2128 5252 2148
rect 6564 1873 6592 4966
rect 6736 2304 6788 2310
rect 6736 2246 6788 2252
rect 6550 1864 6606 1873
rect 6550 1799 6606 1808
rect 4618 54 4844 82
rect 6458 82 6514 480
rect 6748 82 6776 2246
rect 8036 2009 8064 8298
rect 8116 8288 8168 8294
rect 8116 8230 8168 8236
rect 8128 8090 8156 8230
rect 8116 8084 8168 8090
rect 8116 8026 8168 8032
rect 8312 7478 8340 9862
rect 8772 9450 8800 10950
rect 8864 10606 8892 11086
rect 8852 10600 8904 10606
rect 8852 10542 8904 10548
rect 8864 10130 8892 10542
rect 8956 10364 9252 10384
rect 9012 10362 9036 10364
rect 9092 10362 9116 10364
rect 9172 10362 9196 10364
rect 9034 10310 9036 10362
rect 9098 10310 9110 10362
rect 9172 10310 9174 10362
rect 9012 10308 9036 10310
rect 9092 10308 9116 10310
rect 9172 10308 9196 10310
rect 8956 10288 9252 10308
rect 8852 10124 8904 10130
rect 8852 10066 8904 10072
rect 8864 9722 8892 10066
rect 8852 9716 8904 9722
rect 8852 9658 8904 9664
rect 8668 9444 8720 9450
rect 8668 9386 8720 9392
rect 8760 9444 8812 9450
rect 8760 9386 8812 9392
rect 8680 8566 8708 9386
rect 8956 9276 9252 9296
rect 9012 9274 9036 9276
rect 9092 9274 9116 9276
rect 9172 9274 9196 9276
rect 9034 9222 9036 9274
rect 9098 9222 9110 9274
rect 9172 9222 9174 9274
rect 9012 9220 9036 9222
rect 9092 9220 9116 9222
rect 9172 9220 9196 9222
rect 8956 9200 9252 9220
rect 8668 8560 8720 8566
rect 8668 8502 8720 8508
rect 8392 8356 8444 8362
rect 8392 8298 8444 8304
rect 8404 7750 8432 8298
rect 8956 8188 9252 8208
rect 9012 8186 9036 8188
rect 9092 8186 9116 8188
rect 9172 8186 9196 8188
rect 9034 8134 9036 8186
rect 9098 8134 9110 8186
rect 9172 8134 9174 8186
rect 9012 8132 9036 8134
rect 9092 8132 9116 8134
rect 9172 8132 9196 8134
rect 8956 8112 9252 8132
rect 8392 7744 8444 7750
rect 8392 7686 8444 7692
rect 8668 7744 8720 7750
rect 8668 7686 8720 7692
rect 8300 7472 8352 7478
rect 8300 7414 8352 7420
rect 8208 7336 8260 7342
rect 8208 7278 8260 7284
rect 8220 7002 8248 7278
rect 8404 7002 8432 7686
rect 8680 7313 8708 7686
rect 9312 7472 9364 7478
rect 9312 7414 9364 7420
rect 8666 7304 8722 7313
rect 8666 7239 8722 7248
rect 8680 7206 8708 7239
rect 9324 7206 9352 7414
rect 8668 7200 8720 7206
rect 8668 7142 8720 7148
rect 8852 7200 8904 7206
rect 8852 7142 8904 7148
rect 9312 7200 9364 7206
rect 9312 7142 9364 7148
rect 8208 6996 8260 7002
rect 8208 6938 8260 6944
rect 8392 6996 8444 7002
rect 8392 6938 8444 6944
rect 8680 4154 8708 7142
rect 8864 6390 8892 7142
rect 8956 7100 9252 7120
rect 9012 7098 9036 7100
rect 9092 7098 9116 7100
rect 9172 7098 9196 7100
rect 9034 7046 9036 7098
rect 9098 7046 9110 7098
rect 9172 7046 9174 7098
rect 9012 7044 9036 7046
rect 9092 7044 9116 7046
rect 9172 7044 9196 7046
rect 8956 7024 9252 7044
rect 8852 6384 8904 6390
rect 8852 6326 8904 6332
rect 8864 5166 8892 6326
rect 9312 6180 9364 6186
rect 9312 6122 9364 6128
rect 8956 6012 9252 6032
rect 9012 6010 9036 6012
rect 9092 6010 9116 6012
rect 9172 6010 9196 6012
rect 9034 5958 9036 6010
rect 9098 5958 9110 6010
rect 9172 5958 9174 6010
rect 9012 5956 9036 5958
rect 9092 5956 9116 5958
rect 9172 5956 9196 5958
rect 8956 5936 9252 5956
rect 9324 5778 9352 6122
rect 9312 5772 9364 5778
rect 9312 5714 9364 5720
rect 8852 5160 8904 5166
rect 8852 5102 8904 5108
rect 8956 4924 9252 4944
rect 9012 4922 9036 4924
rect 9092 4922 9116 4924
rect 9172 4922 9196 4924
rect 9034 4870 9036 4922
rect 9098 4870 9110 4922
rect 9172 4870 9174 4922
rect 9012 4868 9036 4870
rect 9092 4868 9116 4870
rect 9172 4868 9196 4870
rect 8956 4848 9252 4868
rect 9416 4185 9444 13874
rect 10508 13728 10560 13734
rect 10508 13670 10560 13676
rect 10520 13462 10548 13670
rect 10508 13456 10560 13462
rect 10508 13398 10560 13404
rect 10508 13320 10560 13326
rect 10508 13262 10560 13268
rect 10140 13184 10192 13190
rect 10140 13126 10192 13132
rect 10048 12980 10100 12986
rect 10048 12922 10100 12928
rect 10060 12782 10088 12922
rect 10152 12782 10180 13126
rect 10520 12850 10548 13262
rect 10508 12844 10560 12850
rect 10508 12786 10560 12792
rect 10048 12776 10100 12782
rect 10048 12718 10100 12724
rect 10140 12776 10192 12782
rect 10140 12718 10192 12724
rect 9772 12708 9824 12714
rect 9772 12650 9824 12656
rect 9496 12640 9548 12646
rect 9496 12582 9548 12588
rect 9508 12374 9536 12582
rect 9496 12368 9548 12374
rect 9496 12310 9548 12316
rect 9508 11762 9536 12310
rect 9784 11898 9812 12650
rect 10060 12102 10088 12718
rect 10152 12238 10180 12718
rect 10612 12442 10640 13874
rect 11256 13530 11284 13942
rect 11244 13524 11296 13530
rect 11244 13466 11296 13472
rect 11704 13456 11756 13462
rect 11704 13398 11756 13404
rect 11336 12776 11388 12782
rect 11336 12718 11388 12724
rect 10600 12436 10652 12442
rect 10600 12378 10652 12384
rect 11348 12306 11376 12718
rect 11716 12646 11744 13398
rect 11704 12640 11756 12646
rect 11704 12582 11756 12588
rect 10324 12300 10376 12306
rect 10324 12242 10376 12248
rect 11336 12300 11388 12306
rect 11336 12242 11388 12248
rect 10140 12232 10192 12238
rect 10140 12174 10192 12180
rect 10048 12096 10100 12102
rect 10048 12038 10100 12044
rect 9772 11892 9824 11898
rect 9772 11834 9824 11840
rect 9496 11756 9548 11762
rect 9496 11698 9548 11704
rect 10060 11694 10088 12038
rect 9588 11688 9640 11694
rect 9588 11630 9640 11636
rect 10048 11688 10100 11694
rect 10048 11630 10100 11636
rect 9496 11620 9548 11626
rect 9496 11562 9548 11568
rect 9508 11218 9536 11562
rect 9496 11212 9548 11218
rect 9496 11154 9548 11160
rect 9508 10266 9536 11154
rect 9496 10260 9548 10266
rect 9496 10202 9548 10208
rect 9496 7336 9548 7342
rect 9600 7324 9628 11630
rect 10152 11558 10180 12174
rect 10140 11552 10192 11558
rect 10140 11494 10192 11500
rect 10048 11348 10100 11354
rect 10048 11290 10100 11296
rect 9956 11280 10008 11286
rect 9956 11222 10008 11228
rect 9680 10532 9732 10538
rect 9968 10520 9996 11222
rect 10060 10674 10088 11290
rect 10152 11218 10180 11494
rect 10336 11286 10364 12242
rect 10600 12232 10652 12238
rect 10600 12174 10652 12180
rect 10612 11898 10640 12174
rect 10600 11892 10652 11898
rect 10600 11834 10652 11840
rect 10324 11280 10376 11286
rect 10324 11222 10376 11228
rect 10612 11218 10640 11834
rect 10140 11212 10192 11218
rect 10140 11154 10192 11160
rect 10600 11212 10652 11218
rect 10600 11154 10652 11160
rect 10048 10668 10100 10674
rect 10048 10610 10100 10616
rect 10152 10606 10180 11154
rect 10140 10600 10192 10606
rect 10140 10542 10192 10548
rect 10048 10532 10100 10538
rect 9968 10492 10048 10520
rect 9680 10474 9732 10480
rect 10048 10474 10100 10480
rect 9692 9926 9720 10474
rect 9680 9920 9732 9926
rect 9680 9862 9732 9868
rect 9692 7750 9720 9862
rect 9772 9716 9824 9722
rect 9772 9658 9824 9664
rect 9680 7744 9732 7750
rect 9680 7686 9732 7692
rect 9692 7342 9720 7686
rect 9784 7546 9812 9658
rect 10060 8090 10088 10474
rect 11152 10464 11204 10470
rect 11152 10406 11204 10412
rect 11164 10198 11192 10406
rect 10600 10192 10652 10198
rect 10600 10134 10652 10140
rect 11152 10192 11204 10198
rect 11152 10134 11204 10140
rect 10232 10056 10284 10062
rect 10232 9998 10284 10004
rect 10140 9648 10192 9654
rect 10140 9590 10192 9596
rect 10152 9110 10180 9590
rect 10244 9110 10272 9998
rect 10612 9722 10640 10134
rect 11152 9920 11204 9926
rect 11152 9862 11204 9868
rect 10600 9716 10652 9722
rect 11164 9674 11192 9862
rect 10600 9658 10652 9664
rect 10612 9382 10640 9658
rect 10888 9646 11192 9674
rect 10888 9450 10916 9646
rect 10876 9444 10928 9450
rect 10876 9386 10928 9392
rect 11244 9444 11296 9450
rect 11244 9386 11296 9392
rect 10600 9376 10652 9382
rect 10600 9318 10652 9324
rect 10888 9178 10916 9386
rect 10876 9172 10928 9178
rect 10876 9114 10928 9120
rect 10140 9104 10192 9110
rect 10140 9046 10192 9052
rect 10232 9104 10284 9110
rect 10232 9046 10284 9052
rect 11060 9104 11112 9110
rect 11060 9046 11112 9052
rect 10152 8634 10180 9046
rect 10968 8968 11020 8974
rect 10968 8910 11020 8916
rect 10416 8900 10468 8906
rect 10416 8842 10468 8848
rect 10140 8628 10192 8634
rect 10192 8588 10272 8616
rect 10140 8570 10192 8576
rect 10048 8084 10100 8090
rect 10048 8026 10100 8032
rect 9772 7540 9824 7546
rect 9772 7482 9824 7488
rect 9548 7296 9628 7324
rect 9680 7336 9732 7342
rect 9496 7278 9548 7284
rect 9680 7278 9732 7284
rect 9508 7002 9536 7278
rect 10060 7002 10088 8026
rect 9496 6996 9548 7002
rect 9496 6938 9548 6944
rect 10048 6996 10100 7002
rect 10048 6938 10100 6944
rect 9588 6928 9640 6934
rect 9588 6870 9640 6876
rect 9600 6118 9628 6870
rect 10048 6792 10100 6798
rect 10048 6734 10100 6740
rect 9772 6724 9824 6730
rect 9772 6666 9824 6672
rect 9784 6322 9812 6666
rect 9772 6316 9824 6322
rect 9772 6258 9824 6264
rect 10060 6225 10088 6734
rect 10046 6216 10102 6225
rect 10046 6151 10102 6160
rect 10060 6118 10088 6151
rect 9588 6112 9640 6118
rect 9588 6054 9640 6060
rect 10048 6112 10100 6118
rect 10048 6054 10100 6060
rect 9600 4214 9628 6054
rect 9864 5772 9916 5778
rect 9864 5714 9916 5720
rect 9876 5370 9904 5714
rect 10060 5692 10088 6054
rect 10140 5704 10192 5710
rect 10060 5664 10140 5692
rect 10140 5646 10192 5652
rect 9864 5364 9916 5370
rect 9864 5306 9916 5312
rect 9876 4826 9904 5306
rect 9864 4820 9916 4826
rect 9864 4762 9916 4768
rect 9680 4684 9732 4690
rect 9680 4626 9732 4632
rect 9692 4282 9720 4626
rect 9680 4276 9732 4282
rect 9680 4218 9732 4224
rect 9588 4208 9640 4214
rect 8588 4126 8708 4154
rect 9402 4176 9458 4185
rect 8022 2000 8078 2009
rect 8022 1935 8078 1944
rect 6458 54 6776 82
rect 8298 82 8354 480
rect 8588 82 8616 4126
rect 9588 4150 9640 4156
rect 9772 4208 9824 4214
rect 9772 4150 9824 4156
rect 10244 4154 10272 8588
rect 10428 8362 10456 8842
rect 10692 8832 10744 8838
rect 10692 8774 10744 8780
rect 10704 8498 10732 8774
rect 10980 8634 11008 8910
rect 10968 8628 11020 8634
rect 10968 8570 11020 8576
rect 10692 8492 10744 8498
rect 10692 8434 10744 8440
rect 10416 8356 10468 8362
rect 10416 8298 10468 8304
rect 10428 8022 10456 8298
rect 11072 8294 11100 9046
rect 11256 8974 11284 9386
rect 11244 8968 11296 8974
rect 11244 8910 11296 8916
rect 11060 8288 11112 8294
rect 11060 8230 11112 8236
rect 10416 8016 10468 8022
rect 10416 7958 10468 7964
rect 10876 7744 10928 7750
rect 10876 7686 10928 7692
rect 10888 7410 10916 7686
rect 11060 7540 11112 7546
rect 11060 7482 11112 7488
rect 10876 7404 10928 7410
rect 10876 7346 10928 7352
rect 11072 7002 11100 7482
rect 11060 6996 11112 7002
rect 11060 6938 11112 6944
rect 10416 6860 10468 6866
rect 10416 6802 10468 6808
rect 10428 5778 10456 6802
rect 10600 6656 10652 6662
rect 10600 6598 10652 6604
rect 10692 6656 10744 6662
rect 10692 6598 10744 6604
rect 10612 6322 10640 6598
rect 10704 6458 10732 6598
rect 10692 6452 10744 6458
rect 10692 6394 10744 6400
rect 10600 6316 10652 6322
rect 10600 6258 10652 6264
rect 10416 5772 10468 5778
rect 10416 5714 10468 5720
rect 10416 5568 10468 5574
rect 10416 5510 10468 5516
rect 10428 5166 10456 5510
rect 10704 5370 10732 6394
rect 11244 6248 11296 6254
rect 11244 6190 11296 6196
rect 10876 5704 10928 5710
rect 10876 5646 10928 5652
rect 10692 5364 10744 5370
rect 10692 5306 10744 5312
rect 10888 5302 10916 5646
rect 11256 5642 11284 6190
rect 11348 5846 11376 12242
rect 11520 11688 11572 11694
rect 11520 11630 11572 11636
rect 11532 11286 11560 11630
rect 11520 11280 11572 11286
rect 11520 11222 11572 11228
rect 11716 10470 11744 12582
rect 12440 12096 12492 12102
rect 12440 12038 12492 12044
rect 12348 11552 12400 11558
rect 12348 11494 12400 11500
rect 12360 11014 12388 11494
rect 12452 11082 12480 12038
rect 12440 11076 12492 11082
rect 12440 11018 12492 11024
rect 12348 11008 12400 11014
rect 12348 10950 12400 10956
rect 12360 10538 12388 10950
rect 12348 10532 12400 10538
rect 12348 10474 12400 10480
rect 11704 10464 11756 10470
rect 11704 10406 11756 10412
rect 12360 10130 12388 10474
rect 12348 10124 12400 10130
rect 12348 10066 12400 10072
rect 11888 10056 11940 10062
rect 11888 9998 11940 10004
rect 11900 8566 11928 9998
rect 12360 9722 12388 10066
rect 12348 9716 12400 9722
rect 12348 9658 12400 9664
rect 11888 8560 11940 8566
rect 11888 8502 11940 8508
rect 11520 8288 11572 8294
rect 11520 8230 11572 8236
rect 11532 8022 11560 8230
rect 11520 8016 11572 8022
rect 11520 7958 11572 7964
rect 11532 7546 11560 7958
rect 11900 7886 11928 8502
rect 12636 8498 12664 23582
rect 12898 23520 12954 23582
rect 13912 23588 13964 23594
rect 13912 23530 13964 23536
rect 14922 23588 14978 24000
rect 16946 23610 17002 24000
rect 18878 23610 18934 24000
rect 20902 23610 20958 24000
rect 22926 23610 22982 24000
rect 14922 23536 14924 23588
rect 14976 23536 14978 23588
rect 12956 21788 13252 21808
rect 13012 21786 13036 21788
rect 13092 21786 13116 21788
rect 13172 21786 13196 21788
rect 13034 21734 13036 21786
rect 13098 21734 13110 21786
rect 13172 21734 13174 21786
rect 13012 21732 13036 21734
rect 13092 21732 13116 21734
rect 13172 21732 13196 21734
rect 12956 21712 13252 21732
rect 12956 20700 13252 20720
rect 13012 20698 13036 20700
rect 13092 20698 13116 20700
rect 13172 20698 13196 20700
rect 13034 20646 13036 20698
rect 13098 20646 13110 20698
rect 13172 20646 13174 20698
rect 13012 20644 13036 20646
rect 13092 20644 13116 20646
rect 13172 20644 13196 20646
rect 12956 20624 13252 20644
rect 12956 19612 13252 19632
rect 13012 19610 13036 19612
rect 13092 19610 13116 19612
rect 13172 19610 13196 19612
rect 13034 19558 13036 19610
rect 13098 19558 13110 19610
rect 13172 19558 13174 19610
rect 13012 19556 13036 19558
rect 13092 19556 13116 19558
rect 13172 19556 13196 19558
rect 12956 19536 13252 19556
rect 12956 18524 13252 18544
rect 13012 18522 13036 18524
rect 13092 18522 13116 18524
rect 13172 18522 13196 18524
rect 13034 18470 13036 18522
rect 13098 18470 13110 18522
rect 13172 18470 13174 18522
rect 13012 18468 13036 18470
rect 13092 18468 13116 18470
rect 13172 18468 13196 18470
rect 12956 18448 13252 18468
rect 12956 17436 13252 17456
rect 13012 17434 13036 17436
rect 13092 17434 13116 17436
rect 13172 17434 13196 17436
rect 13034 17382 13036 17434
rect 13098 17382 13110 17434
rect 13172 17382 13174 17434
rect 13012 17380 13036 17382
rect 13092 17380 13116 17382
rect 13172 17380 13196 17382
rect 12956 17360 13252 17380
rect 12956 16348 13252 16368
rect 13012 16346 13036 16348
rect 13092 16346 13116 16348
rect 13172 16346 13196 16348
rect 13034 16294 13036 16346
rect 13098 16294 13110 16346
rect 13172 16294 13174 16346
rect 13012 16292 13036 16294
rect 13092 16292 13116 16294
rect 13172 16292 13196 16294
rect 12956 16272 13252 16292
rect 13544 15564 13596 15570
rect 13544 15506 13596 15512
rect 12956 15260 13252 15280
rect 13012 15258 13036 15260
rect 13092 15258 13116 15260
rect 13172 15258 13196 15260
rect 13034 15206 13036 15258
rect 13098 15206 13110 15258
rect 13172 15206 13174 15258
rect 13012 15204 13036 15206
rect 13092 15204 13116 15206
rect 13172 15204 13196 15206
rect 12956 15184 13252 15204
rect 13556 15094 13584 15506
rect 13544 15088 13596 15094
rect 13544 15030 13596 15036
rect 13556 14822 13584 15030
rect 13544 14816 13596 14822
rect 13544 14758 13596 14764
rect 12956 14172 13252 14192
rect 13012 14170 13036 14172
rect 13092 14170 13116 14172
rect 13172 14170 13196 14172
rect 13034 14118 13036 14170
rect 13098 14118 13110 14170
rect 13172 14118 13174 14170
rect 13012 14116 13036 14118
rect 13092 14116 13116 14118
rect 13172 14116 13196 14118
rect 12956 14096 13252 14116
rect 13360 13184 13412 13190
rect 13360 13126 13412 13132
rect 12956 13084 13252 13104
rect 13012 13082 13036 13084
rect 13092 13082 13116 13084
rect 13172 13082 13196 13084
rect 13034 13030 13036 13082
rect 13098 13030 13110 13082
rect 13172 13030 13174 13082
rect 13012 13028 13036 13030
rect 13092 13028 13116 13030
rect 13172 13028 13196 13030
rect 12956 13008 13252 13028
rect 13372 12918 13400 13126
rect 13360 12912 13412 12918
rect 13360 12854 13412 12860
rect 13268 12776 13320 12782
rect 13268 12718 13320 12724
rect 13372 12764 13400 12854
rect 13452 12776 13504 12782
rect 13372 12736 13452 12764
rect 12808 12708 12860 12714
rect 12808 12650 12860 12656
rect 12820 12442 12848 12650
rect 13280 12646 13308 12718
rect 13268 12640 13320 12646
rect 13268 12582 13320 12588
rect 12808 12436 12860 12442
rect 12808 12378 12860 12384
rect 13280 12238 13308 12582
rect 13372 12306 13400 12736
rect 13452 12718 13504 12724
rect 13360 12300 13412 12306
rect 13360 12242 13412 12248
rect 13268 12232 13320 12238
rect 13268 12174 13320 12180
rect 12956 11996 13252 12016
rect 13012 11994 13036 11996
rect 13092 11994 13116 11996
rect 13172 11994 13196 11996
rect 13034 11942 13036 11994
rect 13098 11942 13110 11994
rect 13172 11942 13174 11994
rect 13012 11940 13036 11942
rect 13092 11940 13116 11942
rect 13172 11940 13196 11942
rect 12956 11920 13252 11940
rect 12808 11892 12860 11898
rect 12808 11834 12860 11840
rect 12820 10810 12848 11834
rect 13280 11778 13308 12174
rect 13372 11898 13400 12242
rect 13360 11892 13412 11898
rect 13412 11852 13492 11880
rect 13360 11834 13412 11840
rect 13188 11750 13308 11778
rect 13084 11620 13136 11626
rect 13188 11608 13216 11750
rect 13268 11688 13320 11694
rect 13320 11648 13400 11676
rect 13268 11630 13320 11636
rect 13136 11580 13216 11608
rect 13084 11562 13136 11568
rect 13188 11132 13216 11580
rect 13268 11144 13320 11150
rect 13188 11104 13268 11132
rect 13268 11086 13320 11092
rect 12956 10908 13252 10928
rect 13012 10906 13036 10908
rect 13092 10906 13116 10908
rect 13172 10906 13196 10908
rect 13034 10854 13036 10906
rect 13098 10854 13110 10906
rect 13172 10854 13174 10906
rect 13012 10852 13036 10854
rect 13092 10852 13116 10854
rect 13172 10852 13196 10854
rect 12956 10832 13252 10852
rect 12808 10804 12860 10810
rect 12808 10746 12860 10752
rect 13176 10736 13228 10742
rect 13176 10678 13228 10684
rect 13188 10470 13216 10678
rect 13176 10464 13228 10470
rect 13176 10406 13228 10412
rect 12956 9820 13252 9840
rect 13012 9818 13036 9820
rect 13092 9818 13116 9820
rect 13172 9818 13196 9820
rect 13034 9766 13036 9818
rect 13098 9766 13110 9818
rect 13172 9766 13174 9818
rect 13012 9764 13036 9766
rect 13092 9764 13116 9766
rect 13172 9764 13196 9766
rect 12956 9744 13252 9764
rect 13280 9382 13308 11086
rect 13372 11014 13400 11648
rect 13360 11008 13412 11014
rect 13360 10950 13412 10956
rect 13372 10606 13400 10950
rect 13360 10600 13412 10606
rect 13360 10542 13412 10548
rect 13464 10198 13492 11852
rect 13452 10192 13504 10198
rect 13452 10134 13504 10140
rect 13452 10056 13504 10062
rect 13452 9998 13504 10004
rect 13464 9518 13492 9998
rect 13452 9512 13504 9518
rect 13452 9454 13504 9460
rect 13268 9376 13320 9382
rect 13268 9318 13320 9324
rect 13280 9042 13308 9318
rect 13464 9042 13492 9454
rect 13268 9036 13320 9042
rect 13268 8978 13320 8984
rect 13452 9036 13504 9042
rect 13452 8978 13504 8984
rect 12808 8968 12860 8974
rect 12808 8910 12860 8916
rect 12624 8492 12676 8498
rect 12624 8434 12676 8440
rect 11796 7880 11848 7886
rect 11796 7822 11848 7828
rect 11888 7880 11940 7886
rect 11888 7822 11940 7828
rect 11808 7546 11836 7822
rect 11520 7540 11572 7546
rect 11520 7482 11572 7488
rect 11796 7540 11848 7546
rect 11796 7482 11848 7488
rect 12532 7200 12584 7206
rect 12532 7142 12584 7148
rect 12544 7002 12572 7142
rect 12532 6996 12584 7002
rect 12532 6938 12584 6944
rect 11520 6724 11572 6730
rect 11520 6666 11572 6672
rect 11336 5840 11388 5846
rect 11336 5782 11388 5788
rect 11244 5636 11296 5642
rect 11244 5578 11296 5584
rect 10876 5296 10928 5302
rect 10876 5238 10928 5244
rect 10416 5160 10468 5166
rect 10416 5102 10468 5108
rect 10428 4622 10456 5102
rect 10888 4826 10916 5238
rect 11532 4826 11560 6666
rect 12072 6112 12124 6118
rect 12072 6054 12124 6060
rect 11888 5772 11940 5778
rect 11888 5714 11940 5720
rect 11796 5704 11848 5710
rect 11796 5646 11848 5652
rect 11808 5030 11836 5646
rect 11900 5642 11928 5714
rect 11888 5636 11940 5642
rect 11888 5578 11940 5584
rect 12084 5234 12112 6054
rect 12164 5772 12216 5778
rect 12164 5714 12216 5720
rect 12176 5370 12204 5714
rect 12164 5364 12216 5370
rect 12164 5306 12216 5312
rect 12072 5228 12124 5234
rect 12072 5170 12124 5176
rect 11980 5092 12032 5098
rect 11980 5034 12032 5040
rect 11796 5024 11848 5030
rect 11796 4966 11848 4972
rect 10692 4820 10744 4826
rect 10692 4762 10744 4768
rect 10876 4820 10928 4826
rect 10876 4762 10928 4768
rect 11520 4820 11572 4826
rect 11520 4762 11572 4768
rect 10416 4616 10468 4622
rect 10416 4558 10468 4564
rect 9402 4111 9458 4120
rect 8956 3836 9252 3856
rect 9012 3834 9036 3836
rect 9092 3834 9116 3836
rect 9172 3834 9196 3836
rect 9034 3782 9036 3834
rect 9098 3782 9110 3834
rect 9172 3782 9174 3834
rect 9012 3780 9036 3782
rect 9092 3780 9116 3782
rect 9172 3780 9196 3782
rect 8956 3760 9252 3780
rect 8956 2748 9252 2768
rect 9012 2746 9036 2748
rect 9092 2746 9116 2748
rect 9172 2746 9196 2748
rect 9034 2694 9036 2746
rect 9098 2694 9110 2746
rect 9172 2694 9174 2746
rect 9012 2692 9036 2694
rect 9092 2692 9116 2694
rect 9172 2692 9196 2694
rect 8956 2672 9252 2692
rect 9784 2514 9812 4150
rect 10152 4126 10272 4154
rect 10152 3126 10180 4126
rect 10704 3602 10732 4762
rect 10888 4282 10916 4762
rect 11612 4684 11664 4690
rect 11612 4626 11664 4632
rect 10876 4276 10928 4282
rect 10876 4218 10928 4224
rect 10888 4154 10916 4218
rect 11624 4154 11652 4626
rect 10888 4126 11008 4154
rect 11532 4146 11652 4154
rect 10980 4078 11008 4126
rect 11520 4140 11652 4146
rect 11572 4126 11652 4140
rect 11520 4082 11572 4088
rect 10968 4072 11020 4078
rect 10968 4014 11020 4020
rect 11532 3738 11560 4082
rect 11520 3732 11572 3738
rect 11520 3674 11572 3680
rect 11808 3602 11836 4966
rect 11888 4616 11940 4622
rect 11888 4558 11940 4564
rect 11900 4282 11928 4558
rect 11888 4276 11940 4282
rect 11888 4218 11940 4224
rect 11992 3670 12020 5034
rect 12084 4690 12112 5170
rect 12544 4690 12572 6938
rect 12636 6934 12664 8434
rect 12820 8294 12848 8910
rect 12956 8732 13252 8752
rect 13012 8730 13036 8732
rect 13092 8730 13116 8732
rect 13172 8730 13196 8732
rect 13034 8678 13036 8730
rect 13098 8678 13110 8730
rect 13172 8678 13174 8730
rect 13012 8676 13036 8678
rect 13092 8676 13116 8678
rect 13172 8676 13196 8678
rect 12956 8656 13252 8676
rect 13280 8362 13308 8978
rect 13464 8634 13492 8978
rect 13452 8628 13504 8634
rect 13452 8570 13504 8576
rect 13268 8356 13320 8362
rect 13268 8298 13320 8304
rect 12808 8288 12860 8294
rect 12808 8230 12860 8236
rect 12716 7744 12768 7750
rect 12716 7686 12768 7692
rect 12728 7342 12756 7686
rect 12716 7336 12768 7342
rect 12716 7278 12768 7284
rect 12624 6928 12676 6934
rect 12624 6870 12676 6876
rect 12728 6866 12756 7278
rect 12716 6860 12768 6866
rect 12716 6802 12768 6808
rect 12728 6662 12756 6802
rect 12716 6656 12768 6662
rect 12716 6598 12768 6604
rect 12728 5574 12756 6598
rect 12820 6390 12848 8230
rect 12956 7644 13252 7664
rect 13012 7642 13036 7644
rect 13092 7642 13116 7644
rect 13172 7642 13196 7644
rect 13034 7590 13036 7642
rect 13098 7590 13110 7642
rect 13172 7590 13174 7642
rect 13012 7588 13036 7590
rect 13092 7588 13116 7590
rect 13172 7588 13196 7590
rect 12956 7568 13252 7588
rect 13452 7200 13504 7206
rect 13452 7142 13504 7148
rect 13464 6866 13492 7142
rect 13452 6860 13504 6866
rect 13452 6802 13504 6808
rect 12956 6556 13252 6576
rect 13012 6554 13036 6556
rect 13092 6554 13116 6556
rect 13172 6554 13196 6556
rect 13034 6502 13036 6554
rect 13098 6502 13110 6554
rect 13172 6502 13174 6554
rect 13012 6500 13036 6502
rect 13092 6500 13116 6502
rect 13172 6500 13196 6502
rect 12956 6480 13252 6500
rect 12808 6384 12860 6390
rect 12808 6326 12860 6332
rect 13268 6384 13320 6390
rect 13268 6326 13320 6332
rect 12716 5568 12768 5574
rect 12716 5510 12768 5516
rect 12728 5302 12756 5510
rect 12956 5468 13252 5488
rect 13012 5466 13036 5468
rect 13092 5466 13116 5468
rect 13172 5466 13196 5468
rect 13034 5414 13036 5466
rect 13098 5414 13110 5466
rect 13172 5414 13174 5466
rect 13012 5412 13036 5414
rect 13092 5412 13116 5414
rect 13172 5412 13196 5414
rect 12956 5392 13252 5412
rect 12716 5296 12768 5302
rect 12716 5238 12768 5244
rect 12072 4684 12124 4690
rect 12072 4626 12124 4632
rect 12532 4684 12584 4690
rect 12532 4626 12584 4632
rect 12544 4282 12572 4626
rect 12716 4548 12768 4554
rect 12716 4490 12768 4496
rect 12532 4276 12584 4282
rect 12532 4218 12584 4224
rect 12440 3936 12492 3942
rect 12440 3878 12492 3884
rect 11980 3664 12032 3670
rect 11980 3606 12032 3612
rect 10692 3596 10744 3602
rect 10692 3538 10744 3544
rect 11796 3596 11848 3602
rect 11796 3538 11848 3544
rect 10704 3194 10732 3538
rect 10692 3188 10744 3194
rect 10692 3130 10744 3136
rect 10140 3120 10192 3126
rect 10140 3062 10192 3068
rect 11808 2854 11836 3538
rect 11612 2848 11664 2854
rect 11612 2790 11664 2796
rect 11796 2848 11848 2854
rect 11796 2790 11848 2796
rect 9772 2508 9824 2514
rect 9772 2450 9824 2456
rect 10232 2304 10284 2310
rect 10232 2246 10284 2252
rect 8298 54 8616 82
rect 10138 82 10194 480
rect 10244 82 10272 2246
rect 10138 54 10272 82
rect 11624 82 11652 2790
rect 11808 1601 11836 2790
rect 12452 2650 12480 3878
rect 12728 3738 12756 4490
rect 12956 4380 13252 4400
rect 13012 4378 13036 4380
rect 13092 4378 13116 4380
rect 13172 4378 13196 4380
rect 13034 4326 13036 4378
rect 13098 4326 13110 4378
rect 13172 4326 13174 4378
rect 13012 4324 13036 4326
rect 13092 4324 13116 4326
rect 13172 4324 13196 4326
rect 12956 4304 13252 4324
rect 13280 4146 13308 6326
rect 13360 6248 13412 6254
rect 13360 6190 13412 6196
rect 13372 5642 13400 6190
rect 13464 6118 13492 6802
rect 13452 6112 13504 6118
rect 13452 6054 13504 6060
rect 13360 5636 13412 5642
rect 13360 5578 13412 5584
rect 13372 5166 13400 5578
rect 13464 5574 13492 6054
rect 13452 5568 13504 5574
rect 13452 5510 13504 5516
rect 13464 5234 13492 5510
rect 13452 5228 13504 5234
rect 13452 5170 13504 5176
rect 13360 5160 13412 5166
rect 13360 5102 13412 5108
rect 13372 4622 13400 5102
rect 13464 4826 13492 5170
rect 13452 4820 13504 4826
rect 13452 4762 13504 4768
rect 13360 4616 13412 4622
rect 13360 4558 13412 4564
rect 13268 4140 13320 4146
rect 13268 4082 13320 4088
rect 13280 3942 13308 4082
rect 13372 4078 13400 4558
rect 13360 4072 13412 4078
rect 13360 4014 13412 4020
rect 13268 3936 13320 3942
rect 13268 3878 13320 3884
rect 12716 3732 12768 3738
rect 12716 3674 12768 3680
rect 12728 3058 12756 3674
rect 13452 3664 13504 3670
rect 13452 3606 13504 3612
rect 12956 3292 13252 3312
rect 13012 3290 13036 3292
rect 13092 3290 13116 3292
rect 13172 3290 13196 3292
rect 13034 3238 13036 3290
rect 13098 3238 13110 3290
rect 13172 3238 13174 3290
rect 13012 3236 13036 3238
rect 13092 3236 13116 3238
rect 13172 3236 13196 3238
rect 12956 3216 13252 3236
rect 12716 3052 12768 3058
rect 12716 2994 12768 3000
rect 13464 2854 13492 3606
rect 13556 2990 13584 14758
rect 13636 12708 13688 12714
rect 13636 12650 13688 12656
rect 13648 11694 13676 12650
rect 13924 12424 13952 23530
rect 14922 23520 14978 23536
rect 16592 23582 17002 23610
rect 14936 23499 14964 23520
rect 15844 20392 15896 20398
rect 15844 20334 15896 20340
rect 14188 17672 14240 17678
rect 14188 17614 14240 17620
rect 13924 12396 14044 12424
rect 13912 12300 13964 12306
rect 13912 12242 13964 12248
rect 13636 11688 13688 11694
rect 13636 11630 13688 11636
rect 13648 9926 13676 11630
rect 13728 11552 13780 11558
rect 13728 11494 13780 11500
rect 13740 11082 13768 11494
rect 13728 11076 13780 11082
rect 13728 11018 13780 11024
rect 13740 10266 13768 11018
rect 13924 10606 13952 12242
rect 14016 11218 14044 12396
rect 14004 11212 14056 11218
rect 14056 11172 14136 11200
rect 14004 11154 14056 11160
rect 13912 10600 13964 10606
rect 13912 10542 13964 10548
rect 13728 10260 13780 10266
rect 13728 10202 13780 10208
rect 13636 9920 13688 9926
rect 13636 9862 13688 9868
rect 13648 9586 13676 9862
rect 13636 9580 13688 9586
rect 13636 9522 13688 9528
rect 13740 9178 13768 10202
rect 13728 9172 13780 9178
rect 13728 9114 13780 9120
rect 13924 9042 13952 10542
rect 14004 9444 14056 9450
rect 14004 9386 14056 9392
rect 14016 9042 14044 9386
rect 13912 9036 13964 9042
rect 13912 8978 13964 8984
rect 14004 9036 14056 9042
rect 14004 8978 14056 8984
rect 13820 8356 13872 8362
rect 13820 8298 13872 8304
rect 13728 7744 13780 7750
rect 13728 7686 13780 7692
rect 13740 7342 13768 7686
rect 13728 7336 13780 7342
rect 13728 7278 13780 7284
rect 13636 7200 13688 7206
rect 13636 7142 13688 7148
rect 13648 7002 13676 7142
rect 13636 6996 13688 7002
rect 13636 6938 13688 6944
rect 13740 6866 13768 7278
rect 13728 6860 13780 6866
rect 13728 6802 13780 6808
rect 13636 6384 13688 6390
rect 13636 6326 13688 6332
rect 13648 6118 13676 6326
rect 13636 6112 13688 6118
rect 13636 6054 13688 6060
rect 13636 4820 13688 4826
rect 13636 4762 13688 4768
rect 13648 4078 13676 4762
rect 13636 4072 13688 4078
rect 13636 4014 13688 4020
rect 13728 3460 13780 3466
rect 13728 3402 13780 3408
rect 13544 2984 13596 2990
rect 13544 2926 13596 2932
rect 12532 2848 12584 2854
rect 12532 2790 12584 2796
rect 13452 2848 13504 2854
rect 13452 2790 13504 2796
rect 12440 2644 12492 2650
rect 12440 2586 12492 2592
rect 12452 2378 12480 2586
rect 12544 2514 12572 2790
rect 13740 2582 13768 3402
rect 13728 2576 13780 2582
rect 13728 2518 13780 2524
rect 12532 2508 12584 2514
rect 12532 2450 12584 2456
rect 12440 2372 12492 2378
rect 12440 2314 12492 2320
rect 12956 2204 13252 2224
rect 13012 2202 13036 2204
rect 13092 2202 13116 2204
rect 13172 2202 13196 2204
rect 13034 2150 13036 2202
rect 13098 2150 13110 2202
rect 13172 2150 13174 2202
rect 13012 2148 13036 2150
rect 13092 2148 13116 2150
rect 13172 2148 13196 2150
rect 12956 2128 13252 2148
rect 11794 1592 11850 1601
rect 11794 1527 11850 1536
rect 13832 1329 13860 8298
rect 14016 8294 14044 8978
rect 14108 8430 14136 11172
rect 14200 8566 14228 17614
rect 14832 15972 14884 15978
rect 14832 15914 14884 15920
rect 14844 15162 14872 15914
rect 15856 15910 15884 20334
rect 15844 15904 15896 15910
rect 15844 15846 15896 15852
rect 15856 15570 15884 15846
rect 15844 15564 15896 15570
rect 15844 15506 15896 15512
rect 15856 15162 15884 15506
rect 16120 15428 16172 15434
rect 16120 15370 16172 15376
rect 16028 15360 16080 15366
rect 16028 15302 16080 15308
rect 14832 15156 14884 15162
rect 14832 15098 14884 15104
rect 15844 15156 15896 15162
rect 15844 15098 15896 15104
rect 14844 14958 14872 15098
rect 14832 14952 14884 14958
rect 14832 14894 14884 14900
rect 16040 14890 16068 15302
rect 16132 15026 16160 15370
rect 16120 15020 16172 15026
rect 16120 14962 16172 14968
rect 16028 14884 16080 14890
rect 16028 14826 16080 14832
rect 15200 14816 15252 14822
rect 15200 14758 15252 14764
rect 15212 14414 15240 14758
rect 15200 14408 15252 14414
rect 15200 14350 15252 14356
rect 15212 14074 15240 14350
rect 15200 14068 15252 14074
rect 15200 14010 15252 14016
rect 16040 13870 16068 14826
rect 16120 14544 16172 14550
rect 16120 14486 16172 14492
rect 16132 13938 16160 14486
rect 16394 13968 16450 13977
rect 16120 13932 16172 13938
rect 16394 13903 16450 13912
rect 16120 13874 16172 13880
rect 16028 13864 16080 13870
rect 16028 13806 16080 13812
rect 15844 13456 15896 13462
rect 15844 13398 15896 13404
rect 15292 13320 15344 13326
rect 15292 13262 15344 13268
rect 14556 13184 14608 13190
rect 14556 13126 14608 13132
rect 14568 12782 14596 13126
rect 15304 12850 15332 13262
rect 15292 12844 15344 12850
rect 15292 12786 15344 12792
rect 14556 12776 14608 12782
rect 14556 12718 14608 12724
rect 14568 12306 14596 12718
rect 15856 12646 15884 13398
rect 15936 12776 15988 12782
rect 15936 12718 15988 12724
rect 15844 12640 15896 12646
rect 15844 12582 15896 12588
rect 15856 12442 15884 12582
rect 15844 12436 15896 12442
rect 15844 12378 15896 12384
rect 14280 12300 14332 12306
rect 14280 12242 14332 12248
rect 14556 12300 14608 12306
rect 14556 12242 14608 12248
rect 14292 11694 14320 12242
rect 15474 12200 15530 12209
rect 15474 12135 15530 12144
rect 14280 11688 14332 11694
rect 14280 11630 14332 11636
rect 15108 11552 15160 11558
rect 15108 11494 15160 11500
rect 15120 10742 15148 11494
rect 15488 11354 15516 12135
rect 15568 11688 15620 11694
rect 15568 11630 15620 11636
rect 15580 11354 15608 11630
rect 15856 11626 15884 12378
rect 15844 11620 15896 11626
rect 15844 11562 15896 11568
rect 15476 11348 15528 11354
rect 15476 11290 15528 11296
rect 15568 11348 15620 11354
rect 15568 11290 15620 11296
rect 15200 11212 15252 11218
rect 15200 11154 15252 11160
rect 15212 10810 15240 11154
rect 15844 11008 15896 11014
rect 15844 10950 15896 10956
rect 15200 10804 15252 10810
rect 15200 10746 15252 10752
rect 15108 10736 15160 10742
rect 15108 10678 15160 10684
rect 14280 10600 14332 10606
rect 14280 10542 14332 10548
rect 14292 10266 14320 10542
rect 15120 10538 15148 10678
rect 15856 10674 15884 10950
rect 15844 10668 15896 10674
rect 15844 10610 15896 10616
rect 15108 10532 15160 10538
rect 15108 10474 15160 10480
rect 15476 10532 15528 10538
rect 15476 10474 15528 10480
rect 14280 10260 14332 10266
rect 14280 10202 14332 10208
rect 14280 9512 14332 9518
rect 14280 9454 14332 9460
rect 14188 8560 14240 8566
rect 14188 8502 14240 8508
rect 14096 8424 14148 8430
rect 14096 8366 14148 8372
rect 14004 8288 14056 8294
rect 14004 8230 14056 8236
rect 14016 5846 14044 8230
rect 14292 7342 14320 9454
rect 15488 9382 15516 10474
rect 15568 9920 15620 9926
rect 15568 9862 15620 9868
rect 15580 9586 15608 9862
rect 15568 9580 15620 9586
rect 15568 9522 15620 9528
rect 15476 9376 15528 9382
rect 15476 9318 15528 9324
rect 15488 9110 15516 9318
rect 15476 9104 15528 9110
rect 15476 9046 15528 9052
rect 15844 9104 15896 9110
rect 15844 9046 15896 9052
rect 14832 8968 14884 8974
rect 14832 8910 14884 8916
rect 14844 8634 14872 8910
rect 14832 8628 14884 8634
rect 14832 8570 14884 8576
rect 15856 8294 15884 9046
rect 15844 8288 15896 8294
rect 15844 8230 15896 8236
rect 15856 8022 15884 8230
rect 15844 8016 15896 8022
rect 15290 7984 15346 7993
rect 15844 7958 15896 7964
rect 15290 7919 15346 7928
rect 14280 7336 14332 7342
rect 14280 7278 14332 7284
rect 15016 7200 15068 7206
rect 15016 7142 15068 7148
rect 15028 6934 15056 7142
rect 15016 6928 15068 6934
rect 15016 6870 15068 6876
rect 15304 6866 15332 7919
rect 15384 7880 15436 7886
rect 15384 7822 15436 7828
rect 15396 7410 15424 7822
rect 15384 7404 15436 7410
rect 15384 7346 15436 7352
rect 15396 7002 15424 7346
rect 15856 7206 15884 7958
rect 15844 7200 15896 7206
rect 15844 7142 15896 7148
rect 15384 6996 15436 7002
rect 15384 6938 15436 6944
rect 14648 6860 14700 6866
rect 14648 6802 14700 6808
rect 15292 6860 15344 6866
rect 15292 6802 15344 6808
rect 14660 6254 14688 6802
rect 15304 6458 15332 6802
rect 15856 6662 15884 7142
rect 15568 6656 15620 6662
rect 15568 6598 15620 6604
rect 15844 6656 15896 6662
rect 15844 6598 15896 6604
rect 15292 6452 15344 6458
rect 15292 6394 15344 6400
rect 14280 6248 14332 6254
rect 14280 6190 14332 6196
rect 14648 6248 14700 6254
rect 14648 6190 14700 6196
rect 14004 5840 14056 5846
rect 14004 5782 14056 5788
rect 14292 5574 14320 6190
rect 14280 5568 14332 5574
rect 14280 5510 14332 5516
rect 14292 5234 14320 5510
rect 14280 5228 14332 5234
rect 14280 5170 14332 5176
rect 14556 5160 14608 5166
rect 14556 5102 14608 5108
rect 14568 4826 14596 5102
rect 15200 5024 15252 5030
rect 15200 4966 15252 4972
rect 14556 4820 14608 4826
rect 14556 4762 14608 4768
rect 14280 4548 14332 4554
rect 14280 4490 14332 4496
rect 14292 4078 14320 4490
rect 14280 4072 14332 4078
rect 14280 4014 14332 4020
rect 14292 3738 14320 4014
rect 14924 4004 14976 4010
rect 14924 3946 14976 3952
rect 14280 3732 14332 3738
rect 14280 3674 14332 3680
rect 14936 3534 14964 3946
rect 15212 3670 15240 4966
rect 15200 3664 15252 3670
rect 15200 3606 15252 3612
rect 14004 3528 14056 3534
rect 14004 3470 14056 3476
rect 14924 3528 14976 3534
rect 14924 3470 14976 3476
rect 14016 3194 14044 3470
rect 14004 3188 14056 3194
rect 14004 3130 14056 3136
rect 15212 2922 15240 3606
rect 15200 2916 15252 2922
rect 15200 2858 15252 2864
rect 14096 2848 14148 2854
rect 14096 2790 14148 2796
rect 13818 1320 13874 1329
rect 13818 1255 13874 1264
rect 11978 82 12034 480
rect 11624 54 12034 82
rect 938 0 994 54
rect 2778 0 2834 54
rect 4618 0 4674 54
rect 6458 0 6514 54
rect 8298 0 8354 54
rect 10138 0 10194 54
rect 11978 0 12034 54
rect 13818 82 13874 480
rect 14108 82 14136 2790
rect 15580 2582 15608 6598
rect 15752 6248 15804 6254
rect 15752 6190 15804 6196
rect 15764 5914 15792 6190
rect 15856 6186 15884 6598
rect 15844 6180 15896 6186
rect 15844 6122 15896 6128
rect 15752 5908 15804 5914
rect 15752 5850 15804 5856
rect 15752 5568 15804 5574
rect 15856 5556 15884 6122
rect 15804 5528 15884 5556
rect 15752 5510 15804 5516
rect 15660 5160 15712 5166
rect 15660 5102 15712 5108
rect 15672 4826 15700 5102
rect 15764 5030 15792 5510
rect 15752 5024 15804 5030
rect 15752 4966 15804 4972
rect 15660 4820 15712 4826
rect 15660 4762 15712 4768
rect 15844 3120 15896 3126
rect 15844 3062 15896 3068
rect 15568 2576 15620 2582
rect 15568 2518 15620 2524
rect 15856 2446 15884 3062
rect 15948 2446 15976 12718
rect 16040 6458 16068 13806
rect 16408 12986 16436 13903
rect 16592 13814 16620 23582
rect 16946 23520 17002 23582
rect 18616 23582 18934 23610
rect 18326 22672 18382 22681
rect 18326 22607 18382 22616
rect 16956 21244 17252 21264
rect 17012 21242 17036 21244
rect 17092 21242 17116 21244
rect 17172 21242 17196 21244
rect 17034 21190 17036 21242
rect 17098 21190 17110 21242
rect 17172 21190 17174 21242
rect 17012 21188 17036 21190
rect 17092 21188 17116 21190
rect 17172 21188 17196 21190
rect 16956 21168 17252 21188
rect 16956 20156 17252 20176
rect 17012 20154 17036 20156
rect 17092 20154 17116 20156
rect 17172 20154 17196 20156
rect 17034 20102 17036 20154
rect 17098 20102 17110 20154
rect 17172 20102 17174 20154
rect 17012 20100 17036 20102
rect 17092 20100 17116 20102
rect 17172 20100 17196 20102
rect 16956 20080 17252 20100
rect 16956 19068 17252 19088
rect 17012 19066 17036 19068
rect 17092 19066 17116 19068
rect 17172 19066 17196 19068
rect 17034 19014 17036 19066
rect 17098 19014 17110 19066
rect 17172 19014 17174 19066
rect 17012 19012 17036 19014
rect 17092 19012 17116 19014
rect 17172 19012 17196 19014
rect 16956 18992 17252 19012
rect 16762 18184 16818 18193
rect 16762 18119 16818 18128
rect 16776 15978 16804 18119
rect 16956 17980 17252 18000
rect 17012 17978 17036 17980
rect 17092 17978 17116 17980
rect 17172 17978 17196 17980
rect 17034 17926 17036 17978
rect 17098 17926 17110 17978
rect 17172 17926 17174 17978
rect 17012 17924 17036 17926
rect 17092 17924 17116 17926
rect 17172 17924 17196 17926
rect 16956 17904 17252 17924
rect 16956 16892 17252 16912
rect 17012 16890 17036 16892
rect 17092 16890 17116 16892
rect 17172 16890 17196 16892
rect 17034 16838 17036 16890
rect 17098 16838 17110 16890
rect 17172 16838 17174 16890
rect 17012 16836 17036 16838
rect 17092 16836 17116 16838
rect 17172 16836 17196 16838
rect 16956 16816 17252 16836
rect 16764 15972 16816 15978
rect 16764 15914 16816 15920
rect 16956 15804 17252 15824
rect 17012 15802 17036 15804
rect 17092 15802 17116 15804
rect 17172 15802 17196 15804
rect 17034 15750 17036 15802
rect 17098 15750 17110 15802
rect 17172 15750 17174 15802
rect 17012 15748 17036 15750
rect 17092 15748 17116 15750
rect 17172 15748 17196 15750
rect 16956 15728 17252 15748
rect 16672 14884 16724 14890
rect 16672 14826 16724 14832
rect 16684 14550 16712 14826
rect 16956 14716 17252 14736
rect 17012 14714 17036 14716
rect 17092 14714 17116 14716
rect 17172 14714 17196 14716
rect 17034 14662 17036 14714
rect 17098 14662 17110 14714
rect 17172 14662 17174 14714
rect 17012 14660 17036 14662
rect 17092 14660 17116 14662
rect 17172 14660 17196 14662
rect 16956 14640 17252 14660
rect 16672 14544 16724 14550
rect 16724 14504 16896 14532
rect 16672 14486 16724 14492
rect 16592 13786 16712 13814
rect 16396 12980 16448 12986
rect 16396 12922 16448 12928
rect 16488 11552 16540 11558
rect 16488 11494 16540 11500
rect 16500 11286 16528 11494
rect 16488 11280 16540 11286
rect 16488 11222 16540 11228
rect 16212 10192 16264 10198
rect 16212 10134 16264 10140
rect 16224 9178 16252 10134
rect 16488 10056 16540 10062
rect 16488 9998 16540 10004
rect 16212 9172 16264 9178
rect 16212 9114 16264 9120
rect 16500 8838 16528 9998
rect 16684 9654 16712 13786
rect 16764 12232 16816 12238
rect 16764 12174 16816 12180
rect 16776 11898 16804 12174
rect 16764 11892 16816 11898
rect 16764 11834 16816 11840
rect 16764 10056 16816 10062
rect 16764 9998 16816 10004
rect 16776 9654 16804 9998
rect 16672 9648 16724 9654
rect 16672 9590 16724 9596
rect 16764 9648 16816 9654
rect 16764 9590 16816 9596
rect 16488 8832 16540 8838
rect 16868 8786 16896 14504
rect 18340 14074 18368 22607
rect 18616 15094 18644 23582
rect 18878 23520 18934 23582
rect 20640 23582 20958 23610
rect 20640 20602 20668 23582
rect 20902 23520 20958 23582
rect 22664 23582 22982 23610
rect 20956 21788 21252 21808
rect 21012 21786 21036 21788
rect 21092 21786 21116 21788
rect 21172 21786 21196 21788
rect 21034 21734 21036 21786
rect 21098 21734 21110 21786
rect 21172 21734 21174 21786
rect 21012 21732 21036 21734
rect 21092 21732 21116 21734
rect 21172 21732 21196 21734
rect 20956 21712 21252 21732
rect 21362 21176 21418 21185
rect 21362 21111 21418 21120
rect 20956 20700 21252 20720
rect 21012 20698 21036 20700
rect 21092 20698 21116 20700
rect 21172 20698 21196 20700
rect 21034 20646 21036 20698
rect 21098 20646 21110 20698
rect 21172 20646 21174 20698
rect 21012 20644 21036 20646
rect 21092 20644 21116 20646
rect 21172 20644 21196 20646
rect 20956 20624 21252 20644
rect 20628 20596 20680 20602
rect 20628 20538 20680 20544
rect 20812 20392 20864 20398
rect 20812 20334 20864 20340
rect 20824 18737 20852 20334
rect 20956 19612 21252 19632
rect 21012 19610 21036 19612
rect 21092 19610 21116 19612
rect 21172 19610 21196 19612
rect 21034 19558 21036 19610
rect 21098 19558 21110 19610
rect 21172 19558 21174 19610
rect 21012 19556 21036 19558
rect 21092 19556 21116 19558
rect 21172 19556 21196 19558
rect 20956 19536 21252 19556
rect 20810 18728 20866 18737
rect 20810 18663 20866 18672
rect 20956 18524 21252 18544
rect 21012 18522 21036 18524
rect 21092 18522 21116 18524
rect 21172 18522 21196 18524
rect 21034 18470 21036 18522
rect 21098 18470 21110 18522
rect 21172 18470 21174 18522
rect 21012 18468 21036 18470
rect 21092 18468 21116 18470
rect 21172 18468 21196 18470
rect 20956 18448 21252 18468
rect 20956 17436 21252 17456
rect 21012 17434 21036 17436
rect 21092 17434 21116 17436
rect 21172 17434 21196 17436
rect 21034 17382 21036 17434
rect 21098 17382 21110 17434
rect 21172 17382 21174 17434
rect 21012 17380 21036 17382
rect 21092 17380 21116 17382
rect 21172 17380 21196 17382
rect 20956 17360 21252 17380
rect 20956 16348 21252 16368
rect 21012 16346 21036 16348
rect 21092 16346 21116 16348
rect 21172 16346 21196 16348
rect 21034 16294 21036 16346
rect 21098 16294 21110 16346
rect 21172 16294 21174 16346
rect 21012 16292 21036 16294
rect 21092 16292 21116 16294
rect 21172 16292 21196 16294
rect 20956 16272 21252 16292
rect 21270 15464 21326 15473
rect 21270 15399 21326 15408
rect 20956 15260 21252 15280
rect 21012 15258 21036 15260
rect 21092 15258 21116 15260
rect 21172 15258 21196 15260
rect 21034 15206 21036 15258
rect 21098 15206 21110 15258
rect 21172 15206 21174 15258
rect 21012 15204 21036 15206
rect 21092 15204 21116 15206
rect 21172 15204 21196 15206
rect 20956 15184 21252 15204
rect 21284 15162 21312 15399
rect 21272 15156 21324 15162
rect 21272 15098 21324 15104
rect 18604 15088 18656 15094
rect 18604 15030 18656 15036
rect 20812 14952 20864 14958
rect 20812 14894 20864 14900
rect 18328 14068 18380 14074
rect 18328 14010 18380 14016
rect 17776 13864 17828 13870
rect 17776 13806 17828 13812
rect 16956 13628 17252 13648
rect 17012 13626 17036 13628
rect 17092 13626 17116 13628
rect 17172 13626 17196 13628
rect 17034 13574 17036 13626
rect 17098 13574 17110 13626
rect 17172 13574 17174 13626
rect 17012 13572 17036 13574
rect 17092 13572 17116 13574
rect 17172 13572 17196 13574
rect 16956 13552 17252 13572
rect 17500 13456 17552 13462
rect 17500 13398 17552 13404
rect 17132 13320 17184 13326
rect 17132 13262 17184 13268
rect 17144 12986 17172 13262
rect 17132 12980 17184 12986
rect 17132 12922 17184 12928
rect 17512 12918 17540 13398
rect 17788 13326 17816 13806
rect 17776 13320 17828 13326
rect 17776 13262 17828 13268
rect 17500 12912 17552 12918
rect 17500 12854 17552 12860
rect 16956 12540 17252 12560
rect 17012 12538 17036 12540
rect 17092 12538 17116 12540
rect 17172 12538 17196 12540
rect 17034 12486 17036 12538
rect 17098 12486 17110 12538
rect 17172 12486 17174 12538
rect 17012 12484 17036 12486
rect 17092 12484 17116 12486
rect 17172 12484 17196 12486
rect 16956 12464 17252 12484
rect 17316 12436 17368 12442
rect 17316 12378 17368 12384
rect 17328 11898 17356 12378
rect 17788 12238 17816 13262
rect 20824 12306 20852 14894
rect 20956 14172 21252 14192
rect 21012 14170 21036 14172
rect 21092 14170 21116 14172
rect 21172 14170 21196 14172
rect 21034 14118 21036 14170
rect 21098 14118 21110 14170
rect 21172 14118 21174 14170
rect 21012 14116 21036 14118
rect 21092 14116 21116 14118
rect 21172 14116 21196 14118
rect 20956 14096 21252 14116
rect 21376 13814 21404 21111
rect 22664 20602 22692 23582
rect 22926 23520 22982 23582
rect 22652 20596 22704 20602
rect 22652 20538 22704 20544
rect 21546 19680 21602 19689
rect 21546 19615 21602 19624
rect 21560 15162 21588 19615
rect 21548 15156 21600 15162
rect 21548 15098 21600 15104
rect 21560 14958 21588 15098
rect 21548 14952 21600 14958
rect 21548 14894 21600 14900
rect 21284 13786 21404 13814
rect 20956 13084 21252 13104
rect 21012 13082 21036 13084
rect 21092 13082 21116 13084
rect 21172 13082 21196 13084
rect 21034 13030 21036 13082
rect 21098 13030 21110 13082
rect 21172 13030 21174 13082
rect 21012 13028 21036 13030
rect 21092 13028 21116 13030
rect 21172 13028 21196 13030
rect 20956 13008 21252 13028
rect 18880 12300 18932 12306
rect 18880 12242 18932 12248
rect 20812 12300 20864 12306
rect 20812 12242 20864 12248
rect 17408 12232 17460 12238
rect 17408 12174 17460 12180
rect 17776 12232 17828 12238
rect 17776 12174 17828 12180
rect 17316 11892 17368 11898
rect 17316 11834 17368 11840
rect 17420 11558 17448 12174
rect 17408 11552 17460 11558
rect 17408 11494 17460 11500
rect 16956 11452 17252 11472
rect 17012 11450 17036 11452
rect 17092 11450 17116 11452
rect 17172 11450 17196 11452
rect 17034 11398 17036 11450
rect 17098 11398 17110 11450
rect 17172 11398 17174 11450
rect 17012 11396 17036 11398
rect 17092 11396 17116 11398
rect 17172 11396 17196 11398
rect 16956 11376 17252 11396
rect 17788 11286 17816 12174
rect 18696 12096 18748 12102
rect 18696 12038 18748 12044
rect 18708 11286 18736 12038
rect 18892 11898 18920 12242
rect 20956 11996 21252 12016
rect 21012 11994 21036 11996
rect 21092 11994 21116 11996
rect 21172 11994 21196 11996
rect 21034 11942 21036 11994
rect 21098 11942 21110 11994
rect 21172 11942 21174 11994
rect 21012 11940 21036 11942
rect 21092 11940 21116 11942
rect 21172 11940 21196 11942
rect 20956 11920 21252 11940
rect 18880 11892 18932 11898
rect 18880 11834 18932 11840
rect 18972 11552 19024 11558
rect 18972 11494 19024 11500
rect 17132 11280 17184 11286
rect 17132 11222 17184 11228
rect 17776 11280 17828 11286
rect 17776 11222 17828 11228
rect 18696 11280 18748 11286
rect 18696 11222 18748 11228
rect 18880 11280 18932 11286
rect 18880 11222 18932 11228
rect 17144 10810 17172 11222
rect 17408 11144 17460 11150
rect 17408 11086 17460 11092
rect 17420 10810 17448 11086
rect 18144 11008 18196 11014
rect 18144 10950 18196 10956
rect 17132 10804 17184 10810
rect 17132 10746 17184 10752
rect 17408 10804 17460 10810
rect 17408 10746 17460 10752
rect 18156 10538 18184 10950
rect 18708 10810 18736 11222
rect 18696 10804 18748 10810
rect 18696 10746 18748 10752
rect 18328 10668 18380 10674
rect 18328 10610 18380 10616
rect 18144 10532 18196 10538
rect 18144 10474 18196 10480
rect 16956 10364 17252 10384
rect 17012 10362 17036 10364
rect 17092 10362 17116 10364
rect 17172 10362 17196 10364
rect 17034 10310 17036 10362
rect 17098 10310 17110 10362
rect 17172 10310 17174 10362
rect 17012 10308 17036 10310
rect 17092 10308 17116 10310
rect 17172 10308 17196 10310
rect 16956 10288 17252 10308
rect 18156 10266 18184 10474
rect 18144 10260 18196 10266
rect 18144 10202 18196 10208
rect 18340 10198 18368 10610
rect 18892 10470 18920 11222
rect 18984 11150 19012 11494
rect 18972 11144 19024 11150
rect 18972 11086 19024 11092
rect 18880 10464 18932 10470
rect 18880 10406 18932 10412
rect 17776 10192 17828 10198
rect 17776 10134 17828 10140
rect 18328 10192 18380 10198
rect 18328 10134 18380 10140
rect 17684 10056 17736 10062
rect 17684 9998 17736 10004
rect 17696 9586 17724 9998
rect 17684 9580 17736 9586
rect 17684 9522 17736 9528
rect 17500 9376 17552 9382
rect 17500 9318 17552 9324
rect 16956 9276 17252 9296
rect 17012 9274 17036 9276
rect 17092 9274 17116 9276
rect 17172 9274 17196 9276
rect 17034 9222 17036 9274
rect 17098 9222 17110 9274
rect 17172 9222 17174 9274
rect 17012 9220 17036 9222
rect 17092 9220 17116 9222
rect 17172 9220 17196 9222
rect 16956 9200 17252 9220
rect 17512 9110 17540 9318
rect 17696 9178 17724 9522
rect 17788 9518 17816 10134
rect 17960 9716 18012 9722
rect 17960 9658 18012 9664
rect 17776 9512 17828 9518
rect 17776 9454 17828 9460
rect 17684 9172 17736 9178
rect 17684 9114 17736 9120
rect 17500 9104 17552 9110
rect 17500 9046 17552 9052
rect 17132 8968 17184 8974
rect 17132 8910 17184 8916
rect 16488 8774 16540 8780
rect 16500 8634 16528 8774
rect 16776 8758 16896 8786
rect 16488 8628 16540 8634
rect 16488 8570 16540 8576
rect 16580 7200 16632 7206
rect 16580 7142 16632 7148
rect 16592 6934 16620 7142
rect 16580 6928 16632 6934
rect 16580 6870 16632 6876
rect 16028 6452 16080 6458
rect 16028 6394 16080 6400
rect 16776 5642 16804 8758
rect 17144 8634 17172 8910
rect 17512 8634 17540 9046
rect 16856 8628 16908 8634
rect 16856 8570 16908 8576
rect 17132 8628 17184 8634
rect 17132 8570 17184 8576
rect 17500 8628 17552 8634
rect 17500 8570 17552 8576
rect 16868 8090 16896 8570
rect 17316 8288 17368 8294
rect 17316 8230 17368 8236
rect 16956 8188 17252 8208
rect 17012 8186 17036 8188
rect 17092 8186 17116 8188
rect 17172 8186 17196 8188
rect 17034 8134 17036 8186
rect 17098 8134 17110 8186
rect 17172 8134 17174 8186
rect 17012 8132 17036 8134
rect 17092 8132 17116 8134
rect 17172 8132 17196 8134
rect 16956 8112 17252 8132
rect 16856 8084 16908 8090
rect 16856 8026 16908 8032
rect 16956 7100 17252 7120
rect 17012 7098 17036 7100
rect 17092 7098 17116 7100
rect 17172 7098 17196 7100
rect 17034 7046 17036 7098
rect 17098 7046 17110 7098
rect 17172 7046 17174 7098
rect 17012 7044 17036 7046
rect 17092 7044 17116 7046
rect 17172 7044 17196 7046
rect 16956 7024 17252 7044
rect 17328 6866 17356 8230
rect 17972 7313 18000 9658
rect 18144 9444 18196 9450
rect 18144 9386 18196 9392
rect 18156 8974 18184 9386
rect 18340 9110 18368 10134
rect 18984 9654 19012 11086
rect 20956 10908 21252 10928
rect 21012 10906 21036 10908
rect 21092 10906 21116 10908
rect 21172 10906 21196 10908
rect 21034 10854 21036 10906
rect 21098 10854 21110 10906
rect 21172 10854 21174 10906
rect 21012 10852 21036 10854
rect 21092 10852 21116 10854
rect 21172 10852 21196 10854
rect 20956 10832 21252 10852
rect 20076 10600 20128 10606
rect 20076 10542 20128 10548
rect 19156 10124 19208 10130
rect 19156 10066 19208 10072
rect 19168 9722 19196 10066
rect 19156 9716 19208 9722
rect 19156 9658 19208 9664
rect 18972 9648 19024 9654
rect 18972 9590 19024 9596
rect 20088 9518 20116 10542
rect 20956 9820 21252 9840
rect 21012 9818 21036 9820
rect 21092 9818 21116 9820
rect 21172 9818 21196 9820
rect 21034 9766 21036 9818
rect 21098 9766 21110 9818
rect 21172 9766 21174 9818
rect 21012 9764 21036 9766
rect 21092 9764 21116 9766
rect 21172 9764 21196 9766
rect 20956 9744 21252 9764
rect 20076 9512 20128 9518
rect 20076 9454 20128 9460
rect 18604 9444 18656 9450
rect 18604 9386 18656 9392
rect 18328 9104 18380 9110
rect 18328 9046 18380 9052
rect 18616 9042 18644 9386
rect 21284 9178 21312 13786
rect 21362 10840 21418 10849
rect 21362 10775 21418 10784
rect 21376 10742 21404 10775
rect 21364 10736 21416 10742
rect 21364 10678 21416 10684
rect 21362 9752 21418 9761
rect 21362 9687 21418 9696
rect 21272 9172 21324 9178
rect 21272 9114 21324 9120
rect 18604 9036 18656 9042
rect 18604 8978 18656 8984
rect 20076 9036 20128 9042
rect 20076 8978 20128 8984
rect 20812 9036 20864 9042
rect 20812 8978 20864 8984
rect 18144 8968 18196 8974
rect 18144 8910 18196 8916
rect 18512 8832 18564 8838
rect 18512 8774 18564 8780
rect 18052 8016 18104 8022
rect 18052 7958 18104 7964
rect 17958 7304 18014 7313
rect 17958 7239 18014 7248
rect 17868 6928 17920 6934
rect 17868 6870 17920 6876
rect 17040 6860 17092 6866
rect 17040 6802 17092 6808
rect 17316 6860 17368 6866
rect 17316 6802 17368 6808
rect 17052 6186 17080 6802
rect 17408 6656 17460 6662
rect 17408 6598 17460 6604
rect 17420 6458 17448 6598
rect 17880 6458 17908 6870
rect 17408 6452 17460 6458
rect 17408 6394 17460 6400
rect 17868 6452 17920 6458
rect 17868 6394 17920 6400
rect 17880 6254 17908 6394
rect 17868 6248 17920 6254
rect 17868 6190 17920 6196
rect 17040 6180 17092 6186
rect 17040 6122 17092 6128
rect 16956 6012 17252 6032
rect 17012 6010 17036 6012
rect 17092 6010 17116 6012
rect 17172 6010 17196 6012
rect 17034 5958 17036 6010
rect 17098 5958 17110 6010
rect 17172 5958 17174 6010
rect 17012 5956 17036 5958
rect 17092 5956 17116 5958
rect 17172 5956 17196 5958
rect 16956 5936 17252 5956
rect 17880 5914 17908 6190
rect 17868 5908 17920 5914
rect 17868 5850 17920 5856
rect 16948 5840 17000 5846
rect 16948 5782 17000 5788
rect 16764 5636 16816 5642
rect 16764 5578 16816 5584
rect 16776 5370 16804 5578
rect 16764 5364 16816 5370
rect 16764 5306 16816 5312
rect 16960 5098 16988 5782
rect 17408 5636 17460 5642
rect 17408 5578 17460 5584
rect 17776 5636 17828 5642
rect 17776 5578 17828 5584
rect 16948 5092 17000 5098
rect 16948 5034 17000 5040
rect 16956 4924 17252 4944
rect 17012 4922 17036 4924
rect 17092 4922 17116 4924
rect 17172 4922 17196 4924
rect 17034 4870 17036 4922
rect 17098 4870 17110 4922
rect 17172 4870 17174 4922
rect 17012 4868 17036 4870
rect 17092 4868 17116 4870
rect 17172 4868 17196 4870
rect 16956 4848 17252 4868
rect 17040 4752 17092 4758
rect 17040 4694 17092 4700
rect 16856 4548 16908 4554
rect 16856 4490 16908 4496
rect 16868 4214 16896 4490
rect 16856 4208 16908 4214
rect 16856 4150 16908 4156
rect 16212 4072 16264 4078
rect 16212 4014 16264 4020
rect 16224 3738 16252 4014
rect 16488 4004 16540 4010
rect 16488 3946 16540 3952
rect 16212 3732 16264 3738
rect 16212 3674 16264 3680
rect 16224 2582 16252 3674
rect 16500 3194 16528 3946
rect 16868 3738 16896 4150
rect 17052 4146 17080 4694
rect 17420 4622 17448 5578
rect 17408 4616 17460 4622
rect 17408 4558 17460 4564
rect 17040 4140 17092 4146
rect 17040 4082 17092 4088
rect 17420 4078 17448 4558
rect 17408 4072 17460 4078
rect 17408 4014 17460 4020
rect 16956 3836 17252 3856
rect 17012 3834 17036 3836
rect 17092 3834 17116 3836
rect 17172 3834 17196 3836
rect 17034 3782 17036 3834
rect 17098 3782 17110 3834
rect 17172 3782 17174 3834
rect 17012 3780 17036 3782
rect 17092 3780 17116 3782
rect 17172 3780 17196 3782
rect 16956 3760 17252 3780
rect 16856 3732 16908 3738
rect 16856 3674 16908 3680
rect 16764 3528 16816 3534
rect 16764 3470 16816 3476
rect 16776 3194 16804 3470
rect 16488 3188 16540 3194
rect 16488 3130 16540 3136
rect 16764 3188 16816 3194
rect 16764 3130 16816 3136
rect 16500 2854 16528 3130
rect 16856 3052 16908 3058
rect 16856 2994 16908 3000
rect 16488 2848 16540 2854
rect 16488 2790 16540 2796
rect 16868 2650 16896 2994
rect 16956 2748 17252 2768
rect 17012 2746 17036 2748
rect 17092 2746 17116 2748
rect 17172 2746 17196 2748
rect 17034 2694 17036 2746
rect 17098 2694 17110 2746
rect 17172 2694 17174 2746
rect 17012 2692 17036 2694
rect 17092 2692 17116 2694
rect 17172 2692 17196 2694
rect 16956 2672 17252 2692
rect 16856 2644 16908 2650
rect 16856 2586 16908 2592
rect 16212 2576 16264 2582
rect 16212 2518 16264 2524
rect 15844 2440 15896 2446
rect 15844 2382 15896 2388
rect 15936 2440 15988 2446
rect 15936 2382 15988 2388
rect 13818 54 14136 82
rect 15658 82 15714 480
rect 15948 82 15976 2382
rect 15658 54 15976 82
rect 17498 82 17554 480
rect 17788 82 17816 5578
rect 17972 2514 18000 7239
rect 18064 7206 18092 7958
rect 18524 7886 18552 8774
rect 18616 8566 18644 8978
rect 20088 8634 20116 8978
rect 20076 8628 20128 8634
rect 20076 8570 20128 8576
rect 18604 8560 18656 8566
rect 18604 8502 18656 8508
rect 19064 8424 19116 8430
rect 19064 8366 19116 8372
rect 18512 7880 18564 7886
rect 18512 7822 18564 7828
rect 18880 7880 18932 7886
rect 18880 7822 18932 7828
rect 18328 7812 18380 7818
rect 18328 7754 18380 7760
rect 18340 7274 18368 7754
rect 18524 7546 18552 7822
rect 18892 7546 18920 7822
rect 19076 7750 19104 8366
rect 20824 8362 20852 8978
rect 20956 8732 21252 8752
rect 21012 8730 21036 8732
rect 21092 8730 21116 8732
rect 21172 8730 21196 8732
rect 21034 8678 21036 8730
rect 21098 8678 21110 8730
rect 21172 8678 21174 8730
rect 21012 8676 21036 8678
rect 21092 8676 21116 8678
rect 21172 8676 21196 8678
rect 20956 8656 21252 8676
rect 21376 8634 21404 9687
rect 21364 8628 21416 8634
rect 21364 8570 21416 8576
rect 21272 8560 21324 8566
rect 21272 8502 21324 8508
rect 19708 8356 19760 8362
rect 19708 8298 19760 8304
rect 20812 8356 20864 8362
rect 20812 8298 20864 8304
rect 19432 8288 19484 8294
rect 19432 8230 19484 8236
rect 19444 8022 19472 8230
rect 19432 8016 19484 8022
rect 19432 7958 19484 7964
rect 19064 7744 19116 7750
rect 19064 7686 19116 7692
rect 18512 7540 18564 7546
rect 18512 7482 18564 7488
rect 18880 7540 18932 7546
rect 18880 7482 18932 7488
rect 18328 7268 18380 7274
rect 18328 7210 18380 7216
rect 19076 7256 19104 7686
rect 19444 7546 19472 7958
rect 19720 7818 19748 8298
rect 19708 7812 19760 7818
rect 19708 7754 19760 7760
rect 19432 7540 19484 7546
rect 19432 7482 19484 7488
rect 19720 7410 19748 7754
rect 20956 7644 21252 7664
rect 21012 7642 21036 7644
rect 21092 7642 21116 7644
rect 21172 7642 21196 7644
rect 21034 7590 21036 7642
rect 21098 7590 21110 7642
rect 21172 7590 21174 7642
rect 21012 7588 21036 7590
rect 21092 7588 21116 7590
rect 21172 7588 21196 7590
rect 20956 7568 21252 7588
rect 19708 7404 19760 7410
rect 19708 7346 19760 7352
rect 19156 7268 19208 7274
rect 19076 7228 19156 7256
rect 18052 7200 18104 7206
rect 18052 7142 18104 7148
rect 18064 6322 18092 7142
rect 18340 6798 18368 7210
rect 19076 7002 19104 7228
rect 19156 7210 19208 7216
rect 19064 6996 19116 7002
rect 19064 6938 19116 6944
rect 18328 6792 18380 6798
rect 18328 6734 18380 6740
rect 20956 6556 21252 6576
rect 21012 6554 21036 6556
rect 21092 6554 21116 6556
rect 21172 6554 21196 6556
rect 21034 6502 21036 6554
rect 21098 6502 21110 6554
rect 21172 6502 21174 6554
rect 21012 6500 21036 6502
rect 21092 6500 21116 6502
rect 21172 6500 21196 6502
rect 20956 6480 21252 6500
rect 18052 6316 18104 6322
rect 18052 6258 18104 6264
rect 18326 6216 18382 6225
rect 18326 6151 18328 6160
rect 18380 6151 18382 6160
rect 18328 6122 18380 6128
rect 18340 5778 18368 6122
rect 18328 5772 18380 5778
rect 18328 5714 18380 5720
rect 18340 5370 18368 5714
rect 20956 5468 21252 5488
rect 21012 5466 21036 5468
rect 21092 5466 21116 5468
rect 21172 5466 21196 5468
rect 21034 5414 21036 5466
rect 21098 5414 21110 5466
rect 21172 5414 21174 5466
rect 21012 5412 21036 5414
rect 21092 5412 21116 5414
rect 21172 5412 21196 5414
rect 20956 5392 21252 5412
rect 18328 5364 18380 5370
rect 18328 5306 18380 5312
rect 18512 5092 18564 5098
rect 18512 5034 18564 5040
rect 18524 4690 18552 5034
rect 18512 4684 18564 4690
rect 18512 4626 18564 4632
rect 18524 4282 18552 4626
rect 20956 4380 21252 4400
rect 21012 4378 21036 4380
rect 21092 4378 21116 4380
rect 21172 4378 21196 4380
rect 21034 4326 21036 4378
rect 21098 4326 21110 4378
rect 21172 4326 21174 4378
rect 21012 4324 21036 4326
rect 21092 4324 21116 4326
rect 21172 4324 21196 4326
rect 20956 4304 21252 4324
rect 18512 4276 18564 4282
rect 18512 4218 18564 4224
rect 20956 3292 21252 3312
rect 21012 3290 21036 3292
rect 21092 3290 21116 3292
rect 21172 3290 21196 3292
rect 21034 3238 21036 3290
rect 21098 3238 21110 3290
rect 21172 3238 21174 3290
rect 21012 3236 21036 3238
rect 21092 3236 21116 3238
rect 21172 3236 21196 3238
rect 20956 3216 21252 3236
rect 17960 2508 18012 2514
rect 17960 2450 18012 2456
rect 19892 2508 19944 2514
rect 19892 2450 19944 2456
rect 19432 2372 19484 2378
rect 19432 2314 19484 2320
rect 17498 54 17816 82
rect 19338 82 19394 480
rect 19444 82 19472 2314
rect 19904 2009 19932 2450
rect 20956 2204 21252 2224
rect 21012 2202 21036 2204
rect 21092 2202 21116 2204
rect 21172 2202 21196 2204
rect 21034 2150 21036 2202
rect 21098 2150 21110 2202
rect 21172 2150 21174 2202
rect 21012 2148 21036 2150
rect 21092 2148 21116 2150
rect 21172 2148 21196 2150
rect 20956 2128 21252 2148
rect 19890 2000 19946 2009
rect 19890 1935 19946 1944
rect 19338 54 19472 82
rect 21178 82 21234 480
rect 21284 82 21312 8502
rect 23570 5264 23626 5273
rect 23570 5199 23626 5208
rect 23584 4185 23612 5199
rect 23570 4176 23626 4185
rect 23570 4111 23626 4120
rect 23572 4004 23624 4010
rect 23572 3946 23624 3952
rect 23584 3777 23612 3946
rect 23570 3768 23626 3777
rect 23570 3703 23626 3712
rect 23112 2372 23164 2378
rect 23112 2314 23164 2320
rect 21178 54 21312 82
rect 23018 82 23074 480
rect 23124 82 23152 2314
rect 23018 54 23152 82
rect 13818 0 13874 54
rect 15658 0 15714 54
rect 17498 0 17554 54
rect 19338 0 19394 54
rect 21178 0 21234 54
rect 23018 0 23074 54
<< via2 >>
rect 110 22480 166 22536
rect 1766 19216 1822 19272
rect 1214 18808 1270 18864
rect 1398 16632 1454 16688
rect 1490 14184 1546 14240
rect 110 11872 166 11928
rect 110 9152 166 9208
rect 4956 21786 5012 21788
rect 5036 21786 5092 21788
rect 5116 21786 5172 21788
rect 5196 21786 5252 21788
rect 4956 21734 4982 21786
rect 4982 21734 5012 21786
rect 5036 21734 5046 21786
rect 5046 21734 5092 21786
rect 5116 21734 5162 21786
rect 5162 21734 5172 21786
rect 5196 21734 5226 21786
rect 5226 21734 5252 21786
rect 4956 21732 5012 21734
rect 5036 21732 5092 21734
rect 5116 21732 5172 21734
rect 5196 21732 5252 21734
rect 4956 20698 5012 20700
rect 5036 20698 5092 20700
rect 5116 20698 5172 20700
rect 5196 20698 5252 20700
rect 4956 20646 4982 20698
rect 4982 20646 5012 20698
rect 5036 20646 5046 20698
rect 5046 20646 5092 20698
rect 5116 20646 5162 20698
rect 5162 20646 5172 20698
rect 5196 20646 5226 20698
rect 5226 20646 5252 20698
rect 4956 20644 5012 20646
rect 5036 20644 5092 20646
rect 5116 20644 5172 20646
rect 5196 20644 5252 20646
rect 4956 19610 5012 19612
rect 5036 19610 5092 19612
rect 5116 19610 5172 19612
rect 5196 19610 5252 19612
rect 4956 19558 4982 19610
rect 4982 19558 5012 19610
rect 5036 19558 5046 19610
rect 5046 19558 5092 19610
rect 5116 19558 5162 19610
rect 5162 19558 5172 19610
rect 5196 19558 5226 19610
rect 5226 19558 5252 19610
rect 4956 19556 5012 19558
rect 5036 19556 5092 19558
rect 5116 19556 5172 19558
rect 5196 19556 5252 19558
rect 4956 18522 5012 18524
rect 5036 18522 5092 18524
rect 5116 18522 5172 18524
rect 5196 18522 5252 18524
rect 4956 18470 4982 18522
rect 4982 18470 5012 18522
rect 5036 18470 5046 18522
rect 5046 18470 5092 18522
rect 5116 18470 5162 18522
rect 5162 18470 5172 18522
rect 5196 18470 5226 18522
rect 5226 18470 5252 18522
rect 4956 18468 5012 18470
rect 5036 18468 5092 18470
rect 5116 18468 5172 18470
rect 5196 18468 5252 18470
rect 4956 17434 5012 17436
rect 5036 17434 5092 17436
rect 5116 17434 5172 17436
rect 5196 17434 5252 17436
rect 4956 17382 4982 17434
rect 4982 17382 5012 17434
rect 5036 17382 5046 17434
rect 5046 17382 5092 17434
rect 5116 17382 5162 17434
rect 5162 17382 5172 17434
rect 5196 17382 5226 17434
rect 5226 17382 5252 17434
rect 4956 17380 5012 17382
rect 5036 17380 5092 17382
rect 5116 17380 5172 17382
rect 5196 17380 5252 17382
rect 8956 21242 9012 21244
rect 9036 21242 9092 21244
rect 9116 21242 9172 21244
rect 9196 21242 9252 21244
rect 8956 21190 8982 21242
rect 8982 21190 9012 21242
rect 9036 21190 9046 21242
rect 9046 21190 9092 21242
rect 9116 21190 9162 21242
rect 9162 21190 9172 21242
rect 9196 21190 9226 21242
rect 9226 21190 9252 21242
rect 8956 21188 9012 21190
rect 9036 21188 9092 21190
rect 9116 21188 9172 21190
rect 9196 21188 9252 21190
rect 8956 20154 9012 20156
rect 9036 20154 9092 20156
rect 9116 20154 9172 20156
rect 9196 20154 9252 20156
rect 8956 20102 8982 20154
rect 8982 20102 9012 20154
rect 9036 20102 9046 20154
rect 9046 20102 9092 20154
rect 9116 20102 9162 20154
rect 9162 20102 9172 20154
rect 9196 20102 9226 20154
rect 9226 20102 9252 20154
rect 8956 20100 9012 20102
rect 9036 20100 9092 20102
rect 9116 20100 9172 20102
rect 9196 20100 9252 20102
rect 8956 19066 9012 19068
rect 9036 19066 9092 19068
rect 9116 19066 9172 19068
rect 9196 19066 9252 19068
rect 8956 19014 8982 19066
rect 8982 19014 9012 19066
rect 9036 19014 9046 19066
rect 9046 19014 9092 19066
rect 9116 19014 9162 19066
rect 9162 19014 9172 19066
rect 9196 19014 9226 19066
rect 9226 19014 9252 19066
rect 8956 19012 9012 19014
rect 9036 19012 9092 19014
rect 9116 19012 9172 19014
rect 9196 19012 9252 19014
rect 8390 18672 8446 18728
rect 8956 17978 9012 17980
rect 9036 17978 9092 17980
rect 9116 17978 9172 17980
rect 9196 17978 9252 17980
rect 8956 17926 8982 17978
rect 8982 17926 9012 17978
rect 9036 17926 9046 17978
rect 9046 17926 9092 17978
rect 9116 17926 9162 17978
rect 9162 17926 9172 17978
rect 9196 17926 9226 17978
rect 9226 17926 9252 17978
rect 8956 17924 9012 17926
rect 9036 17924 9092 17926
rect 9116 17924 9172 17926
rect 9196 17924 9252 17926
rect 8956 16890 9012 16892
rect 9036 16890 9092 16892
rect 9116 16890 9172 16892
rect 9196 16890 9252 16892
rect 8956 16838 8982 16890
rect 8982 16838 9012 16890
rect 9036 16838 9046 16890
rect 9046 16838 9092 16890
rect 9116 16838 9162 16890
rect 9162 16838 9172 16890
rect 9196 16838 9226 16890
rect 9226 16838 9252 16890
rect 8956 16836 9012 16838
rect 9036 16836 9092 16838
rect 9116 16836 9172 16838
rect 9196 16836 9252 16838
rect 7746 16652 7802 16688
rect 7746 16632 7748 16652
rect 7748 16632 7800 16652
rect 7800 16632 7802 16652
rect 4956 16346 5012 16348
rect 5036 16346 5092 16348
rect 5116 16346 5172 16348
rect 5196 16346 5252 16348
rect 4956 16294 4982 16346
rect 4982 16294 5012 16346
rect 5036 16294 5046 16346
rect 5046 16294 5092 16346
rect 5116 16294 5162 16346
rect 5162 16294 5172 16346
rect 5196 16294 5226 16346
rect 5226 16294 5252 16346
rect 4956 16292 5012 16294
rect 5036 16292 5092 16294
rect 5116 16292 5172 16294
rect 5196 16292 5252 16294
rect 4956 15258 5012 15260
rect 5036 15258 5092 15260
rect 5116 15258 5172 15260
rect 5196 15258 5252 15260
rect 4956 15206 4982 15258
rect 4982 15206 5012 15258
rect 5036 15206 5046 15258
rect 5046 15206 5092 15258
rect 5116 15206 5162 15258
rect 5162 15206 5172 15258
rect 5196 15206 5226 15258
rect 5226 15206 5252 15258
rect 4956 15204 5012 15206
rect 5036 15204 5092 15206
rect 5116 15204 5172 15206
rect 5196 15204 5252 15206
rect 11426 18808 11482 18864
rect 8956 15802 9012 15804
rect 9036 15802 9092 15804
rect 9116 15802 9172 15804
rect 9196 15802 9252 15804
rect 8956 15750 8982 15802
rect 8982 15750 9012 15802
rect 9036 15750 9046 15802
rect 9046 15750 9092 15802
rect 9116 15750 9162 15802
rect 9162 15750 9172 15802
rect 9196 15750 9226 15802
rect 9226 15750 9252 15802
rect 8956 15748 9012 15750
rect 9036 15748 9092 15750
rect 9116 15748 9172 15750
rect 9196 15748 9252 15750
rect 4956 14170 5012 14172
rect 5036 14170 5092 14172
rect 5116 14170 5172 14172
rect 5196 14170 5252 14172
rect 4956 14118 4982 14170
rect 4982 14118 5012 14170
rect 5036 14118 5046 14170
rect 5046 14118 5092 14170
rect 5116 14118 5162 14170
rect 5162 14118 5172 14170
rect 5196 14118 5226 14170
rect 5226 14118 5252 14170
rect 4956 14116 5012 14118
rect 5036 14116 5092 14118
rect 5116 14116 5172 14118
rect 5196 14116 5252 14118
rect 4956 13082 5012 13084
rect 5036 13082 5092 13084
rect 5116 13082 5172 13084
rect 5196 13082 5252 13084
rect 4956 13030 4982 13082
rect 4982 13030 5012 13082
rect 5036 13030 5046 13082
rect 5046 13030 5092 13082
rect 5116 13030 5162 13082
rect 5162 13030 5172 13082
rect 5196 13030 5226 13082
rect 5226 13030 5252 13082
rect 4956 13028 5012 13030
rect 5036 13028 5092 13030
rect 5116 13028 5172 13030
rect 5196 13028 5252 13030
rect 4956 11994 5012 11996
rect 5036 11994 5092 11996
rect 5116 11994 5172 11996
rect 5196 11994 5252 11996
rect 4956 11942 4982 11994
rect 4982 11942 5012 11994
rect 5036 11942 5046 11994
rect 5046 11942 5092 11994
rect 5116 11942 5162 11994
rect 5162 11942 5172 11994
rect 5196 11942 5226 11994
rect 5226 11942 5252 11994
rect 4956 11940 5012 11942
rect 5036 11940 5092 11942
rect 5116 11940 5172 11942
rect 5196 11940 5252 11942
rect 4956 10906 5012 10908
rect 5036 10906 5092 10908
rect 5116 10906 5172 10908
rect 5196 10906 5252 10908
rect 4956 10854 4982 10906
rect 4982 10854 5012 10906
rect 5036 10854 5046 10906
rect 5046 10854 5092 10906
rect 5116 10854 5162 10906
rect 5162 10854 5172 10906
rect 5196 10854 5226 10906
rect 5226 10854 5252 10906
rect 4956 10852 5012 10854
rect 5036 10852 5092 10854
rect 5116 10852 5172 10854
rect 5196 10852 5252 10854
rect 4956 9818 5012 9820
rect 5036 9818 5092 9820
rect 5116 9818 5172 9820
rect 5196 9818 5252 9820
rect 4956 9766 4982 9818
rect 4982 9766 5012 9818
rect 5036 9766 5046 9818
rect 5046 9766 5092 9818
rect 5116 9766 5162 9818
rect 5162 9766 5172 9818
rect 5196 9766 5226 9818
rect 5226 9766 5252 9818
rect 4956 9764 5012 9766
rect 5036 9764 5092 9766
rect 5116 9764 5172 9766
rect 5196 9764 5252 9766
rect 8956 14714 9012 14716
rect 9036 14714 9092 14716
rect 9116 14714 9172 14716
rect 9196 14714 9252 14716
rect 8956 14662 8982 14714
rect 8982 14662 9012 14714
rect 9036 14662 9046 14714
rect 9046 14662 9092 14714
rect 9116 14662 9162 14714
rect 9162 14662 9172 14714
rect 9196 14662 9226 14714
rect 9226 14662 9252 14714
rect 8956 14660 9012 14662
rect 9036 14660 9092 14662
rect 9116 14660 9172 14662
rect 9196 14660 9252 14662
rect 8956 13626 9012 13628
rect 9036 13626 9092 13628
rect 9116 13626 9172 13628
rect 9196 13626 9252 13628
rect 8956 13574 8982 13626
rect 8982 13574 9012 13626
rect 9036 13574 9046 13626
rect 9046 13574 9092 13626
rect 9116 13574 9162 13626
rect 9162 13574 9172 13626
rect 9196 13574 9226 13626
rect 9226 13574 9252 13626
rect 8956 13572 9012 13574
rect 9036 13572 9092 13574
rect 9116 13572 9172 13574
rect 9196 13572 9252 13574
rect 8956 12538 9012 12540
rect 9036 12538 9092 12540
rect 9116 12538 9172 12540
rect 9196 12538 9252 12540
rect 8956 12486 8982 12538
rect 8982 12486 9012 12538
rect 9036 12486 9046 12538
rect 9046 12486 9092 12538
rect 9116 12486 9162 12538
rect 9162 12486 9172 12538
rect 9196 12486 9226 12538
rect 9226 12486 9252 12538
rect 8956 12484 9012 12486
rect 9036 12484 9092 12486
rect 9116 12484 9172 12486
rect 9196 12484 9252 12486
rect 8956 11450 9012 11452
rect 9036 11450 9092 11452
rect 9116 11450 9172 11452
rect 9196 11450 9252 11452
rect 8956 11398 8982 11450
rect 8982 11398 9012 11450
rect 9036 11398 9046 11450
rect 9046 11398 9092 11450
rect 9116 11398 9162 11450
rect 9162 11398 9172 11450
rect 9196 11398 9226 11450
rect 9226 11398 9252 11450
rect 8956 11396 9012 11398
rect 9036 11396 9092 11398
rect 9116 11396 9172 11398
rect 9196 11396 9252 11398
rect 4956 8730 5012 8732
rect 5036 8730 5092 8732
rect 5116 8730 5172 8732
rect 5196 8730 5252 8732
rect 4956 8678 4982 8730
rect 4982 8678 5012 8730
rect 5036 8678 5046 8730
rect 5046 8678 5092 8730
rect 5116 8678 5162 8730
rect 5162 8678 5172 8730
rect 5196 8678 5226 8730
rect 5226 8678 5252 8730
rect 4956 8676 5012 8678
rect 5036 8676 5092 8678
rect 5116 8676 5172 8678
rect 5196 8676 5252 8678
rect 2042 7928 2098 7984
rect 4956 7642 5012 7644
rect 5036 7642 5092 7644
rect 5116 7642 5172 7644
rect 5196 7642 5252 7644
rect 4956 7590 4982 7642
rect 4982 7590 5012 7642
rect 5036 7590 5046 7642
rect 5046 7590 5092 7642
rect 5116 7590 5162 7642
rect 5162 7590 5172 7642
rect 5196 7590 5226 7642
rect 5226 7590 5252 7642
rect 4956 7588 5012 7590
rect 5036 7588 5092 7590
rect 5116 7588 5172 7590
rect 5196 7588 5252 7590
rect 110 3848 166 3904
rect 4956 6554 5012 6556
rect 5036 6554 5092 6556
rect 5116 6554 5172 6556
rect 5196 6554 5252 6556
rect 4956 6502 4982 6554
rect 4982 6502 5012 6554
rect 5036 6502 5046 6554
rect 5046 6502 5092 6554
rect 5116 6502 5162 6554
rect 5162 6502 5172 6554
rect 5196 6502 5226 6554
rect 5226 6502 5252 6554
rect 4956 6500 5012 6502
rect 5036 6500 5092 6502
rect 5116 6500 5172 6502
rect 5196 6500 5252 6502
rect 4956 5466 5012 5468
rect 5036 5466 5092 5468
rect 5116 5466 5172 5468
rect 5196 5466 5252 5468
rect 4956 5414 4982 5466
rect 4982 5414 5012 5466
rect 5036 5414 5046 5466
rect 5046 5414 5092 5466
rect 5116 5414 5162 5466
rect 5162 5414 5172 5466
rect 5196 5414 5226 5466
rect 5226 5414 5252 5466
rect 4956 5412 5012 5414
rect 5036 5412 5092 5414
rect 5116 5412 5172 5414
rect 5196 5412 5252 5414
rect 4956 4378 5012 4380
rect 5036 4378 5092 4380
rect 5116 4378 5172 4380
rect 5196 4378 5252 4380
rect 4956 4326 4982 4378
rect 4982 4326 5012 4378
rect 5036 4326 5046 4378
rect 5046 4326 5092 4378
rect 5116 4326 5162 4378
rect 5162 4326 5172 4378
rect 5196 4326 5226 4378
rect 5226 4326 5252 4378
rect 4956 4324 5012 4326
rect 5036 4324 5092 4326
rect 5116 4324 5172 4326
rect 5196 4324 5252 4326
rect 4956 3290 5012 3292
rect 5036 3290 5092 3292
rect 5116 3290 5172 3292
rect 5196 3290 5252 3292
rect 4956 3238 4982 3290
rect 4982 3238 5012 3290
rect 5036 3238 5046 3290
rect 5046 3238 5092 3290
rect 5116 3238 5162 3290
rect 5162 3238 5172 3290
rect 5196 3238 5226 3290
rect 5226 3238 5252 3290
rect 4956 3236 5012 3238
rect 5036 3236 5092 3238
rect 5116 3236 5172 3238
rect 5196 3236 5252 3238
rect 4956 2202 5012 2204
rect 5036 2202 5092 2204
rect 5116 2202 5172 2204
rect 5196 2202 5252 2204
rect 4956 2150 4982 2202
rect 4982 2150 5012 2202
rect 5036 2150 5046 2202
rect 5046 2150 5092 2202
rect 5116 2150 5162 2202
rect 5162 2150 5172 2202
rect 5196 2150 5226 2202
rect 5226 2150 5252 2202
rect 4956 2148 5012 2150
rect 5036 2148 5092 2150
rect 5116 2148 5172 2150
rect 5196 2148 5252 2150
rect 6550 1808 6606 1864
rect 8956 10362 9012 10364
rect 9036 10362 9092 10364
rect 9116 10362 9172 10364
rect 9196 10362 9252 10364
rect 8956 10310 8982 10362
rect 8982 10310 9012 10362
rect 9036 10310 9046 10362
rect 9046 10310 9092 10362
rect 9116 10310 9162 10362
rect 9162 10310 9172 10362
rect 9196 10310 9226 10362
rect 9226 10310 9252 10362
rect 8956 10308 9012 10310
rect 9036 10308 9092 10310
rect 9116 10308 9172 10310
rect 9196 10308 9252 10310
rect 8956 9274 9012 9276
rect 9036 9274 9092 9276
rect 9116 9274 9172 9276
rect 9196 9274 9252 9276
rect 8956 9222 8982 9274
rect 8982 9222 9012 9274
rect 9036 9222 9046 9274
rect 9046 9222 9092 9274
rect 9116 9222 9162 9274
rect 9162 9222 9172 9274
rect 9196 9222 9226 9274
rect 9226 9222 9252 9274
rect 8956 9220 9012 9222
rect 9036 9220 9092 9222
rect 9116 9220 9172 9222
rect 9196 9220 9252 9222
rect 8956 8186 9012 8188
rect 9036 8186 9092 8188
rect 9116 8186 9172 8188
rect 9196 8186 9252 8188
rect 8956 8134 8982 8186
rect 8982 8134 9012 8186
rect 9036 8134 9046 8186
rect 9046 8134 9092 8186
rect 9116 8134 9162 8186
rect 9162 8134 9172 8186
rect 9196 8134 9226 8186
rect 9226 8134 9252 8186
rect 8956 8132 9012 8134
rect 9036 8132 9092 8134
rect 9116 8132 9172 8134
rect 9196 8132 9252 8134
rect 8666 7248 8722 7304
rect 8956 7098 9012 7100
rect 9036 7098 9092 7100
rect 9116 7098 9172 7100
rect 9196 7098 9252 7100
rect 8956 7046 8982 7098
rect 8982 7046 9012 7098
rect 9036 7046 9046 7098
rect 9046 7046 9092 7098
rect 9116 7046 9162 7098
rect 9162 7046 9172 7098
rect 9196 7046 9226 7098
rect 9226 7046 9252 7098
rect 8956 7044 9012 7046
rect 9036 7044 9092 7046
rect 9116 7044 9172 7046
rect 9196 7044 9252 7046
rect 8956 6010 9012 6012
rect 9036 6010 9092 6012
rect 9116 6010 9172 6012
rect 9196 6010 9252 6012
rect 8956 5958 8982 6010
rect 8982 5958 9012 6010
rect 9036 5958 9046 6010
rect 9046 5958 9092 6010
rect 9116 5958 9162 6010
rect 9162 5958 9172 6010
rect 9196 5958 9226 6010
rect 9226 5958 9252 6010
rect 8956 5956 9012 5958
rect 9036 5956 9092 5958
rect 9116 5956 9172 5958
rect 9196 5956 9252 5958
rect 8956 4922 9012 4924
rect 9036 4922 9092 4924
rect 9116 4922 9172 4924
rect 9196 4922 9252 4924
rect 8956 4870 8982 4922
rect 8982 4870 9012 4922
rect 9036 4870 9046 4922
rect 9046 4870 9092 4922
rect 9116 4870 9162 4922
rect 9162 4870 9172 4922
rect 9196 4870 9226 4922
rect 9226 4870 9252 4922
rect 8956 4868 9012 4870
rect 9036 4868 9092 4870
rect 9116 4868 9172 4870
rect 9196 4868 9252 4870
rect 10046 6160 10102 6216
rect 8022 1944 8078 2000
rect 9402 4120 9458 4176
rect 12956 21786 13012 21788
rect 13036 21786 13092 21788
rect 13116 21786 13172 21788
rect 13196 21786 13252 21788
rect 12956 21734 12982 21786
rect 12982 21734 13012 21786
rect 13036 21734 13046 21786
rect 13046 21734 13092 21786
rect 13116 21734 13162 21786
rect 13162 21734 13172 21786
rect 13196 21734 13226 21786
rect 13226 21734 13252 21786
rect 12956 21732 13012 21734
rect 13036 21732 13092 21734
rect 13116 21732 13172 21734
rect 13196 21732 13252 21734
rect 12956 20698 13012 20700
rect 13036 20698 13092 20700
rect 13116 20698 13172 20700
rect 13196 20698 13252 20700
rect 12956 20646 12982 20698
rect 12982 20646 13012 20698
rect 13036 20646 13046 20698
rect 13046 20646 13092 20698
rect 13116 20646 13162 20698
rect 13162 20646 13172 20698
rect 13196 20646 13226 20698
rect 13226 20646 13252 20698
rect 12956 20644 13012 20646
rect 13036 20644 13092 20646
rect 13116 20644 13172 20646
rect 13196 20644 13252 20646
rect 12956 19610 13012 19612
rect 13036 19610 13092 19612
rect 13116 19610 13172 19612
rect 13196 19610 13252 19612
rect 12956 19558 12982 19610
rect 12982 19558 13012 19610
rect 13036 19558 13046 19610
rect 13046 19558 13092 19610
rect 13116 19558 13162 19610
rect 13162 19558 13172 19610
rect 13196 19558 13226 19610
rect 13226 19558 13252 19610
rect 12956 19556 13012 19558
rect 13036 19556 13092 19558
rect 13116 19556 13172 19558
rect 13196 19556 13252 19558
rect 12956 18522 13012 18524
rect 13036 18522 13092 18524
rect 13116 18522 13172 18524
rect 13196 18522 13252 18524
rect 12956 18470 12982 18522
rect 12982 18470 13012 18522
rect 13036 18470 13046 18522
rect 13046 18470 13092 18522
rect 13116 18470 13162 18522
rect 13162 18470 13172 18522
rect 13196 18470 13226 18522
rect 13226 18470 13252 18522
rect 12956 18468 13012 18470
rect 13036 18468 13092 18470
rect 13116 18468 13172 18470
rect 13196 18468 13252 18470
rect 12956 17434 13012 17436
rect 13036 17434 13092 17436
rect 13116 17434 13172 17436
rect 13196 17434 13252 17436
rect 12956 17382 12982 17434
rect 12982 17382 13012 17434
rect 13036 17382 13046 17434
rect 13046 17382 13092 17434
rect 13116 17382 13162 17434
rect 13162 17382 13172 17434
rect 13196 17382 13226 17434
rect 13226 17382 13252 17434
rect 12956 17380 13012 17382
rect 13036 17380 13092 17382
rect 13116 17380 13172 17382
rect 13196 17380 13252 17382
rect 12956 16346 13012 16348
rect 13036 16346 13092 16348
rect 13116 16346 13172 16348
rect 13196 16346 13252 16348
rect 12956 16294 12982 16346
rect 12982 16294 13012 16346
rect 13036 16294 13046 16346
rect 13046 16294 13092 16346
rect 13116 16294 13162 16346
rect 13162 16294 13172 16346
rect 13196 16294 13226 16346
rect 13226 16294 13252 16346
rect 12956 16292 13012 16294
rect 13036 16292 13092 16294
rect 13116 16292 13172 16294
rect 13196 16292 13252 16294
rect 12956 15258 13012 15260
rect 13036 15258 13092 15260
rect 13116 15258 13172 15260
rect 13196 15258 13252 15260
rect 12956 15206 12982 15258
rect 12982 15206 13012 15258
rect 13036 15206 13046 15258
rect 13046 15206 13092 15258
rect 13116 15206 13162 15258
rect 13162 15206 13172 15258
rect 13196 15206 13226 15258
rect 13226 15206 13252 15258
rect 12956 15204 13012 15206
rect 13036 15204 13092 15206
rect 13116 15204 13172 15206
rect 13196 15204 13252 15206
rect 12956 14170 13012 14172
rect 13036 14170 13092 14172
rect 13116 14170 13172 14172
rect 13196 14170 13252 14172
rect 12956 14118 12982 14170
rect 12982 14118 13012 14170
rect 13036 14118 13046 14170
rect 13046 14118 13092 14170
rect 13116 14118 13162 14170
rect 13162 14118 13172 14170
rect 13196 14118 13226 14170
rect 13226 14118 13252 14170
rect 12956 14116 13012 14118
rect 13036 14116 13092 14118
rect 13116 14116 13172 14118
rect 13196 14116 13252 14118
rect 12956 13082 13012 13084
rect 13036 13082 13092 13084
rect 13116 13082 13172 13084
rect 13196 13082 13252 13084
rect 12956 13030 12982 13082
rect 12982 13030 13012 13082
rect 13036 13030 13046 13082
rect 13046 13030 13092 13082
rect 13116 13030 13162 13082
rect 13162 13030 13172 13082
rect 13196 13030 13226 13082
rect 13226 13030 13252 13082
rect 12956 13028 13012 13030
rect 13036 13028 13092 13030
rect 13116 13028 13172 13030
rect 13196 13028 13252 13030
rect 12956 11994 13012 11996
rect 13036 11994 13092 11996
rect 13116 11994 13172 11996
rect 13196 11994 13252 11996
rect 12956 11942 12982 11994
rect 12982 11942 13012 11994
rect 13036 11942 13046 11994
rect 13046 11942 13092 11994
rect 13116 11942 13162 11994
rect 13162 11942 13172 11994
rect 13196 11942 13226 11994
rect 13226 11942 13252 11994
rect 12956 11940 13012 11942
rect 13036 11940 13092 11942
rect 13116 11940 13172 11942
rect 13196 11940 13252 11942
rect 12956 10906 13012 10908
rect 13036 10906 13092 10908
rect 13116 10906 13172 10908
rect 13196 10906 13252 10908
rect 12956 10854 12982 10906
rect 12982 10854 13012 10906
rect 13036 10854 13046 10906
rect 13046 10854 13092 10906
rect 13116 10854 13162 10906
rect 13162 10854 13172 10906
rect 13196 10854 13226 10906
rect 13226 10854 13252 10906
rect 12956 10852 13012 10854
rect 13036 10852 13092 10854
rect 13116 10852 13172 10854
rect 13196 10852 13252 10854
rect 12956 9818 13012 9820
rect 13036 9818 13092 9820
rect 13116 9818 13172 9820
rect 13196 9818 13252 9820
rect 12956 9766 12982 9818
rect 12982 9766 13012 9818
rect 13036 9766 13046 9818
rect 13046 9766 13092 9818
rect 13116 9766 13162 9818
rect 13162 9766 13172 9818
rect 13196 9766 13226 9818
rect 13226 9766 13252 9818
rect 12956 9764 13012 9766
rect 13036 9764 13092 9766
rect 13116 9764 13172 9766
rect 13196 9764 13252 9766
rect 8956 3834 9012 3836
rect 9036 3834 9092 3836
rect 9116 3834 9172 3836
rect 9196 3834 9252 3836
rect 8956 3782 8982 3834
rect 8982 3782 9012 3834
rect 9036 3782 9046 3834
rect 9046 3782 9092 3834
rect 9116 3782 9162 3834
rect 9162 3782 9172 3834
rect 9196 3782 9226 3834
rect 9226 3782 9252 3834
rect 8956 3780 9012 3782
rect 9036 3780 9092 3782
rect 9116 3780 9172 3782
rect 9196 3780 9252 3782
rect 8956 2746 9012 2748
rect 9036 2746 9092 2748
rect 9116 2746 9172 2748
rect 9196 2746 9252 2748
rect 8956 2694 8982 2746
rect 8982 2694 9012 2746
rect 9036 2694 9046 2746
rect 9046 2694 9092 2746
rect 9116 2694 9162 2746
rect 9162 2694 9172 2746
rect 9196 2694 9226 2746
rect 9226 2694 9252 2746
rect 8956 2692 9012 2694
rect 9036 2692 9092 2694
rect 9116 2692 9172 2694
rect 9196 2692 9252 2694
rect 12956 8730 13012 8732
rect 13036 8730 13092 8732
rect 13116 8730 13172 8732
rect 13196 8730 13252 8732
rect 12956 8678 12982 8730
rect 12982 8678 13012 8730
rect 13036 8678 13046 8730
rect 13046 8678 13092 8730
rect 13116 8678 13162 8730
rect 13162 8678 13172 8730
rect 13196 8678 13226 8730
rect 13226 8678 13252 8730
rect 12956 8676 13012 8678
rect 13036 8676 13092 8678
rect 13116 8676 13172 8678
rect 13196 8676 13252 8678
rect 12956 7642 13012 7644
rect 13036 7642 13092 7644
rect 13116 7642 13172 7644
rect 13196 7642 13252 7644
rect 12956 7590 12982 7642
rect 12982 7590 13012 7642
rect 13036 7590 13046 7642
rect 13046 7590 13092 7642
rect 13116 7590 13162 7642
rect 13162 7590 13172 7642
rect 13196 7590 13226 7642
rect 13226 7590 13252 7642
rect 12956 7588 13012 7590
rect 13036 7588 13092 7590
rect 13116 7588 13172 7590
rect 13196 7588 13252 7590
rect 12956 6554 13012 6556
rect 13036 6554 13092 6556
rect 13116 6554 13172 6556
rect 13196 6554 13252 6556
rect 12956 6502 12982 6554
rect 12982 6502 13012 6554
rect 13036 6502 13046 6554
rect 13046 6502 13092 6554
rect 13116 6502 13162 6554
rect 13162 6502 13172 6554
rect 13196 6502 13226 6554
rect 13226 6502 13252 6554
rect 12956 6500 13012 6502
rect 13036 6500 13092 6502
rect 13116 6500 13172 6502
rect 13196 6500 13252 6502
rect 12956 5466 13012 5468
rect 13036 5466 13092 5468
rect 13116 5466 13172 5468
rect 13196 5466 13252 5468
rect 12956 5414 12982 5466
rect 12982 5414 13012 5466
rect 13036 5414 13046 5466
rect 13046 5414 13092 5466
rect 13116 5414 13162 5466
rect 13162 5414 13172 5466
rect 13196 5414 13226 5466
rect 13226 5414 13252 5466
rect 12956 5412 13012 5414
rect 13036 5412 13092 5414
rect 13116 5412 13172 5414
rect 13196 5412 13252 5414
rect 12956 4378 13012 4380
rect 13036 4378 13092 4380
rect 13116 4378 13172 4380
rect 13196 4378 13252 4380
rect 12956 4326 12982 4378
rect 12982 4326 13012 4378
rect 13036 4326 13046 4378
rect 13046 4326 13092 4378
rect 13116 4326 13162 4378
rect 13162 4326 13172 4378
rect 13196 4326 13226 4378
rect 13226 4326 13252 4378
rect 12956 4324 13012 4326
rect 13036 4324 13092 4326
rect 13116 4324 13172 4326
rect 13196 4324 13252 4326
rect 12956 3290 13012 3292
rect 13036 3290 13092 3292
rect 13116 3290 13172 3292
rect 13196 3290 13252 3292
rect 12956 3238 12982 3290
rect 12982 3238 13012 3290
rect 13036 3238 13046 3290
rect 13046 3238 13092 3290
rect 13116 3238 13162 3290
rect 13162 3238 13172 3290
rect 13196 3238 13226 3290
rect 13226 3238 13252 3290
rect 12956 3236 13012 3238
rect 13036 3236 13092 3238
rect 13116 3236 13172 3238
rect 13196 3236 13252 3238
rect 12956 2202 13012 2204
rect 13036 2202 13092 2204
rect 13116 2202 13172 2204
rect 13196 2202 13252 2204
rect 12956 2150 12982 2202
rect 12982 2150 13012 2202
rect 13036 2150 13046 2202
rect 13046 2150 13092 2202
rect 13116 2150 13162 2202
rect 13162 2150 13172 2202
rect 13196 2150 13226 2202
rect 13226 2150 13252 2202
rect 12956 2148 13012 2150
rect 13036 2148 13092 2150
rect 13116 2148 13172 2150
rect 13196 2148 13252 2150
rect 11794 1536 11850 1592
rect 16394 13912 16450 13968
rect 15474 12144 15530 12200
rect 15290 7928 15346 7984
rect 13818 1264 13874 1320
rect 18326 22616 18382 22672
rect 16956 21242 17012 21244
rect 17036 21242 17092 21244
rect 17116 21242 17172 21244
rect 17196 21242 17252 21244
rect 16956 21190 16982 21242
rect 16982 21190 17012 21242
rect 17036 21190 17046 21242
rect 17046 21190 17092 21242
rect 17116 21190 17162 21242
rect 17162 21190 17172 21242
rect 17196 21190 17226 21242
rect 17226 21190 17252 21242
rect 16956 21188 17012 21190
rect 17036 21188 17092 21190
rect 17116 21188 17172 21190
rect 17196 21188 17252 21190
rect 16956 20154 17012 20156
rect 17036 20154 17092 20156
rect 17116 20154 17172 20156
rect 17196 20154 17252 20156
rect 16956 20102 16982 20154
rect 16982 20102 17012 20154
rect 17036 20102 17046 20154
rect 17046 20102 17092 20154
rect 17116 20102 17162 20154
rect 17162 20102 17172 20154
rect 17196 20102 17226 20154
rect 17226 20102 17252 20154
rect 16956 20100 17012 20102
rect 17036 20100 17092 20102
rect 17116 20100 17172 20102
rect 17196 20100 17252 20102
rect 16956 19066 17012 19068
rect 17036 19066 17092 19068
rect 17116 19066 17172 19068
rect 17196 19066 17252 19068
rect 16956 19014 16982 19066
rect 16982 19014 17012 19066
rect 17036 19014 17046 19066
rect 17046 19014 17092 19066
rect 17116 19014 17162 19066
rect 17162 19014 17172 19066
rect 17196 19014 17226 19066
rect 17226 19014 17252 19066
rect 16956 19012 17012 19014
rect 17036 19012 17092 19014
rect 17116 19012 17172 19014
rect 17196 19012 17252 19014
rect 16762 18128 16818 18184
rect 16956 17978 17012 17980
rect 17036 17978 17092 17980
rect 17116 17978 17172 17980
rect 17196 17978 17252 17980
rect 16956 17926 16982 17978
rect 16982 17926 17012 17978
rect 17036 17926 17046 17978
rect 17046 17926 17092 17978
rect 17116 17926 17162 17978
rect 17162 17926 17172 17978
rect 17196 17926 17226 17978
rect 17226 17926 17252 17978
rect 16956 17924 17012 17926
rect 17036 17924 17092 17926
rect 17116 17924 17172 17926
rect 17196 17924 17252 17926
rect 16956 16890 17012 16892
rect 17036 16890 17092 16892
rect 17116 16890 17172 16892
rect 17196 16890 17252 16892
rect 16956 16838 16982 16890
rect 16982 16838 17012 16890
rect 17036 16838 17046 16890
rect 17046 16838 17092 16890
rect 17116 16838 17162 16890
rect 17162 16838 17172 16890
rect 17196 16838 17226 16890
rect 17226 16838 17252 16890
rect 16956 16836 17012 16838
rect 17036 16836 17092 16838
rect 17116 16836 17172 16838
rect 17196 16836 17252 16838
rect 16956 15802 17012 15804
rect 17036 15802 17092 15804
rect 17116 15802 17172 15804
rect 17196 15802 17252 15804
rect 16956 15750 16982 15802
rect 16982 15750 17012 15802
rect 17036 15750 17046 15802
rect 17046 15750 17092 15802
rect 17116 15750 17162 15802
rect 17162 15750 17172 15802
rect 17196 15750 17226 15802
rect 17226 15750 17252 15802
rect 16956 15748 17012 15750
rect 17036 15748 17092 15750
rect 17116 15748 17172 15750
rect 17196 15748 17252 15750
rect 16956 14714 17012 14716
rect 17036 14714 17092 14716
rect 17116 14714 17172 14716
rect 17196 14714 17252 14716
rect 16956 14662 16982 14714
rect 16982 14662 17012 14714
rect 17036 14662 17046 14714
rect 17046 14662 17092 14714
rect 17116 14662 17162 14714
rect 17162 14662 17172 14714
rect 17196 14662 17226 14714
rect 17226 14662 17252 14714
rect 16956 14660 17012 14662
rect 17036 14660 17092 14662
rect 17116 14660 17172 14662
rect 17196 14660 17252 14662
rect 20956 21786 21012 21788
rect 21036 21786 21092 21788
rect 21116 21786 21172 21788
rect 21196 21786 21252 21788
rect 20956 21734 20982 21786
rect 20982 21734 21012 21786
rect 21036 21734 21046 21786
rect 21046 21734 21092 21786
rect 21116 21734 21162 21786
rect 21162 21734 21172 21786
rect 21196 21734 21226 21786
rect 21226 21734 21252 21786
rect 20956 21732 21012 21734
rect 21036 21732 21092 21734
rect 21116 21732 21172 21734
rect 21196 21732 21252 21734
rect 21362 21120 21418 21176
rect 20956 20698 21012 20700
rect 21036 20698 21092 20700
rect 21116 20698 21172 20700
rect 21196 20698 21252 20700
rect 20956 20646 20982 20698
rect 20982 20646 21012 20698
rect 21036 20646 21046 20698
rect 21046 20646 21092 20698
rect 21116 20646 21162 20698
rect 21162 20646 21172 20698
rect 21196 20646 21226 20698
rect 21226 20646 21252 20698
rect 20956 20644 21012 20646
rect 21036 20644 21092 20646
rect 21116 20644 21172 20646
rect 21196 20644 21252 20646
rect 20956 19610 21012 19612
rect 21036 19610 21092 19612
rect 21116 19610 21172 19612
rect 21196 19610 21252 19612
rect 20956 19558 20982 19610
rect 20982 19558 21012 19610
rect 21036 19558 21046 19610
rect 21046 19558 21092 19610
rect 21116 19558 21162 19610
rect 21162 19558 21172 19610
rect 21196 19558 21226 19610
rect 21226 19558 21252 19610
rect 20956 19556 21012 19558
rect 21036 19556 21092 19558
rect 21116 19556 21172 19558
rect 21196 19556 21252 19558
rect 20810 18672 20866 18728
rect 20956 18522 21012 18524
rect 21036 18522 21092 18524
rect 21116 18522 21172 18524
rect 21196 18522 21252 18524
rect 20956 18470 20982 18522
rect 20982 18470 21012 18522
rect 21036 18470 21046 18522
rect 21046 18470 21092 18522
rect 21116 18470 21162 18522
rect 21162 18470 21172 18522
rect 21196 18470 21226 18522
rect 21226 18470 21252 18522
rect 20956 18468 21012 18470
rect 21036 18468 21092 18470
rect 21116 18468 21172 18470
rect 21196 18468 21252 18470
rect 20956 17434 21012 17436
rect 21036 17434 21092 17436
rect 21116 17434 21172 17436
rect 21196 17434 21252 17436
rect 20956 17382 20982 17434
rect 20982 17382 21012 17434
rect 21036 17382 21046 17434
rect 21046 17382 21092 17434
rect 21116 17382 21162 17434
rect 21162 17382 21172 17434
rect 21196 17382 21226 17434
rect 21226 17382 21252 17434
rect 20956 17380 21012 17382
rect 21036 17380 21092 17382
rect 21116 17380 21172 17382
rect 21196 17380 21252 17382
rect 20956 16346 21012 16348
rect 21036 16346 21092 16348
rect 21116 16346 21172 16348
rect 21196 16346 21252 16348
rect 20956 16294 20982 16346
rect 20982 16294 21012 16346
rect 21036 16294 21046 16346
rect 21046 16294 21092 16346
rect 21116 16294 21162 16346
rect 21162 16294 21172 16346
rect 21196 16294 21226 16346
rect 21226 16294 21252 16346
rect 20956 16292 21012 16294
rect 21036 16292 21092 16294
rect 21116 16292 21172 16294
rect 21196 16292 21252 16294
rect 21270 15408 21326 15464
rect 20956 15258 21012 15260
rect 21036 15258 21092 15260
rect 21116 15258 21172 15260
rect 21196 15258 21252 15260
rect 20956 15206 20982 15258
rect 20982 15206 21012 15258
rect 21036 15206 21046 15258
rect 21046 15206 21092 15258
rect 21116 15206 21162 15258
rect 21162 15206 21172 15258
rect 21196 15206 21226 15258
rect 21226 15206 21252 15258
rect 20956 15204 21012 15206
rect 21036 15204 21092 15206
rect 21116 15204 21172 15206
rect 21196 15204 21252 15206
rect 16956 13626 17012 13628
rect 17036 13626 17092 13628
rect 17116 13626 17172 13628
rect 17196 13626 17252 13628
rect 16956 13574 16982 13626
rect 16982 13574 17012 13626
rect 17036 13574 17046 13626
rect 17046 13574 17092 13626
rect 17116 13574 17162 13626
rect 17162 13574 17172 13626
rect 17196 13574 17226 13626
rect 17226 13574 17252 13626
rect 16956 13572 17012 13574
rect 17036 13572 17092 13574
rect 17116 13572 17172 13574
rect 17196 13572 17252 13574
rect 16956 12538 17012 12540
rect 17036 12538 17092 12540
rect 17116 12538 17172 12540
rect 17196 12538 17252 12540
rect 16956 12486 16982 12538
rect 16982 12486 17012 12538
rect 17036 12486 17046 12538
rect 17046 12486 17092 12538
rect 17116 12486 17162 12538
rect 17162 12486 17172 12538
rect 17196 12486 17226 12538
rect 17226 12486 17252 12538
rect 16956 12484 17012 12486
rect 17036 12484 17092 12486
rect 17116 12484 17172 12486
rect 17196 12484 17252 12486
rect 20956 14170 21012 14172
rect 21036 14170 21092 14172
rect 21116 14170 21172 14172
rect 21196 14170 21252 14172
rect 20956 14118 20982 14170
rect 20982 14118 21012 14170
rect 21036 14118 21046 14170
rect 21046 14118 21092 14170
rect 21116 14118 21162 14170
rect 21162 14118 21172 14170
rect 21196 14118 21226 14170
rect 21226 14118 21252 14170
rect 20956 14116 21012 14118
rect 21036 14116 21092 14118
rect 21116 14116 21172 14118
rect 21196 14116 21252 14118
rect 21546 19624 21602 19680
rect 20956 13082 21012 13084
rect 21036 13082 21092 13084
rect 21116 13082 21172 13084
rect 21196 13082 21252 13084
rect 20956 13030 20982 13082
rect 20982 13030 21012 13082
rect 21036 13030 21046 13082
rect 21046 13030 21092 13082
rect 21116 13030 21162 13082
rect 21162 13030 21172 13082
rect 21196 13030 21226 13082
rect 21226 13030 21252 13082
rect 20956 13028 21012 13030
rect 21036 13028 21092 13030
rect 21116 13028 21172 13030
rect 21196 13028 21252 13030
rect 16956 11450 17012 11452
rect 17036 11450 17092 11452
rect 17116 11450 17172 11452
rect 17196 11450 17252 11452
rect 16956 11398 16982 11450
rect 16982 11398 17012 11450
rect 17036 11398 17046 11450
rect 17046 11398 17092 11450
rect 17116 11398 17162 11450
rect 17162 11398 17172 11450
rect 17196 11398 17226 11450
rect 17226 11398 17252 11450
rect 16956 11396 17012 11398
rect 17036 11396 17092 11398
rect 17116 11396 17172 11398
rect 17196 11396 17252 11398
rect 20956 11994 21012 11996
rect 21036 11994 21092 11996
rect 21116 11994 21172 11996
rect 21196 11994 21252 11996
rect 20956 11942 20982 11994
rect 20982 11942 21012 11994
rect 21036 11942 21046 11994
rect 21046 11942 21092 11994
rect 21116 11942 21162 11994
rect 21162 11942 21172 11994
rect 21196 11942 21226 11994
rect 21226 11942 21252 11994
rect 20956 11940 21012 11942
rect 21036 11940 21092 11942
rect 21116 11940 21172 11942
rect 21196 11940 21252 11942
rect 16956 10362 17012 10364
rect 17036 10362 17092 10364
rect 17116 10362 17172 10364
rect 17196 10362 17252 10364
rect 16956 10310 16982 10362
rect 16982 10310 17012 10362
rect 17036 10310 17046 10362
rect 17046 10310 17092 10362
rect 17116 10310 17162 10362
rect 17162 10310 17172 10362
rect 17196 10310 17226 10362
rect 17226 10310 17252 10362
rect 16956 10308 17012 10310
rect 17036 10308 17092 10310
rect 17116 10308 17172 10310
rect 17196 10308 17252 10310
rect 16956 9274 17012 9276
rect 17036 9274 17092 9276
rect 17116 9274 17172 9276
rect 17196 9274 17252 9276
rect 16956 9222 16982 9274
rect 16982 9222 17012 9274
rect 17036 9222 17046 9274
rect 17046 9222 17092 9274
rect 17116 9222 17162 9274
rect 17162 9222 17172 9274
rect 17196 9222 17226 9274
rect 17226 9222 17252 9274
rect 16956 9220 17012 9222
rect 17036 9220 17092 9222
rect 17116 9220 17172 9222
rect 17196 9220 17252 9222
rect 16956 8186 17012 8188
rect 17036 8186 17092 8188
rect 17116 8186 17172 8188
rect 17196 8186 17252 8188
rect 16956 8134 16982 8186
rect 16982 8134 17012 8186
rect 17036 8134 17046 8186
rect 17046 8134 17092 8186
rect 17116 8134 17162 8186
rect 17162 8134 17172 8186
rect 17196 8134 17226 8186
rect 17226 8134 17252 8186
rect 16956 8132 17012 8134
rect 17036 8132 17092 8134
rect 17116 8132 17172 8134
rect 17196 8132 17252 8134
rect 16956 7098 17012 7100
rect 17036 7098 17092 7100
rect 17116 7098 17172 7100
rect 17196 7098 17252 7100
rect 16956 7046 16982 7098
rect 16982 7046 17012 7098
rect 17036 7046 17046 7098
rect 17046 7046 17092 7098
rect 17116 7046 17162 7098
rect 17162 7046 17172 7098
rect 17196 7046 17226 7098
rect 17226 7046 17252 7098
rect 16956 7044 17012 7046
rect 17036 7044 17092 7046
rect 17116 7044 17172 7046
rect 17196 7044 17252 7046
rect 20956 10906 21012 10908
rect 21036 10906 21092 10908
rect 21116 10906 21172 10908
rect 21196 10906 21252 10908
rect 20956 10854 20982 10906
rect 20982 10854 21012 10906
rect 21036 10854 21046 10906
rect 21046 10854 21092 10906
rect 21116 10854 21162 10906
rect 21162 10854 21172 10906
rect 21196 10854 21226 10906
rect 21226 10854 21252 10906
rect 20956 10852 21012 10854
rect 21036 10852 21092 10854
rect 21116 10852 21172 10854
rect 21196 10852 21252 10854
rect 20956 9818 21012 9820
rect 21036 9818 21092 9820
rect 21116 9818 21172 9820
rect 21196 9818 21252 9820
rect 20956 9766 20982 9818
rect 20982 9766 21012 9818
rect 21036 9766 21046 9818
rect 21046 9766 21092 9818
rect 21116 9766 21162 9818
rect 21162 9766 21172 9818
rect 21196 9766 21226 9818
rect 21226 9766 21252 9818
rect 20956 9764 21012 9766
rect 21036 9764 21092 9766
rect 21116 9764 21172 9766
rect 21196 9764 21252 9766
rect 21362 10784 21418 10840
rect 21362 9696 21418 9752
rect 17958 7248 18014 7304
rect 16956 6010 17012 6012
rect 17036 6010 17092 6012
rect 17116 6010 17172 6012
rect 17196 6010 17252 6012
rect 16956 5958 16982 6010
rect 16982 5958 17012 6010
rect 17036 5958 17046 6010
rect 17046 5958 17092 6010
rect 17116 5958 17162 6010
rect 17162 5958 17172 6010
rect 17196 5958 17226 6010
rect 17226 5958 17252 6010
rect 16956 5956 17012 5958
rect 17036 5956 17092 5958
rect 17116 5956 17172 5958
rect 17196 5956 17252 5958
rect 16956 4922 17012 4924
rect 17036 4922 17092 4924
rect 17116 4922 17172 4924
rect 17196 4922 17252 4924
rect 16956 4870 16982 4922
rect 16982 4870 17012 4922
rect 17036 4870 17046 4922
rect 17046 4870 17092 4922
rect 17116 4870 17162 4922
rect 17162 4870 17172 4922
rect 17196 4870 17226 4922
rect 17226 4870 17252 4922
rect 16956 4868 17012 4870
rect 17036 4868 17092 4870
rect 17116 4868 17172 4870
rect 17196 4868 17252 4870
rect 16956 3834 17012 3836
rect 17036 3834 17092 3836
rect 17116 3834 17172 3836
rect 17196 3834 17252 3836
rect 16956 3782 16982 3834
rect 16982 3782 17012 3834
rect 17036 3782 17046 3834
rect 17046 3782 17092 3834
rect 17116 3782 17162 3834
rect 17162 3782 17172 3834
rect 17196 3782 17226 3834
rect 17226 3782 17252 3834
rect 16956 3780 17012 3782
rect 17036 3780 17092 3782
rect 17116 3780 17172 3782
rect 17196 3780 17252 3782
rect 16956 2746 17012 2748
rect 17036 2746 17092 2748
rect 17116 2746 17172 2748
rect 17196 2746 17252 2748
rect 16956 2694 16982 2746
rect 16982 2694 17012 2746
rect 17036 2694 17046 2746
rect 17046 2694 17092 2746
rect 17116 2694 17162 2746
rect 17162 2694 17172 2746
rect 17196 2694 17226 2746
rect 17226 2694 17252 2746
rect 16956 2692 17012 2694
rect 17036 2692 17092 2694
rect 17116 2692 17172 2694
rect 17196 2692 17252 2694
rect 20956 8730 21012 8732
rect 21036 8730 21092 8732
rect 21116 8730 21172 8732
rect 21196 8730 21252 8732
rect 20956 8678 20982 8730
rect 20982 8678 21012 8730
rect 21036 8678 21046 8730
rect 21046 8678 21092 8730
rect 21116 8678 21162 8730
rect 21162 8678 21172 8730
rect 21196 8678 21226 8730
rect 21226 8678 21252 8730
rect 20956 8676 21012 8678
rect 21036 8676 21092 8678
rect 21116 8676 21172 8678
rect 21196 8676 21252 8678
rect 20956 7642 21012 7644
rect 21036 7642 21092 7644
rect 21116 7642 21172 7644
rect 21196 7642 21252 7644
rect 20956 7590 20982 7642
rect 20982 7590 21012 7642
rect 21036 7590 21046 7642
rect 21046 7590 21092 7642
rect 21116 7590 21162 7642
rect 21162 7590 21172 7642
rect 21196 7590 21226 7642
rect 21226 7590 21252 7642
rect 20956 7588 21012 7590
rect 21036 7588 21092 7590
rect 21116 7588 21172 7590
rect 21196 7588 21252 7590
rect 20956 6554 21012 6556
rect 21036 6554 21092 6556
rect 21116 6554 21172 6556
rect 21196 6554 21252 6556
rect 20956 6502 20982 6554
rect 20982 6502 21012 6554
rect 21036 6502 21046 6554
rect 21046 6502 21092 6554
rect 21116 6502 21162 6554
rect 21162 6502 21172 6554
rect 21196 6502 21226 6554
rect 21226 6502 21252 6554
rect 20956 6500 21012 6502
rect 21036 6500 21092 6502
rect 21116 6500 21172 6502
rect 21196 6500 21252 6502
rect 18326 6180 18382 6216
rect 18326 6160 18328 6180
rect 18328 6160 18380 6180
rect 18380 6160 18382 6180
rect 20956 5466 21012 5468
rect 21036 5466 21092 5468
rect 21116 5466 21172 5468
rect 21196 5466 21252 5468
rect 20956 5414 20982 5466
rect 20982 5414 21012 5466
rect 21036 5414 21046 5466
rect 21046 5414 21092 5466
rect 21116 5414 21162 5466
rect 21162 5414 21172 5466
rect 21196 5414 21226 5466
rect 21226 5414 21252 5466
rect 20956 5412 21012 5414
rect 21036 5412 21092 5414
rect 21116 5412 21172 5414
rect 21196 5412 21252 5414
rect 20956 4378 21012 4380
rect 21036 4378 21092 4380
rect 21116 4378 21172 4380
rect 21196 4378 21252 4380
rect 20956 4326 20982 4378
rect 20982 4326 21012 4378
rect 21036 4326 21046 4378
rect 21046 4326 21092 4378
rect 21116 4326 21162 4378
rect 21162 4326 21172 4378
rect 21196 4326 21226 4378
rect 21226 4326 21252 4378
rect 20956 4324 21012 4326
rect 21036 4324 21092 4326
rect 21116 4324 21172 4326
rect 21196 4324 21252 4326
rect 20956 3290 21012 3292
rect 21036 3290 21092 3292
rect 21116 3290 21172 3292
rect 21196 3290 21252 3292
rect 20956 3238 20982 3290
rect 20982 3238 21012 3290
rect 21036 3238 21046 3290
rect 21046 3238 21092 3290
rect 21116 3238 21162 3290
rect 21162 3238 21172 3290
rect 21196 3238 21226 3290
rect 21226 3238 21252 3290
rect 20956 3236 21012 3238
rect 21036 3236 21092 3238
rect 21116 3236 21172 3238
rect 21196 3236 21252 3238
rect 20956 2202 21012 2204
rect 21036 2202 21092 2204
rect 21116 2202 21172 2204
rect 21196 2202 21252 2204
rect 20956 2150 20982 2202
rect 20982 2150 21012 2202
rect 21036 2150 21046 2202
rect 21046 2150 21092 2202
rect 21116 2150 21162 2202
rect 21162 2150 21172 2202
rect 21196 2150 21226 2202
rect 21226 2150 21252 2202
rect 20956 2148 21012 2150
rect 21036 2148 21092 2150
rect 21116 2148 21172 2150
rect 21196 2148 21252 2150
rect 19890 1944 19946 2000
rect 23570 5208 23626 5264
rect 23570 4120 23626 4176
rect 23570 3712 23626 3768
<< metal3 >>
rect 23520 23128 24000 23248
rect 18321 22674 18387 22677
rect 23614 22674 23674 23128
rect 18321 22672 23674 22674
rect 18321 22616 18326 22672
rect 18382 22616 23674 22672
rect 18321 22614 23674 22616
rect 18321 22611 18387 22614
rect 0 22536 480 22568
rect 0 22480 110 22536
rect 166 22480 480 22536
rect 0 22448 480 22480
rect 4944 21792 5264 21793
rect 4944 21728 4952 21792
rect 5016 21728 5032 21792
rect 5096 21728 5112 21792
rect 5176 21728 5192 21792
rect 5256 21728 5264 21792
rect 4944 21727 5264 21728
rect 12944 21792 13264 21793
rect 12944 21728 12952 21792
rect 13016 21728 13032 21792
rect 13096 21728 13112 21792
rect 13176 21728 13192 21792
rect 13256 21728 13264 21792
rect 12944 21727 13264 21728
rect 20944 21792 21264 21793
rect 20944 21728 20952 21792
rect 21016 21728 21032 21792
rect 21096 21728 21112 21792
rect 21176 21728 21192 21792
rect 21256 21728 21264 21792
rect 20944 21727 21264 21728
rect 23520 21632 24000 21752
rect 8944 21248 9264 21249
rect 8944 21184 8952 21248
rect 9016 21184 9032 21248
rect 9096 21184 9112 21248
rect 9176 21184 9192 21248
rect 9256 21184 9264 21248
rect 8944 21183 9264 21184
rect 16944 21248 17264 21249
rect 16944 21184 16952 21248
rect 17016 21184 17032 21248
rect 17096 21184 17112 21248
rect 17176 21184 17192 21248
rect 17256 21184 17264 21248
rect 16944 21183 17264 21184
rect 21357 21178 21423 21181
rect 23614 21178 23674 21632
rect 21357 21176 23674 21178
rect 21357 21120 21362 21176
rect 21418 21120 23674 21176
rect 21357 21118 23674 21120
rect 21357 21115 21423 21118
rect 4944 20704 5264 20705
rect 4944 20640 4952 20704
rect 5016 20640 5032 20704
rect 5096 20640 5112 20704
rect 5176 20640 5192 20704
rect 5256 20640 5264 20704
rect 4944 20639 5264 20640
rect 12944 20704 13264 20705
rect 12944 20640 12952 20704
rect 13016 20640 13032 20704
rect 13096 20640 13112 20704
rect 13176 20640 13192 20704
rect 13256 20640 13264 20704
rect 12944 20639 13264 20640
rect 20944 20704 21264 20705
rect 20944 20640 20952 20704
rect 21016 20640 21032 20704
rect 21096 20640 21112 20704
rect 21176 20640 21192 20704
rect 21256 20640 21264 20704
rect 20944 20639 21264 20640
rect 8944 20160 9264 20161
rect 8944 20096 8952 20160
rect 9016 20096 9032 20160
rect 9096 20096 9112 20160
rect 9176 20096 9192 20160
rect 9256 20096 9264 20160
rect 8944 20095 9264 20096
rect 16944 20160 17264 20161
rect 16944 20096 16952 20160
rect 17016 20096 17032 20160
rect 17096 20096 17112 20160
rect 17176 20096 17192 20160
rect 17256 20096 17264 20160
rect 23520 20136 24000 20256
rect 16944 20095 17264 20096
rect 0 19728 480 19848
rect 62 19274 122 19728
rect 21541 19682 21607 19685
rect 23614 19682 23674 20136
rect 21541 19680 23674 19682
rect 21541 19624 21546 19680
rect 21602 19624 23674 19680
rect 21541 19622 23674 19624
rect 21541 19619 21607 19622
rect 4944 19616 5264 19617
rect 4944 19552 4952 19616
rect 5016 19552 5032 19616
rect 5096 19552 5112 19616
rect 5176 19552 5192 19616
rect 5256 19552 5264 19616
rect 4944 19551 5264 19552
rect 12944 19616 13264 19617
rect 12944 19552 12952 19616
rect 13016 19552 13032 19616
rect 13096 19552 13112 19616
rect 13176 19552 13192 19616
rect 13256 19552 13264 19616
rect 12944 19551 13264 19552
rect 20944 19616 21264 19617
rect 20944 19552 20952 19616
rect 21016 19552 21032 19616
rect 21096 19552 21112 19616
rect 21176 19552 21192 19616
rect 21256 19552 21264 19616
rect 20944 19551 21264 19552
rect 1761 19274 1827 19277
rect 62 19272 1827 19274
rect 62 19216 1766 19272
rect 1822 19216 1827 19272
rect 62 19214 1827 19216
rect 1761 19211 1827 19214
rect 8944 19072 9264 19073
rect 8944 19008 8952 19072
rect 9016 19008 9032 19072
rect 9096 19008 9112 19072
rect 9176 19008 9192 19072
rect 9256 19008 9264 19072
rect 8944 19007 9264 19008
rect 16944 19072 17264 19073
rect 16944 19008 16952 19072
rect 17016 19008 17032 19072
rect 17096 19008 17112 19072
rect 17176 19008 17192 19072
rect 17256 19008 17264 19072
rect 16944 19007 17264 19008
rect 1209 18866 1275 18869
rect 11421 18866 11487 18869
rect 1209 18864 11487 18866
rect 1209 18808 1214 18864
rect 1270 18808 11426 18864
rect 11482 18808 11487 18864
rect 1209 18806 11487 18808
rect 1209 18803 1275 18806
rect 11421 18803 11487 18806
rect 8385 18730 8451 18733
rect 20805 18730 20871 18733
rect 8385 18728 20871 18730
rect 8385 18672 8390 18728
rect 8446 18672 20810 18728
rect 20866 18672 20871 18728
rect 8385 18670 20871 18672
rect 8385 18667 8451 18670
rect 20805 18667 20871 18670
rect 23520 18640 24000 18760
rect 4944 18528 5264 18529
rect 4944 18464 4952 18528
rect 5016 18464 5032 18528
rect 5096 18464 5112 18528
rect 5176 18464 5192 18528
rect 5256 18464 5264 18528
rect 4944 18463 5264 18464
rect 12944 18528 13264 18529
rect 12944 18464 12952 18528
rect 13016 18464 13032 18528
rect 13096 18464 13112 18528
rect 13176 18464 13192 18528
rect 13256 18464 13264 18528
rect 12944 18463 13264 18464
rect 20944 18528 21264 18529
rect 20944 18464 20952 18528
rect 21016 18464 21032 18528
rect 21096 18464 21112 18528
rect 21176 18464 21192 18528
rect 21256 18464 21264 18528
rect 20944 18463 21264 18464
rect 16757 18186 16823 18189
rect 23614 18186 23674 18640
rect 16757 18184 23674 18186
rect 16757 18128 16762 18184
rect 16818 18128 23674 18184
rect 16757 18126 23674 18128
rect 16757 18123 16823 18126
rect 8944 17984 9264 17985
rect 8944 17920 8952 17984
rect 9016 17920 9032 17984
rect 9096 17920 9112 17984
rect 9176 17920 9192 17984
rect 9256 17920 9264 17984
rect 8944 17919 9264 17920
rect 16944 17984 17264 17985
rect 16944 17920 16952 17984
rect 17016 17920 17032 17984
rect 17096 17920 17112 17984
rect 17176 17920 17192 17984
rect 17256 17920 17264 17984
rect 16944 17919 17264 17920
rect 4944 17440 5264 17441
rect 4944 17376 4952 17440
rect 5016 17376 5032 17440
rect 5096 17376 5112 17440
rect 5176 17376 5192 17440
rect 5256 17376 5264 17440
rect 4944 17375 5264 17376
rect 12944 17440 13264 17441
rect 12944 17376 12952 17440
rect 13016 17376 13032 17440
rect 13096 17376 13112 17440
rect 13176 17376 13192 17440
rect 13256 17376 13264 17440
rect 12944 17375 13264 17376
rect 20944 17440 21264 17441
rect 20944 17376 20952 17440
rect 21016 17376 21032 17440
rect 21096 17376 21112 17440
rect 21176 17376 21192 17440
rect 21256 17376 21264 17440
rect 20944 17375 21264 17376
rect 0 17144 480 17264
rect 23520 17144 24000 17264
rect 62 16690 122 17144
rect 8944 16896 9264 16897
rect 8944 16832 8952 16896
rect 9016 16832 9032 16896
rect 9096 16832 9112 16896
rect 9176 16832 9192 16896
rect 9256 16832 9264 16896
rect 8944 16831 9264 16832
rect 16944 16896 17264 16897
rect 16944 16832 16952 16896
rect 17016 16832 17032 16896
rect 17096 16832 17112 16896
rect 17176 16832 17192 16896
rect 17256 16832 17264 16896
rect 16944 16831 17264 16832
rect 1393 16690 1459 16693
rect 62 16688 1459 16690
rect 62 16632 1398 16688
rect 1454 16632 1459 16688
rect 62 16630 1459 16632
rect 1393 16627 1459 16630
rect 7741 16690 7807 16693
rect 23614 16690 23674 17144
rect 7741 16688 23674 16690
rect 7741 16632 7746 16688
rect 7802 16632 23674 16688
rect 7741 16630 23674 16632
rect 7741 16627 7807 16630
rect 4944 16352 5264 16353
rect 4944 16288 4952 16352
rect 5016 16288 5032 16352
rect 5096 16288 5112 16352
rect 5176 16288 5192 16352
rect 5256 16288 5264 16352
rect 4944 16287 5264 16288
rect 12944 16352 13264 16353
rect 12944 16288 12952 16352
rect 13016 16288 13032 16352
rect 13096 16288 13112 16352
rect 13176 16288 13192 16352
rect 13256 16288 13264 16352
rect 12944 16287 13264 16288
rect 20944 16352 21264 16353
rect 20944 16288 20952 16352
rect 21016 16288 21032 16352
rect 21096 16288 21112 16352
rect 21176 16288 21192 16352
rect 21256 16288 21264 16352
rect 20944 16287 21264 16288
rect 8944 15808 9264 15809
rect 8944 15744 8952 15808
rect 9016 15744 9032 15808
rect 9096 15744 9112 15808
rect 9176 15744 9192 15808
rect 9256 15744 9264 15808
rect 8944 15743 9264 15744
rect 16944 15808 17264 15809
rect 16944 15744 16952 15808
rect 17016 15744 17032 15808
rect 17096 15744 17112 15808
rect 17176 15744 17192 15808
rect 17256 15744 17264 15808
rect 16944 15743 17264 15744
rect 23520 15648 24000 15768
rect 21265 15466 21331 15469
rect 23614 15466 23674 15648
rect 21265 15464 23674 15466
rect 21265 15408 21270 15464
rect 21326 15408 23674 15464
rect 21265 15406 23674 15408
rect 21265 15403 21331 15406
rect 4944 15264 5264 15265
rect 4944 15200 4952 15264
rect 5016 15200 5032 15264
rect 5096 15200 5112 15264
rect 5176 15200 5192 15264
rect 5256 15200 5264 15264
rect 4944 15199 5264 15200
rect 12944 15264 13264 15265
rect 12944 15200 12952 15264
rect 13016 15200 13032 15264
rect 13096 15200 13112 15264
rect 13176 15200 13192 15264
rect 13256 15200 13264 15264
rect 12944 15199 13264 15200
rect 20944 15264 21264 15265
rect 20944 15200 20952 15264
rect 21016 15200 21032 15264
rect 21096 15200 21112 15264
rect 21176 15200 21192 15264
rect 21256 15200 21264 15264
rect 20944 15199 21264 15200
rect 8944 14720 9264 14721
rect 8944 14656 8952 14720
rect 9016 14656 9032 14720
rect 9096 14656 9112 14720
rect 9176 14656 9192 14720
rect 9256 14656 9264 14720
rect 8944 14655 9264 14656
rect 16944 14720 17264 14721
rect 16944 14656 16952 14720
rect 17016 14656 17032 14720
rect 17096 14656 17112 14720
rect 17176 14656 17192 14720
rect 17256 14656 17264 14720
rect 16944 14655 17264 14656
rect 0 14424 480 14544
rect 62 14242 122 14424
rect 1485 14242 1551 14245
rect 62 14240 1551 14242
rect 62 14184 1490 14240
rect 1546 14184 1551 14240
rect 62 14182 1551 14184
rect 1485 14179 1551 14182
rect 4944 14176 5264 14177
rect 4944 14112 4952 14176
rect 5016 14112 5032 14176
rect 5096 14112 5112 14176
rect 5176 14112 5192 14176
rect 5256 14112 5264 14176
rect 4944 14111 5264 14112
rect 12944 14176 13264 14177
rect 12944 14112 12952 14176
rect 13016 14112 13032 14176
rect 13096 14112 13112 14176
rect 13176 14112 13192 14176
rect 13256 14112 13264 14176
rect 12944 14111 13264 14112
rect 20944 14176 21264 14177
rect 20944 14112 20952 14176
rect 21016 14112 21032 14176
rect 21096 14112 21112 14176
rect 21176 14112 21192 14176
rect 21256 14112 21264 14176
rect 23520 14152 24000 14272
rect 20944 14111 21264 14112
rect 16389 13970 16455 13973
rect 23614 13970 23674 14152
rect 16389 13968 23674 13970
rect 16389 13912 16394 13968
rect 16450 13912 23674 13968
rect 16389 13910 23674 13912
rect 16389 13907 16455 13910
rect 8944 13632 9264 13633
rect 8944 13568 8952 13632
rect 9016 13568 9032 13632
rect 9096 13568 9112 13632
rect 9176 13568 9192 13632
rect 9256 13568 9264 13632
rect 8944 13567 9264 13568
rect 16944 13632 17264 13633
rect 16944 13568 16952 13632
rect 17016 13568 17032 13632
rect 17096 13568 17112 13632
rect 17176 13568 17192 13632
rect 17256 13568 17264 13632
rect 16944 13567 17264 13568
rect 4944 13088 5264 13089
rect 4944 13024 4952 13088
rect 5016 13024 5032 13088
rect 5096 13024 5112 13088
rect 5176 13024 5192 13088
rect 5256 13024 5264 13088
rect 4944 13023 5264 13024
rect 12944 13088 13264 13089
rect 12944 13024 12952 13088
rect 13016 13024 13032 13088
rect 13096 13024 13112 13088
rect 13176 13024 13192 13088
rect 13256 13024 13264 13088
rect 12944 13023 13264 13024
rect 20944 13088 21264 13089
rect 20944 13024 20952 13088
rect 21016 13024 21032 13088
rect 21096 13024 21112 13088
rect 21176 13024 21192 13088
rect 21256 13024 21264 13088
rect 20944 13023 21264 13024
rect 23520 12656 24000 12776
rect 8944 12544 9264 12545
rect 8944 12480 8952 12544
rect 9016 12480 9032 12544
rect 9096 12480 9112 12544
rect 9176 12480 9192 12544
rect 9256 12480 9264 12544
rect 8944 12479 9264 12480
rect 16944 12544 17264 12545
rect 16944 12480 16952 12544
rect 17016 12480 17032 12544
rect 17096 12480 17112 12544
rect 17176 12480 17192 12544
rect 17256 12480 17264 12544
rect 16944 12479 17264 12480
rect 15469 12202 15535 12205
rect 23614 12202 23674 12656
rect 15469 12200 23674 12202
rect 15469 12144 15474 12200
rect 15530 12144 23674 12200
rect 15469 12142 23674 12144
rect 15469 12139 15535 12142
rect 4944 12000 5264 12001
rect 0 11928 480 11960
rect 4944 11936 4952 12000
rect 5016 11936 5032 12000
rect 5096 11936 5112 12000
rect 5176 11936 5192 12000
rect 5256 11936 5264 12000
rect 4944 11935 5264 11936
rect 12944 12000 13264 12001
rect 12944 11936 12952 12000
rect 13016 11936 13032 12000
rect 13096 11936 13112 12000
rect 13176 11936 13192 12000
rect 13256 11936 13264 12000
rect 12944 11935 13264 11936
rect 20944 12000 21264 12001
rect 20944 11936 20952 12000
rect 21016 11936 21032 12000
rect 21096 11936 21112 12000
rect 21176 11936 21192 12000
rect 21256 11936 21264 12000
rect 20944 11935 21264 11936
rect 0 11872 110 11928
rect 166 11872 480 11928
rect 0 11840 480 11872
rect 8944 11456 9264 11457
rect 8944 11392 8952 11456
rect 9016 11392 9032 11456
rect 9096 11392 9112 11456
rect 9176 11392 9192 11456
rect 9256 11392 9264 11456
rect 8944 11391 9264 11392
rect 16944 11456 17264 11457
rect 16944 11392 16952 11456
rect 17016 11392 17032 11456
rect 17096 11392 17112 11456
rect 17176 11392 17192 11456
rect 17256 11392 17264 11456
rect 16944 11391 17264 11392
rect 23520 11160 24000 11280
rect 4944 10912 5264 10913
rect 4944 10848 4952 10912
rect 5016 10848 5032 10912
rect 5096 10848 5112 10912
rect 5176 10848 5192 10912
rect 5256 10848 5264 10912
rect 4944 10847 5264 10848
rect 12944 10912 13264 10913
rect 12944 10848 12952 10912
rect 13016 10848 13032 10912
rect 13096 10848 13112 10912
rect 13176 10848 13192 10912
rect 13256 10848 13264 10912
rect 12944 10847 13264 10848
rect 20944 10912 21264 10913
rect 20944 10848 20952 10912
rect 21016 10848 21032 10912
rect 21096 10848 21112 10912
rect 21176 10848 21192 10912
rect 21256 10848 21264 10912
rect 20944 10847 21264 10848
rect 21357 10842 21423 10845
rect 23614 10842 23674 11160
rect 21357 10840 23674 10842
rect 21357 10784 21362 10840
rect 21418 10784 23674 10840
rect 21357 10782 23674 10784
rect 21357 10779 21423 10782
rect 8944 10368 9264 10369
rect 8944 10304 8952 10368
rect 9016 10304 9032 10368
rect 9096 10304 9112 10368
rect 9176 10304 9192 10368
rect 9256 10304 9264 10368
rect 8944 10303 9264 10304
rect 16944 10368 17264 10369
rect 16944 10304 16952 10368
rect 17016 10304 17032 10368
rect 17096 10304 17112 10368
rect 17176 10304 17192 10368
rect 17256 10304 17264 10368
rect 16944 10303 17264 10304
rect 4944 9824 5264 9825
rect 4944 9760 4952 9824
rect 5016 9760 5032 9824
rect 5096 9760 5112 9824
rect 5176 9760 5192 9824
rect 5256 9760 5264 9824
rect 4944 9759 5264 9760
rect 12944 9824 13264 9825
rect 12944 9760 12952 9824
rect 13016 9760 13032 9824
rect 13096 9760 13112 9824
rect 13176 9760 13192 9824
rect 13256 9760 13264 9824
rect 12944 9759 13264 9760
rect 20944 9824 21264 9825
rect 20944 9760 20952 9824
rect 21016 9760 21032 9824
rect 21096 9760 21112 9824
rect 21176 9760 21192 9824
rect 21256 9760 21264 9824
rect 20944 9759 21264 9760
rect 21357 9754 21423 9757
rect 23520 9754 24000 9784
rect 21357 9752 24000 9754
rect 21357 9696 21362 9752
rect 21418 9696 24000 9752
rect 21357 9694 24000 9696
rect 21357 9691 21423 9694
rect 23520 9664 24000 9694
rect 8944 9280 9264 9281
rect 0 9208 480 9240
rect 8944 9216 8952 9280
rect 9016 9216 9032 9280
rect 9096 9216 9112 9280
rect 9176 9216 9192 9280
rect 9256 9216 9264 9280
rect 8944 9215 9264 9216
rect 16944 9280 17264 9281
rect 16944 9216 16952 9280
rect 17016 9216 17032 9280
rect 17096 9216 17112 9280
rect 17176 9216 17192 9280
rect 17256 9216 17264 9280
rect 16944 9215 17264 9216
rect 0 9152 110 9208
rect 166 9152 480 9208
rect 0 9120 480 9152
rect 4944 8736 5264 8737
rect 4944 8672 4952 8736
rect 5016 8672 5032 8736
rect 5096 8672 5112 8736
rect 5176 8672 5192 8736
rect 5256 8672 5264 8736
rect 4944 8671 5264 8672
rect 12944 8736 13264 8737
rect 12944 8672 12952 8736
rect 13016 8672 13032 8736
rect 13096 8672 13112 8736
rect 13176 8672 13192 8736
rect 13256 8672 13264 8736
rect 12944 8671 13264 8672
rect 20944 8736 21264 8737
rect 20944 8672 20952 8736
rect 21016 8672 21032 8736
rect 21096 8672 21112 8736
rect 21176 8672 21192 8736
rect 21256 8672 21264 8736
rect 20944 8671 21264 8672
rect 8944 8192 9264 8193
rect 8944 8128 8952 8192
rect 9016 8128 9032 8192
rect 9096 8128 9112 8192
rect 9176 8128 9192 8192
rect 9256 8128 9264 8192
rect 8944 8127 9264 8128
rect 16944 8192 17264 8193
rect 16944 8128 16952 8192
rect 17016 8128 17032 8192
rect 17096 8128 17112 8192
rect 17176 8128 17192 8192
rect 17256 8128 17264 8192
rect 23520 8168 24000 8288
rect 16944 8127 17264 8128
rect 2037 7986 2103 7989
rect 15285 7986 15351 7989
rect 23614 7986 23674 8168
rect 2037 7984 23674 7986
rect 2037 7928 2042 7984
rect 2098 7928 15290 7984
rect 15346 7928 23674 7984
rect 2037 7926 23674 7928
rect 2037 7923 2103 7926
rect 15285 7923 15351 7926
rect 4944 7648 5264 7649
rect 4944 7584 4952 7648
rect 5016 7584 5032 7648
rect 5096 7584 5112 7648
rect 5176 7584 5192 7648
rect 5256 7584 5264 7648
rect 4944 7583 5264 7584
rect 12944 7648 13264 7649
rect 12944 7584 12952 7648
rect 13016 7584 13032 7648
rect 13096 7584 13112 7648
rect 13176 7584 13192 7648
rect 13256 7584 13264 7648
rect 12944 7583 13264 7584
rect 20944 7648 21264 7649
rect 20944 7584 20952 7648
rect 21016 7584 21032 7648
rect 21096 7584 21112 7648
rect 21176 7584 21192 7648
rect 21256 7584 21264 7648
rect 20944 7583 21264 7584
rect 8661 7306 8727 7309
rect 17953 7306 18019 7309
rect 8661 7304 18019 7306
rect 8661 7248 8666 7304
rect 8722 7248 17958 7304
rect 18014 7248 18019 7304
rect 8661 7246 18019 7248
rect 8661 7243 8727 7246
rect 17953 7243 18019 7246
rect 8944 7104 9264 7105
rect 8944 7040 8952 7104
rect 9016 7040 9032 7104
rect 9096 7040 9112 7104
rect 9176 7040 9192 7104
rect 9256 7040 9264 7104
rect 8944 7039 9264 7040
rect 16944 7104 17264 7105
rect 16944 7040 16952 7104
rect 17016 7040 17032 7104
rect 17096 7040 17112 7104
rect 17176 7040 17192 7104
rect 17256 7040 17264 7104
rect 16944 7039 17264 7040
rect 23520 6672 24000 6792
rect 0 6536 480 6656
rect 4944 6560 5264 6561
rect 62 6218 122 6536
rect 4944 6496 4952 6560
rect 5016 6496 5032 6560
rect 5096 6496 5112 6560
rect 5176 6496 5192 6560
rect 5256 6496 5264 6560
rect 4944 6495 5264 6496
rect 12944 6560 13264 6561
rect 12944 6496 12952 6560
rect 13016 6496 13032 6560
rect 13096 6496 13112 6560
rect 13176 6496 13192 6560
rect 13256 6496 13264 6560
rect 12944 6495 13264 6496
rect 20944 6560 21264 6561
rect 20944 6496 20952 6560
rect 21016 6496 21032 6560
rect 21096 6496 21112 6560
rect 21176 6496 21192 6560
rect 21256 6496 21264 6560
rect 20944 6495 21264 6496
rect 10041 6218 10107 6221
rect 62 6216 10107 6218
rect 62 6160 10046 6216
rect 10102 6160 10107 6216
rect 62 6158 10107 6160
rect 10041 6155 10107 6158
rect 18321 6218 18387 6221
rect 23614 6218 23674 6672
rect 18321 6216 23674 6218
rect 18321 6160 18326 6216
rect 18382 6160 23674 6216
rect 18321 6158 23674 6160
rect 18321 6155 18387 6158
rect 8944 6016 9264 6017
rect 8944 5952 8952 6016
rect 9016 5952 9032 6016
rect 9096 5952 9112 6016
rect 9176 5952 9192 6016
rect 9256 5952 9264 6016
rect 8944 5951 9264 5952
rect 16944 6016 17264 6017
rect 16944 5952 16952 6016
rect 17016 5952 17032 6016
rect 17096 5952 17112 6016
rect 17176 5952 17192 6016
rect 17256 5952 17264 6016
rect 16944 5951 17264 5952
rect 4944 5472 5264 5473
rect 4944 5408 4952 5472
rect 5016 5408 5032 5472
rect 5096 5408 5112 5472
rect 5176 5408 5192 5472
rect 5256 5408 5264 5472
rect 4944 5407 5264 5408
rect 12944 5472 13264 5473
rect 12944 5408 12952 5472
rect 13016 5408 13032 5472
rect 13096 5408 13112 5472
rect 13176 5408 13192 5472
rect 13256 5408 13264 5472
rect 12944 5407 13264 5408
rect 20944 5472 21264 5473
rect 20944 5408 20952 5472
rect 21016 5408 21032 5472
rect 21096 5408 21112 5472
rect 21176 5408 21192 5472
rect 21256 5408 21264 5472
rect 20944 5407 21264 5408
rect 23520 5266 24000 5296
rect 23484 5264 24000 5266
rect 23484 5208 23570 5264
rect 23626 5208 24000 5264
rect 23484 5206 24000 5208
rect 23520 5176 24000 5206
rect 8944 4928 9264 4929
rect 8944 4864 8952 4928
rect 9016 4864 9032 4928
rect 9096 4864 9112 4928
rect 9176 4864 9192 4928
rect 9256 4864 9264 4928
rect 8944 4863 9264 4864
rect 16944 4928 17264 4929
rect 16944 4864 16952 4928
rect 17016 4864 17032 4928
rect 17096 4864 17112 4928
rect 17176 4864 17192 4928
rect 17256 4864 17264 4928
rect 16944 4863 17264 4864
rect 4944 4384 5264 4385
rect 4944 4320 4952 4384
rect 5016 4320 5032 4384
rect 5096 4320 5112 4384
rect 5176 4320 5192 4384
rect 5256 4320 5264 4384
rect 4944 4319 5264 4320
rect 12944 4384 13264 4385
rect 12944 4320 12952 4384
rect 13016 4320 13032 4384
rect 13096 4320 13112 4384
rect 13176 4320 13192 4384
rect 13256 4320 13264 4384
rect 12944 4319 13264 4320
rect 20944 4384 21264 4385
rect 20944 4320 20952 4384
rect 21016 4320 21032 4384
rect 21096 4320 21112 4384
rect 21176 4320 21192 4384
rect 21256 4320 21264 4384
rect 20944 4319 21264 4320
rect 9397 4178 9463 4181
rect 23565 4178 23631 4181
rect 9397 4176 23631 4178
rect 9397 4120 9402 4176
rect 9458 4120 23570 4176
rect 23626 4120 23631 4176
rect 9397 4118 23631 4120
rect 9397 4115 9463 4118
rect 23565 4115 23631 4118
rect 0 3904 480 3936
rect 0 3848 110 3904
rect 166 3848 480 3904
rect 0 3816 480 3848
rect 8944 3840 9264 3841
rect 8944 3776 8952 3840
rect 9016 3776 9032 3840
rect 9096 3776 9112 3840
rect 9176 3776 9192 3840
rect 9256 3776 9264 3840
rect 8944 3775 9264 3776
rect 16944 3840 17264 3841
rect 16944 3776 16952 3840
rect 17016 3776 17032 3840
rect 17096 3776 17112 3840
rect 17176 3776 17192 3840
rect 17256 3776 17264 3840
rect 16944 3775 17264 3776
rect 23520 3770 24000 3800
rect 23484 3768 24000 3770
rect 23484 3712 23570 3768
rect 23626 3712 24000 3768
rect 23484 3710 24000 3712
rect 23520 3680 24000 3710
rect 4944 3296 5264 3297
rect 4944 3232 4952 3296
rect 5016 3232 5032 3296
rect 5096 3232 5112 3296
rect 5176 3232 5192 3296
rect 5256 3232 5264 3296
rect 4944 3231 5264 3232
rect 12944 3296 13264 3297
rect 12944 3232 12952 3296
rect 13016 3232 13032 3296
rect 13096 3232 13112 3296
rect 13176 3232 13192 3296
rect 13256 3232 13264 3296
rect 12944 3231 13264 3232
rect 20944 3296 21264 3297
rect 20944 3232 20952 3296
rect 21016 3232 21032 3296
rect 21096 3232 21112 3296
rect 21176 3232 21192 3296
rect 21256 3232 21264 3296
rect 20944 3231 21264 3232
rect 8944 2752 9264 2753
rect 8944 2688 8952 2752
rect 9016 2688 9032 2752
rect 9096 2688 9112 2752
rect 9176 2688 9192 2752
rect 9256 2688 9264 2752
rect 8944 2687 9264 2688
rect 16944 2752 17264 2753
rect 16944 2688 16952 2752
rect 17016 2688 17032 2752
rect 17096 2688 17112 2752
rect 17176 2688 17192 2752
rect 17256 2688 17264 2752
rect 16944 2687 17264 2688
rect 4944 2208 5264 2209
rect 4944 2144 4952 2208
rect 5016 2144 5032 2208
rect 5096 2144 5112 2208
rect 5176 2144 5192 2208
rect 5256 2144 5264 2208
rect 4944 2143 5264 2144
rect 12944 2208 13264 2209
rect 12944 2144 12952 2208
rect 13016 2144 13032 2208
rect 13096 2144 13112 2208
rect 13176 2144 13192 2208
rect 13256 2144 13264 2208
rect 12944 2143 13264 2144
rect 20944 2208 21264 2209
rect 20944 2144 20952 2208
rect 21016 2144 21032 2208
rect 21096 2144 21112 2208
rect 21176 2144 21192 2208
rect 21256 2144 21264 2208
rect 23520 2184 24000 2304
rect 20944 2143 21264 2144
rect 8017 2002 8083 2005
rect 19885 2002 19951 2005
rect 8017 2000 19951 2002
rect 8017 1944 8022 2000
rect 8078 1944 19890 2000
rect 19946 1944 19951 2000
rect 8017 1942 19951 1944
rect 8017 1939 8083 1942
rect 19885 1939 19951 1942
rect 6545 1866 6611 1869
rect 62 1864 6611 1866
rect 62 1808 6550 1864
rect 6606 1808 6611 1864
rect 62 1806 6611 1808
rect 62 1352 122 1806
rect 6545 1803 6611 1806
rect 11789 1594 11855 1597
rect 23614 1594 23674 2184
rect 11789 1592 23674 1594
rect 11789 1536 11794 1592
rect 11850 1536 23674 1592
rect 11789 1534 23674 1536
rect 11789 1531 11855 1534
rect 0 1232 480 1352
rect 13813 1322 13879 1325
rect 13813 1320 23674 1322
rect 13813 1264 13818 1320
rect 13874 1264 23674 1320
rect 13813 1262 23674 1264
rect 13813 1259 13879 1262
rect 23614 808 23674 1262
rect 23520 688 24000 808
<< via3 >>
rect 4952 21788 5016 21792
rect 4952 21732 4956 21788
rect 4956 21732 5012 21788
rect 5012 21732 5016 21788
rect 4952 21728 5016 21732
rect 5032 21788 5096 21792
rect 5032 21732 5036 21788
rect 5036 21732 5092 21788
rect 5092 21732 5096 21788
rect 5032 21728 5096 21732
rect 5112 21788 5176 21792
rect 5112 21732 5116 21788
rect 5116 21732 5172 21788
rect 5172 21732 5176 21788
rect 5112 21728 5176 21732
rect 5192 21788 5256 21792
rect 5192 21732 5196 21788
rect 5196 21732 5252 21788
rect 5252 21732 5256 21788
rect 5192 21728 5256 21732
rect 12952 21788 13016 21792
rect 12952 21732 12956 21788
rect 12956 21732 13012 21788
rect 13012 21732 13016 21788
rect 12952 21728 13016 21732
rect 13032 21788 13096 21792
rect 13032 21732 13036 21788
rect 13036 21732 13092 21788
rect 13092 21732 13096 21788
rect 13032 21728 13096 21732
rect 13112 21788 13176 21792
rect 13112 21732 13116 21788
rect 13116 21732 13172 21788
rect 13172 21732 13176 21788
rect 13112 21728 13176 21732
rect 13192 21788 13256 21792
rect 13192 21732 13196 21788
rect 13196 21732 13252 21788
rect 13252 21732 13256 21788
rect 13192 21728 13256 21732
rect 20952 21788 21016 21792
rect 20952 21732 20956 21788
rect 20956 21732 21012 21788
rect 21012 21732 21016 21788
rect 20952 21728 21016 21732
rect 21032 21788 21096 21792
rect 21032 21732 21036 21788
rect 21036 21732 21092 21788
rect 21092 21732 21096 21788
rect 21032 21728 21096 21732
rect 21112 21788 21176 21792
rect 21112 21732 21116 21788
rect 21116 21732 21172 21788
rect 21172 21732 21176 21788
rect 21112 21728 21176 21732
rect 21192 21788 21256 21792
rect 21192 21732 21196 21788
rect 21196 21732 21252 21788
rect 21252 21732 21256 21788
rect 21192 21728 21256 21732
rect 8952 21244 9016 21248
rect 8952 21188 8956 21244
rect 8956 21188 9012 21244
rect 9012 21188 9016 21244
rect 8952 21184 9016 21188
rect 9032 21244 9096 21248
rect 9032 21188 9036 21244
rect 9036 21188 9092 21244
rect 9092 21188 9096 21244
rect 9032 21184 9096 21188
rect 9112 21244 9176 21248
rect 9112 21188 9116 21244
rect 9116 21188 9172 21244
rect 9172 21188 9176 21244
rect 9112 21184 9176 21188
rect 9192 21244 9256 21248
rect 9192 21188 9196 21244
rect 9196 21188 9252 21244
rect 9252 21188 9256 21244
rect 9192 21184 9256 21188
rect 16952 21244 17016 21248
rect 16952 21188 16956 21244
rect 16956 21188 17012 21244
rect 17012 21188 17016 21244
rect 16952 21184 17016 21188
rect 17032 21244 17096 21248
rect 17032 21188 17036 21244
rect 17036 21188 17092 21244
rect 17092 21188 17096 21244
rect 17032 21184 17096 21188
rect 17112 21244 17176 21248
rect 17112 21188 17116 21244
rect 17116 21188 17172 21244
rect 17172 21188 17176 21244
rect 17112 21184 17176 21188
rect 17192 21244 17256 21248
rect 17192 21188 17196 21244
rect 17196 21188 17252 21244
rect 17252 21188 17256 21244
rect 17192 21184 17256 21188
rect 4952 20700 5016 20704
rect 4952 20644 4956 20700
rect 4956 20644 5012 20700
rect 5012 20644 5016 20700
rect 4952 20640 5016 20644
rect 5032 20700 5096 20704
rect 5032 20644 5036 20700
rect 5036 20644 5092 20700
rect 5092 20644 5096 20700
rect 5032 20640 5096 20644
rect 5112 20700 5176 20704
rect 5112 20644 5116 20700
rect 5116 20644 5172 20700
rect 5172 20644 5176 20700
rect 5112 20640 5176 20644
rect 5192 20700 5256 20704
rect 5192 20644 5196 20700
rect 5196 20644 5252 20700
rect 5252 20644 5256 20700
rect 5192 20640 5256 20644
rect 12952 20700 13016 20704
rect 12952 20644 12956 20700
rect 12956 20644 13012 20700
rect 13012 20644 13016 20700
rect 12952 20640 13016 20644
rect 13032 20700 13096 20704
rect 13032 20644 13036 20700
rect 13036 20644 13092 20700
rect 13092 20644 13096 20700
rect 13032 20640 13096 20644
rect 13112 20700 13176 20704
rect 13112 20644 13116 20700
rect 13116 20644 13172 20700
rect 13172 20644 13176 20700
rect 13112 20640 13176 20644
rect 13192 20700 13256 20704
rect 13192 20644 13196 20700
rect 13196 20644 13252 20700
rect 13252 20644 13256 20700
rect 13192 20640 13256 20644
rect 20952 20700 21016 20704
rect 20952 20644 20956 20700
rect 20956 20644 21012 20700
rect 21012 20644 21016 20700
rect 20952 20640 21016 20644
rect 21032 20700 21096 20704
rect 21032 20644 21036 20700
rect 21036 20644 21092 20700
rect 21092 20644 21096 20700
rect 21032 20640 21096 20644
rect 21112 20700 21176 20704
rect 21112 20644 21116 20700
rect 21116 20644 21172 20700
rect 21172 20644 21176 20700
rect 21112 20640 21176 20644
rect 21192 20700 21256 20704
rect 21192 20644 21196 20700
rect 21196 20644 21252 20700
rect 21252 20644 21256 20700
rect 21192 20640 21256 20644
rect 8952 20156 9016 20160
rect 8952 20100 8956 20156
rect 8956 20100 9012 20156
rect 9012 20100 9016 20156
rect 8952 20096 9016 20100
rect 9032 20156 9096 20160
rect 9032 20100 9036 20156
rect 9036 20100 9092 20156
rect 9092 20100 9096 20156
rect 9032 20096 9096 20100
rect 9112 20156 9176 20160
rect 9112 20100 9116 20156
rect 9116 20100 9172 20156
rect 9172 20100 9176 20156
rect 9112 20096 9176 20100
rect 9192 20156 9256 20160
rect 9192 20100 9196 20156
rect 9196 20100 9252 20156
rect 9252 20100 9256 20156
rect 9192 20096 9256 20100
rect 16952 20156 17016 20160
rect 16952 20100 16956 20156
rect 16956 20100 17012 20156
rect 17012 20100 17016 20156
rect 16952 20096 17016 20100
rect 17032 20156 17096 20160
rect 17032 20100 17036 20156
rect 17036 20100 17092 20156
rect 17092 20100 17096 20156
rect 17032 20096 17096 20100
rect 17112 20156 17176 20160
rect 17112 20100 17116 20156
rect 17116 20100 17172 20156
rect 17172 20100 17176 20156
rect 17112 20096 17176 20100
rect 17192 20156 17256 20160
rect 17192 20100 17196 20156
rect 17196 20100 17252 20156
rect 17252 20100 17256 20156
rect 17192 20096 17256 20100
rect 4952 19612 5016 19616
rect 4952 19556 4956 19612
rect 4956 19556 5012 19612
rect 5012 19556 5016 19612
rect 4952 19552 5016 19556
rect 5032 19612 5096 19616
rect 5032 19556 5036 19612
rect 5036 19556 5092 19612
rect 5092 19556 5096 19612
rect 5032 19552 5096 19556
rect 5112 19612 5176 19616
rect 5112 19556 5116 19612
rect 5116 19556 5172 19612
rect 5172 19556 5176 19612
rect 5112 19552 5176 19556
rect 5192 19612 5256 19616
rect 5192 19556 5196 19612
rect 5196 19556 5252 19612
rect 5252 19556 5256 19612
rect 5192 19552 5256 19556
rect 12952 19612 13016 19616
rect 12952 19556 12956 19612
rect 12956 19556 13012 19612
rect 13012 19556 13016 19612
rect 12952 19552 13016 19556
rect 13032 19612 13096 19616
rect 13032 19556 13036 19612
rect 13036 19556 13092 19612
rect 13092 19556 13096 19612
rect 13032 19552 13096 19556
rect 13112 19612 13176 19616
rect 13112 19556 13116 19612
rect 13116 19556 13172 19612
rect 13172 19556 13176 19612
rect 13112 19552 13176 19556
rect 13192 19612 13256 19616
rect 13192 19556 13196 19612
rect 13196 19556 13252 19612
rect 13252 19556 13256 19612
rect 13192 19552 13256 19556
rect 20952 19612 21016 19616
rect 20952 19556 20956 19612
rect 20956 19556 21012 19612
rect 21012 19556 21016 19612
rect 20952 19552 21016 19556
rect 21032 19612 21096 19616
rect 21032 19556 21036 19612
rect 21036 19556 21092 19612
rect 21092 19556 21096 19612
rect 21032 19552 21096 19556
rect 21112 19612 21176 19616
rect 21112 19556 21116 19612
rect 21116 19556 21172 19612
rect 21172 19556 21176 19612
rect 21112 19552 21176 19556
rect 21192 19612 21256 19616
rect 21192 19556 21196 19612
rect 21196 19556 21252 19612
rect 21252 19556 21256 19612
rect 21192 19552 21256 19556
rect 8952 19068 9016 19072
rect 8952 19012 8956 19068
rect 8956 19012 9012 19068
rect 9012 19012 9016 19068
rect 8952 19008 9016 19012
rect 9032 19068 9096 19072
rect 9032 19012 9036 19068
rect 9036 19012 9092 19068
rect 9092 19012 9096 19068
rect 9032 19008 9096 19012
rect 9112 19068 9176 19072
rect 9112 19012 9116 19068
rect 9116 19012 9172 19068
rect 9172 19012 9176 19068
rect 9112 19008 9176 19012
rect 9192 19068 9256 19072
rect 9192 19012 9196 19068
rect 9196 19012 9252 19068
rect 9252 19012 9256 19068
rect 9192 19008 9256 19012
rect 16952 19068 17016 19072
rect 16952 19012 16956 19068
rect 16956 19012 17012 19068
rect 17012 19012 17016 19068
rect 16952 19008 17016 19012
rect 17032 19068 17096 19072
rect 17032 19012 17036 19068
rect 17036 19012 17092 19068
rect 17092 19012 17096 19068
rect 17032 19008 17096 19012
rect 17112 19068 17176 19072
rect 17112 19012 17116 19068
rect 17116 19012 17172 19068
rect 17172 19012 17176 19068
rect 17112 19008 17176 19012
rect 17192 19068 17256 19072
rect 17192 19012 17196 19068
rect 17196 19012 17252 19068
rect 17252 19012 17256 19068
rect 17192 19008 17256 19012
rect 4952 18524 5016 18528
rect 4952 18468 4956 18524
rect 4956 18468 5012 18524
rect 5012 18468 5016 18524
rect 4952 18464 5016 18468
rect 5032 18524 5096 18528
rect 5032 18468 5036 18524
rect 5036 18468 5092 18524
rect 5092 18468 5096 18524
rect 5032 18464 5096 18468
rect 5112 18524 5176 18528
rect 5112 18468 5116 18524
rect 5116 18468 5172 18524
rect 5172 18468 5176 18524
rect 5112 18464 5176 18468
rect 5192 18524 5256 18528
rect 5192 18468 5196 18524
rect 5196 18468 5252 18524
rect 5252 18468 5256 18524
rect 5192 18464 5256 18468
rect 12952 18524 13016 18528
rect 12952 18468 12956 18524
rect 12956 18468 13012 18524
rect 13012 18468 13016 18524
rect 12952 18464 13016 18468
rect 13032 18524 13096 18528
rect 13032 18468 13036 18524
rect 13036 18468 13092 18524
rect 13092 18468 13096 18524
rect 13032 18464 13096 18468
rect 13112 18524 13176 18528
rect 13112 18468 13116 18524
rect 13116 18468 13172 18524
rect 13172 18468 13176 18524
rect 13112 18464 13176 18468
rect 13192 18524 13256 18528
rect 13192 18468 13196 18524
rect 13196 18468 13252 18524
rect 13252 18468 13256 18524
rect 13192 18464 13256 18468
rect 20952 18524 21016 18528
rect 20952 18468 20956 18524
rect 20956 18468 21012 18524
rect 21012 18468 21016 18524
rect 20952 18464 21016 18468
rect 21032 18524 21096 18528
rect 21032 18468 21036 18524
rect 21036 18468 21092 18524
rect 21092 18468 21096 18524
rect 21032 18464 21096 18468
rect 21112 18524 21176 18528
rect 21112 18468 21116 18524
rect 21116 18468 21172 18524
rect 21172 18468 21176 18524
rect 21112 18464 21176 18468
rect 21192 18524 21256 18528
rect 21192 18468 21196 18524
rect 21196 18468 21252 18524
rect 21252 18468 21256 18524
rect 21192 18464 21256 18468
rect 8952 17980 9016 17984
rect 8952 17924 8956 17980
rect 8956 17924 9012 17980
rect 9012 17924 9016 17980
rect 8952 17920 9016 17924
rect 9032 17980 9096 17984
rect 9032 17924 9036 17980
rect 9036 17924 9092 17980
rect 9092 17924 9096 17980
rect 9032 17920 9096 17924
rect 9112 17980 9176 17984
rect 9112 17924 9116 17980
rect 9116 17924 9172 17980
rect 9172 17924 9176 17980
rect 9112 17920 9176 17924
rect 9192 17980 9256 17984
rect 9192 17924 9196 17980
rect 9196 17924 9252 17980
rect 9252 17924 9256 17980
rect 9192 17920 9256 17924
rect 16952 17980 17016 17984
rect 16952 17924 16956 17980
rect 16956 17924 17012 17980
rect 17012 17924 17016 17980
rect 16952 17920 17016 17924
rect 17032 17980 17096 17984
rect 17032 17924 17036 17980
rect 17036 17924 17092 17980
rect 17092 17924 17096 17980
rect 17032 17920 17096 17924
rect 17112 17980 17176 17984
rect 17112 17924 17116 17980
rect 17116 17924 17172 17980
rect 17172 17924 17176 17980
rect 17112 17920 17176 17924
rect 17192 17980 17256 17984
rect 17192 17924 17196 17980
rect 17196 17924 17252 17980
rect 17252 17924 17256 17980
rect 17192 17920 17256 17924
rect 4952 17436 5016 17440
rect 4952 17380 4956 17436
rect 4956 17380 5012 17436
rect 5012 17380 5016 17436
rect 4952 17376 5016 17380
rect 5032 17436 5096 17440
rect 5032 17380 5036 17436
rect 5036 17380 5092 17436
rect 5092 17380 5096 17436
rect 5032 17376 5096 17380
rect 5112 17436 5176 17440
rect 5112 17380 5116 17436
rect 5116 17380 5172 17436
rect 5172 17380 5176 17436
rect 5112 17376 5176 17380
rect 5192 17436 5256 17440
rect 5192 17380 5196 17436
rect 5196 17380 5252 17436
rect 5252 17380 5256 17436
rect 5192 17376 5256 17380
rect 12952 17436 13016 17440
rect 12952 17380 12956 17436
rect 12956 17380 13012 17436
rect 13012 17380 13016 17436
rect 12952 17376 13016 17380
rect 13032 17436 13096 17440
rect 13032 17380 13036 17436
rect 13036 17380 13092 17436
rect 13092 17380 13096 17436
rect 13032 17376 13096 17380
rect 13112 17436 13176 17440
rect 13112 17380 13116 17436
rect 13116 17380 13172 17436
rect 13172 17380 13176 17436
rect 13112 17376 13176 17380
rect 13192 17436 13256 17440
rect 13192 17380 13196 17436
rect 13196 17380 13252 17436
rect 13252 17380 13256 17436
rect 13192 17376 13256 17380
rect 20952 17436 21016 17440
rect 20952 17380 20956 17436
rect 20956 17380 21012 17436
rect 21012 17380 21016 17436
rect 20952 17376 21016 17380
rect 21032 17436 21096 17440
rect 21032 17380 21036 17436
rect 21036 17380 21092 17436
rect 21092 17380 21096 17436
rect 21032 17376 21096 17380
rect 21112 17436 21176 17440
rect 21112 17380 21116 17436
rect 21116 17380 21172 17436
rect 21172 17380 21176 17436
rect 21112 17376 21176 17380
rect 21192 17436 21256 17440
rect 21192 17380 21196 17436
rect 21196 17380 21252 17436
rect 21252 17380 21256 17436
rect 21192 17376 21256 17380
rect 8952 16892 9016 16896
rect 8952 16836 8956 16892
rect 8956 16836 9012 16892
rect 9012 16836 9016 16892
rect 8952 16832 9016 16836
rect 9032 16892 9096 16896
rect 9032 16836 9036 16892
rect 9036 16836 9092 16892
rect 9092 16836 9096 16892
rect 9032 16832 9096 16836
rect 9112 16892 9176 16896
rect 9112 16836 9116 16892
rect 9116 16836 9172 16892
rect 9172 16836 9176 16892
rect 9112 16832 9176 16836
rect 9192 16892 9256 16896
rect 9192 16836 9196 16892
rect 9196 16836 9252 16892
rect 9252 16836 9256 16892
rect 9192 16832 9256 16836
rect 16952 16892 17016 16896
rect 16952 16836 16956 16892
rect 16956 16836 17012 16892
rect 17012 16836 17016 16892
rect 16952 16832 17016 16836
rect 17032 16892 17096 16896
rect 17032 16836 17036 16892
rect 17036 16836 17092 16892
rect 17092 16836 17096 16892
rect 17032 16832 17096 16836
rect 17112 16892 17176 16896
rect 17112 16836 17116 16892
rect 17116 16836 17172 16892
rect 17172 16836 17176 16892
rect 17112 16832 17176 16836
rect 17192 16892 17256 16896
rect 17192 16836 17196 16892
rect 17196 16836 17252 16892
rect 17252 16836 17256 16892
rect 17192 16832 17256 16836
rect 4952 16348 5016 16352
rect 4952 16292 4956 16348
rect 4956 16292 5012 16348
rect 5012 16292 5016 16348
rect 4952 16288 5016 16292
rect 5032 16348 5096 16352
rect 5032 16292 5036 16348
rect 5036 16292 5092 16348
rect 5092 16292 5096 16348
rect 5032 16288 5096 16292
rect 5112 16348 5176 16352
rect 5112 16292 5116 16348
rect 5116 16292 5172 16348
rect 5172 16292 5176 16348
rect 5112 16288 5176 16292
rect 5192 16348 5256 16352
rect 5192 16292 5196 16348
rect 5196 16292 5252 16348
rect 5252 16292 5256 16348
rect 5192 16288 5256 16292
rect 12952 16348 13016 16352
rect 12952 16292 12956 16348
rect 12956 16292 13012 16348
rect 13012 16292 13016 16348
rect 12952 16288 13016 16292
rect 13032 16348 13096 16352
rect 13032 16292 13036 16348
rect 13036 16292 13092 16348
rect 13092 16292 13096 16348
rect 13032 16288 13096 16292
rect 13112 16348 13176 16352
rect 13112 16292 13116 16348
rect 13116 16292 13172 16348
rect 13172 16292 13176 16348
rect 13112 16288 13176 16292
rect 13192 16348 13256 16352
rect 13192 16292 13196 16348
rect 13196 16292 13252 16348
rect 13252 16292 13256 16348
rect 13192 16288 13256 16292
rect 20952 16348 21016 16352
rect 20952 16292 20956 16348
rect 20956 16292 21012 16348
rect 21012 16292 21016 16348
rect 20952 16288 21016 16292
rect 21032 16348 21096 16352
rect 21032 16292 21036 16348
rect 21036 16292 21092 16348
rect 21092 16292 21096 16348
rect 21032 16288 21096 16292
rect 21112 16348 21176 16352
rect 21112 16292 21116 16348
rect 21116 16292 21172 16348
rect 21172 16292 21176 16348
rect 21112 16288 21176 16292
rect 21192 16348 21256 16352
rect 21192 16292 21196 16348
rect 21196 16292 21252 16348
rect 21252 16292 21256 16348
rect 21192 16288 21256 16292
rect 8952 15804 9016 15808
rect 8952 15748 8956 15804
rect 8956 15748 9012 15804
rect 9012 15748 9016 15804
rect 8952 15744 9016 15748
rect 9032 15804 9096 15808
rect 9032 15748 9036 15804
rect 9036 15748 9092 15804
rect 9092 15748 9096 15804
rect 9032 15744 9096 15748
rect 9112 15804 9176 15808
rect 9112 15748 9116 15804
rect 9116 15748 9172 15804
rect 9172 15748 9176 15804
rect 9112 15744 9176 15748
rect 9192 15804 9256 15808
rect 9192 15748 9196 15804
rect 9196 15748 9252 15804
rect 9252 15748 9256 15804
rect 9192 15744 9256 15748
rect 16952 15804 17016 15808
rect 16952 15748 16956 15804
rect 16956 15748 17012 15804
rect 17012 15748 17016 15804
rect 16952 15744 17016 15748
rect 17032 15804 17096 15808
rect 17032 15748 17036 15804
rect 17036 15748 17092 15804
rect 17092 15748 17096 15804
rect 17032 15744 17096 15748
rect 17112 15804 17176 15808
rect 17112 15748 17116 15804
rect 17116 15748 17172 15804
rect 17172 15748 17176 15804
rect 17112 15744 17176 15748
rect 17192 15804 17256 15808
rect 17192 15748 17196 15804
rect 17196 15748 17252 15804
rect 17252 15748 17256 15804
rect 17192 15744 17256 15748
rect 4952 15260 5016 15264
rect 4952 15204 4956 15260
rect 4956 15204 5012 15260
rect 5012 15204 5016 15260
rect 4952 15200 5016 15204
rect 5032 15260 5096 15264
rect 5032 15204 5036 15260
rect 5036 15204 5092 15260
rect 5092 15204 5096 15260
rect 5032 15200 5096 15204
rect 5112 15260 5176 15264
rect 5112 15204 5116 15260
rect 5116 15204 5172 15260
rect 5172 15204 5176 15260
rect 5112 15200 5176 15204
rect 5192 15260 5256 15264
rect 5192 15204 5196 15260
rect 5196 15204 5252 15260
rect 5252 15204 5256 15260
rect 5192 15200 5256 15204
rect 12952 15260 13016 15264
rect 12952 15204 12956 15260
rect 12956 15204 13012 15260
rect 13012 15204 13016 15260
rect 12952 15200 13016 15204
rect 13032 15260 13096 15264
rect 13032 15204 13036 15260
rect 13036 15204 13092 15260
rect 13092 15204 13096 15260
rect 13032 15200 13096 15204
rect 13112 15260 13176 15264
rect 13112 15204 13116 15260
rect 13116 15204 13172 15260
rect 13172 15204 13176 15260
rect 13112 15200 13176 15204
rect 13192 15260 13256 15264
rect 13192 15204 13196 15260
rect 13196 15204 13252 15260
rect 13252 15204 13256 15260
rect 13192 15200 13256 15204
rect 20952 15260 21016 15264
rect 20952 15204 20956 15260
rect 20956 15204 21012 15260
rect 21012 15204 21016 15260
rect 20952 15200 21016 15204
rect 21032 15260 21096 15264
rect 21032 15204 21036 15260
rect 21036 15204 21092 15260
rect 21092 15204 21096 15260
rect 21032 15200 21096 15204
rect 21112 15260 21176 15264
rect 21112 15204 21116 15260
rect 21116 15204 21172 15260
rect 21172 15204 21176 15260
rect 21112 15200 21176 15204
rect 21192 15260 21256 15264
rect 21192 15204 21196 15260
rect 21196 15204 21252 15260
rect 21252 15204 21256 15260
rect 21192 15200 21256 15204
rect 8952 14716 9016 14720
rect 8952 14660 8956 14716
rect 8956 14660 9012 14716
rect 9012 14660 9016 14716
rect 8952 14656 9016 14660
rect 9032 14716 9096 14720
rect 9032 14660 9036 14716
rect 9036 14660 9092 14716
rect 9092 14660 9096 14716
rect 9032 14656 9096 14660
rect 9112 14716 9176 14720
rect 9112 14660 9116 14716
rect 9116 14660 9172 14716
rect 9172 14660 9176 14716
rect 9112 14656 9176 14660
rect 9192 14716 9256 14720
rect 9192 14660 9196 14716
rect 9196 14660 9252 14716
rect 9252 14660 9256 14716
rect 9192 14656 9256 14660
rect 16952 14716 17016 14720
rect 16952 14660 16956 14716
rect 16956 14660 17012 14716
rect 17012 14660 17016 14716
rect 16952 14656 17016 14660
rect 17032 14716 17096 14720
rect 17032 14660 17036 14716
rect 17036 14660 17092 14716
rect 17092 14660 17096 14716
rect 17032 14656 17096 14660
rect 17112 14716 17176 14720
rect 17112 14660 17116 14716
rect 17116 14660 17172 14716
rect 17172 14660 17176 14716
rect 17112 14656 17176 14660
rect 17192 14716 17256 14720
rect 17192 14660 17196 14716
rect 17196 14660 17252 14716
rect 17252 14660 17256 14716
rect 17192 14656 17256 14660
rect 4952 14172 5016 14176
rect 4952 14116 4956 14172
rect 4956 14116 5012 14172
rect 5012 14116 5016 14172
rect 4952 14112 5016 14116
rect 5032 14172 5096 14176
rect 5032 14116 5036 14172
rect 5036 14116 5092 14172
rect 5092 14116 5096 14172
rect 5032 14112 5096 14116
rect 5112 14172 5176 14176
rect 5112 14116 5116 14172
rect 5116 14116 5172 14172
rect 5172 14116 5176 14172
rect 5112 14112 5176 14116
rect 5192 14172 5256 14176
rect 5192 14116 5196 14172
rect 5196 14116 5252 14172
rect 5252 14116 5256 14172
rect 5192 14112 5256 14116
rect 12952 14172 13016 14176
rect 12952 14116 12956 14172
rect 12956 14116 13012 14172
rect 13012 14116 13016 14172
rect 12952 14112 13016 14116
rect 13032 14172 13096 14176
rect 13032 14116 13036 14172
rect 13036 14116 13092 14172
rect 13092 14116 13096 14172
rect 13032 14112 13096 14116
rect 13112 14172 13176 14176
rect 13112 14116 13116 14172
rect 13116 14116 13172 14172
rect 13172 14116 13176 14172
rect 13112 14112 13176 14116
rect 13192 14172 13256 14176
rect 13192 14116 13196 14172
rect 13196 14116 13252 14172
rect 13252 14116 13256 14172
rect 13192 14112 13256 14116
rect 20952 14172 21016 14176
rect 20952 14116 20956 14172
rect 20956 14116 21012 14172
rect 21012 14116 21016 14172
rect 20952 14112 21016 14116
rect 21032 14172 21096 14176
rect 21032 14116 21036 14172
rect 21036 14116 21092 14172
rect 21092 14116 21096 14172
rect 21032 14112 21096 14116
rect 21112 14172 21176 14176
rect 21112 14116 21116 14172
rect 21116 14116 21172 14172
rect 21172 14116 21176 14172
rect 21112 14112 21176 14116
rect 21192 14172 21256 14176
rect 21192 14116 21196 14172
rect 21196 14116 21252 14172
rect 21252 14116 21256 14172
rect 21192 14112 21256 14116
rect 8952 13628 9016 13632
rect 8952 13572 8956 13628
rect 8956 13572 9012 13628
rect 9012 13572 9016 13628
rect 8952 13568 9016 13572
rect 9032 13628 9096 13632
rect 9032 13572 9036 13628
rect 9036 13572 9092 13628
rect 9092 13572 9096 13628
rect 9032 13568 9096 13572
rect 9112 13628 9176 13632
rect 9112 13572 9116 13628
rect 9116 13572 9172 13628
rect 9172 13572 9176 13628
rect 9112 13568 9176 13572
rect 9192 13628 9256 13632
rect 9192 13572 9196 13628
rect 9196 13572 9252 13628
rect 9252 13572 9256 13628
rect 9192 13568 9256 13572
rect 16952 13628 17016 13632
rect 16952 13572 16956 13628
rect 16956 13572 17012 13628
rect 17012 13572 17016 13628
rect 16952 13568 17016 13572
rect 17032 13628 17096 13632
rect 17032 13572 17036 13628
rect 17036 13572 17092 13628
rect 17092 13572 17096 13628
rect 17032 13568 17096 13572
rect 17112 13628 17176 13632
rect 17112 13572 17116 13628
rect 17116 13572 17172 13628
rect 17172 13572 17176 13628
rect 17112 13568 17176 13572
rect 17192 13628 17256 13632
rect 17192 13572 17196 13628
rect 17196 13572 17252 13628
rect 17252 13572 17256 13628
rect 17192 13568 17256 13572
rect 4952 13084 5016 13088
rect 4952 13028 4956 13084
rect 4956 13028 5012 13084
rect 5012 13028 5016 13084
rect 4952 13024 5016 13028
rect 5032 13084 5096 13088
rect 5032 13028 5036 13084
rect 5036 13028 5092 13084
rect 5092 13028 5096 13084
rect 5032 13024 5096 13028
rect 5112 13084 5176 13088
rect 5112 13028 5116 13084
rect 5116 13028 5172 13084
rect 5172 13028 5176 13084
rect 5112 13024 5176 13028
rect 5192 13084 5256 13088
rect 5192 13028 5196 13084
rect 5196 13028 5252 13084
rect 5252 13028 5256 13084
rect 5192 13024 5256 13028
rect 12952 13084 13016 13088
rect 12952 13028 12956 13084
rect 12956 13028 13012 13084
rect 13012 13028 13016 13084
rect 12952 13024 13016 13028
rect 13032 13084 13096 13088
rect 13032 13028 13036 13084
rect 13036 13028 13092 13084
rect 13092 13028 13096 13084
rect 13032 13024 13096 13028
rect 13112 13084 13176 13088
rect 13112 13028 13116 13084
rect 13116 13028 13172 13084
rect 13172 13028 13176 13084
rect 13112 13024 13176 13028
rect 13192 13084 13256 13088
rect 13192 13028 13196 13084
rect 13196 13028 13252 13084
rect 13252 13028 13256 13084
rect 13192 13024 13256 13028
rect 20952 13084 21016 13088
rect 20952 13028 20956 13084
rect 20956 13028 21012 13084
rect 21012 13028 21016 13084
rect 20952 13024 21016 13028
rect 21032 13084 21096 13088
rect 21032 13028 21036 13084
rect 21036 13028 21092 13084
rect 21092 13028 21096 13084
rect 21032 13024 21096 13028
rect 21112 13084 21176 13088
rect 21112 13028 21116 13084
rect 21116 13028 21172 13084
rect 21172 13028 21176 13084
rect 21112 13024 21176 13028
rect 21192 13084 21256 13088
rect 21192 13028 21196 13084
rect 21196 13028 21252 13084
rect 21252 13028 21256 13084
rect 21192 13024 21256 13028
rect 8952 12540 9016 12544
rect 8952 12484 8956 12540
rect 8956 12484 9012 12540
rect 9012 12484 9016 12540
rect 8952 12480 9016 12484
rect 9032 12540 9096 12544
rect 9032 12484 9036 12540
rect 9036 12484 9092 12540
rect 9092 12484 9096 12540
rect 9032 12480 9096 12484
rect 9112 12540 9176 12544
rect 9112 12484 9116 12540
rect 9116 12484 9172 12540
rect 9172 12484 9176 12540
rect 9112 12480 9176 12484
rect 9192 12540 9256 12544
rect 9192 12484 9196 12540
rect 9196 12484 9252 12540
rect 9252 12484 9256 12540
rect 9192 12480 9256 12484
rect 16952 12540 17016 12544
rect 16952 12484 16956 12540
rect 16956 12484 17012 12540
rect 17012 12484 17016 12540
rect 16952 12480 17016 12484
rect 17032 12540 17096 12544
rect 17032 12484 17036 12540
rect 17036 12484 17092 12540
rect 17092 12484 17096 12540
rect 17032 12480 17096 12484
rect 17112 12540 17176 12544
rect 17112 12484 17116 12540
rect 17116 12484 17172 12540
rect 17172 12484 17176 12540
rect 17112 12480 17176 12484
rect 17192 12540 17256 12544
rect 17192 12484 17196 12540
rect 17196 12484 17252 12540
rect 17252 12484 17256 12540
rect 17192 12480 17256 12484
rect 4952 11996 5016 12000
rect 4952 11940 4956 11996
rect 4956 11940 5012 11996
rect 5012 11940 5016 11996
rect 4952 11936 5016 11940
rect 5032 11996 5096 12000
rect 5032 11940 5036 11996
rect 5036 11940 5092 11996
rect 5092 11940 5096 11996
rect 5032 11936 5096 11940
rect 5112 11996 5176 12000
rect 5112 11940 5116 11996
rect 5116 11940 5172 11996
rect 5172 11940 5176 11996
rect 5112 11936 5176 11940
rect 5192 11996 5256 12000
rect 5192 11940 5196 11996
rect 5196 11940 5252 11996
rect 5252 11940 5256 11996
rect 5192 11936 5256 11940
rect 12952 11996 13016 12000
rect 12952 11940 12956 11996
rect 12956 11940 13012 11996
rect 13012 11940 13016 11996
rect 12952 11936 13016 11940
rect 13032 11996 13096 12000
rect 13032 11940 13036 11996
rect 13036 11940 13092 11996
rect 13092 11940 13096 11996
rect 13032 11936 13096 11940
rect 13112 11996 13176 12000
rect 13112 11940 13116 11996
rect 13116 11940 13172 11996
rect 13172 11940 13176 11996
rect 13112 11936 13176 11940
rect 13192 11996 13256 12000
rect 13192 11940 13196 11996
rect 13196 11940 13252 11996
rect 13252 11940 13256 11996
rect 13192 11936 13256 11940
rect 20952 11996 21016 12000
rect 20952 11940 20956 11996
rect 20956 11940 21012 11996
rect 21012 11940 21016 11996
rect 20952 11936 21016 11940
rect 21032 11996 21096 12000
rect 21032 11940 21036 11996
rect 21036 11940 21092 11996
rect 21092 11940 21096 11996
rect 21032 11936 21096 11940
rect 21112 11996 21176 12000
rect 21112 11940 21116 11996
rect 21116 11940 21172 11996
rect 21172 11940 21176 11996
rect 21112 11936 21176 11940
rect 21192 11996 21256 12000
rect 21192 11940 21196 11996
rect 21196 11940 21252 11996
rect 21252 11940 21256 11996
rect 21192 11936 21256 11940
rect 8952 11452 9016 11456
rect 8952 11396 8956 11452
rect 8956 11396 9012 11452
rect 9012 11396 9016 11452
rect 8952 11392 9016 11396
rect 9032 11452 9096 11456
rect 9032 11396 9036 11452
rect 9036 11396 9092 11452
rect 9092 11396 9096 11452
rect 9032 11392 9096 11396
rect 9112 11452 9176 11456
rect 9112 11396 9116 11452
rect 9116 11396 9172 11452
rect 9172 11396 9176 11452
rect 9112 11392 9176 11396
rect 9192 11452 9256 11456
rect 9192 11396 9196 11452
rect 9196 11396 9252 11452
rect 9252 11396 9256 11452
rect 9192 11392 9256 11396
rect 16952 11452 17016 11456
rect 16952 11396 16956 11452
rect 16956 11396 17012 11452
rect 17012 11396 17016 11452
rect 16952 11392 17016 11396
rect 17032 11452 17096 11456
rect 17032 11396 17036 11452
rect 17036 11396 17092 11452
rect 17092 11396 17096 11452
rect 17032 11392 17096 11396
rect 17112 11452 17176 11456
rect 17112 11396 17116 11452
rect 17116 11396 17172 11452
rect 17172 11396 17176 11452
rect 17112 11392 17176 11396
rect 17192 11452 17256 11456
rect 17192 11396 17196 11452
rect 17196 11396 17252 11452
rect 17252 11396 17256 11452
rect 17192 11392 17256 11396
rect 4952 10908 5016 10912
rect 4952 10852 4956 10908
rect 4956 10852 5012 10908
rect 5012 10852 5016 10908
rect 4952 10848 5016 10852
rect 5032 10908 5096 10912
rect 5032 10852 5036 10908
rect 5036 10852 5092 10908
rect 5092 10852 5096 10908
rect 5032 10848 5096 10852
rect 5112 10908 5176 10912
rect 5112 10852 5116 10908
rect 5116 10852 5172 10908
rect 5172 10852 5176 10908
rect 5112 10848 5176 10852
rect 5192 10908 5256 10912
rect 5192 10852 5196 10908
rect 5196 10852 5252 10908
rect 5252 10852 5256 10908
rect 5192 10848 5256 10852
rect 12952 10908 13016 10912
rect 12952 10852 12956 10908
rect 12956 10852 13012 10908
rect 13012 10852 13016 10908
rect 12952 10848 13016 10852
rect 13032 10908 13096 10912
rect 13032 10852 13036 10908
rect 13036 10852 13092 10908
rect 13092 10852 13096 10908
rect 13032 10848 13096 10852
rect 13112 10908 13176 10912
rect 13112 10852 13116 10908
rect 13116 10852 13172 10908
rect 13172 10852 13176 10908
rect 13112 10848 13176 10852
rect 13192 10908 13256 10912
rect 13192 10852 13196 10908
rect 13196 10852 13252 10908
rect 13252 10852 13256 10908
rect 13192 10848 13256 10852
rect 20952 10908 21016 10912
rect 20952 10852 20956 10908
rect 20956 10852 21012 10908
rect 21012 10852 21016 10908
rect 20952 10848 21016 10852
rect 21032 10908 21096 10912
rect 21032 10852 21036 10908
rect 21036 10852 21092 10908
rect 21092 10852 21096 10908
rect 21032 10848 21096 10852
rect 21112 10908 21176 10912
rect 21112 10852 21116 10908
rect 21116 10852 21172 10908
rect 21172 10852 21176 10908
rect 21112 10848 21176 10852
rect 21192 10908 21256 10912
rect 21192 10852 21196 10908
rect 21196 10852 21252 10908
rect 21252 10852 21256 10908
rect 21192 10848 21256 10852
rect 8952 10364 9016 10368
rect 8952 10308 8956 10364
rect 8956 10308 9012 10364
rect 9012 10308 9016 10364
rect 8952 10304 9016 10308
rect 9032 10364 9096 10368
rect 9032 10308 9036 10364
rect 9036 10308 9092 10364
rect 9092 10308 9096 10364
rect 9032 10304 9096 10308
rect 9112 10364 9176 10368
rect 9112 10308 9116 10364
rect 9116 10308 9172 10364
rect 9172 10308 9176 10364
rect 9112 10304 9176 10308
rect 9192 10364 9256 10368
rect 9192 10308 9196 10364
rect 9196 10308 9252 10364
rect 9252 10308 9256 10364
rect 9192 10304 9256 10308
rect 16952 10364 17016 10368
rect 16952 10308 16956 10364
rect 16956 10308 17012 10364
rect 17012 10308 17016 10364
rect 16952 10304 17016 10308
rect 17032 10364 17096 10368
rect 17032 10308 17036 10364
rect 17036 10308 17092 10364
rect 17092 10308 17096 10364
rect 17032 10304 17096 10308
rect 17112 10364 17176 10368
rect 17112 10308 17116 10364
rect 17116 10308 17172 10364
rect 17172 10308 17176 10364
rect 17112 10304 17176 10308
rect 17192 10364 17256 10368
rect 17192 10308 17196 10364
rect 17196 10308 17252 10364
rect 17252 10308 17256 10364
rect 17192 10304 17256 10308
rect 4952 9820 5016 9824
rect 4952 9764 4956 9820
rect 4956 9764 5012 9820
rect 5012 9764 5016 9820
rect 4952 9760 5016 9764
rect 5032 9820 5096 9824
rect 5032 9764 5036 9820
rect 5036 9764 5092 9820
rect 5092 9764 5096 9820
rect 5032 9760 5096 9764
rect 5112 9820 5176 9824
rect 5112 9764 5116 9820
rect 5116 9764 5172 9820
rect 5172 9764 5176 9820
rect 5112 9760 5176 9764
rect 5192 9820 5256 9824
rect 5192 9764 5196 9820
rect 5196 9764 5252 9820
rect 5252 9764 5256 9820
rect 5192 9760 5256 9764
rect 12952 9820 13016 9824
rect 12952 9764 12956 9820
rect 12956 9764 13012 9820
rect 13012 9764 13016 9820
rect 12952 9760 13016 9764
rect 13032 9820 13096 9824
rect 13032 9764 13036 9820
rect 13036 9764 13092 9820
rect 13092 9764 13096 9820
rect 13032 9760 13096 9764
rect 13112 9820 13176 9824
rect 13112 9764 13116 9820
rect 13116 9764 13172 9820
rect 13172 9764 13176 9820
rect 13112 9760 13176 9764
rect 13192 9820 13256 9824
rect 13192 9764 13196 9820
rect 13196 9764 13252 9820
rect 13252 9764 13256 9820
rect 13192 9760 13256 9764
rect 20952 9820 21016 9824
rect 20952 9764 20956 9820
rect 20956 9764 21012 9820
rect 21012 9764 21016 9820
rect 20952 9760 21016 9764
rect 21032 9820 21096 9824
rect 21032 9764 21036 9820
rect 21036 9764 21092 9820
rect 21092 9764 21096 9820
rect 21032 9760 21096 9764
rect 21112 9820 21176 9824
rect 21112 9764 21116 9820
rect 21116 9764 21172 9820
rect 21172 9764 21176 9820
rect 21112 9760 21176 9764
rect 21192 9820 21256 9824
rect 21192 9764 21196 9820
rect 21196 9764 21252 9820
rect 21252 9764 21256 9820
rect 21192 9760 21256 9764
rect 8952 9276 9016 9280
rect 8952 9220 8956 9276
rect 8956 9220 9012 9276
rect 9012 9220 9016 9276
rect 8952 9216 9016 9220
rect 9032 9276 9096 9280
rect 9032 9220 9036 9276
rect 9036 9220 9092 9276
rect 9092 9220 9096 9276
rect 9032 9216 9096 9220
rect 9112 9276 9176 9280
rect 9112 9220 9116 9276
rect 9116 9220 9172 9276
rect 9172 9220 9176 9276
rect 9112 9216 9176 9220
rect 9192 9276 9256 9280
rect 9192 9220 9196 9276
rect 9196 9220 9252 9276
rect 9252 9220 9256 9276
rect 9192 9216 9256 9220
rect 16952 9276 17016 9280
rect 16952 9220 16956 9276
rect 16956 9220 17012 9276
rect 17012 9220 17016 9276
rect 16952 9216 17016 9220
rect 17032 9276 17096 9280
rect 17032 9220 17036 9276
rect 17036 9220 17092 9276
rect 17092 9220 17096 9276
rect 17032 9216 17096 9220
rect 17112 9276 17176 9280
rect 17112 9220 17116 9276
rect 17116 9220 17172 9276
rect 17172 9220 17176 9276
rect 17112 9216 17176 9220
rect 17192 9276 17256 9280
rect 17192 9220 17196 9276
rect 17196 9220 17252 9276
rect 17252 9220 17256 9276
rect 17192 9216 17256 9220
rect 4952 8732 5016 8736
rect 4952 8676 4956 8732
rect 4956 8676 5012 8732
rect 5012 8676 5016 8732
rect 4952 8672 5016 8676
rect 5032 8732 5096 8736
rect 5032 8676 5036 8732
rect 5036 8676 5092 8732
rect 5092 8676 5096 8732
rect 5032 8672 5096 8676
rect 5112 8732 5176 8736
rect 5112 8676 5116 8732
rect 5116 8676 5172 8732
rect 5172 8676 5176 8732
rect 5112 8672 5176 8676
rect 5192 8732 5256 8736
rect 5192 8676 5196 8732
rect 5196 8676 5252 8732
rect 5252 8676 5256 8732
rect 5192 8672 5256 8676
rect 12952 8732 13016 8736
rect 12952 8676 12956 8732
rect 12956 8676 13012 8732
rect 13012 8676 13016 8732
rect 12952 8672 13016 8676
rect 13032 8732 13096 8736
rect 13032 8676 13036 8732
rect 13036 8676 13092 8732
rect 13092 8676 13096 8732
rect 13032 8672 13096 8676
rect 13112 8732 13176 8736
rect 13112 8676 13116 8732
rect 13116 8676 13172 8732
rect 13172 8676 13176 8732
rect 13112 8672 13176 8676
rect 13192 8732 13256 8736
rect 13192 8676 13196 8732
rect 13196 8676 13252 8732
rect 13252 8676 13256 8732
rect 13192 8672 13256 8676
rect 20952 8732 21016 8736
rect 20952 8676 20956 8732
rect 20956 8676 21012 8732
rect 21012 8676 21016 8732
rect 20952 8672 21016 8676
rect 21032 8732 21096 8736
rect 21032 8676 21036 8732
rect 21036 8676 21092 8732
rect 21092 8676 21096 8732
rect 21032 8672 21096 8676
rect 21112 8732 21176 8736
rect 21112 8676 21116 8732
rect 21116 8676 21172 8732
rect 21172 8676 21176 8732
rect 21112 8672 21176 8676
rect 21192 8732 21256 8736
rect 21192 8676 21196 8732
rect 21196 8676 21252 8732
rect 21252 8676 21256 8732
rect 21192 8672 21256 8676
rect 8952 8188 9016 8192
rect 8952 8132 8956 8188
rect 8956 8132 9012 8188
rect 9012 8132 9016 8188
rect 8952 8128 9016 8132
rect 9032 8188 9096 8192
rect 9032 8132 9036 8188
rect 9036 8132 9092 8188
rect 9092 8132 9096 8188
rect 9032 8128 9096 8132
rect 9112 8188 9176 8192
rect 9112 8132 9116 8188
rect 9116 8132 9172 8188
rect 9172 8132 9176 8188
rect 9112 8128 9176 8132
rect 9192 8188 9256 8192
rect 9192 8132 9196 8188
rect 9196 8132 9252 8188
rect 9252 8132 9256 8188
rect 9192 8128 9256 8132
rect 16952 8188 17016 8192
rect 16952 8132 16956 8188
rect 16956 8132 17012 8188
rect 17012 8132 17016 8188
rect 16952 8128 17016 8132
rect 17032 8188 17096 8192
rect 17032 8132 17036 8188
rect 17036 8132 17092 8188
rect 17092 8132 17096 8188
rect 17032 8128 17096 8132
rect 17112 8188 17176 8192
rect 17112 8132 17116 8188
rect 17116 8132 17172 8188
rect 17172 8132 17176 8188
rect 17112 8128 17176 8132
rect 17192 8188 17256 8192
rect 17192 8132 17196 8188
rect 17196 8132 17252 8188
rect 17252 8132 17256 8188
rect 17192 8128 17256 8132
rect 4952 7644 5016 7648
rect 4952 7588 4956 7644
rect 4956 7588 5012 7644
rect 5012 7588 5016 7644
rect 4952 7584 5016 7588
rect 5032 7644 5096 7648
rect 5032 7588 5036 7644
rect 5036 7588 5092 7644
rect 5092 7588 5096 7644
rect 5032 7584 5096 7588
rect 5112 7644 5176 7648
rect 5112 7588 5116 7644
rect 5116 7588 5172 7644
rect 5172 7588 5176 7644
rect 5112 7584 5176 7588
rect 5192 7644 5256 7648
rect 5192 7588 5196 7644
rect 5196 7588 5252 7644
rect 5252 7588 5256 7644
rect 5192 7584 5256 7588
rect 12952 7644 13016 7648
rect 12952 7588 12956 7644
rect 12956 7588 13012 7644
rect 13012 7588 13016 7644
rect 12952 7584 13016 7588
rect 13032 7644 13096 7648
rect 13032 7588 13036 7644
rect 13036 7588 13092 7644
rect 13092 7588 13096 7644
rect 13032 7584 13096 7588
rect 13112 7644 13176 7648
rect 13112 7588 13116 7644
rect 13116 7588 13172 7644
rect 13172 7588 13176 7644
rect 13112 7584 13176 7588
rect 13192 7644 13256 7648
rect 13192 7588 13196 7644
rect 13196 7588 13252 7644
rect 13252 7588 13256 7644
rect 13192 7584 13256 7588
rect 20952 7644 21016 7648
rect 20952 7588 20956 7644
rect 20956 7588 21012 7644
rect 21012 7588 21016 7644
rect 20952 7584 21016 7588
rect 21032 7644 21096 7648
rect 21032 7588 21036 7644
rect 21036 7588 21092 7644
rect 21092 7588 21096 7644
rect 21032 7584 21096 7588
rect 21112 7644 21176 7648
rect 21112 7588 21116 7644
rect 21116 7588 21172 7644
rect 21172 7588 21176 7644
rect 21112 7584 21176 7588
rect 21192 7644 21256 7648
rect 21192 7588 21196 7644
rect 21196 7588 21252 7644
rect 21252 7588 21256 7644
rect 21192 7584 21256 7588
rect 8952 7100 9016 7104
rect 8952 7044 8956 7100
rect 8956 7044 9012 7100
rect 9012 7044 9016 7100
rect 8952 7040 9016 7044
rect 9032 7100 9096 7104
rect 9032 7044 9036 7100
rect 9036 7044 9092 7100
rect 9092 7044 9096 7100
rect 9032 7040 9096 7044
rect 9112 7100 9176 7104
rect 9112 7044 9116 7100
rect 9116 7044 9172 7100
rect 9172 7044 9176 7100
rect 9112 7040 9176 7044
rect 9192 7100 9256 7104
rect 9192 7044 9196 7100
rect 9196 7044 9252 7100
rect 9252 7044 9256 7100
rect 9192 7040 9256 7044
rect 16952 7100 17016 7104
rect 16952 7044 16956 7100
rect 16956 7044 17012 7100
rect 17012 7044 17016 7100
rect 16952 7040 17016 7044
rect 17032 7100 17096 7104
rect 17032 7044 17036 7100
rect 17036 7044 17092 7100
rect 17092 7044 17096 7100
rect 17032 7040 17096 7044
rect 17112 7100 17176 7104
rect 17112 7044 17116 7100
rect 17116 7044 17172 7100
rect 17172 7044 17176 7100
rect 17112 7040 17176 7044
rect 17192 7100 17256 7104
rect 17192 7044 17196 7100
rect 17196 7044 17252 7100
rect 17252 7044 17256 7100
rect 17192 7040 17256 7044
rect 4952 6556 5016 6560
rect 4952 6500 4956 6556
rect 4956 6500 5012 6556
rect 5012 6500 5016 6556
rect 4952 6496 5016 6500
rect 5032 6556 5096 6560
rect 5032 6500 5036 6556
rect 5036 6500 5092 6556
rect 5092 6500 5096 6556
rect 5032 6496 5096 6500
rect 5112 6556 5176 6560
rect 5112 6500 5116 6556
rect 5116 6500 5172 6556
rect 5172 6500 5176 6556
rect 5112 6496 5176 6500
rect 5192 6556 5256 6560
rect 5192 6500 5196 6556
rect 5196 6500 5252 6556
rect 5252 6500 5256 6556
rect 5192 6496 5256 6500
rect 12952 6556 13016 6560
rect 12952 6500 12956 6556
rect 12956 6500 13012 6556
rect 13012 6500 13016 6556
rect 12952 6496 13016 6500
rect 13032 6556 13096 6560
rect 13032 6500 13036 6556
rect 13036 6500 13092 6556
rect 13092 6500 13096 6556
rect 13032 6496 13096 6500
rect 13112 6556 13176 6560
rect 13112 6500 13116 6556
rect 13116 6500 13172 6556
rect 13172 6500 13176 6556
rect 13112 6496 13176 6500
rect 13192 6556 13256 6560
rect 13192 6500 13196 6556
rect 13196 6500 13252 6556
rect 13252 6500 13256 6556
rect 13192 6496 13256 6500
rect 20952 6556 21016 6560
rect 20952 6500 20956 6556
rect 20956 6500 21012 6556
rect 21012 6500 21016 6556
rect 20952 6496 21016 6500
rect 21032 6556 21096 6560
rect 21032 6500 21036 6556
rect 21036 6500 21092 6556
rect 21092 6500 21096 6556
rect 21032 6496 21096 6500
rect 21112 6556 21176 6560
rect 21112 6500 21116 6556
rect 21116 6500 21172 6556
rect 21172 6500 21176 6556
rect 21112 6496 21176 6500
rect 21192 6556 21256 6560
rect 21192 6500 21196 6556
rect 21196 6500 21252 6556
rect 21252 6500 21256 6556
rect 21192 6496 21256 6500
rect 8952 6012 9016 6016
rect 8952 5956 8956 6012
rect 8956 5956 9012 6012
rect 9012 5956 9016 6012
rect 8952 5952 9016 5956
rect 9032 6012 9096 6016
rect 9032 5956 9036 6012
rect 9036 5956 9092 6012
rect 9092 5956 9096 6012
rect 9032 5952 9096 5956
rect 9112 6012 9176 6016
rect 9112 5956 9116 6012
rect 9116 5956 9172 6012
rect 9172 5956 9176 6012
rect 9112 5952 9176 5956
rect 9192 6012 9256 6016
rect 9192 5956 9196 6012
rect 9196 5956 9252 6012
rect 9252 5956 9256 6012
rect 9192 5952 9256 5956
rect 16952 6012 17016 6016
rect 16952 5956 16956 6012
rect 16956 5956 17012 6012
rect 17012 5956 17016 6012
rect 16952 5952 17016 5956
rect 17032 6012 17096 6016
rect 17032 5956 17036 6012
rect 17036 5956 17092 6012
rect 17092 5956 17096 6012
rect 17032 5952 17096 5956
rect 17112 6012 17176 6016
rect 17112 5956 17116 6012
rect 17116 5956 17172 6012
rect 17172 5956 17176 6012
rect 17112 5952 17176 5956
rect 17192 6012 17256 6016
rect 17192 5956 17196 6012
rect 17196 5956 17252 6012
rect 17252 5956 17256 6012
rect 17192 5952 17256 5956
rect 4952 5468 5016 5472
rect 4952 5412 4956 5468
rect 4956 5412 5012 5468
rect 5012 5412 5016 5468
rect 4952 5408 5016 5412
rect 5032 5468 5096 5472
rect 5032 5412 5036 5468
rect 5036 5412 5092 5468
rect 5092 5412 5096 5468
rect 5032 5408 5096 5412
rect 5112 5468 5176 5472
rect 5112 5412 5116 5468
rect 5116 5412 5172 5468
rect 5172 5412 5176 5468
rect 5112 5408 5176 5412
rect 5192 5468 5256 5472
rect 5192 5412 5196 5468
rect 5196 5412 5252 5468
rect 5252 5412 5256 5468
rect 5192 5408 5256 5412
rect 12952 5468 13016 5472
rect 12952 5412 12956 5468
rect 12956 5412 13012 5468
rect 13012 5412 13016 5468
rect 12952 5408 13016 5412
rect 13032 5468 13096 5472
rect 13032 5412 13036 5468
rect 13036 5412 13092 5468
rect 13092 5412 13096 5468
rect 13032 5408 13096 5412
rect 13112 5468 13176 5472
rect 13112 5412 13116 5468
rect 13116 5412 13172 5468
rect 13172 5412 13176 5468
rect 13112 5408 13176 5412
rect 13192 5468 13256 5472
rect 13192 5412 13196 5468
rect 13196 5412 13252 5468
rect 13252 5412 13256 5468
rect 13192 5408 13256 5412
rect 20952 5468 21016 5472
rect 20952 5412 20956 5468
rect 20956 5412 21012 5468
rect 21012 5412 21016 5468
rect 20952 5408 21016 5412
rect 21032 5468 21096 5472
rect 21032 5412 21036 5468
rect 21036 5412 21092 5468
rect 21092 5412 21096 5468
rect 21032 5408 21096 5412
rect 21112 5468 21176 5472
rect 21112 5412 21116 5468
rect 21116 5412 21172 5468
rect 21172 5412 21176 5468
rect 21112 5408 21176 5412
rect 21192 5468 21256 5472
rect 21192 5412 21196 5468
rect 21196 5412 21252 5468
rect 21252 5412 21256 5468
rect 21192 5408 21256 5412
rect 8952 4924 9016 4928
rect 8952 4868 8956 4924
rect 8956 4868 9012 4924
rect 9012 4868 9016 4924
rect 8952 4864 9016 4868
rect 9032 4924 9096 4928
rect 9032 4868 9036 4924
rect 9036 4868 9092 4924
rect 9092 4868 9096 4924
rect 9032 4864 9096 4868
rect 9112 4924 9176 4928
rect 9112 4868 9116 4924
rect 9116 4868 9172 4924
rect 9172 4868 9176 4924
rect 9112 4864 9176 4868
rect 9192 4924 9256 4928
rect 9192 4868 9196 4924
rect 9196 4868 9252 4924
rect 9252 4868 9256 4924
rect 9192 4864 9256 4868
rect 16952 4924 17016 4928
rect 16952 4868 16956 4924
rect 16956 4868 17012 4924
rect 17012 4868 17016 4924
rect 16952 4864 17016 4868
rect 17032 4924 17096 4928
rect 17032 4868 17036 4924
rect 17036 4868 17092 4924
rect 17092 4868 17096 4924
rect 17032 4864 17096 4868
rect 17112 4924 17176 4928
rect 17112 4868 17116 4924
rect 17116 4868 17172 4924
rect 17172 4868 17176 4924
rect 17112 4864 17176 4868
rect 17192 4924 17256 4928
rect 17192 4868 17196 4924
rect 17196 4868 17252 4924
rect 17252 4868 17256 4924
rect 17192 4864 17256 4868
rect 4952 4380 5016 4384
rect 4952 4324 4956 4380
rect 4956 4324 5012 4380
rect 5012 4324 5016 4380
rect 4952 4320 5016 4324
rect 5032 4380 5096 4384
rect 5032 4324 5036 4380
rect 5036 4324 5092 4380
rect 5092 4324 5096 4380
rect 5032 4320 5096 4324
rect 5112 4380 5176 4384
rect 5112 4324 5116 4380
rect 5116 4324 5172 4380
rect 5172 4324 5176 4380
rect 5112 4320 5176 4324
rect 5192 4380 5256 4384
rect 5192 4324 5196 4380
rect 5196 4324 5252 4380
rect 5252 4324 5256 4380
rect 5192 4320 5256 4324
rect 12952 4380 13016 4384
rect 12952 4324 12956 4380
rect 12956 4324 13012 4380
rect 13012 4324 13016 4380
rect 12952 4320 13016 4324
rect 13032 4380 13096 4384
rect 13032 4324 13036 4380
rect 13036 4324 13092 4380
rect 13092 4324 13096 4380
rect 13032 4320 13096 4324
rect 13112 4380 13176 4384
rect 13112 4324 13116 4380
rect 13116 4324 13172 4380
rect 13172 4324 13176 4380
rect 13112 4320 13176 4324
rect 13192 4380 13256 4384
rect 13192 4324 13196 4380
rect 13196 4324 13252 4380
rect 13252 4324 13256 4380
rect 13192 4320 13256 4324
rect 20952 4380 21016 4384
rect 20952 4324 20956 4380
rect 20956 4324 21012 4380
rect 21012 4324 21016 4380
rect 20952 4320 21016 4324
rect 21032 4380 21096 4384
rect 21032 4324 21036 4380
rect 21036 4324 21092 4380
rect 21092 4324 21096 4380
rect 21032 4320 21096 4324
rect 21112 4380 21176 4384
rect 21112 4324 21116 4380
rect 21116 4324 21172 4380
rect 21172 4324 21176 4380
rect 21112 4320 21176 4324
rect 21192 4380 21256 4384
rect 21192 4324 21196 4380
rect 21196 4324 21252 4380
rect 21252 4324 21256 4380
rect 21192 4320 21256 4324
rect 8952 3836 9016 3840
rect 8952 3780 8956 3836
rect 8956 3780 9012 3836
rect 9012 3780 9016 3836
rect 8952 3776 9016 3780
rect 9032 3836 9096 3840
rect 9032 3780 9036 3836
rect 9036 3780 9092 3836
rect 9092 3780 9096 3836
rect 9032 3776 9096 3780
rect 9112 3836 9176 3840
rect 9112 3780 9116 3836
rect 9116 3780 9172 3836
rect 9172 3780 9176 3836
rect 9112 3776 9176 3780
rect 9192 3836 9256 3840
rect 9192 3780 9196 3836
rect 9196 3780 9252 3836
rect 9252 3780 9256 3836
rect 9192 3776 9256 3780
rect 16952 3836 17016 3840
rect 16952 3780 16956 3836
rect 16956 3780 17012 3836
rect 17012 3780 17016 3836
rect 16952 3776 17016 3780
rect 17032 3836 17096 3840
rect 17032 3780 17036 3836
rect 17036 3780 17092 3836
rect 17092 3780 17096 3836
rect 17032 3776 17096 3780
rect 17112 3836 17176 3840
rect 17112 3780 17116 3836
rect 17116 3780 17172 3836
rect 17172 3780 17176 3836
rect 17112 3776 17176 3780
rect 17192 3836 17256 3840
rect 17192 3780 17196 3836
rect 17196 3780 17252 3836
rect 17252 3780 17256 3836
rect 17192 3776 17256 3780
rect 4952 3292 5016 3296
rect 4952 3236 4956 3292
rect 4956 3236 5012 3292
rect 5012 3236 5016 3292
rect 4952 3232 5016 3236
rect 5032 3292 5096 3296
rect 5032 3236 5036 3292
rect 5036 3236 5092 3292
rect 5092 3236 5096 3292
rect 5032 3232 5096 3236
rect 5112 3292 5176 3296
rect 5112 3236 5116 3292
rect 5116 3236 5172 3292
rect 5172 3236 5176 3292
rect 5112 3232 5176 3236
rect 5192 3292 5256 3296
rect 5192 3236 5196 3292
rect 5196 3236 5252 3292
rect 5252 3236 5256 3292
rect 5192 3232 5256 3236
rect 12952 3292 13016 3296
rect 12952 3236 12956 3292
rect 12956 3236 13012 3292
rect 13012 3236 13016 3292
rect 12952 3232 13016 3236
rect 13032 3292 13096 3296
rect 13032 3236 13036 3292
rect 13036 3236 13092 3292
rect 13092 3236 13096 3292
rect 13032 3232 13096 3236
rect 13112 3292 13176 3296
rect 13112 3236 13116 3292
rect 13116 3236 13172 3292
rect 13172 3236 13176 3292
rect 13112 3232 13176 3236
rect 13192 3292 13256 3296
rect 13192 3236 13196 3292
rect 13196 3236 13252 3292
rect 13252 3236 13256 3292
rect 13192 3232 13256 3236
rect 20952 3292 21016 3296
rect 20952 3236 20956 3292
rect 20956 3236 21012 3292
rect 21012 3236 21016 3292
rect 20952 3232 21016 3236
rect 21032 3292 21096 3296
rect 21032 3236 21036 3292
rect 21036 3236 21092 3292
rect 21092 3236 21096 3292
rect 21032 3232 21096 3236
rect 21112 3292 21176 3296
rect 21112 3236 21116 3292
rect 21116 3236 21172 3292
rect 21172 3236 21176 3292
rect 21112 3232 21176 3236
rect 21192 3292 21256 3296
rect 21192 3236 21196 3292
rect 21196 3236 21252 3292
rect 21252 3236 21256 3292
rect 21192 3232 21256 3236
rect 8952 2748 9016 2752
rect 8952 2692 8956 2748
rect 8956 2692 9012 2748
rect 9012 2692 9016 2748
rect 8952 2688 9016 2692
rect 9032 2748 9096 2752
rect 9032 2692 9036 2748
rect 9036 2692 9092 2748
rect 9092 2692 9096 2748
rect 9032 2688 9096 2692
rect 9112 2748 9176 2752
rect 9112 2692 9116 2748
rect 9116 2692 9172 2748
rect 9172 2692 9176 2748
rect 9112 2688 9176 2692
rect 9192 2748 9256 2752
rect 9192 2692 9196 2748
rect 9196 2692 9252 2748
rect 9252 2692 9256 2748
rect 9192 2688 9256 2692
rect 16952 2748 17016 2752
rect 16952 2692 16956 2748
rect 16956 2692 17012 2748
rect 17012 2692 17016 2748
rect 16952 2688 17016 2692
rect 17032 2748 17096 2752
rect 17032 2692 17036 2748
rect 17036 2692 17092 2748
rect 17092 2692 17096 2748
rect 17032 2688 17096 2692
rect 17112 2748 17176 2752
rect 17112 2692 17116 2748
rect 17116 2692 17172 2748
rect 17172 2692 17176 2748
rect 17112 2688 17176 2692
rect 17192 2748 17256 2752
rect 17192 2692 17196 2748
rect 17196 2692 17252 2748
rect 17252 2692 17256 2748
rect 17192 2688 17256 2692
rect 4952 2204 5016 2208
rect 4952 2148 4956 2204
rect 4956 2148 5012 2204
rect 5012 2148 5016 2204
rect 4952 2144 5016 2148
rect 5032 2204 5096 2208
rect 5032 2148 5036 2204
rect 5036 2148 5092 2204
rect 5092 2148 5096 2204
rect 5032 2144 5096 2148
rect 5112 2204 5176 2208
rect 5112 2148 5116 2204
rect 5116 2148 5172 2204
rect 5172 2148 5176 2204
rect 5112 2144 5176 2148
rect 5192 2204 5256 2208
rect 5192 2148 5196 2204
rect 5196 2148 5252 2204
rect 5252 2148 5256 2204
rect 5192 2144 5256 2148
rect 12952 2204 13016 2208
rect 12952 2148 12956 2204
rect 12956 2148 13012 2204
rect 13012 2148 13016 2204
rect 12952 2144 13016 2148
rect 13032 2204 13096 2208
rect 13032 2148 13036 2204
rect 13036 2148 13092 2204
rect 13092 2148 13096 2204
rect 13032 2144 13096 2148
rect 13112 2204 13176 2208
rect 13112 2148 13116 2204
rect 13116 2148 13172 2204
rect 13172 2148 13176 2204
rect 13112 2144 13176 2148
rect 13192 2204 13256 2208
rect 13192 2148 13196 2204
rect 13196 2148 13252 2204
rect 13252 2148 13256 2204
rect 13192 2144 13256 2148
rect 20952 2204 21016 2208
rect 20952 2148 20956 2204
rect 20956 2148 21012 2204
rect 21012 2148 21016 2204
rect 20952 2144 21016 2148
rect 21032 2204 21096 2208
rect 21032 2148 21036 2204
rect 21036 2148 21092 2204
rect 21092 2148 21096 2204
rect 21032 2144 21096 2148
rect 21112 2204 21176 2208
rect 21112 2148 21116 2204
rect 21116 2148 21172 2204
rect 21172 2148 21176 2204
rect 21112 2144 21176 2148
rect 21192 2204 21256 2208
rect 21192 2148 21196 2204
rect 21196 2148 21252 2204
rect 21252 2148 21256 2204
rect 21192 2144 21256 2148
<< metal4 >>
rect 4944 21792 5264 21808
rect 4944 21728 4952 21792
rect 5016 21728 5032 21792
rect 5096 21728 5112 21792
rect 5176 21728 5192 21792
rect 5256 21728 5264 21792
rect 4944 20704 5264 21728
rect 4944 20640 4952 20704
rect 5016 20640 5032 20704
rect 5096 20640 5112 20704
rect 5176 20640 5192 20704
rect 5256 20640 5264 20704
rect 4944 19616 5264 20640
rect 4944 19552 4952 19616
rect 5016 19552 5032 19616
rect 5096 19552 5112 19616
rect 5176 19552 5192 19616
rect 5256 19552 5264 19616
rect 4944 18528 5264 19552
rect 4944 18464 4952 18528
rect 5016 18464 5032 18528
rect 5096 18464 5112 18528
rect 5176 18464 5192 18528
rect 5256 18464 5264 18528
rect 4944 17440 5264 18464
rect 4944 17376 4952 17440
rect 5016 17376 5032 17440
rect 5096 17376 5112 17440
rect 5176 17376 5192 17440
rect 5256 17376 5264 17440
rect 4944 16352 5264 17376
rect 4944 16288 4952 16352
rect 5016 16288 5032 16352
rect 5096 16288 5112 16352
rect 5176 16288 5192 16352
rect 5256 16288 5264 16352
rect 4944 15264 5264 16288
rect 4944 15200 4952 15264
rect 5016 15200 5032 15264
rect 5096 15200 5112 15264
rect 5176 15200 5192 15264
rect 5256 15200 5264 15264
rect 4944 14176 5264 15200
rect 4944 14112 4952 14176
rect 5016 14112 5032 14176
rect 5096 14112 5112 14176
rect 5176 14112 5192 14176
rect 5256 14112 5264 14176
rect 4944 13088 5264 14112
rect 4944 13024 4952 13088
rect 5016 13024 5032 13088
rect 5096 13024 5112 13088
rect 5176 13024 5192 13088
rect 5256 13024 5264 13088
rect 4944 12000 5264 13024
rect 4944 11936 4952 12000
rect 5016 11936 5032 12000
rect 5096 11936 5112 12000
rect 5176 11936 5192 12000
rect 5256 11936 5264 12000
rect 4944 10912 5264 11936
rect 4944 10848 4952 10912
rect 5016 10848 5032 10912
rect 5096 10848 5112 10912
rect 5176 10848 5192 10912
rect 5256 10848 5264 10912
rect 4944 9824 5264 10848
rect 4944 9760 4952 9824
rect 5016 9760 5032 9824
rect 5096 9760 5112 9824
rect 5176 9760 5192 9824
rect 5256 9760 5264 9824
rect 4944 8736 5264 9760
rect 4944 8672 4952 8736
rect 5016 8672 5032 8736
rect 5096 8672 5112 8736
rect 5176 8672 5192 8736
rect 5256 8672 5264 8736
rect 4944 7648 5264 8672
rect 4944 7584 4952 7648
rect 5016 7584 5032 7648
rect 5096 7584 5112 7648
rect 5176 7584 5192 7648
rect 5256 7584 5264 7648
rect 4944 6560 5264 7584
rect 4944 6496 4952 6560
rect 5016 6496 5032 6560
rect 5096 6496 5112 6560
rect 5176 6496 5192 6560
rect 5256 6496 5264 6560
rect 4944 5472 5264 6496
rect 4944 5408 4952 5472
rect 5016 5408 5032 5472
rect 5096 5408 5112 5472
rect 5176 5408 5192 5472
rect 5256 5408 5264 5472
rect 4944 4384 5264 5408
rect 4944 4320 4952 4384
rect 5016 4320 5032 4384
rect 5096 4320 5112 4384
rect 5176 4320 5192 4384
rect 5256 4320 5264 4384
rect 4944 3296 5264 4320
rect 4944 3232 4952 3296
rect 5016 3232 5032 3296
rect 5096 3232 5112 3296
rect 5176 3232 5192 3296
rect 5256 3232 5264 3296
rect 4944 2208 5264 3232
rect 4944 2144 4952 2208
rect 5016 2144 5032 2208
rect 5096 2144 5112 2208
rect 5176 2144 5192 2208
rect 5256 2144 5264 2208
rect 4944 2128 5264 2144
rect 8944 21248 9264 21808
rect 8944 21184 8952 21248
rect 9016 21184 9032 21248
rect 9096 21184 9112 21248
rect 9176 21184 9192 21248
rect 9256 21184 9264 21248
rect 8944 20160 9264 21184
rect 8944 20096 8952 20160
rect 9016 20096 9032 20160
rect 9096 20096 9112 20160
rect 9176 20096 9192 20160
rect 9256 20096 9264 20160
rect 8944 19072 9264 20096
rect 8944 19008 8952 19072
rect 9016 19008 9032 19072
rect 9096 19008 9112 19072
rect 9176 19008 9192 19072
rect 9256 19008 9264 19072
rect 8944 17984 9264 19008
rect 8944 17920 8952 17984
rect 9016 17920 9032 17984
rect 9096 17920 9112 17984
rect 9176 17920 9192 17984
rect 9256 17920 9264 17984
rect 8944 16896 9264 17920
rect 8944 16832 8952 16896
rect 9016 16832 9032 16896
rect 9096 16832 9112 16896
rect 9176 16832 9192 16896
rect 9256 16832 9264 16896
rect 8944 15808 9264 16832
rect 8944 15744 8952 15808
rect 9016 15744 9032 15808
rect 9096 15744 9112 15808
rect 9176 15744 9192 15808
rect 9256 15744 9264 15808
rect 8944 14720 9264 15744
rect 8944 14656 8952 14720
rect 9016 14656 9032 14720
rect 9096 14656 9112 14720
rect 9176 14656 9192 14720
rect 9256 14656 9264 14720
rect 8944 13632 9264 14656
rect 8944 13568 8952 13632
rect 9016 13568 9032 13632
rect 9096 13568 9112 13632
rect 9176 13568 9192 13632
rect 9256 13568 9264 13632
rect 8944 12544 9264 13568
rect 8944 12480 8952 12544
rect 9016 12480 9032 12544
rect 9096 12480 9112 12544
rect 9176 12480 9192 12544
rect 9256 12480 9264 12544
rect 8944 11456 9264 12480
rect 8944 11392 8952 11456
rect 9016 11392 9032 11456
rect 9096 11392 9112 11456
rect 9176 11392 9192 11456
rect 9256 11392 9264 11456
rect 8944 10368 9264 11392
rect 8944 10304 8952 10368
rect 9016 10304 9032 10368
rect 9096 10304 9112 10368
rect 9176 10304 9192 10368
rect 9256 10304 9264 10368
rect 8944 9280 9264 10304
rect 8944 9216 8952 9280
rect 9016 9216 9032 9280
rect 9096 9216 9112 9280
rect 9176 9216 9192 9280
rect 9256 9216 9264 9280
rect 8944 8192 9264 9216
rect 8944 8128 8952 8192
rect 9016 8128 9032 8192
rect 9096 8128 9112 8192
rect 9176 8128 9192 8192
rect 9256 8128 9264 8192
rect 8944 7104 9264 8128
rect 8944 7040 8952 7104
rect 9016 7040 9032 7104
rect 9096 7040 9112 7104
rect 9176 7040 9192 7104
rect 9256 7040 9264 7104
rect 8944 6016 9264 7040
rect 8944 5952 8952 6016
rect 9016 5952 9032 6016
rect 9096 5952 9112 6016
rect 9176 5952 9192 6016
rect 9256 5952 9264 6016
rect 8944 4928 9264 5952
rect 8944 4864 8952 4928
rect 9016 4864 9032 4928
rect 9096 4864 9112 4928
rect 9176 4864 9192 4928
rect 9256 4864 9264 4928
rect 8944 3840 9264 4864
rect 8944 3776 8952 3840
rect 9016 3776 9032 3840
rect 9096 3776 9112 3840
rect 9176 3776 9192 3840
rect 9256 3776 9264 3840
rect 8944 2752 9264 3776
rect 8944 2688 8952 2752
rect 9016 2688 9032 2752
rect 9096 2688 9112 2752
rect 9176 2688 9192 2752
rect 9256 2688 9264 2752
rect 8944 2128 9264 2688
rect 12944 21792 13264 21808
rect 12944 21728 12952 21792
rect 13016 21728 13032 21792
rect 13096 21728 13112 21792
rect 13176 21728 13192 21792
rect 13256 21728 13264 21792
rect 12944 20704 13264 21728
rect 12944 20640 12952 20704
rect 13016 20640 13032 20704
rect 13096 20640 13112 20704
rect 13176 20640 13192 20704
rect 13256 20640 13264 20704
rect 12944 19616 13264 20640
rect 12944 19552 12952 19616
rect 13016 19552 13032 19616
rect 13096 19552 13112 19616
rect 13176 19552 13192 19616
rect 13256 19552 13264 19616
rect 12944 18528 13264 19552
rect 12944 18464 12952 18528
rect 13016 18464 13032 18528
rect 13096 18464 13112 18528
rect 13176 18464 13192 18528
rect 13256 18464 13264 18528
rect 12944 17440 13264 18464
rect 12944 17376 12952 17440
rect 13016 17376 13032 17440
rect 13096 17376 13112 17440
rect 13176 17376 13192 17440
rect 13256 17376 13264 17440
rect 12944 16352 13264 17376
rect 12944 16288 12952 16352
rect 13016 16288 13032 16352
rect 13096 16288 13112 16352
rect 13176 16288 13192 16352
rect 13256 16288 13264 16352
rect 12944 15264 13264 16288
rect 12944 15200 12952 15264
rect 13016 15200 13032 15264
rect 13096 15200 13112 15264
rect 13176 15200 13192 15264
rect 13256 15200 13264 15264
rect 12944 14176 13264 15200
rect 12944 14112 12952 14176
rect 13016 14112 13032 14176
rect 13096 14112 13112 14176
rect 13176 14112 13192 14176
rect 13256 14112 13264 14176
rect 12944 13088 13264 14112
rect 12944 13024 12952 13088
rect 13016 13024 13032 13088
rect 13096 13024 13112 13088
rect 13176 13024 13192 13088
rect 13256 13024 13264 13088
rect 12944 12000 13264 13024
rect 12944 11936 12952 12000
rect 13016 11936 13032 12000
rect 13096 11936 13112 12000
rect 13176 11936 13192 12000
rect 13256 11936 13264 12000
rect 12944 10912 13264 11936
rect 12944 10848 12952 10912
rect 13016 10848 13032 10912
rect 13096 10848 13112 10912
rect 13176 10848 13192 10912
rect 13256 10848 13264 10912
rect 12944 9824 13264 10848
rect 12944 9760 12952 9824
rect 13016 9760 13032 9824
rect 13096 9760 13112 9824
rect 13176 9760 13192 9824
rect 13256 9760 13264 9824
rect 12944 8736 13264 9760
rect 12944 8672 12952 8736
rect 13016 8672 13032 8736
rect 13096 8672 13112 8736
rect 13176 8672 13192 8736
rect 13256 8672 13264 8736
rect 12944 7648 13264 8672
rect 12944 7584 12952 7648
rect 13016 7584 13032 7648
rect 13096 7584 13112 7648
rect 13176 7584 13192 7648
rect 13256 7584 13264 7648
rect 12944 6560 13264 7584
rect 12944 6496 12952 6560
rect 13016 6496 13032 6560
rect 13096 6496 13112 6560
rect 13176 6496 13192 6560
rect 13256 6496 13264 6560
rect 12944 5472 13264 6496
rect 12944 5408 12952 5472
rect 13016 5408 13032 5472
rect 13096 5408 13112 5472
rect 13176 5408 13192 5472
rect 13256 5408 13264 5472
rect 12944 4384 13264 5408
rect 12944 4320 12952 4384
rect 13016 4320 13032 4384
rect 13096 4320 13112 4384
rect 13176 4320 13192 4384
rect 13256 4320 13264 4384
rect 12944 3296 13264 4320
rect 12944 3232 12952 3296
rect 13016 3232 13032 3296
rect 13096 3232 13112 3296
rect 13176 3232 13192 3296
rect 13256 3232 13264 3296
rect 12944 2208 13264 3232
rect 12944 2144 12952 2208
rect 13016 2144 13032 2208
rect 13096 2144 13112 2208
rect 13176 2144 13192 2208
rect 13256 2144 13264 2208
rect 12944 2128 13264 2144
rect 16944 21248 17264 21808
rect 16944 21184 16952 21248
rect 17016 21184 17032 21248
rect 17096 21184 17112 21248
rect 17176 21184 17192 21248
rect 17256 21184 17264 21248
rect 16944 20160 17264 21184
rect 16944 20096 16952 20160
rect 17016 20096 17032 20160
rect 17096 20096 17112 20160
rect 17176 20096 17192 20160
rect 17256 20096 17264 20160
rect 16944 19072 17264 20096
rect 16944 19008 16952 19072
rect 17016 19008 17032 19072
rect 17096 19008 17112 19072
rect 17176 19008 17192 19072
rect 17256 19008 17264 19072
rect 16944 17984 17264 19008
rect 16944 17920 16952 17984
rect 17016 17920 17032 17984
rect 17096 17920 17112 17984
rect 17176 17920 17192 17984
rect 17256 17920 17264 17984
rect 16944 16896 17264 17920
rect 16944 16832 16952 16896
rect 17016 16832 17032 16896
rect 17096 16832 17112 16896
rect 17176 16832 17192 16896
rect 17256 16832 17264 16896
rect 16944 15808 17264 16832
rect 16944 15744 16952 15808
rect 17016 15744 17032 15808
rect 17096 15744 17112 15808
rect 17176 15744 17192 15808
rect 17256 15744 17264 15808
rect 16944 14720 17264 15744
rect 16944 14656 16952 14720
rect 17016 14656 17032 14720
rect 17096 14656 17112 14720
rect 17176 14656 17192 14720
rect 17256 14656 17264 14720
rect 16944 13632 17264 14656
rect 16944 13568 16952 13632
rect 17016 13568 17032 13632
rect 17096 13568 17112 13632
rect 17176 13568 17192 13632
rect 17256 13568 17264 13632
rect 16944 12544 17264 13568
rect 16944 12480 16952 12544
rect 17016 12480 17032 12544
rect 17096 12480 17112 12544
rect 17176 12480 17192 12544
rect 17256 12480 17264 12544
rect 16944 11456 17264 12480
rect 16944 11392 16952 11456
rect 17016 11392 17032 11456
rect 17096 11392 17112 11456
rect 17176 11392 17192 11456
rect 17256 11392 17264 11456
rect 16944 10368 17264 11392
rect 16944 10304 16952 10368
rect 17016 10304 17032 10368
rect 17096 10304 17112 10368
rect 17176 10304 17192 10368
rect 17256 10304 17264 10368
rect 16944 9280 17264 10304
rect 16944 9216 16952 9280
rect 17016 9216 17032 9280
rect 17096 9216 17112 9280
rect 17176 9216 17192 9280
rect 17256 9216 17264 9280
rect 16944 8192 17264 9216
rect 16944 8128 16952 8192
rect 17016 8128 17032 8192
rect 17096 8128 17112 8192
rect 17176 8128 17192 8192
rect 17256 8128 17264 8192
rect 16944 7104 17264 8128
rect 16944 7040 16952 7104
rect 17016 7040 17032 7104
rect 17096 7040 17112 7104
rect 17176 7040 17192 7104
rect 17256 7040 17264 7104
rect 16944 6016 17264 7040
rect 16944 5952 16952 6016
rect 17016 5952 17032 6016
rect 17096 5952 17112 6016
rect 17176 5952 17192 6016
rect 17256 5952 17264 6016
rect 16944 4928 17264 5952
rect 16944 4864 16952 4928
rect 17016 4864 17032 4928
rect 17096 4864 17112 4928
rect 17176 4864 17192 4928
rect 17256 4864 17264 4928
rect 16944 3840 17264 4864
rect 16944 3776 16952 3840
rect 17016 3776 17032 3840
rect 17096 3776 17112 3840
rect 17176 3776 17192 3840
rect 17256 3776 17264 3840
rect 16944 2752 17264 3776
rect 16944 2688 16952 2752
rect 17016 2688 17032 2752
rect 17096 2688 17112 2752
rect 17176 2688 17192 2752
rect 17256 2688 17264 2752
rect 16944 2128 17264 2688
rect 20944 21792 21264 21808
rect 20944 21728 20952 21792
rect 21016 21728 21032 21792
rect 21096 21728 21112 21792
rect 21176 21728 21192 21792
rect 21256 21728 21264 21792
rect 20944 20704 21264 21728
rect 20944 20640 20952 20704
rect 21016 20640 21032 20704
rect 21096 20640 21112 20704
rect 21176 20640 21192 20704
rect 21256 20640 21264 20704
rect 20944 19616 21264 20640
rect 20944 19552 20952 19616
rect 21016 19552 21032 19616
rect 21096 19552 21112 19616
rect 21176 19552 21192 19616
rect 21256 19552 21264 19616
rect 20944 18528 21264 19552
rect 20944 18464 20952 18528
rect 21016 18464 21032 18528
rect 21096 18464 21112 18528
rect 21176 18464 21192 18528
rect 21256 18464 21264 18528
rect 20944 17440 21264 18464
rect 20944 17376 20952 17440
rect 21016 17376 21032 17440
rect 21096 17376 21112 17440
rect 21176 17376 21192 17440
rect 21256 17376 21264 17440
rect 20944 16352 21264 17376
rect 20944 16288 20952 16352
rect 21016 16288 21032 16352
rect 21096 16288 21112 16352
rect 21176 16288 21192 16352
rect 21256 16288 21264 16352
rect 20944 15264 21264 16288
rect 20944 15200 20952 15264
rect 21016 15200 21032 15264
rect 21096 15200 21112 15264
rect 21176 15200 21192 15264
rect 21256 15200 21264 15264
rect 20944 14176 21264 15200
rect 20944 14112 20952 14176
rect 21016 14112 21032 14176
rect 21096 14112 21112 14176
rect 21176 14112 21192 14176
rect 21256 14112 21264 14176
rect 20944 13088 21264 14112
rect 20944 13024 20952 13088
rect 21016 13024 21032 13088
rect 21096 13024 21112 13088
rect 21176 13024 21192 13088
rect 21256 13024 21264 13088
rect 20944 12000 21264 13024
rect 20944 11936 20952 12000
rect 21016 11936 21032 12000
rect 21096 11936 21112 12000
rect 21176 11936 21192 12000
rect 21256 11936 21264 12000
rect 20944 10912 21264 11936
rect 20944 10848 20952 10912
rect 21016 10848 21032 10912
rect 21096 10848 21112 10912
rect 21176 10848 21192 10912
rect 21256 10848 21264 10912
rect 20944 9824 21264 10848
rect 20944 9760 20952 9824
rect 21016 9760 21032 9824
rect 21096 9760 21112 9824
rect 21176 9760 21192 9824
rect 21256 9760 21264 9824
rect 20944 8736 21264 9760
rect 20944 8672 20952 8736
rect 21016 8672 21032 8736
rect 21096 8672 21112 8736
rect 21176 8672 21192 8736
rect 21256 8672 21264 8736
rect 20944 7648 21264 8672
rect 20944 7584 20952 7648
rect 21016 7584 21032 7648
rect 21096 7584 21112 7648
rect 21176 7584 21192 7648
rect 21256 7584 21264 7648
rect 20944 6560 21264 7584
rect 20944 6496 20952 6560
rect 21016 6496 21032 6560
rect 21096 6496 21112 6560
rect 21176 6496 21192 6560
rect 21256 6496 21264 6560
rect 20944 5472 21264 6496
rect 20944 5408 20952 5472
rect 21016 5408 21032 5472
rect 21096 5408 21112 5472
rect 21176 5408 21192 5472
rect 21256 5408 21264 5472
rect 20944 4384 21264 5408
rect 20944 4320 20952 4384
rect 21016 4320 21032 4384
rect 21096 4320 21112 4384
rect 21176 4320 21192 4384
rect 21256 4320 21264 4384
rect 20944 3296 21264 4320
rect 20944 3232 20952 3296
rect 21016 3232 21032 3296
rect 21096 3232 21112 3296
rect 21176 3232 21192 3296
rect 21256 3232 21264 3296
rect 20944 2208 21264 3232
rect 20944 2144 20952 2208
rect 21016 2144 21032 2208
rect 21096 2144 21112 2208
rect 21176 2144 21192 2208
rect 21256 2144 21264 2208
rect 20944 2128 21264 2144
use scs8hd_decap_3  PHY_0 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1104 0 -1 2720
box -38 -48 314 592
use scs8hd_decap_3  PHY_2
timestamp 1586364061
transform 1 0 1104 0 1 2720
box -38 -48 314 592
use scs8hd_decap_12  FILLER_0_3 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1380 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_15
timestamp 1586364061
transform 1 0 2484 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_3
timestamp 1586364061
transform 1 0 1380 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_15
timestamp 1586364061
transform 1 0 2484 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_72 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 3956 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_4  FILLER_0_27 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 3588 0 -1 2720
box -38 -48 406 592
use scs8hd_decap_12  FILLER_0_32
timestamp 1586364061
transform 1 0 4048 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_27
timestamp 1586364061
transform 1 0 3588 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_44
timestamp 1586364061
transform 1 0 5152 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_39
timestamp 1586364061
transform 1 0 4692 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_1_51 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 5796 0 1 2720
box -38 -48 774 592
use scs8hd_inv_1  mux_top_ipin_2.tap_buf4_0_.scs8hd_inv_1 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 6900 0 -1 2720
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_73
timestamp 1586364061
transform 1 0 6808 0 -1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_79
timestamp 1586364061
transform 1 0 6716 0 1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_2.tap_buf4_0_.scs8hd_inv_1_A tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 7360 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_6  FILLER_0_56 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 6256 0 -1 2720
box -38 -48 590 592
use scs8hd_fill_2  FILLER_0_66 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 7176 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_12  FILLER_0_70
timestamp 1586364061
transform 1 0 7544 0 -1 2720
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_1_59
timestamp 1586364061
transform 1 0 6532 0 1 2720
box -38 -48 222 592
use scs8hd_decap_12  FILLER_1_62
timestamp 1586364061
transform 1 0 6808 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_0_82
timestamp 1586364061
transform 1 0 8648 0 -1 2720
box -38 -48 774 592
use scs8hd_decap_12  FILLER_1_74
timestamp 1586364061
transform 1 0 7912 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_86
timestamp 1586364061
transform 1 0 9016 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_1_98
timestamp 1586364061
transform 1 0 10120 0 1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_0_98
timestamp 1586364061
transform 1 0 10120 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_3  FILLER_0_90
timestamp 1586364061
transform 1 0 9384 0 -1 2720
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_74
timestamp 1586364061
transform 1 0 9660 0 -1 2720
box -38 -48 130 592
use scs8hd_buf_2  _78_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 9752 0 -1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_1_105
timestamp 1586364061
transform 1 0 10764 0 1 2720
box -38 -48 222 592
use scs8hd_fill_1  FILLER_1_102 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 10488 0 1 2720
box -38 -48 130 592
use scs8hd_decap_3  FILLER_0_102
timestamp 1586364061
transform 1 0 10488 0 -1 2720
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__35__A
timestamp 1586364061
transform 1 0 10764 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__37__B
timestamp 1586364061
transform 1 0 10580 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__73__A
timestamp 1586364061
transform 1 0 10948 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__78__A
timestamp 1586364061
transform 1 0 10304 0 -1 2720
box -38 -48 222 592
use scs8hd_inv_8  _35_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 10948 0 -1 2720
box -38 -48 866 592
use scs8hd_fill_2  FILLER_1_113
timestamp 1586364061
transform 1 0 11500 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__37__A
timestamp 1586364061
transform 1 0 11684 0 1 2720
box -38 -48 222 592
use scs8hd_buf_2  _73_
timestamp 1586364061
transform 1 0 11132 0 1 2720
box -38 -48 406 592
use scs8hd_decap_3  FILLER_1_117
timestamp 1586364061
transform 1 0 11868 0 1 2720
box -38 -48 314 592
use scs8hd_decap_6  FILLER_0_116
timestamp 1586364061
transform 1 0 11776 0 -1 2720
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 12328 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_2.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 12144 0 1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_80
timestamp 1586364061
transform 1 0 12328 0 1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_75
timestamp 1586364061
transform 1 0 12512 0 -1 2720
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  mem_top_ipin_2.LATCH_1_.latch tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 12420 0 1 2720
box -38 -48 1050 592
use scs8hd_buf_2  _72_
timestamp 1586364061
transform 1 0 14168 0 1 2720
box -38 -48 406 592
use scs8hd_ebufn_2  mux_top_ipin_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 12972 0 -1 2720
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 12788 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 13616 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 13984 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_125
timestamp 1586364061
transform 1 0 12604 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_8  FILLER_0_138
timestamp 1586364061
transform 1 0 13800 0 -1 2720
box -38 -48 774 592
use scs8hd_fill_2  FILLER_1_134
timestamp 1586364061
transform 1 0 13432 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_138
timestamp 1586364061
transform 1 0 13800 0 1 2720
box -38 -48 222 592
use scs8hd_decap_3  FILLER_1_150
timestamp 1586364061
transform 1 0 14904 0 1 2720
box -38 -48 314 592
use scs8hd_fill_2  FILLER_1_146
timestamp 1586364061
transform 1 0 14536 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_151
timestamp 1586364061
transform 1 0 14996 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_3  FILLER_0_146
timestamp 1586364061
transform 1 0 14536 0 -1 2720
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14812 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__72__A
timestamp 1586364061
transform 1 0 14720 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 15180 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_2.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 15180 0 1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_76
timestamp 1586364061
transform 1 0 15364 0 -1 2720
box -38 -48 130 592
use scs8hd_ebufn_2  mux_top_ipin_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15364 0 1 2720
box -38 -48 866 592
use scs8hd_ebufn_2  mux_top_ipin_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15456 0 -1 2720
box -38 -48 866 592
use scs8hd_fill_2  FILLER_1_168
timestamp 1586364061
transform 1 0 16560 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_164
timestamp 1586364061
transform 1 0 16192 0 1 2720
box -38 -48 222 592
use scs8hd_decap_8  FILLER_0_165
timestamp 1586364061
transform 1 0 16284 0 -1 2720
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 16376 0 1 2720
box -38 -48 222 592
use scs8hd_decap_6  FILLER_1_176
timestamp 1586364061
transform 1 0 17296 0 1 2720
box -38 -48 590 592
use scs8hd_fill_2  FILLER_1_172
timestamp 1586364061
transform 1 0 16928 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_176
timestamp 1586364061
transform 1 0 17296 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 17112 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_2.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 16744 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_2.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 17480 0 -1 2720
box -38 -48 222 592
use scs8hd_inv_1  mux_top_ipin_2.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 17020 0 -1 2720
box -38 -48 314 592
use scs8hd_fill_1  FILLER_1_182
timestamp 1586364061
transform 1 0 17848 0 1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_180
timestamp 1586364061
transform 1 0 17664 0 -1 2720
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_81
timestamp 1586364061
transform 1 0 17940 0 1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_77
timestamp 1586364061
transform 1 0 18216 0 -1 2720
box -38 -48 130 592
use scs8hd_buf_2  _87_
timestamp 1586364061
transform 1 0 18308 0 -1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_0_191
timestamp 1586364061
transform 1 0 18676 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__87__A
timestamp 1586364061
transform 1 0 18860 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_12  FILLER_1_196
timestamp 1586364061
transform 1 0 19136 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_184
timestamp 1586364061
transform 1 0 18032 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_195
timestamp 1586364061
transform 1 0 19044 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_0_207
timestamp 1586364061
transform 1 0 20148 0 -1 2720
box -38 -48 774 592
use scs8hd_decap_12  FILLER_1_208
timestamp 1586364061
transform 1 0 20240 0 1 2720
box -38 -48 1142 592
use scs8hd_buf_2  _82_
timestamp 1586364061
transform 1 0 21160 0 -1 2720
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_78
timestamp 1586364061
transform 1 0 21068 0 -1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__82__A
timestamp 1586364061
transform 1 0 21712 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_215
timestamp 1586364061
transform 1 0 20884 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_222
timestamp 1586364061
transform 1 0 21528 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_6  FILLER_0_226
timestamp 1586364061
transform 1 0 21896 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_1_220
timestamp 1586364061
transform 1 0 21344 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_3  PHY_1
timestamp 1586364061
transform -1 0 22816 0 -1 2720
box -38 -48 314 592
use scs8hd_decap_3  PHY_3
timestamp 1586364061
transform -1 0 22816 0 1 2720
box -38 -48 314 592
use scs8hd_fill_1  FILLER_0_232
timestamp 1586364061
transform 1 0 22448 0 -1 2720
box -38 -48 130 592
use scs8hd_fill_1  FILLER_1_232
timestamp 1586364061
transform 1 0 22448 0 1 2720
box -38 -48 130 592
use scs8hd_decap_3  PHY_4
timestamp 1586364061
transform 1 0 1104 0 -1 3808
box -38 -48 314 592
use scs8hd_decap_12  FILLER_2_3
timestamp 1586364061
transform 1 0 1380 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_15
timestamp 1586364061
transform 1 0 2484 0 -1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_82
timestamp 1586364061
transform 1 0 3956 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_4  FILLER_2_27
timestamp 1586364061
transform 1 0 3588 0 -1 3808
box -38 -48 406 592
use scs8hd_decap_12  FILLER_2_32
timestamp 1586364061
transform 1 0 4048 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_44
timestamp 1586364061
transform 1 0 5152 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_56
timestamp 1586364061
transform 1 0 6256 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_68
timestamp 1586364061
transform 1 0 7360 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_80
timestamp 1586364061
transform 1 0 8464 0 -1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_83
timestamp 1586364061
transform 1 0 9568 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_2_93
timestamp 1586364061
transform 1 0 9660 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_2_105
timestamp 1586364061
transform 1 0 10764 0 -1 3808
box -38 -48 590 592
use scs8hd_or2_4  _37_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 11408 0 -1 3808
box -38 -48 682 592
use scs8hd_diode_2  ANTENNA__64__A
timestamp 1586364061
transform 1 0 12236 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_1  FILLER_2_111
timestamp 1586364061
transform 1 0 11316 0 -1 3808
box -38 -48 130 592
use scs8hd_fill_2  FILLER_2_119
timestamp 1586364061
transform 1 0 12052 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_123
timestamp 1586364061
transform 1 0 12420 0 -1 3808
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_ipin_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 13248 0 -1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_2.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 12604 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_2_127
timestamp 1586364061
transform 1 0 12788 0 -1 3808
box -38 -48 406 592
use scs8hd_fill_1  FILLER_2_131
timestamp 1586364061
transform 1 0 13156 0 -1 3808
box -38 -48 130 592
use scs8hd_fill_2  FILLER_2_141
timestamp 1586364061
transform 1 0 14076 0 -1 3808
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_top_ipin_2.LATCH_0_.latch
timestamp 1586364061
transform 1 0 15272 0 -1 3808
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_84
timestamp 1586364061
transform 1 0 15180 0 -1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__65__C
timestamp 1586364061
transform 1 0 14260 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_8  FILLER_2_145
timestamp 1586364061
transform 1 0 14444 0 -1 3808
box -38 -48 774 592
use scs8hd_conb_1  _70_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 17112 0 -1 3808
box -38 -48 314 592
use scs8hd_decap_8  FILLER_2_165
timestamp 1586364061
transform 1 0 16284 0 -1 3808
box -38 -48 774 592
use scs8hd_fill_1  FILLER_2_173
timestamp 1586364061
transform 1 0 17020 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_2_177
timestamp 1586364061
transform 1 0 17388 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_189
timestamp 1586364061
transform 1 0 18492 0 -1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_85
timestamp 1586364061
transform 1 0 20792 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_2_201
timestamp 1586364061
transform 1 0 19596 0 -1 3808
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_2_213
timestamp 1586364061
transform 1 0 20700 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_2_215
timestamp 1586364061
transform 1 0 20884 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_2_227
timestamp 1586364061
transform 1 0 21988 0 -1 3808
box -38 -48 590 592
use scs8hd_decap_3  PHY_5
timestamp 1586364061
transform -1 0 22816 0 -1 3808
box -38 -48 314 592
use scs8hd_decap_3  PHY_6
timestamp 1586364061
transform 1 0 1104 0 1 3808
box -38 -48 314 592
use scs8hd_decap_12  FILLER_3_3
timestamp 1586364061
transform 1 0 1380 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_15
timestamp 1586364061
transform 1 0 2484 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_27
timestamp 1586364061
transform 1 0 3588 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_39
timestamp 1586364061
transform 1 0 4692 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_3_51
timestamp 1586364061
transform 1 0 5796 0 1 3808
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_86
timestamp 1586364061
transform 1 0 6716 0 1 3808
box -38 -48 130 592
use scs8hd_fill_2  FILLER_3_59
timestamp 1586364061
transform 1 0 6532 0 1 3808
box -38 -48 222 592
use scs8hd_decap_12  FILLER_3_62
timestamp 1586364061
transform 1 0 6808 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_74
timestamp 1586364061
transform 1 0 7912 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_3_86
timestamp 1586364061
transform 1 0 9016 0 1 3808
box -38 -48 590 592
use scs8hd_inv_8  _27_
timestamp 1586364061
transform 1 0 10764 0 1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__27__A
timestamp 1586364061
transform 1 0 10580 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__30__A
timestamp 1586364061
transform 1 0 9660 0 1 3808
box -38 -48 222 592
use scs8hd_fill_1  FILLER_3_92
timestamp 1586364061
transform 1 0 9568 0 1 3808
box -38 -48 130 592
use scs8hd_decap_8  FILLER_3_95
timestamp 1586364061
transform 1 0 9844 0 1 3808
box -38 -48 774 592
use scs8hd_conb_1  _71_
timestamp 1586364061
transform 1 0 12420 0 1 3808
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_87
timestamp 1586364061
transform 1 0 12328 0 1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__64__B
timestamp 1586364061
transform 1 0 11776 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__64__D
timestamp 1586364061
transform 1 0 12144 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_114
timestamp 1586364061
transform 1 0 11592 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_118
timestamp 1586364061
transform 1 0 11960 0 1 3808
box -38 -48 222 592
use scs8hd_nor4_4  _65_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 13432 0 1 3808
box -38 -48 1602 592
use scs8hd_diode_2  ANTENNA__65__D
timestamp 1586364061
transform 1 0 13248 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__65__A
timestamp 1586364061
transform 1 0 12880 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_126
timestamp 1586364061
transform 1 0 12696 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_130
timestamp 1586364061
transform 1 0 13064 0 1 3808
box -38 -48 222 592
use scs8hd_inv_8  _36_
timestamp 1586364061
transform 1 0 15732 0 1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__36__A
timestamp 1586364061
transform 1 0 15548 0 1 3808
box -38 -48 222 592
use scs8hd_decap_6  FILLER_3_151
timestamp 1586364061
transform 1 0 14996 0 1 3808
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 16836 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 17204 0 1 3808
box -38 -48 222 592
use scs8hd_decap_3  FILLER_3_168
timestamp 1586364061
transform 1 0 16560 0 1 3808
box -38 -48 314 592
use scs8hd_fill_2  FILLER_3_173
timestamp 1586364061
transform 1 0 17020 0 1 3808
box -38 -48 222 592
use scs8hd_decap_6  FILLER_3_177
timestamp 1586364061
transform 1 0 17388 0 1 3808
box -38 -48 590 592
use scs8hd_inv_1  mux_top_ipin_1.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 18032 0 1 3808
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_88
timestamp 1586364061
transform 1 0 17940 0 1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__33__A
timestamp 1586364061
transform 1 0 18492 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_1.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 18860 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_187
timestamp 1586364061
transform 1 0 18308 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_191
timestamp 1586364061
transform 1 0 18676 0 1 3808
box -38 -48 222 592
use scs8hd_decap_12  FILLER_3_195
timestamp 1586364061
transform 1 0 19044 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_207
timestamp 1586364061
transform 1 0 20148 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_219
timestamp 1586364061
transform 1 0 21252 0 1 3808
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_3_231
timestamp 1586364061
transform 1 0 22356 0 1 3808
box -38 -48 222 592
use scs8hd_decap_3  PHY_7
timestamp 1586364061
transform -1 0 22816 0 1 3808
box -38 -48 314 592
use scs8hd_decap_3  PHY_8
timestamp 1586364061
transform 1 0 1104 0 -1 4896
box -38 -48 314 592
use scs8hd_decap_12  FILLER_4_3
timestamp 1586364061
transform 1 0 1380 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_15
timestamp 1586364061
transform 1 0 2484 0 -1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_89
timestamp 1586364061
transform 1 0 3956 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_4  FILLER_4_27
timestamp 1586364061
transform 1 0 3588 0 -1 4896
box -38 -48 406 592
use scs8hd_decap_12  FILLER_4_32
timestamp 1586364061
transform 1 0 4048 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_44
timestamp 1586364061
transform 1 0 5152 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_56
timestamp 1586364061
transform 1 0 6256 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_68
timestamp 1586364061
transform 1 0 7360 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_80
timestamp 1586364061
transform 1 0 8464 0 -1 4896
box -38 -48 1142 592
use scs8hd_inv_8  _30_
timestamp 1586364061
transform 1 0 9660 0 -1 4896
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_90
timestamp 1586364061
transform 1 0 9568 0 -1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__38__A
timestamp 1586364061
transform 1 0 10672 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_102
timestamp 1586364061
transform 1 0 10488 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_6  FILLER_4_106
timestamp 1586364061
transform 1 0 10856 0 -1 4896
box -38 -48 590 592
use scs8hd_nor4_4  _64_
timestamp 1586364061
transform 1 0 11592 0 -1 4896
box -38 -48 1602 592
use scs8hd_diode_2  ANTENNA__64__C
timestamp 1586364061
transform 1 0 11408 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__65__B
timestamp 1586364061
transform 1 0 13432 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__62__D
timestamp 1586364061
transform 1 0 13800 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__62__A
timestamp 1586364061
transform 1 0 14168 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_3  FILLER_4_131
timestamp 1586364061
transform 1 0 13156 0 -1 4896
box -38 -48 314 592
use scs8hd_fill_2  FILLER_4_136
timestamp 1586364061
transform 1 0 13616 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_140
timestamp 1586364061
transform 1 0 13984 0 -1 4896
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_91
timestamp 1586364061
transform 1 0 15180 0 -1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_1.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 15640 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_8  FILLER_4_144
timestamp 1586364061
transform 1 0 14352 0 -1 4896
box -38 -48 774 592
use scs8hd_fill_1  FILLER_4_152
timestamp 1586364061
transform 1 0 15088 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_4  FILLER_4_154
timestamp 1586364061
transform 1 0 15272 0 -1 4896
box -38 -48 406 592
use scs8hd_decap_8  FILLER_4_160
timestamp 1586364061
transform 1 0 15824 0 -1 4896
box -38 -48 774 592
use scs8hd_ebufn_2  mux_top_ipin_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 16836 0 -1 4896
box -38 -48 866 592
use scs8hd_decap_3  FILLER_4_168
timestamp 1586364061
transform 1 0 16560 0 -1 4896
box -38 -48 314 592
use scs8hd_inv_8  _33_
timestamp 1586364061
transform 1 0 18400 0 -1 4896
box -38 -48 866 592
use scs8hd_decap_8  FILLER_4_180
timestamp 1586364061
transform 1 0 17664 0 -1 4896
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_92
timestamp 1586364061
transform 1 0 20792 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_4_197
timestamp 1586364061
transform 1 0 19228 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_4_209
timestamp 1586364061
transform 1 0 20332 0 -1 4896
box -38 -48 406 592
use scs8hd_fill_1  FILLER_4_213
timestamp 1586364061
transform 1 0 20700 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_4_215
timestamp 1586364061
transform 1 0 20884 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_4_227
timestamp 1586364061
transform 1 0 21988 0 -1 4896
box -38 -48 590 592
use scs8hd_decap_3  PHY_9
timestamp 1586364061
transform -1 0 22816 0 -1 4896
box -38 -48 314 592
use scs8hd_decap_3  PHY_10
timestamp 1586364061
transform 1 0 1104 0 1 4896
box -38 -48 314 592
use scs8hd_decap_12  FILLER_5_3
timestamp 1586364061
transform 1 0 1380 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_15
timestamp 1586364061
transform 1 0 2484 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_27
timestamp 1586364061
transform 1 0 3588 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_39
timestamp 1586364061
transform 1 0 4692 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_5_51
timestamp 1586364061
transform 1 0 5796 0 1 4896
box -38 -48 774 592
use scs8hd_inv_8  _26_
timestamp 1586364061
transform 1 0 6900 0 1 4896
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_93
timestamp 1586364061
transform 1 0 6716 0 1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__26__A
timestamp 1586364061
transform 1 0 6532 0 1 4896
box -38 -48 222 592
use scs8hd_fill_1  FILLER_5_62
timestamp 1586364061
transform 1 0 6808 0 1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_5_72
timestamp 1586364061
transform 1 0 7728 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_5_84
timestamp 1586364061
transform 1 0 8832 0 1 4896
box -38 -48 774 592
use scs8hd_inv_8  _28_
timestamp 1586364061
transform 1 0 10304 0 1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__38__B
timestamp 1586364061
transform 1 0 10120 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__38__D
timestamp 1586364061
transform 1 0 9752 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_92
timestamp 1586364061
transform 1 0 9568 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_96
timestamp 1586364061
transform 1 0 9936 0 1 4896
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_94
timestamp 1586364061
transform 1 0 12328 0 1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__45__A
timestamp 1586364061
transform 1 0 12144 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__38__C
timestamp 1586364061
transform 1 0 11316 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__45__D
timestamp 1586364061
transform 1 0 11776 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_109
timestamp 1586364061
transform 1 0 11132 0 1 4896
box -38 -48 222 592
use scs8hd_decap_3  FILLER_5_113
timestamp 1586364061
transform 1 0 11500 0 1 4896
box -38 -48 314 592
use scs8hd_fill_2  FILLER_5_118
timestamp 1586364061
transform 1 0 11960 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_123
timestamp 1586364061
transform 1 0 12420 0 1 4896
box -38 -48 222 592
use scs8hd_nor4_4  _62_
timestamp 1586364061
transform 1 0 13340 0 1 4896
box -38 -48 1602 592
use scs8hd_diode_2  ANTENNA__62__B
timestamp 1586364061
transform 1 0 13156 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__45__C
timestamp 1586364061
transform 1 0 12604 0 1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_5_127
timestamp 1586364061
transform 1 0 12788 0 1 4896
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_top_ipin_1.LATCH_1_.latch
timestamp 1586364061
transform 1 0 15640 0 1 4896
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_1.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 15456 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__62__C
timestamp 1586364061
transform 1 0 15088 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_150
timestamp 1586364061
transform 1 0 14904 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_154
timestamp 1586364061
transform 1 0 15272 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 16836 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 17204 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_169
timestamp 1586364061
transform 1 0 16652 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_173
timestamp 1586364061
transform 1 0 17020 0 1 4896
box -38 -48 222 592
use scs8hd_decap_6  FILLER_5_177
timestamp 1586364061
transform 1 0 17388 0 1 4896
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_95
timestamp 1586364061
transform 1 0 17940 0 1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__88__A
timestamp 1586364061
transform 1 0 18308 0 1 4896
box -38 -48 222 592
use scs8hd_decap_3  FILLER_5_184
timestamp 1586364061
transform 1 0 18032 0 1 4896
box -38 -48 314 592
use scs8hd_decap_12  FILLER_5_189
timestamp 1586364061
transform 1 0 18492 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_201
timestamp 1586364061
transform 1 0 19596 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_213
timestamp 1586364061
transform 1 0 20700 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_5_225
timestamp 1586364061
transform 1 0 21804 0 1 4896
box -38 -48 774 592
use scs8hd_decap_3  PHY_11
timestamp 1586364061
transform -1 0 22816 0 1 4896
box -38 -48 314 592
use scs8hd_decap_3  PHY_12
timestamp 1586364061
transform 1 0 1104 0 -1 5984
box -38 -48 314 592
use scs8hd_decap_3  PHY_14
timestamp 1586364061
transform 1 0 1104 0 1 5984
box -38 -48 314 592
use scs8hd_decap_12  FILLER_6_3
timestamp 1586364061
transform 1 0 1380 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_15
timestamp 1586364061
transform 1 0 2484 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_3
timestamp 1586364061
transform 1 0 1380 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_15
timestamp 1586364061
transform 1 0 2484 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_96
timestamp 1586364061
transform 1 0 3956 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_4  FILLER_6_27
timestamp 1586364061
transform 1 0 3588 0 -1 5984
box -38 -48 406 592
use scs8hd_decap_12  FILLER_6_32
timestamp 1586364061
transform 1 0 4048 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_27
timestamp 1586364061
transform 1 0 3588 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_44
timestamp 1586364061
transform 1 0 5152 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_39
timestamp 1586364061
transform 1 0 4692 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_7_51
timestamp 1586364061
transform 1 0 5796 0 1 5984
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_100
timestamp 1586364061
transform 1 0 6716 0 1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_56
timestamp 1586364061
transform 1 0 6256 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_68
timestamp 1586364061
transform 1 0 7360 0 -1 5984
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_7_59
timestamp 1586364061
transform 1 0 6532 0 1 5984
box -38 -48 222 592
use scs8hd_decap_12  FILLER_7_62
timestamp 1586364061
transform 1 0 6808 0 1 5984
box -38 -48 1142 592
use scs8hd_or2_4  _52_
timestamp 1586364061
transform 1 0 9200 0 1 5984
box -38 -48 682 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 8464 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__52__A
timestamp 1586364061
transform 1 0 9016 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__52__B
timestamp 1586364061
transform 1 0 9200 0 -1 5984
box -38 -48 222 592
use scs8hd_decap_8  FILLER_6_80
timestamp 1586364061
transform 1 0 8464 0 -1 5984
box -38 -48 774 592
use scs8hd_decap_6  FILLER_7_74
timestamp 1586364061
transform 1 0 7912 0 1 5984
box -38 -48 590 592
use scs8hd_decap_4  FILLER_7_82
timestamp 1586364061
transform 1 0 8648 0 1 5984
box -38 -48 406 592
use scs8hd_fill_2  FILLER_7_95
timestamp 1586364061
transform 1 0 9844 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_98
timestamp 1586364061
transform 1 0 10120 0 -1 5984
box -38 -48 222 592
use scs8hd_decap_3  FILLER_6_93
timestamp 1586364061
transform 1 0 9660 0 -1 5984
box -38 -48 314 592
use scs8hd_fill_2  FILLER_6_90
timestamp 1586364061
transform 1 0 9384 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__53__D
timestamp 1586364061
transform 1 0 9936 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__53__A
timestamp 1586364061
transform 1 0 10028 0 1 5984
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_97
timestamp 1586364061
transform 1 0 9568 0 -1 5984
box -38 -48 130 592
use scs8hd_fill_2  FILLER_7_99
timestamp 1586364061
transform 1 0 10212 0 1 5984
box -38 -48 222 592
use scs8hd_fill_1  FILLER_6_102
timestamp 1586364061
transform 1 0 10488 0 -1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__28__A
timestamp 1586364061
transform 1 0 10304 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__29__A
timestamp 1586364061
transform 1 0 10396 0 1 5984
box -38 -48 222 592
use scs8hd_or4_4  _38_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 10580 0 -1 5984
box -38 -48 866 592
use scs8hd_inv_8  _29_
timestamp 1586364061
transform 1 0 10580 0 1 5984
box -38 -48 866 592
use scs8hd_or4_4  _45_
timestamp 1586364061
transform 1 0 12144 0 -1 5984
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_101
timestamp 1586364061
transform 1 0 12328 0 1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__61__B
timestamp 1586364061
transform 1 0 12144 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__53__B
timestamp 1586364061
transform 1 0 11592 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__45__B
timestamp 1586364061
transform 1 0 11960 0 -1 5984
box -38 -48 222 592
use scs8hd_decap_6  FILLER_6_112
timestamp 1586364061
transform 1 0 11408 0 -1 5984
box -38 -48 590 592
use scs8hd_fill_2  FILLER_7_112
timestamp 1586364061
transform 1 0 11408 0 1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_7_116
timestamp 1586364061
transform 1 0 11776 0 1 5984
box -38 -48 406 592
use scs8hd_decap_4  FILLER_7_123
timestamp 1586364061
transform 1 0 12420 0 1 5984
box -38 -48 406 592
use scs8hd_fill_2  FILLER_7_130
timestamp 1586364061
transform 1 0 13064 0 1 5984
box -38 -48 222 592
use scs8hd_fill_1  FILLER_7_127
timestamp 1586364061
transform 1 0 12788 0 1 5984
box -38 -48 130 592
use scs8hd_fill_1  FILLER_6_133
timestamp 1586364061
transform 1 0 13340 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_4  FILLER_6_129
timestamp 1586364061
transform 1 0 12972 0 -1 5984
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__61__D
timestamp 1586364061
transform 1 0 12880 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__63__D
timestamp 1586364061
transform 1 0 13248 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_140
timestamp 1586364061
transform 1 0 13984 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_136
timestamp 1586364061
transform 1 0 13616 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__63__C
timestamp 1586364061
transform 1 0 14168 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__63__A
timestamp 1586364061
transform 1 0 13800 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__63__B
timestamp 1586364061
transform 1 0 13432 0 -1 5984
box -38 -48 222 592
use scs8hd_nor4_4  _63_
timestamp 1586364061
transform 1 0 13432 0 1 5984
box -38 -48 1602 592
use scs8hd_decap_3  FILLER_7_151
timestamp 1586364061
transform 1 0 14996 0 1 5984
box -38 -48 314 592
use scs8hd_decap_8  FILLER_6_144
timestamp 1586364061
transform 1 0 14352 0 -1 5984
box -38 -48 774 592
use scs8hd_decap_3  FILLER_7_156
timestamp 1586364061
transform 1 0 15456 0 1 5984
box -38 -48 314 592
use scs8hd_fill_1  FILLER_6_158
timestamp 1586364061
transform 1 0 15640 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_4  FILLER_6_154
timestamp 1586364061
transform 1 0 15272 0 -1 5984
box -38 -48 406 592
use scs8hd_fill_1  FILLER_6_152
timestamp 1586364061
transform 1 0 15088 0 -1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_1.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 15732 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_2.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 15272 0 1 5984
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_98
timestamp 1586364061
transform 1 0 15180 0 -1 5984
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  mem_top_ipin_1.LATCH_0_.latch
timestamp 1586364061
transform 1 0 15732 0 1 5984
box -38 -48 1050 592
use scs8hd_ebufn_2  mux_top_ipin_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 16744 0 -1 5984
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 16928 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_1.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 16100 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 17388 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_161
timestamp 1586364061
transform 1 0 15916 0 -1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_6_165
timestamp 1586364061
transform 1 0 16284 0 -1 5984
box -38 -48 406 592
use scs8hd_fill_1  FILLER_6_169
timestamp 1586364061
transform 1 0 16652 0 -1 5984
box -38 -48 130 592
use scs8hd_fill_2  FILLER_7_170
timestamp 1586364061
transform 1 0 16744 0 1 5984
box -38 -48 222 592
use scs8hd_decap_3  FILLER_7_174
timestamp 1586364061
transform 1 0 17112 0 1 5984
box -38 -48 314 592
use scs8hd_fill_2  FILLER_7_179
timestamp 1586364061
transform 1 0 17572 0 1 5984
box -38 -48 222 592
use scs8hd_fill_1  FILLER_6_186
timestamp 1586364061
transform 1 0 18216 0 -1 5984
box -38 -48 130 592
use scs8hd_fill_1  FILLER_6_183
timestamp 1586364061
transform 1 0 17940 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_4  FILLER_6_179
timestamp 1586364061
transform 1 0 17572 0 -1 5984
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__32__A
timestamp 1586364061
transform 1 0 18032 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 17756 0 1 5984
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_102
timestamp 1586364061
transform 1 0 17940 0 1 5984
box -38 -48 130 592
use scs8hd_buf_2  _88_
timestamp 1586364061
transform 1 0 18308 0 -1 5984
box -38 -48 406 592
use scs8hd_decap_12  FILLER_7_193
timestamp 1586364061
transform 1 0 18860 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_191
timestamp 1586364061
transform 1 0 18676 0 -1 5984
box -38 -48 1142 592
use scs8hd_inv_8  _32_
timestamp 1586364061
transform 1 0 18032 0 1 5984
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_99
timestamp 1586364061
transform 1 0 20792 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_8  FILLER_6_203
timestamp 1586364061
transform 1 0 19780 0 -1 5984
box -38 -48 774 592
use scs8hd_decap_3  FILLER_6_211
timestamp 1586364061
transform 1 0 20516 0 -1 5984
box -38 -48 314 592
use scs8hd_decap_12  FILLER_7_205
timestamp 1586364061
transform 1 0 19964 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_215
timestamp 1586364061
transform 1 0 20884 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_6_227
timestamp 1586364061
transform 1 0 21988 0 -1 5984
box -38 -48 590 592
use scs8hd_decap_12  FILLER_7_217
timestamp 1586364061
transform 1 0 21068 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_7_229
timestamp 1586364061
transform 1 0 22172 0 1 5984
box -38 -48 406 592
use scs8hd_decap_3  PHY_13
timestamp 1586364061
transform -1 0 22816 0 -1 5984
box -38 -48 314 592
use scs8hd_decap_3  PHY_15
timestamp 1586364061
transform -1 0 22816 0 1 5984
box -38 -48 314 592
use scs8hd_decap_3  PHY_16
timestamp 1586364061
transform 1 0 1104 0 -1 7072
box -38 -48 314 592
use scs8hd_decap_12  FILLER_8_3
timestamp 1586364061
transform 1 0 1380 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_15
timestamp 1586364061
transform 1 0 2484 0 -1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_103
timestamp 1586364061
transform 1 0 3956 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_4  FILLER_8_27
timestamp 1586364061
transform 1 0 3588 0 -1 7072
box -38 -48 406 592
use scs8hd_decap_12  FILLER_8_32
timestamp 1586364061
transform 1 0 4048 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_44
timestamp 1586364061
transform 1 0 5152 0 -1 7072
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA__58__B
timestamp 1586364061
transform 1 0 6808 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__58__C
timestamp 1586364061
transform 1 0 7176 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__58__D
timestamp 1586364061
transform 1 0 7544 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_6  FILLER_8_56
timestamp 1586364061
transform 1 0 6256 0 -1 7072
box -38 -48 590 592
use scs8hd_fill_2  FILLER_8_64
timestamp 1586364061
transform 1 0 6992 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_68
timestamp 1586364061
transform 1 0 7360 0 -1 7072
box -38 -48 222 592
use scs8hd_inv_1  mux_top_ipin_0.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 8464 0 -1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__59__A
timestamp 1586364061
transform 1 0 9108 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_8  FILLER_8_72
timestamp 1586364061
transform 1 0 7728 0 -1 7072
box -38 -48 774 592
use scs8hd_decap_4  FILLER_8_83
timestamp 1586364061
transform 1 0 8740 0 -1 7072
box -38 -48 406 592
use scs8hd_decap_3  FILLER_8_89
timestamp 1586364061
transform 1 0 9292 0 -1 7072
box -38 -48 314 592
use scs8hd_or4_4  _53_
timestamp 1586364061
transform 1 0 10396 0 -1 7072
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_104
timestamp 1586364061
transform 1 0 9568 0 -1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_0.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 9844 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__53__C
timestamp 1586364061
transform 1 0 10212 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_93
timestamp 1586364061
transform 1 0 9660 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_97
timestamp 1586364061
transform 1 0 10028 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__61__C
timestamp 1586364061
transform 1 0 12328 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_12  FILLER_8_110
timestamp 1586364061
transform 1 0 11224 0 -1 7072
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_8_124
timestamp 1586364061
transform 1 0 12512 0 -1 7072
box -38 -48 222 592
use scs8hd_nor4_4  _61_
timestamp 1586364061
transform 1 0 12880 0 -1 7072
box -38 -48 1602 592
use scs8hd_diode_2  ANTENNA__61__A
timestamp 1586364061
transform 1 0 12696 0 -1 7072
box -38 -48 222 592
use scs8hd_inv_1  mux_top_ipin_2.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 15272 0 -1 7072
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_105
timestamp 1586364061
transform 1 0 15180 0 -1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_1.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 15732 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_8  FILLER_8_145
timestamp 1586364061
transform 1 0 14444 0 -1 7072
box -38 -48 774 592
use scs8hd_fill_2  FILLER_8_157
timestamp 1586364061
transform 1 0 15548 0 -1 7072
box -38 -48 222 592
use scs8hd_inv_1  mux_bottom_ipin_1.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 16744 0 -1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_1.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 16100 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_161
timestamp 1586364061
transform 1 0 15916 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_8_165
timestamp 1586364061
transform 1 0 16284 0 -1 7072
box -38 -48 406 592
use scs8hd_fill_1  FILLER_8_169
timestamp 1586364061
transform 1 0 16652 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_8  FILLER_8_173
timestamp 1586364061
transform 1 0 17020 0 -1 7072
box -38 -48 774 592
use scs8hd_ebufn_2  mux_bottom_ipin_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 17756 0 -1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 18952 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_8_190
timestamp 1586364061
transform 1 0 18584 0 -1 7072
box -38 -48 406 592
use scs8hd_fill_2  FILLER_8_196
timestamp 1586364061
transform 1 0 19136 0 -1 7072
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_106
timestamp 1586364061
transform 1 0 20792 0 -1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 19320 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_12  FILLER_8_200
timestamp 1586364061
transform 1 0 19504 0 -1 7072
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_8_212
timestamp 1586364061
transform 1 0 20608 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_12  FILLER_8_215
timestamp 1586364061
transform 1 0 20884 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_8_227
timestamp 1586364061
transform 1 0 21988 0 -1 7072
box -38 -48 590 592
use scs8hd_decap_3  PHY_17
timestamp 1586364061
transform -1 0 22816 0 -1 7072
box -38 -48 314 592
use scs8hd_decap_3  PHY_18
timestamp 1586364061
transform 1 0 1104 0 1 7072
box -38 -48 314 592
use scs8hd_decap_12  FILLER_9_3
timestamp 1586364061
transform 1 0 1380 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_15
timestamp 1586364061
transform 1 0 2484 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_27
timestamp 1586364061
transform 1 0 3588 0 1 7072
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_0.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 5796 0 1 7072
box -38 -48 222 592
use scs8hd_decap_12  FILLER_9_39
timestamp 1586364061
transform 1 0 4692 0 1 7072
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_9_53
timestamp 1586364061
transform 1 0 5980 0 1 7072
box -38 -48 222 592
use scs8hd_nor4_4  _58_
timestamp 1586364061
transform 1 0 6808 0 1 7072
box -38 -48 1602 592
use scs8hd_tapvpwrvgnd_1  PHY_107
timestamp 1586364061
transform 1 0 6716 0 1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__58__A
timestamp 1586364061
transform 1 0 6532 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_0.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 6164 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_57
timestamp 1586364061
transform 1 0 6348 0 1 7072
box -38 -48 222 592
use scs8hd_nor4_4  _59_
timestamp 1586364061
transform 1 0 9108 0 1 7072
box -38 -48 1602 592
use scs8hd_diode_2  ANTENNA__59__C
timestamp 1586364061
transform 1 0 8924 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 8556 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_79
timestamp 1586364061
transform 1 0 8372 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_83
timestamp 1586364061
transform 1 0 8740 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__59__D
timestamp 1586364061
transform 1 0 10856 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_104
timestamp 1586364061
transform 1 0 10672 0 1 7072
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_108
timestamp 1586364061
transform 1 0 12328 0 1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 11408 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11776 0 1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_9_108
timestamp 1586364061
transform 1 0 11040 0 1 7072
box -38 -48 406 592
use scs8hd_fill_2  FILLER_9_114
timestamp 1586364061
transform 1 0 11592 0 1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_9_118
timestamp 1586364061
transform 1 0 11960 0 1 7072
box -38 -48 406 592
use scs8hd_fill_2  FILLER_9_123
timestamp 1586364061
transform 1 0 12420 0 1 7072
box -38 -48 222 592
use scs8hd_nor4_4  _60_
timestamp 1586364061
transform 1 0 13156 0 1 7072
box -38 -48 1602 592
use scs8hd_diode_2  ANTENNA__60__B
timestamp 1586364061
transform 1 0 12972 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__60__D
timestamp 1586364061
transform 1 0 12604 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_127
timestamp 1586364061
transform 1 0 12788 0 1 7072
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_1.LATCH_0_.latch
timestamp 1586364061
transform 1 0 15640 0 1 7072
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_1.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 15364 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_1.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 14996 0 1 7072
box -38 -48 222 592
use scs8hd_decap_3  FILLER_9_148
timestamp 1586364061
transform 1 0 14720 0 1 7072
box -38 -48 314 592
use scs8hd_fill_2  FILLER_9_153
timestamp 1586364061
transform 1 0 15180 0 1 7072
box -38 -48 222 592
use scs8hd_fill_1  FILLER_9_157
timestamp 1586364061
transform 1 0 15548 0 1 7072
box -38 -48 130 592
use scs8hd_decap_8  FILLER_9_169
timestamp 1586364061
transform 1 0 16652 0 1 7072
box -38 -48 774 592
use scs8hd_decap_3  FILLER_9_177
timestamp 1586364061
transform 1 0 17388 0 1 7072
box -38 -48 314 592
use scs8hd_ebufn_2  mux_bottom_ipin_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18952 0 1 7072
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_109
timestamp 1586364061
transform 1 0 17940 0 1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 17664 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 18768 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 18216 0 1 7072
box -38 -48 222 592
use scs8hd_fill_1  FILLER_9_182
timestamp 1586364061
transform 1 0 17848 0 1 7072
box -38 -48 130 592
use scs8hd_fill_2  FILLER_9_184
timestamp 1586364061
transform 1 0 18032 0 1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_9_188
timestamp 1586364061
transform 1 0 18400 0 1 7072
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 19964 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_203
timestamp 1586364061
transform 1 0 19780 0 1 7072
box -38 -48 222 592
use scs8hd_decap_12  FILLER_9_207
timestamp 1586364061
transform 1 0 20148 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_219
timestamp 1586364061
transform 1 0 21252 0 1 7072
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_9_231
timestamp 1586364061
transform 1 0 22356 0 1 7072
box -38 -48 222 592
use scs8hd_decap_3  PHY_19
timestamp 1586364061
transform -1 0 22816 0 1 7072
box -38 -48 314 592
use scs8hd_decap_3  PHY_20
timestamp 1586364061
transform 1 0 1104 0 -1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 1564 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_3
timestamp 1586364061
transform 1 0 1380 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_12  FILLER_10_7
timestamp 1586364061
transform 1 0 1748 0 -1 8160
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_110
timestamp 1586364061
transform 1 0 3956 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_12  FILLER_10_19
timestamp 1586364061
transform 1 0 2852 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_32
timestamp 1586364061
transform 1 0 4048 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_44
timestamp 1586364061
transform 1 0 5152 0 -1 8160
box -38 -48 1142 592
use scs8hd_lpflow_inputisolatch_1  mem_top_ipin_0.LATCH_1_.latch
timestamp 1586364061
transform 1 0 6716 0 -1 8160
box -38 -48 1050 592
use scs8hd_decap_4  FILLER_10_56
timestamp 1586364061
transform 1 0 6256 0 -1 8160
box -38 -48 406 592
use scs8hd_fill_1  FILLER_10_60
timestamp 1586364061
transform 1 0 6624 0 -1 8160
box -38 -48 130 592
use scs8hd_inv_1  mux_top_ipin_0.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 8556 0 -1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__59__B
timestamp 1586364061
transform 1 0 9108 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 8280 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 7912 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_72
timestamp 1586364061
transform 1 0 7728 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_76
timestamp 1586364061
transform 1 0 8096 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_1  FILLER_10_80
timestamp 1586364061
transform 1 0 8464 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_3  FILLER_10_84
timestamp 1586364061
transform 1 0 8832 0 -1 8160
box -38 -48 314 592
use scs8hd_decap_3  FILLER_10_89
timestamp 1586364061
transform 1 0 9292 0 -1 8160
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_top_ipin_0.LATCH_0_.latch
timestamp 1586364061
transform 1 0 9660 0 -1 8160
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_111
timestamp 1586364061
transform 1 0 9568 0 -1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_0.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 10856 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_104
timestamp 1586364061
transform 1 0 10672 0 -1 8160
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_ipin_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 11408 0 -1 8160
box -38 -48 866 592
use scs8hd_decap_4  FILLER_10_108
timestamp 1586364061
transform 1 0 11040 0 -1 8160
box -38 -48 406 592
use scs8hd_decap_8  FILLER_10_121
timestamp 1586364061
transform 1 0 12236 0 -1 8160
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA__60__A
timestamp 1586364061
transform 1 0 13156 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__60__C
timestamp 1586364061
transform 1 0 13524 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_129
timestamp 1586364061
transform 1 0 12972 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_133
timestamp 1586364061
transform 1 0 13340 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_12  FILLER_10_137
timestamp 1586364061
transform 1 0 13708 0 -1 8160
box -38 -48 1142 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_1.LATCH_1_.latch
timestamp 1586364061
transform 1 0 15364 0 -1 8160
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_112
timestamp 1586364061
transform 1 0 15180 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_4  FILLER_10_149
timestamp 1586364061
transform 1 0 14812 0 -1 8160
box -38 -48 406 592
use scs8hd_fill_1  FILLER_10_154
timestamp 1586364061
transform 1 0 15272 0 -1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 17020 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_6  FILLER_10_166
timestamp 1586364061
transform 1 0 16376 0 -1 8160
box -38 -48 590 592
use scs8hd_fill_1  FILLER_10_172
timestamp 1586364061
transform 1 0 16928 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_4  FILLER_10_175
timestamp 1586364061
transform 1 0 17204 0 -1 8160
box -38 -48 406 592
use scs8hd_ebufn_2  mux_bottom_ipin_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 17664 0 -1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__31__A
timestamp 1586364061
transform 1 0 18952 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_1  FILLER_10_179
timestamp 1586364061
transform 1 0 17572 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_4  FILLER_10_189
timestamp 1586364061
transform 1 0 18492 0 -1 8160
box -38 -48 406 592
use scs8hd_fill_1  FILLER_10_193
timestamp 1586364061
transform 1 0 18860 0 -1 8160
box -38 -48 130 592
use scs8hd_fill_1  FILLER_10_196
timestamp 1586364061
transform 1 0 19136 0 -1 8160
box -38 -48 130 592
use scs8hd_ebufn_2  mux_bottom_ipin_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 19228 0 -1 8160
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_113
timestamp 1586364061
transform 1 0 20792 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_8  FILLER_10_206
timestamp 1586364061
transform 1 0 20056 0 -1 8160
box -38 -48 774 592
use scs8hd_conb_1  _67_
timestamp 1586364061
transform 1 0 20884 0 -1 8160
box -38 -48 314 592
use scs8hd_decap_12  FILLER_10_218
timestamp 1586364061
transform 1 0 21160 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_10_230
timestamp 1586364061
transform 1 0 22264 0 -1 8160
box -38 -48 314 592
use scs8hd_decap_3  PHY_21
timestamp 1586364061
transform -1 0 22816 0 -1 8160
box -38 -48 314 592
use scs8hd_buf_2  _84_
timestamp 1586364061
transform 1 0 1380 0 1 8160
box -38 -48 406 592
use scs8hd_decap_3  PHY_22
timestamp 1586364061
transform 1 0 1104 0 1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__84__A
timestamp 1586364061
transform 1 0 1932 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_7
timestamp 1586364061
transform 1 0 1748 0 1 8160
box -38 -48 222 592
use scs8hd_decap_12  FILLER_11_11
timestamp 1586364061
transform 1 0 2116 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_23
timestamp 1586364061
transform 1 0 3220 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_35
timestamp 1586364061
transform 1 0 4324 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_47
timestamp 1586364061
transform 1 0 5428 0 1 8160
box -38 -48 1142 592
use scs8hd_inv_1  mux_top_ipin_0.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 7268 0 1 8160
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_114
timestamp 1586364061
transform 1 0 6716 0 1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 7084 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_59
timestamp 1586364061
transform 1 0 6532 0 1 8160
box -38 -48 222 592
use scs8hd_decap_3  FILLER_11_62
timestamp 1586364061
transform 1 0 6808 0 1 8160
box -38 -48 314 592
use scs8hd_fill_2  FILLER_11_70
timestamp 1586364061
transform 1 0 7544 0 1 8160
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_ipin_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 8280 0 1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 7728 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 9292 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 8096 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_74
timestamp 1586364061
transform 1 0 7912 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_87
timestamp 1586364061
transform 1 0 9108 0 1 8160
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_ipin_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9844 0 1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 9660 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10856 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_91
timestamp 1586364061
transform 1 0 9476 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_104
timestamp 1586364061
transform 1 0 10672 0 1 8160
box -38 -48 222 592
use scs8hd_inv_1  mux_top_ipin_0.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 12420 0 1 8160
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_115
timestamp 1586364061
transform 1 0 12328 0 1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 12144 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11224 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_108
timestamp 1586364061
transform 1 0 11040 0 1 8160
box -38 -48 222 592
use scs8hd_decap_8  FILLER_11_112
timestamp 1586364061
transform 1 0 11408 0 1 8160
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA__51__C
timestamp 1586364061
transform 1 0 12880 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__51__A
timestamp 1586364061
transform 1 0 13248 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__51__B
timestamp 1586364061
transform 1 0 13616 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__51__D
timestamp 1586364061
transform 1 0 13984 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_126
timestamp 1586364061
transform 1 0 12696 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_130
timestamp 1586364061
transform 1 0 13064 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_134
timestamp 1586364061
transform 1 0 13432 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_138
timestamp 1586364061
transform 1 0 13800 0 1 8160
box -38 -48 222 592
use scs8hd_decap_6  FILLER_11_142
timestamp 1586364061
transform 1 0 14168 0 1 8160
box -38 -48 590 592
use scs8hd_inv_1  mux_bottom_ipin_2.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 14996 0 1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 15456 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_2.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 15824 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_2.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 14812 0 1 8160
box -38 -48 222 592
use scs8hd_fill_1  FILLER_11_148
timestamp 1586364061
transform 1 0 14720 0 1 8160
box -38 -48 130 592
use scs8hd_fill_2  FILLER_11_154
timestamp 1586364061
transform 1 0 15272 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_158
timestamp 1586364061
transform 1 0 15640 0 1 8160
box -38 -48 222 592
use scs8hd_inv_1  mux_bottom_ipin_2.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 16652 0 1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 17112 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 17480 0 1 8160
box -38 -48 222 592
use scs8hd_decap_6  FILLER_11_162
timestamp 1586364061
transform 1 0 16008 0 1 8160
box -38 -48 590 592
use scs8hd_fill_1  FILLER_11_168
timestamp 1586364061
transform 1 0 16560 0 1 8160
box -38 -48 130 592
use scs8hd_fill_2  FILLER_11_172
timestamp 1586364061
transform 1 0 16928 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_176
timestamp 1586364061
transform 1 0 17296 0 1 8160
box -38 -48 222 592
use scs8hd_inv_8  _31_
timestamp 1586364061
transform 1 0 18952 0 1 8160
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_116
timestamp 1586364061
transform 1 0 17940 0 1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 18584 0 1 8160
box -38 -48 222 592
use scs8hd_decap_3  FILLER_11_180
timestamp 1586364061
transform 1 0 17664 0 1 8160
box -38 -48 314 592
use scs8hd_decap_6  FILLER_11_184
timestamp 1586364061
transform 1 0 18032 0 1 8160
box -38 -48 590 592
use scs8hd_fill_2  FILLER_11_192
timestamp 1586364061
transform 1 0 18768 0 1 8160
box -38 -48 222 592
use scs8hd_buf_2  _83_
timestamp 1586364061
transform 1 0 20516 0 1 8160
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 19964 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_203
timestamp 1586364061
transform 1 0 19780 0 1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_11_207
timestamp 1586364061
transform 1 0 20148 0 1 8160
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__83__A
timestamp 1586364061
transform 1 0 21068 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 21436 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_215
timestamp 1586364061
transform 1 0 20884 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_219
timestamp 1586364061
transform 1 0 21252 0 1 8160
box -38 -48 222 592
use scs8hd_decap_8  FILLER_11_223
timestamp 1586364061
transform 1 0 21620 0 1 8160
box -38 -48 774 592
use scs8hd_fill_2  FILLER_11_231
timestamp 1586364061
transform 1 0 22356 0 1 8160
box -38 -48 222 592
use scs8hd_decap_3  PHY_23
timestamp 1586364061
transform -1 0 22816 0 1 8160
box -38 -48 314 592
use scs8hd_inv_1  mux_top_ipin_0.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1380 0 -1 9248
box -38 -48 314 592
use scs8hd_decap_3  PHY_24
timestamp 1586364061
transform 1 0 1104 0 -1 9248
box -38 -48 314 592
use scs8hd_decap_12  FILLER_12_6
timestamp 1586364061
transform 1 0 1656 0 -1 9248
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_117
timestamp 1586364061
transform 1 0 3956 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_12  FILLER_12_18
timestamp 1586364061
transform 1 0 2760 0 -1 9248
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_12_30
timestamp 1586364061
transform 1 0 3864 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_6  FILLER_12_32
timestamp 1586364061
transform 1 0 4048 0 -1 9248
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA__55__B
timestamp 1586364061
transform 1 0 5796 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 4692 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_1  FILLER_12_38
timestamp 1586364061
transform 1 0 4600 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_8  FILLER_12_41
timestamp 1586364061
transform 1 0 4876 0 -1 9248
box -38 -48 774 592
use scs8hd_fill_2  FILLER_12_49
timestamp 1586364061
transform 1 0 5612 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_53
timestamp 1586364061
transform 1 0 5980 0 -1 9248
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_ipin_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 7636 0 -1 9248
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__55__D
timestamp 1586364061
transform 1 0 6164 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_0.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 6808 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_12_57
timestamp 1586364061
transform 1 0 6348 0 -1 9248
box -38 -48 406 592
use scs8hd_fill_1  FILLER_12_61
timestamp 1586364061
transform 1 0 6716 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_6  FILLER_12_64
timestamp 1586364061
transform 1 0 6992 0 -1 9248
box -38 -48 590 592
use scs8hd_fill_1  FILLER_12_70
timestamp 1586364061
transform 1 0 7544 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_12  FILLER_12_80
timestamp 1586364061
transform 1 0 8464 0 -1 9248
box -38 -48 1142 592
use scs8hd_inv_1  mux_top_ipin_0.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 9844 0 -1 9248
box -38 -48 314 592
use scs8hd_ebufn_2  mux_top_ipin_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10856 0 -1 9248
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_118
timestamp 1586364061
transform 1 0 9568 0 -1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10304 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10672 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_93
timestamp 1586364061
transform 1 0 9660 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_98
timestamp 1586364061
transform 1 0 10120 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_102
timestamp 1586364061
transform 1 0 10488 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_12  FILLER_12_115
timestamp 1586364061
transform 1 0 11684 0 -1 9248
box -38 -48 1142 592
use scs8hd_nor4_4  _51_
timestamp 1586364061
transform 1 0 12880 0 -1 9248
box -38 -48 1602 592
use scs8hd_fill_1  FILLER_12_127
timestamp 1586364061
transform 1 0 12788 0 -1 9248
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_2.LATCH_0_.latch
timestamp 1586364061
transform 1 0 15272 0 -1 9248
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_119
timestamp 1586364061
transform 1 0 15180 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_8  FILLER_12_145
timestamp 1586364061
transform 1 0 14444 0 -1 9248
box -38 -48 774 592
use scs8hd_ebufn_2  mux_bottom_ipin_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 17020 0 -1 9248
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 16468 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_165
timestamp 1586364061
transform 1 0 16284 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_12_169
timestamp 1586364061
transform 1 0 16652 0 -1 9248
box -38 -48 406 592
use scs8hd_inv_1  mux_bottom_ipin_1.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 18584 0 -1 9248
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 18032 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 18400 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_182
timestamp 1586364061
transform 1 0 17848 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_186
timestamp 1586364061
transform 1 0 18216 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_8  FILLER_12_193
timestamp 1586364061
transform 1 0 18860 0 -1 9248
box -38 -48 774 592
use scs8hd_inv_1  mux_bottom_ipin_2.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 19596 0 -1 9248
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_120
timestamp 1586364061
transform 1 0 20792 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_8  FILLER_12_204
timestamp 1586364061
transform 1 0 19872 0 -1 9248
box -38 -48 774 592
use scs8hd_fill_2  FILLER_12_212
timestamp 1586364061
transform 1 0 20608 0 -1 9248
box -38 -48 222 592
use scs8hd_inv_1  mux_bottom_ipin_1.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 20884 0 -1 9248
box -38 -48 314 592
use scs8hd_decap_12  FILLER_12_218
timestamp 1586364061
transform 1 0 21160 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_12_230
timestamp 1586364061
transform 1 0 22264 0 -1 9248
box -38 -48 314 592
use scs8hd_decap_3  PHY_25
timestamp 1586364061
transform -1 0 22816 0 -1 9248
box -38 -48 314 592
use scs8hd_decap_3  PHY_26
timestamp 1586364061
transform 1 0 1104 0 1 9248
box -38 -48 314 592
use scs8hd_decap_3  PHY_28
timestamp 1586364061
transform 1 0 1104 0 -1 10336
box -38 -48 314 592
use scs8hd_decap_12  FILLER_13_3
timestamp 1586364061
transform 1 0 1380 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_15
timestamp 1586364061
transform 1 0 2484 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_3
timestamp 1586364061
transform 1 0 1380 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_15
timestamp 1586364061
transform 1 0 2484 0 -1 10336
box -38 -48 1142 592
use scs8hd_lpflow_inputisolatch_1  mem_top_ipin_0.LATCH_5_.latch
timestamp 1586364061
transform 1 0 4048 0 -1 10336
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_124
timestamp 1586364061
transform 1 0 3956 0 -1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_0.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 4048 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_0.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 3680 0 1 9248
box -38 -48 222 592
use scs8hd_fill_1  FILLER_13_27
timestamp 1586364061
transform 1 0 3588 0 1 9248
box -38 -48 130 592
use scs8hd_fill_2  FILLER_13_30
timestamp 1586364061
transform 1 0 3864 0 1 9248
box -38 -48 222 592
use scs8hd_decap_3  FILLER_13_34
timestamp 1586364061
transform 1 0 4232 0 1 9248
box -38 -48 314 592
use scs8hd_decap_4  FILLER_14_27
timestamp 1586364061
transform 1 0 3588 0 -1 10336
box -38 -48 406 592
use scs8hd_nor4_4  _55_
timestamp 1586364061
transform 1 0 5796 0 -1 10336
box -38 -48 1602 592
use scs8hd_ebufn_2  mux_top_ipin_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 4692 0 1 9248
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__55__C
timestamp 1586364061
transform 1 0 5796 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 4508 0 1 9248
box -38 -48 222 592
use scs8hd_decap_3  FILLER_13_48
timestamp 1586364061
transform 1 0 5520 0 1 9248
box -38 -48 314 592
use scs8hd_fill_2  FILLER_13_53
timestamp 1586364061
transform 1 0 5980 0 1 9248
box -38 -48 222 592
use scs8hd_decap_8  FILLER_14_43
timestamp 1586364061
transform 1 0 5060 0 -1 10336
box -38 -48 774 592
use scs8hd_lpflow_inputisolatch_1  mem_top_ipin_0.LATCH_4_.latch
timestamp 1586364061
transform 1 0 6808 0 1 9248
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_121
timestamp 1586364061
transform 1 0 6716 0 1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__55__A
timestamp 1586364061
transform 1 0 6164 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_0.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 6532 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_57
timestamp 1586364061
transform 1 0 6348 0 1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_14_68
timestamp 1586364061
transform 1 0 7360 0 -1 10336
box -38 -48 406 592
use scs8hd_fill_2  FILLER_14_79
timestamp 1586364061
transform 1 0 8372 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_75
timestamp 1586364061
transform 1 0 8004 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_1  FILLER_14_72
timestamp 1586364061
transform 1 0 7728 0 -1 10336
box -38 -48 130 592
use scs8hd_fill_2  FILLER_13_77
timestamp 1586364061
transform 1 0 8188 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_73
timestamp 1586364061
transform 1 0 7820 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 8004 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 8372 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__56__C
timestamp 1586364061
transform 1 0 8188 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_0.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 7820 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_1  FILLER_14_89
timestamp 1586364061
transform 1 0 9292 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_6  FILLER_14_83
timestamp 1586364061
transform 1 0 8740 0 -1 10336
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA__56__D
timestamp 1586364061
transform 1 0 8556 0 -1 10336
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_ipin_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 8556 0 1 9248
box -38 -48 866 592
use scs8hd_fill_1  FILLER_14_97
timestamp 1586364061
transform 1 0 10028 0 -1 10336
box -38 -48 130 592
use scs8hd_fill_2  FILLER_14_93
timestamp 1586364061
transform 1 0 9660 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_96
timestamp 1586364061
transform 1 0 9936 0 1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_13_90
timestamp 1586364061
transform 1 0 9384 0 1 9248
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10120 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__57__D
timestamp 1586364061
transform 1 0 9752 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__57__A
timestamp 1586364061
transform 1 0 9384 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__57__B
timestamp 1586364061
transform 1 0 9844 0 -1 10336
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_125
timestamp 1586364061
transform 1 0 9568 0 -1 10336
box -38 -48 130 592
use scs8hd_fill_2  FILLER_14_107
timestamp 1586364061
transform 1 0 10948 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_3  FILLER_13_100
timestamp 1586364061
transform 1 0 10304 0 1 9248
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10580 0 1 9248
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_ipin_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10764 0 1 9248
box -38 -48 866 592
use scs8hd_ebufn_2  mux_top_ipin_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10120 0 -1 10336
box -38 -48 866 592
use scs8hd_inv_8  _25_
timestamp 1586364061
transform 1 0 12236 0 -1 10336
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_122
timestamp 1586364061
transform 1 0 12328 0 1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11132 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_8  FILLER_13_114
timestamp 1586364061
transform 1 0 11592 0 1 9248
box -38 -48 774 592
use scs8hd_fill_2  FILLER_13_123
timestamp 1586364061
transform 1 0 12420 0 1 9248
box -38 -48 222 592
use scs8hd_decap_8  FILLER_14_111
timestamp 1586364061
transform 1 0 11316 0 -1 10336
box -38 -48 774 592
use scs8hd_fill_2  FILLER_14_119
timestamp 1586364061
transform 1 0 12052 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_130
timestamp 1586364061
transform 1 0 13064 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_3  FILLER_13_127
timestamp 1586364061
transform 1 0 12788 0 1 9248
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__25__A
timestamp 1586364061
transform 1 0 12604 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__50__B
timestamp 1586364061
transform 1 0 13248 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__50__A
timestamp 1586364061
transform 1 0 13064 0 1 9248
box -38 -48 222 592
use scs8hd_decap_8  FILLER_14_142
timestamp 1586364061
transform 1 0 14168 0 -1 10336
box -38 -48 774 592
use scs8hd_fill_2  FILLER_14_138
timestamp 1586364061
transform 1 0 13800 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_134
timestamp 1586364061
transform 1 0 13432 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__50__D
timestamp 1586364061
transform 1 0 13984 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__50__C
timestamp 1586364061
transform 1 0 13616 0 -1 10336
box -38 -48 222 592
use scs8hd_nor4_4  _50_
timestamp 1586364061
transform 1 0 13248 0 1 9248
box -38 -48 1602 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_2.LATCH_1_.latch
timestamp 1586364061
transform 1 0 15548 0 1 9248
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_126
timestamp 1586364061
transform 1 0 15180 0 -1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_2.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 15364 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_2.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 15548 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_6  FILLER_13_149
timestamp 1586364061
transform 1 0 14812 0 1 9248
box -38 -48 590 592
use scs8hd_decap_3  FILLER_14_150
timestamp 1586364061
transform 1 0 14904 0 -1 10336
box -38 -48 314 592
use scs8hd_decap_3  FILLER_14_154
timestamp 1586364061
transform 1 0 15272 0 -1 10336
box -38 -48 314 592
use scs8hd_decap_3  FILLER_14_159
timestamp 1586364061
transform 1 0 15732 0 -1 10336
box -38 -48 314 592
use scs8hd_ebufn_2  mux_bottom_ipin_2.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 16008 0 -1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 16744 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 17388 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_168
timestamp 1586364061
transform 1 0 16560 0 1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_13_172
timestamp 1586364061
transform 1 0 16928 0 1 9248
box -38 -48 406 592
use scs8hd_fill_1  FILLER_13_176
timestamp 1586364061
transform 1 0 17296 0 1 9248
box -38 -48 130 592
use scs8hd_decap_8  FILLER_14_171
timestamp 1586364061
transform 1 0 16836 0 -1 10336
box -38 -48 774 592
use scs8hd_inv_1  mux_bottom_ipin_2.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 19136 0 -1 10336
box -38 -48 314 592
use scs8hd_ebufn_2  mux_bottom_ipin_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 17572 0 -1 10336
box -38 -48 866 592
use scs8hd_ebufn_2  mux_bottom_ipin_2.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18032 0 1 9248
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_123
timestamp 1586364061
transform 1 0 17940 0 1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 19136 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 17756 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_179
timestamp 1586364061
transform 1 0 17572 0 1 9248
box -38 -48 222 592
use scs8hd_decap_3  FILLER_13_193
timestamp 1586364061
transform 1 0 18860 0 1 9248
box -38 -48 314 592
use scs8hd_decap_8  FILLER_14_188
timestamp 1586364061
transform 1 0 18400 0 -1 10336
box -38 -48 774 592
use scs8hd_inv_1  mux_bottom_ipin_2.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 19596 0 1 9248
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_127
timestamp 1586364061
transform 1 0 20792 0 -1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 20056 0 1 9248
box -38 -48 222 592
use scs8hd_decap_3  FILLER_13_198
timestamp 1586364061
transform 1 0 19320 0 1 9248
box -38 -48 314 592
use scs8hd_fill_2  FILLER_13_204
timestamp 1586364061
transform 1 0 19872 0 1 9248
box -38 -48 222 592
use scs8hd_decap_12  FILLER_13_208
timestamp 1586364061
transform 1 0 20240 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_199
timestamp 1586364061
transform 1 0 19412 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_14_211
timestamp 1586364061
transform 1 0 20516 0 -1 10336
box -38 -48 314 592
use scs8hd_decap_12  FILLER_13_220
timestamp 1586364061
transform 1 0 21344 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_215
timestamp 1586364061
transform 1 0 20884 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_14_227
timestamp 1586364061
transform 1 0 21988 0 -1 10336
box -38 -48 590 592
use scs8hd_decap_3  PHY_27
timestamp 1586364061
transform -1 0 22816 0 1 9248
box -38 -48 314 592
use scs8hd_decap_3  PHY_29
timestamp 1586364061
transform -1 0 22816 0 -1 10336
box -38 -48 314 592
use scs8hd_fill_1  FILLER_13_232
timestamp 1586364061
transform 1 0 22448 0 1 9248
box -38 -48 130 592
use scs8hd_inv_1  mux_top_ipin_0.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1472 0 1 10336
box -38 -48 314 592
use scs8hd_decap_3  PHY_30
timestamp 1586364061
transform 1 0 1104 0 1 10336
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 1932 0 1 10336
box -38 -48 222 592
use scs8hd_fill_1  FILLER_15_3
timestamp 1586364061
transform 1 0 1380 0 1 10336
box -38 -48 130 592
use scs8hd_fill_2  FILLER_15_7
timestamp 1586364061
transform 1 0 1748 0 1 10336
box -38 -48 222 592
use scs8hd_decap_12  FILLER_15_11
timestamp 1586364061
transform 1 0 2116 0 1 10336
box -38 -48 1142 592
use scs8hd_conb_1  _69_
timestamp 1586364061
transform 1 0 4324 0 1 10336
box -38 -48 314 592
use scs8hd_decap_12  FILLER_15_23
timestamp 1586364061
transform 1 0 3220 0 1 10336
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA__54__A
timestamp 1586364061
transform 1 0 5428 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__54__B
timestamp 1586364061
transform 1 0 5796 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__54__D
timestamp 1586364061
transform 1 0 5060 0 1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_15_38
timestamp 1586364061
transform 1 0 4600 0 1 10336
box -38 -48 406 592
use scs8hd_fill_1  FILLER_15_42
timestamp 1586364061
transform 1 0 4968 0 1 10336
box -38 -48 130 592
use scs8hd_fill_2  FILLER_15_45
timestamp 1586364061
transform 1 0 5244 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_49
timestamp 1586364061
transform 1 0 5612 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_53
timestamp 1586364061
transform 1 0 5980 0 1 10336
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_128
timestamp 1586364061
transform 1 0 6716 0 1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__56__B
timestamp 1586364061
transform 1 0 7636 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__56__A
timestamp 1586364061
transform 1 0 7268 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__54__C
timestamp 1586364061
transform 1 0 6164 0 1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_15_57
timestamp 1586364061
transform 1 0 6348 0 1 10336
box -38 -48 406 592
use scs8hd_decap_4  FILLER_15_62
timestamp 1586364061
transform 1 0 6808 0 1 10336
box -38 -48 406 592
use scs8hd_fill_1  FILLER_15_66
timestamp 1586364061
transform 1 0 7176 0 1 10336
box -38 -48 130 592
use scs8hd_fill_2  FILLER_15_69
timestamp 1586364061
transform 1 0 7452 0 1 10336
box -38 -48 222 592
use scs8hd_nor4_4  _56_
timestamp 1586364061
transform 1 0 7820 0 1 10336
box -38 -48 1602 592
use scs8hd_lpflow_inputisolatch_1  mem_top_ipin_0.LATCH_2_.latch
timestamp 1586364061
transform 1 0 10212 0 1 10336
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA__57__C
timestamp 1586364061
transform 1 0 9752 0 1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_15_90
timestamp 1586364061
transform 1 0 9384 0 1 10336
box -38 -48 406 592
use scs8hd_decap_3  FILLER_15_96
timestamp 1586364061
transform 1 0 9936 0 1 10336
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_129
timestamp 1586364061
transform 1 0 12328 0 1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_0.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 11408 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__49__A
timestamp 1586364061
transform 1 0 12144 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_0.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 11776 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_110
timestamp 1586364061
transform 1 0 11224 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_114
timestamp 1586364061
transform 1 0 11592 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_118
timestamp 1586364061
transform 1 0 11960 0 1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_15_123
timestamp 1586364061
transform 1 0 12420 0 1 10336
box -38 -48 406 592
use scs8hd_nor4_4  _49_
timestamp 1586364061
transform 1 0 13064 0 1 10336
box -38 -48 1602 592
use scs8hd_diode_2  ANTENNA__49__C
timestamp 1586364061
transform 1 0 12880 0 1 10336
box -38 -48 222 592
use scs8hd_fill_1  FILLER_15_127
timestamp 1586364061
transform 1 0 12788 0 1 10336
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_2.LATCH_2_.latch
timestamp 1586364061
transform 1 0 15364 0 1 10336
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA__77__A
timestamp 1586364061
transform 1 0 15180 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_2.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 14812 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_147
timestamp 1586364061
transform 1 0 14628 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_151
timestamp 1586364061
transform 1 0 14996 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 17020 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 17388 0 1 10336
box -38 -48 222 592
use scs8hd_decap_6  FILLER_15_166
timestamp 1586364061
transform 1 0 16376 0 1 10336
box -38 -48 590 592
use scs8hd_fill_1  FILLER_15_172
timestamp 1586364061
transform 1 0 16928 0 1 10336
box -38 -48 130 592
use scs8hd_fill_2  FILLER_15_175
timestamp 1586364061
transform 1 0 17204 0 1 10336
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_ipin_2.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18032 0 1 10336
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_130
timestamp 1586364061
transform 1 0 17940 0 1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 19044 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 17756 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_179
timestamp 1586364061
transform 1 0 17572 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_193
timestamp 1586364061
transform 1 0 18860 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 19412 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_197
timestamp 1586364061
transform 1 0 19228 0 1 10336
box -38 -48 222 592
use scs8hd_decap_12  FILLER_15_201
timestamp 1586364061
transform 1 0 19596 0 1 10336
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_15_213
timestamp 1586364061
transform 1 0 20700 0 1 10336
box -38 -48 222 592
use scs8hd_buf_2  _79_
timestamp 1586364061
transform 1 0 20884 0 1 10336
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__79__A
timestamp 1586364061
transform 1 0 21436 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_219
timestamp 1586364061
transform 1 0 21252 0 1 10336
box -38 -48 222 592
use scs8hd_decap_8  FILLER_15_223
timestamp 1586364061
transform 1 0 21620 0 1 10336
box -38 -48 774 592
use scs8hd_fill_2  FILLER_15_231
timestamp 1586364061
transform 1 0 22356 0 1 10336
box -38 -48 222 592
use scs8hd_decap_3  PHY_31
timestamp 1586364061
transform -1 0 22816 0 1 10336
box -38 -48 314 592
use scs8hd_decap_3  PHY_32
timestamp 1586364061
transform 1 0 1104 0 -1 11424
box -38 -48 314 592
use scs8hd_decap_12  FILLER_16_3
timestamp 1586364061
transform 1 0 1380 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_15
timestamp 1586364061
transform 1 0 2484 0 -1 11424
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_131
timestamp 1586364061
transform 1 0 3956 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_4  FILLER_16_27
timestamp 1586364061
transform 1 0 3588 0 -1 11424
box -38 -48 406 592
use scs8hd_decap_12  FILLER_16_32
timestamp 1586364061
transform 1 0 4048 0 -1 11424
box -38 -48 1142 592
use scs8hd_nor4_4  _54_
timestamp 1586364061
transform 1 0 5428 0 -1 11424
box -38 -48 1602 592
use scs8hd_decap_3  FILLER_16_44
timestamp 1586364061
transform 1 0 5152 0 -1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_0.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 7636 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_6  FILLER_16_64
timestamp 1586364061
transform 1 0 6992 0 -1 11424
box -38 -48 590 592
use scs8hd_fill_1  FILLER_16_70
timestamp 1586364061
transform 1 0 7544 0 -1 11424
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  mem_top_ipin_0.LATCH_3_.latch
timestamp 1586364061
transform 1 0 7820 0 -1 11424
box -38 -48 1050 592
use scs8hd_decap_6  FILLER_16_84
timestamp 1586364061
transform 1 0 8832 0 -1 11424
box -38 -48 590 592
use scs8hd_nor4_4  _57_
timestamp 1586364061
transform 1 0 9752 0 -1 11424
box -38 -48 1602 592
use scs8hd_tapvpwrvgnd_1  PHY_132
timestamp 1586364061
transform 1 0 9568 0 -1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__42__A
timestamp 1586364061
transform 1 0 9384 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_1  FILLER_16_93
timestamp 1586364061
transform 1 0 9660 0 -1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__49__D
timestamp 1586364061
transform 1 0 12512 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__47__D
timestamp 1586364061
transform 1 0 12144 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_8  FILLER_16_111
timestamp 1586364061
transform 1 0 11316 0 -1 11424
box -38 -48 774 592
use scs8hd_fill_1  FILLER_16_119
timestamp 1586364061
transform 1 0 12052 0 -1 11424
box -38 -48 130 592
use scs8hd_fill_2  FILLER_16_122
timestamp 1586364061
transform 1 0 12328 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__47__A
timestamp 1586364061
transform 1 0 12880 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__49__B
timestamp 1586364061
transform 1 0 13248 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__48__A
timestamp 1586364061
transform 1 0 13616 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_126
timestamp 1586364061
transform 1 0 12696 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_130
timestamp 1586364061
transform 1 0 13064 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_134
timestamp 1586364061
transform 1 0 13432 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_12  FILLER_16_138
timestamp 1586364061
transform 1 0 13800 0 -1 11424
box -38 -48 1142 592
use scs8hd_buf_2  _77_
timestamp 1586364061
transform 1 0 15272 0 -1 11424
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_133
timestamp 1586364061
transform 1 0 15180 0 -1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_2.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 15824 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_3  FILLER_16_150
timestamp 1586364061
transform 1 0 14904 0 -1 11424
box -38 -48 314 592
use scs8hd_fill_2  FILLER_16_158
timestamp 1586364061
transform 1 0 15640 0 -1 11424
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_ipin_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 17020 0 -1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_2.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 16192 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_162
timestamp 1586364061
transform 1 0 16008 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_6  FILLER_16_166
timestamp 1586364061
transform 1 0 16376 0 -1 11424
box -38 -48 590 592
use scs8hd_fill_1  FILLER_16_172
timestamp 1586364061
transform 1 0 16928 0 -1 11424
box -38 -48 130 592
use scs8hd_ebufn_2  mux_bottom_ipin_2.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18584 0 -1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 18032 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_182
timestamp 1586364061
transform 1 0 17848 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_16_186
timestamp 1586364061
transform 1 0 18216 0 -1 11424
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_134
timestamp 1586364061
transform 1 0 20792 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_12  FILLER_16_199
timestamp 1586364061
transform 1 0 19412 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_16_211
timestamp 1586364061
transform 1 0 20516 0 -1 11424
box -38 -48 314 592
use scs8hd_decap_12  FILLER_16_215
timestamp 1586364061
transform 1 0 20884 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_16_227
timestamp 1586364061
transform 1 0 21988 0 -1 11424
box -38 -48 590 592
use scs8hd_decap_3  PHY_33
timestamp 1586364061
transform -1 0 22816 0 -1 11424
box -38 -48 314 592
use scs8hd_buf_2  _86_
timestamp 1586364061
transform 1 0 1380 0 1 11424
box -38 -48 406 592
use scs8hd_decap_3  PHY_34
timestamp 1586364061
transform 1 0 1104 0 1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__86__A
timestamp 1586364061
transform 1 0 1932 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_7
timestamp 1586364061
transform 1 0 1748 0 1 11424
box -38 -48 222 592
use scs8hd_decap_12  FILLER_17_11
timestamp 1586364061
transform 1 0 2116 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_23
timestamp 1586364061
transform 1 0 3220 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_35
timestamp 1586364061
transform 1 0 4324 0 1 11424
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA__43__A
timestamp 1586364061
transform 1 0 5796 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__43__D
timestamp 1586364061
transform 1 0 5428 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_49
timestamp 1586364061
transform 1 0 5612 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_53
timestamp 1586364061
transform 1 0 5980 0 1 11424
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_135
timestamp 1586364061
transform 1 0 6716 0 1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__43__B
timestamp 1586364061
transform 1 0 6164 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__43__C
timestamp 1586364061
transform 1 0 6532 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__41__C
timestamp 1586364061
transform 1 0 7452 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_57
timestamp 1586364061
transform 1 0 6348 0 1 11424
box -38 -48 222 592
use scs8hd_decap_6  FILLER_17_62
timestamp 1586364061
transform 1 0 6808 0 1 11424
box -38 -48 590 592
use scs8hd_fill_1  FILLER_17_68
timestamp 1586364061
transform 1 0 7360 0 1 11424
box -38 -48 130 592
use scs8hd_fill_2  FILLER_17_71
timestamp 1586364061
transform 1 0 7636 0 1 11424
box -38 -48 222 592
use scs8hd_nor4_4  _41_
timestamp 1586364061
transform 1 0 8004 0 1 11424
box -38 -48 1602 592
use scs8hd_diode_2  ANTENNA__41__B
timestamp 1586364061
transform 1 0 7820 0 1 11424
box -38 -48 222 592
use scs8hd_inv_8  _24_
timestamp 1586364061
transform 1 0 10764 0 1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__42__C
timestamp 1586364061
transform 1 0 10304 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__24__A
timestamp 1586364061
transform 1 0 9936 0 1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_17_92
timestamp 1586364061
transform 1 0 9568 0 1 11424
box -38 -48 406 592
use scs8hd_fill_2  FILLER_17_98
timestamp 1586364061
transform 1 0 10120 0 1 11424
box -38 -48 222 592
use scs8hd_decap_3  FILLER_17_102
timestamp 1586364061
transform 1 0 10488 0 1 11424
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_136
timestamp 1586364061
transform 1 0 12328 0 1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__48__B
timestamp 1586364061
transform 1 0 12144 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__42__B
timestamp 1586364061
transform 1 0 11776 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_114
timestamp 1586364061
transform 1 0 11592 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_118
timestamp 1586364061
transform 1 0 11960 0 1 11424
box -38 -48 222 592
use scs8hd_decap_3  FILLER_17_123
timestamp 1586364061
transform 1 0 12420 0 1 11424
box -38 -48 314 592
use scs8hd_nor4_4  _48_
timestamp 1586364061
transform 1 0 12880 0 1 11424
box -38 -48 1602 592
use scs8hd_diode_2  ANTENNA__47__C
timestamp 1586364061
transform 1 0 12696 0 1 11424
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_2.LATCH_3_.latch
timestamp 1586364061
transform 1 0 15548 0 1 11424
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_2.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 15364 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_2.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 14996 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__47__B
timestamp 1586364061
transform 1 0 14628 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_145
timestamp 1586364061
transform 1 0 14444 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_149
timestamp 1586364061
transform 1 0 14812 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_153
timestamp 1586364061
transform 1 0 15180 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 17204 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_2.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 16744 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_168
timestamp 1586364061
transform 1 0 16560 0 1 11424
box -38 -48 222 592
use scs8hd_decap_3  FILLER_17_172
timestamp 1586364061
transform 1 0 16928 0 1 11424
box -38 -48 314 592
use scs8hd_fill_2  FILLER_17_177
timestamp 1586364061
transform 1 0 17388 0 1 11424
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_137
timestamp 1586364061
transform 1 0 17940 0 1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 18768 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 17572 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_181
timestamp 1586364061
transform 1 0 17756 0 1 11424
box -38 -48 222 592
use scs8hd_decap_8  FILLER_17_184
timestamp 1586364061
transform 1 0 18032 0 1 11424
box -38 -48 774 592
use scs8hd_decap_12  FILLER_17_194
timestamp 1586364061
transform 1 0 18952 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_206
timestamp 1586364061
transform 1 0 20056 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_218
timestamp 1586364061
transform 1 0 21160 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_17_230
timestamp 1586364061
transform 1 0 22264 0 1 11424
box -38 -48 314 592
use scs8hd_decap_3  PHY_35
timestamp 1586364061
transform -1 0 22816 0 1 11424
box -38 -48 314 592
use scs8hd_decap_3  PHY_36
timestamp 1586364061
transform 1 0 1104 0 -1 12512
box -38 -48 314 592
use scs8hd_decap_12  FILLER_18_3
timestamp 1586364061
transform 1 0 1380 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_15
timestamp 1586364061
transform 1 0 2484 0 -1 12512
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_138
timestamp 1586364061
transform 1 0 3956 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_4  FILLER_18_27
timestamp 1586364061
transform 1 0 3588 0 -1 12512
box -38 -48 406 592
use scs8hd_decap_12  FILLER_18_32
timestamp 1586364061
transform 1 0 4048 0 -1 12512
box -38 -48 1142 592
use scs8hd_nor4_4  _43_
timestamp 1586364061
transform 1 0 5796 0 -1 12512
box -38 -48 1602 592
use scs8hd_diode_2  ANTENNA__39__C
timestamp 1586364061
transform 1 0 5520 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_18_44
timestamp 1586364061
transform 1 0 5152 0 -1 12512
box -38 -48 406 592
use scs8hd_fill_1  FILLER_18_50
timestamp 1586364061
transform 1 0 5704 0 -1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__40__D
timestamp 1586364061
transform 1 0 7544 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_68
timestamp 1586364061
transform 1 0 7360 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__41__A
timestamp 1586364061
transform 1 0 8004 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__41__D
timestamp 1586364061
transform 1 0 8372 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_3  FILLER_18_72
timestamp 1586364061
transform 1 0 7728 0 -1 12512
box -38 -48 314 592
use scs8hd_fill_2  FILLER_18_77
timestamp 1586364061
transform 1 0 8188 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_8  FILLER_18_81
timestamp 1586364061
transform 1 0 8556 0 -1 12512
box -38 -48 774 592
use scs8hd_fill_1  FILLER_18_89
timestamp 1586364061
transform 1 0 9292 0 -1 12512
box -38 -48 130 592
use scs8hd_nor4_4  _42_
timestamp 1586364061
transform 1 0 10304 0 -1 12512
box -38 -48 1602 592
use scs8hd_tapvpwrvgnd_1  PHY_139
timestamp 1586364061
transform 1 0 9568 0 -1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__44__A
timestamp 1586364061
transform 1 0 9936 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__42__D
timestamp 1586364061
transform 1 0 9384 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_3  FILLER_18_93
timestamp 1586364061
transform 1 0 9660 0 -1 12512
box -38 -48 314 592
use scs8hd_fill_2  FILLER_18_98
timestamp 1586364061
transform 1 0 10120 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__48__D
timestamp 1586364061
transform 1 0 12328 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_18_117
timestamp 1586364061
transform 1 0 11868 0 -1 12512
box -38 -48 406 592
use scs8hd_fill_1  FILLER_18_121
timestamp 1586364061
transform 1 0 12236 0 -1 12512
box -38 -48 130 592
use scs8hd_fill_2  FILLER_18_124
timestamp 1586364061
transform 1 0 12512 0 -1 12512
box -38 -48 222 592
use scs8hd_nor4_4  _47_
timestamp 1586364061
transform 1 0 12880 0 -1 12512
box -38 -48 1602 592
use scs8hd_diode_2  ANTENNA__48__C
timestamp 1586364061
transform 1 0 12696 0 -1 12512
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_2.LATCH_4_.latch
timestamp 1586364061
transform 1 0 15456 0 -1 12512
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_140
timestamp 1586364061
transform 1 0 15180 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_8  FILLER_18_145
timestamp 1586364061
transform 1 0 14444 0 -1 12512
box -38 -48 774 592
use scs8hd_fill_2  FILLER_18_154
timestamp 1586364061
transform 1 0 15272 0 -1 12512
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_ipin_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 17204 0 -1 12512
box -38 -48 866 592
use scs8hd_decap_8  FILLER_18_167
timestamp 1586364061
transform 1 0 16468 0 -1 12512
box -38 -48 774 592
use scs8hd_inv_1  mux_bottom_ipin_2.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 18768 0 -1 12512
box -38 -48 314 592
use scs8hd_decap_8  FILLER_18_184
timestamp 1586364061
transform 1 0 18032 0 -1 12512
box -38 -48 774 592
use scs8hd_decap_12  FILLER_18_195
timestamp 1586364061
transform 1 0 19044 0 -1 12512
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_141
timestamp 1586364061
transform 1 0 20792 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_6  FILLER_18_207
timestamp 1586364061
transform 1 0 20148 0 -1 12512
box -38 -48 590 592
use scs8hd_fill_1  FILLER_18_213
timestamp 1586364061
transform 1 0 20700 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_12  FILLER_18_215
timestamp 1586364061
transform 1 0 20884 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_18_227
timestamp 1586364061
transform 1 0 21988 0 -1 12512
box -38 -48 590 592
use scs8hd_decap_3  PHY_37
timestamp 1586364061
transform -1 0 22816 0 -1 12512
box -38 -48 314 592
use scs8hd_decap_3  PHY_38
timestamp 1586364061
transform 1 0 1104 0 1 12512
box -38 -48 314 592
use scs8hd_decap_3  PHY_40
timestamp 1586364061
transform 1 0 1104 0 -1 13600
box -38 -48 314 592
use scs8hd_decap_12  FILLER_19_3
timestamp 1586364061
transform 1 0 1380 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_15
timestamp 1586364061
transform 1 0 2484 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_3
timestamp 1586364061
transform 1 0 1380 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_15
timestamp 1586364061
transform 1 0 2484 0 -1 13600
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_145
timestamp 1586364061
transform 1 0 3956 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_12  FILLER_19_27
timestamp 1586364061
transform 1 0 3588 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_20_27
timestamp 1586364061
transform 1 0 3588 0 -1 13600
box -38 -48 406 592
use scs8hd_decap_8  FILLER_20_32
timestamp 1586364061
transform 1 0 4048 0 -1 13600
box -38 -48 774 592
use scs8hd_decap_4  FILLER_20_44
timestamp 1586364061
transform 1 0 5152 0 -1 13600
box -38 -48 406 592
use scs8hd_fill_2  FILLER_20_40
timestamp 1586364061
transform 1 0 4784 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_42
timestamp 1586364061
transform 1 0 4968 0 1 12512
box -38 -48 222 592
use scs8hd_fill_1  FILLER_19_39
timestamp 1586364061
transform 1 0 4692 0 1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_0.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 4968 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__39__D
timestamp 1586364061
transform 1 0 4784 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__39__B
timestamp 1586364061
transform 1 0 5152 0 1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_19_50
timestamp 1586364061
transform 1 0 5704 0 1 12512
box -38 -48 406 592
use scs8hd_fill_2  FILLER_19_46
timestamp 1586364061
transform 1 0 5336 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__39__A
timestamp 1586364061
transform 1 0 5520 0 1 12512
box -38 -48 222 592
use scs8hd_nor4_4  _39_
timestamp 1586364061
transform 1 0 5520 0 -1 13600
box -38 -48 1602 592
use scs8hd_nor4_4  _40_
timestamp 1586364061
transform 1 0 6808 0 1 12512
box -38 -48 1602 592
use scs8hd_tapvpwrvgnd_1  PHY_142
timestamp 1586364061
transform 1 0 6716 0 1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__40__C
timestamp 1586364061
transform 1 0 6532 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__40__A
timestamp 1586364061
transform 1 0 6164 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__40__B
timestamp 1586364061
transform 1 0 7268 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_1  FILLER_19_54
timestamp 1586364061
transform 1 0 6072 0 1 12512
box -38 -48 130 592
use scs8hd_fill_2  FILLER_19_57
timestamp 1586364061
transform 1 0 6348 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_65
timestamp 1586364061
transform 1 0 7084 0 -1 13600
box -38 -48 222 592
use scs8hd_decap_8  FILLER_20_69
timestamp 1586364061
transform 1 0 7452 0 -1 13600
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_0.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 8280 0 -1 13600
box -38 -48 222 592
use scs8hd_decap_8  FILLER_19_79
timestamp 1586364061
transform 1 0 8372 0 1 12512
box -38 -48 774 592
use scs8hd_decap_3  FILLER_19_87
timestamp 1586364061
transform 1 0 9108 0 1 12512
box -38 -48 314 592
use scs8hd_fill_1  FILLER_20_77
timestamp 1586364061
transform 1 0 8188 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_12  FILLER_20_80
timestamp 1586364061
transform 1 0 8464 0 -1 13600
box -38 -48 1142 592
use scs8hd_nor4_4  _44_
timestamp 1586364061
transform 1 0 9936 0 1 12512
box -38 -48 1602 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_0.LATCH_0_.latch
timestamp 1586364061
transform 1 0 10488 0 -1 13600
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_146
timestamp 1586364061
transform 1 0 9568 0 -1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__44__C
timestamp 1586364061
transform 1 0 9752 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__44__B
timestamp 1586364061
transform 1 0 9936 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__44__D
timestamp 1586364061
transform 1 0 9384 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_92
timestamp 1586364061
transform 1 0 9568 0 1 12512
box -38 -48 222 592
use scs8hd_decap_3  FILLER_20_93
timestamp 1586364061
transform 1 0 9660 0 -1 13600
box -38 -48 314 592
use scs8hd_decap_4  FILLER_20_98
timestamp 1586364061
transform 1 0 10120 0 -1 13600
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_143
timestamp 1586364061
transform 1 0 12328 0 1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_0.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 11684 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_0.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 12052 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_113
timestamp 1586364061
transform 1 0 11500 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_117
timestamp 1586364061
transform 1 0 11868 0 1 12512
box -38 -48 222 592
use scs8hd_fill_1  FILLER_19_121
timestamp 1586364061
transform 1 0 12236 0 1 12512
box -38 -48 130 592
use scs8hd_decap_4  FILLER_19_123
timestamp 1586364061
transform 1 0 12420 0 1 12512
box -38 -48 406 592
use scs8hd_decap_12  FILLER_20_113
timestamp 1586364061
transform 1 0 11500 0 -1 13600
box -38 -48 1142 592
use scs8hd_nor4_4  _46_
timestamp 1586364061
transform 1 0 13340 0 1 12512
box -38 -48 1602 592
use scs8hd_diode_2  ANTENNA__46__A
timestamp 1586364061
transform 1 0 13156 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__46__B
timestamp 1586364061
transform 1 0 13340 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__46__C
timestamp 1586364061
transform 1 0 12788 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__46__D
timestamp 1586364061
transform 1 0 13708 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_129
timestamp 1586364061
transform 1 0 12972 0 1 12512
box -38 -48 222 592
use scs8hd_decap_8  FILLER_20_125
timestamp 1586364061
transform 1 0 12604 0 -1 13600
box -38 -48 774 592
use scs8hd_fill_2  FILLER_20_135
timestamp 1586364061
transform 1 0 13524 0 -1 13600
box -38 -48 222 592
use scs8hd_decap_12  FILLER_20_139
timestamp 1586364061
transform 1 0 13892 0 -1 13600
box -38 -48 1142 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_2.LATCH_5_.latch
timestamp 1586364061
transform 1 0 15272 0 -1 13600
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_147
timestamp 1586364061
transform 1 0 15180 0 -1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_2.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 15272 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_2.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 15640 0 1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_19_150
timestamp 1586364061
transform 1 0 14904 0 1 12512
box -38 -48 406 592
use scs8hd_fill_2  FILLER_19_156
timestamp 1586364061
transform 1 0 15456 0 1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_19_160
timestamp 1586364061
transform 1 0 15824 0 1 12512
box -38 -48 406 592
use scs8hd_fill_2  FILLER_20_151
timestamp 1586364061
transform 1 0 14996 0 -1 13600
box -38 -48 222 592
use scs8hd_buf_2  _75_
timestamp 1586364061
transform 1 0 16192 0 1 12512
box -38 -48 406 592
use scs8hd_ebufn_2  mux_bottom_ipin_2.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 17020 0 -1 13600
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__75__A
timestamp 1586364061
transform 1 0 16744 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 17112 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 17480 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_168
timestamp 1586364061
transform 1 0 16560 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_172
timestamp 1586364061
transform 1 0 16928 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_176
timestamp 1586364061
transform 1 0 17296 0 1 12512
box -38 -48 222 592
use scs8hd_decap_8  FILLER_20_165
timestamp 1586364061
transform 1 0 16284 0 -1 13600
box -38 -48 774 592
use scs8hd_conb_1  _68_
timestamp 1586364061
transform 1 0 18032 0 1 12512
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_144
timestamp 1586364061
transform 1 0 17940 0 1 12512
box -38 -48 130 592
use scs8hd_decap_3  FILLER_19_180
timestamp 1586364061
transform 1 0 17664 0 1 12512
box -38 -48 314 592
use scs8hd_decap_12  FILLER_19_187
timestamp 1586364061
transform 1 0 18308 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_182
timestamp 1586364061
transform 1 0 17848 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_194
timestamp 1586364061
transform 1 0 18952 0 -1 13600
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_148
timestamp 1586364061
transform 1 0 20792 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_12  FILLER_19_199
timestamp 1586364061
transform 1 0 19412 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_211
timestamp 1586364061
transform 1 0 20516 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_20_206
timestamp 1586364061
transform 1 0 20056 0 -1 13600
box -38 -48 774 592
use scs8hd_decap_8  FILLER_19_223
timestamp 1586364061
transform 1 0 21620 0 1 12512
box -38 -48 774 592
use scs8hd_fill_2  FILLER_19_231
timestamp 1586364061
transform 1 0 22356 0 1 12512
box -38 -48 222 592
use scs8hd_decap_12  FILLER_20_215
timestamp 1586364061
transform 1 0 20884 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_20_227
timestamp 1586364061
transform 1 0 21988 0 -1 13600
box -38 -48 590 592
use scs8hd_decap_3  PHY_39
timestamp 1586364061
transform -1 0 22816 0 1 12512
box -38 -48 314 592
use scs8hd_decap_3  PHY_41
timestamp 1586364061
transform -1 0 22816 0 -1 13600
box -38 -48 314 592
use scs8hd_buf_2  _89_
timestamp 1586364061
transform 1 0 1380 0 1 13600
box -38 -48 406 592
use scs8hd_decap_3  PHY_42
timestamp 1586364061
transform 1 0 1104 0 1 13600
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__89__A
timestamp 1586364061
transform 1 0 1932 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_7
timestamp 1586364061
transform 1 0 1748 0 1 13600
box -38 -48 222 592
use scs8hd_decap_12  FILLER_21_11
timestamp 1586364061
transform 1 0 2116 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_21_23
timestamp 1586364061
transform 1 0 3220 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_21_35
timestamp 1586364061
transform 1 0 4324 0 1 13600
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_0.LATCH_5_.latch
timestamp 1586364061
transform 1 0 4968 0 1 13600
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_0.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 4784 0 1 13600
box -38 -48 222 592
use scs8hd_fill_1  FILLER_21_39
timestamp 1586364061
transform 1 0 4692 0 1 13600
box -38 -48 130 592
use scs8hd_fill_2  FILLER_21_53
timestamp 1586364061
transform 1 0 5980 0 1 13600
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_149
timestamp 1586364061
transform 1 0 6716 0 1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_0.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 7452 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 6164 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_0.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 7084 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 6532 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_57
timestamp 1586364061
transform 1 0 6348 0 1 13600
box -38 -48 222 592
use scs8hd_decap_3  FILLER_21_62
timestamp 1586364061
transform 1 0 6808 0 1 13600
box -38 -48 314 592
use scs8hd_fill_2  FILLER_21_67
timestamp 1586364061
transform 1 0 7268 0 1 13600
box -38 -48 222 592
use scs8hd_decap_4  FILLER_21_71
timestamp 1586364061
transform 1 0 7636 0 1 13600
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_0.LATCH_3_.latch
timestamp 1586364061
transform 1 0 8280 0 1 13600
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_0.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 8096 0 1 13600
box -38 -48 222 592
use scs8hd_fill_1  FILLER_21_75
timestamp 1586364061
transform 1 0 8004 0 1 13600
box -38 -48 130 592
use scs8hd_decap_8  FILLER_21_89
timestamp 1586364061
transform 1 0 9292 0 1 13600
box -38 -48 774 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_0.LATCH_2_.latch
timestamp 1586364061
transform 1 0 10580 0 1 13600
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 10028 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_0.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 10396 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_99
timestamp 1586364061
transform 1 0 10212 0 1 13600
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_150
timestamp 1586364061
transform 1 0 12328 0 1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 11776 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 12144 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_114
timestamp 1586364061
transform 1 0 11592 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_118
timestamp 1586364061
transform 1 0 11960 0 1 13600
box -38 -48 222 592
use scs8hd_decap_12  FILLER_21_123
timestamp 1586364061
transform 1 0 12420 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_21_135
timestamp 1586364061
transform 1 0 13524 0 1 13600
box -38 -48 1142 592
use scs8hd_inv_8  _34_
timestamp 1586364061
transform 1 0 15640 0 1 13600
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__34__A
timestamp 1586364061
transform 1 0 15456 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 15088 0 1 13600
box -38 -48 222 592
use scs8hd_decap_4  FILLER_21_147
timestamp 1586364061
transform 1 0 14628 0 1 13600
box -38 -48 406 592
use scs8hd_fill_1  FILLER_21_151
timestamp 1586364061
transform 1 0 14996 0 1 13600
box -38 -48 130 592
use scs8hd_fill_2  FILLER_21_154
timestamp 1586364061
transform 1 0 15272 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 16652 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_167
timestamp 1586364061
transform 1 0 16468 0 1 13600
box -38 -48 222 592
use scs8hd_decap_12  FILLER_21_171
timestamp 1586364061
transform 1 0 16836 0 1 13600
box -38 -48 1142 592
use scs8hd_inv_1  mux_bottom_ipin_2.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 18032 0 1 13600
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_151
timestamp 1586364061
transform 1 0 17940 0 1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 18492 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_187
timestamp 1586364061
transform 1 0 18308 0 1 13600
box -38 -48 222 592
use scs8hd_decap_12  FILLER_21_191
timestamp 1586364061
transform 1 0 18676 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_21_203
timestamp 1586364061
transform 1 0 19780 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_21_215
timestamp 1586364061
transform 1 0 20884 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_21_227
timestamp 1586364061
transform 1 0 21988 0 1 13600
box -38 -48 590 592
use scs8hd_decap_3  PHY_43
timestamp 1586364061
transform -1 0 22816 0 1 13600
box -38 -48 314 592
use scs8hd_decap_3  PHY_44
timestamp 1586364061
transform 1 0 1104 0 -1 14688
box -38 -48 314 592
use scs8hd_decap_12  FILLER_22_3
timestamp 1586364061
transform 1 0 1380 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_15
timestamp 1586364061
transform 1 0 2484 0 -1 14688
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_152
timestamp 1586364061
transform 1 0 3956 0 -1 14688
box -38 -48 130 592
use scs8hd_decap_4  FILLER_22_27
timestamp 1586364061
transform 1 0 3588 0 -1 14688
box -38 -48 406 592
use scs8hd_decap_12  FILLER_22_32
timestamp 1586364061
transform 1 0 4048 0 -1 14688
box -38 -48 1142 592
use scs8hd_ebufn_2  mux_bottom_ipin_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 5520 0 -1 14688
box -38 -48 866 592
use scs8hd_decap_4  FILLER_22_44
timestamp 1586364061
transform 1 0 5152 0 -1 14688
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_0.LATCH_4_.latch
timestamp 1586364061
transform 1 0 7452 0 -1 14688
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_0.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 6808 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_22_57
timestamp 1586364061
transform 1 0 6348 0 -1 14688
box -38 -48 406 592
use scs8hd_fill_1  FILLER_22_61
timestamp 1586364061
transform 1 0 6716 0 -1 14688
box -38 -48 130 592
use scs8hd_decap_4  FILLER_22_64
timestamp 1586364061
transform 1 0 6992 0 -1 14688
box -38 -48 406 592
use scs8hd_fill_1  FILLER_22_68
timestamp 1586364061
transform 1 0 7360 0 -1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 8648 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9016 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_80
timestamp 1586364061
transform 1 0 8464 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_84
timestamp 1586364061
transform 1 0 8832 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_22_88
timestamp 1586364061
transform 1 0 9200 0 -1 14688
box -38 -48 406 592
use scs8hd_inv_1  mux_bottom_ipin_0.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 10028 0 -1 14688
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_153
timestamp 1586364061
transform 1 0 9568 0 -1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_0.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 10580 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_22_93
timestamp 1586364061
transform 1 0 9660 0 -1 14688
box -38 -48 406 592
use scs8hd_decap_3  FILLER_22_100
timestamp 1586364061
transform 1 0 10304 0 -1 14688
box -38 -48 314 592
use scs8hd_decap_3  FILLER_22_105
timestamp 1586364061
transform 1 0 10764 0 -1 14688
box -38 -48 314 592
use scs8hd_ebufn_2  mux_bottom_ipin_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 11040 0 -1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 12052 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 12420 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_117
timestamp 1586364061
transform 1 0 11868 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_121
timestamp 1586364061
transform 1 0 12236 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_12  FILLER_22_125
timestamp 1586364061
transform 1 0 12604 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_137
timestamp 1586364061
transform 1 0 13708 0 -1 14688
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_154
timestamp 1586364061
transform 1 0 15180 0 -1 14688
box -38 -48 130 592
use scs8hd_decap_4  FILLER_22_149
timestamp 1586364061
transform 1 0 14812 0 -1 14688
box -38 -48 406 592
use scs8hd_decap_6  FILLER_22_154
timestamp 1586364061
transform 1 0 15272 0 -1 14688
box -38 -48 590 592
use scs8hd_fill_1  FILLER_22_160
timestamp 1586364061
transform 1 0 15824 0 -1 14688
box -38 -48 130 592
use scs8hd_ebufn_2  mux_top_ipin_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15916 0 -1 14688
box -38 -48 866 592
use scs8hd_decap_12  FILLER_22_170
timestamp 1586364061
transform 1 0 16744 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_182
timestamp 1586364061
transform 1 0 17848 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_194
timestamp 1586364061
transform 1 0 18952 0 -1 14688
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_155
timestamp 1586364061
transform 1 0 20792 0 -1 14688
box -38 -48 130 592
use scs8hd_decap_8  FILLER_22_206
timestamp 1586364061
transform 1 0 20056 0 -1 14688
box -38 -48 774 592
use scs8hd_decap_12  FILLER_22_215
timestamp 1586364061
transform 1 0 20884 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_22_227
timestamp 1586364061
transform 1 0 21988 0 -1 14688
box -38 -48 590 592
use scs8hd_decap_3  PHY_45
timestamp 1586364061
transform -1 0 22816 0 -1 14688
box -38 -48 314 592
use scs8hd_decap_3  PHY_46
timestamp 1586364061
transform 1 0 1104 0 1 14688
box -38 -48 314 592
use scs8hd_decap_12  FILLER_23_3
timestamp 1586364061
transform 1 0 1380 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_15
timestamp 1586364061
transform 1 0 2484 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_27
timestamp 1586364061
transform 1 0 3588 0 1 14688
box -38 -48 1142 592
use scs8hd_conb_1  _66_
timestamp 1586364061
transform 1 0 5520 0 1 14688
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 5152 0 1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_23_39
timestamp 1586364061
transform 1 0 4692 0 1 14688
box -38 -48 406 592
use scs8hd_fill_1  FILLER_23_43
timestamp 1586364061
transform 1 0 5060 0 1 14688
box -38 -48 130 592
use scs8hd_fill_2  FILLER_23_46
timestamp 1586364061
transform 1 0 5336 0 1 14688
box -38 -48 222 592
use scs8hd_decap_8  FILLER_23_51
timestamp 1586364061
transform 1 0 5796 0 1 14688
box -38 -48 774 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_0.LATCH_1_.latch
timestamp 1586364061
transform 1 0 6808 0 1 14688
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_156
timestamp 1586364061
transform 1 0 6716 0 1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_0.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 6532 0 1 14688
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_ipin_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 8740 0 1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 8004 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 8556 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_73
timestamp 1586364061
transform 1 0 7820 0 1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_23_77
timestamp 1586364061
transform 1 0 8188 0 1 14688
box -38 -48 406 592
use scs8hd_ebufn_2  mux_bottom_ipin_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10764 0 1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10580 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 9752 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10120 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_92
timestamp 1586364061
transform 1 0 9568 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_96
timestamp 1586364061
transform 1 0 9936 0 1 14688
box -38 -48 222 592
use scs8hd_decap_3  FILLER_23_100
timestamp 1586364061
transform 1 0 10304 0 1 14688
box -38 -48 314 592
use scs8hd_ebufn_2  mux_bottom_ipin_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12420 0 1 14688
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_157
timestamp 1586364061
transform 1 0 12328 0 1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 12144 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 11776 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_114
timestamp 1586364061
transform 1 0 11592 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_118
timestamp 1586364061
transform 1 0 11960 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 13432 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_132
timestamp 1586364061
transform 1 0 13248 0 1 14688
box -38 -48 222 592
use scs8hd_decap_12  FILLER_23_136
timestamp 1586364061
transform 1 0 13616 0 1 14688
box -38 -48 1142 592
use scs8hd_inv_1  mux_top_ipin_1.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 14904 0 1 14688
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_1.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 15548 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_1.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 14720 0 1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_23_153
timestamp 1586364061
transform 1 0 15180 0 1 14688
box -38 -48 406 592
use scs8hd_fill_2  FILLER_23_159
timestamp 1586364061
transform 1 0 15732 0 1 14688
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_ipin_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15916 0 1 14688
box -38 -48 866 592
use scs8hd_decap_12  FILLER_23_170
timestamp 1586364061
transform 1 0 16744 0 1 14688
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_158
timestamp 1586364061
transform 1 0 17940 0 1 14688
box -38 -48 130 592
use scs8hd_fill_1  FILLER_23_182
timestamp 1586364061
transform 1 0 17848 0 1 14688
box -38 -48 130 592
use scs8hd_decap_12  FILLER_23_184
timestamp 1586364061
transform 1 0 18032 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_196
timestamp 1586364061
transform 1 0 19136 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_23_208
timestamp 1586364061
transform 1 0 20240 0 1 14688
box -38 -48 590 592
use scs8hd_fill_1  FILLER_23_214
timestamp 1586364061
transform 1 0 20792 0 1 14688
box -38 -48 130 592
use scs8hd_buf_2  _74_
timestamp 1586364061
transform 1 0 20884 0 1 14688
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__74__A
timestamp 1586364061
transform 1 0 21436 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_219
timestamp 1586364061
transform 1 0 21252 0 1 14688
box -38 -48 222 592
use scs8hd_decap_8  FILLER_23_223
timestamp 1586364061
transform 1 0 21620 0 1 14688
box -38 -48 774 592
use scs8hd_fill_2  FILLER_23_231
timestamp 1586364061
transform 1 0 22356 0 1 14688
box -38 -48 222 592
use scs8hd_decap_3  PHY_47
timestamp 1586364061
transform -1 0 22816 0 1 14688
box -38 -48 314 592
use scs8hd_decap_3  PHY_48
timestamp 1586364061
transform 1 0 1104 0 -1 15776
box -38 -48 314 592
use scs8hd_decap_12  FILLER_24_3
timestamp 1586364061
transform 1 0 1380 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_15
timestamp 1586364061
transform 1 0 2484 0 -1 15776
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_159
timestamp 1586364061
transform 1 0 3956 0 -1 15776
box -38 -48 130 592
use scs8hd_decap_4  FILLER_24_27
timestamp 1586364061
transform 1 0 3588 0 -1 15776
box -38 -48 406 592
use scs8hd_decap_12  FILLER_24_32
timestamp 1586364061
transform 1 0 4048 0 -1 15776
box -38 -48 1142 592
use scs8hd_inv_1  mux_bottom_ipin_0.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 5152 0 -1 15776
box -38 -48 314 592
use scs8hd_decap_12  FILLER_24_47
timestamp 1586364061
transform 1 0 5428 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_59
timestamp 1586364061
transform 1 0 6532 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_24_71
timestamp 1586364061
transform 1 0 7636 0 -1 15776
box -38 -48 406 592
use scs8hd_ebufn_2  mux_bottom_ipin_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 8004 0 -1 15776
box -38 -48 866 592
use scs8hd_decap_8  FILLER_24_84
timestamp 1586364061
transform 1 0 8832 0 -1 15776
box -38 -48 774 592
use scs8hd_ebufn_2  mux_bottom_ipin_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9660 0 -1 15776
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_160
timestamp 1586364061
transform 1 0 9568 0 -1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10764 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_3  FILLER_24_102
timestamp 1586364061
transform 1 0 10488 0 -1 15776
box -38 -48 314 592
use scs8hd_decap_3  FILLER_24_107
timestamp 1586364061
transform 1 0 10948 0 -1 15776
box -38 -48 314 592
use scs8hd_ebufn_2  mux_bottom_ipin_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 11224 0 -1 15776
box -38 -48 866 592
use scs8hd_decap_8  FILLER_24_119
timestamp 1586364061
transform 1 0 12052 0 -1 15776
box -38 -48 774 592
use scs8hd_inv_1  mux_bottom_ipin_0.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 12788 0 -1 15776
box -38 -48 314 592
use scs8hd_decap_12  FILLER_24_130
timestamp 1586364061
transform 1 0 13064 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_24_142
timestamp 1586364061
transform 1 0 14168 0 -1 15776
box -38 -48 774 592
use scs8hd_inv_1  mux_top_ipin_1.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 15548 0 -1 15776
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_161
timestamp 1586364061
transform 1 0 15180 0 -1 15776
box -38 -48 130 592
use scs8hd_decap_3  FILLER_24_150
timestamp 1586364061
transform 1 0 14904 0 -1 15776
box -38 -48 314 592
use scs8hd_decap_3  FILLER_24_154
timestamp 1586364061
transform 1 0 15272 0 -1 15776
box -38 -48 314 592
use scs8hd_fill_2  FILLER_24_160
timestamp 1586364061
transform 1 0 15824 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 16008 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 16376 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_164
timestamp 1586364061
transform 1 0 16192 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_12  FILLER_24_168
timestamp 1586364061
transform 1 0 16560 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_180
timestamp 1586364061
transform 1 0 17664 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_192
timestamp 1586364061
transform 1 0 18768 0 -1 15776
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_162
timestamp 1586364061
transform 1 0 20792 0 -1 15776
box -38 -48 130 592
use scs8hd_decap_8  FILLER_24_204
timestamp 1586364061
transform 1 0 19872 0 -1 15776
box -38 -48 774 592
use scs8hd_fill_2  FILLER_24_212
timestamp 1586364061
transform 1 0 20608 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_12  FILLER_24_215
timestamp 1586364061
transform 1 0 20884 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_24_227
timestamp 1586364061
transform 1 0 21988 0 -1 15776
box -38 -48 590 592
use scs8hd_decap_3  PHY_49
timestamp 1586364061
transform -1 0 22816 0 -1 15776
box -38 -48 314 592
use scs8hd_decap_3  PHY_50
timestamp 1586364061
transform 1 0 1104 0 1 15776
box -38 -48 314 592
use scs8hd_decap_12  FILLER_25_3
timestamp 1586364061
transform 1 0 1380 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_15
timestamp 1586364061
transform 1 0 2484 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_27
timestamp 1586364061
transform 1 0 3588 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_39
timestamp 1586364061
transform 1 0 4692 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_25_51
timestamp 1586364061
transform 1 0 5796 0 1 15776
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_163
timestamp 1586364061
transform 1 0 6716 0 1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 7636 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 7268 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_59
timestamp 1586364061
transform 1 0 6532 0 1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_25_62
timestamp 1586364061
transform 1 0 6808 0 1 15776
box -38 -48 406 592
use scs8hd_fill_1  FILLER_25_66
timestamp 1586364061
transform 1 0 7176 0 1 15776
box -38 -48 130 592
use scs8hd_fill_2  FILLER_25_69
timestamp 1586364061
transform 1 0 7452 0 1 15776
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_ipin_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 7912 0 1 15776
box -38 -48 866 592
use scs8hd_fill_1  FILLER_25_73
timestamp 1586364061
transform 1 0 7820 0 1 15776
box -38 -48 130 592
use scs8hd_decap_12  FILLER_25_83
timestamp 1586364061
transform 1 0 8740 0 1 15776
box -38 -48 1142 592
use scs8hd_inv_1  mux_bottom_ipin_0.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 10948 0 1 15776
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 10672 0 1 15776
box -38 -48 222 592
use scs8hd_decap_8  FILLER_25_95
timestamp 1586364061
transform 1 0 9844 0 1 15776
box -38 -48 774 592
use scs8hd_fill_1  FILLER_25_103
timestamp 1586364061
transform 1 0 10580 0 1 15776
box -38 -48 130 592
use scs8hd_fill_1  FILLER_25_106
timestamp 1586364061
transform 1 0 10856 0 1 15776
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_164
timestamp 1586364061
transform 1 0 12328 0 1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 11408 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_110
timestamp 1586364061
transform 1 0 11224 0 1 15776
box -38 -48 222 592
use scs8hd_decap_8  FILLER_25_114
timestamp 1586364061
transform 1 0 11592 0 1 15776
box -38 -48 774 592
use scs8hd_decap_12  FILLER_25_123
timestamp 1586364061
transform 1 0 12420 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_135
timestamp 1586364061
transform 1 0 13524 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_147
timestamp 1586364061
transform 1 0 14628 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_159
timestamp 1586364061
transform 1 0 15732 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_171
timestamp 1586364061
transform 1 0 16836 0 1 15776
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_165
timestamp 1586364061
transform 1 0 17940 0 1 15776
box -38 -48 130 592
use scs8hd_decap_12  FILLER_25_184
timestamp 1586364061
transform 1 0 18032 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_196
timestamp 1586364061
transform 1 0 19136 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_208
timestamp 1586364061
transform 1 0 20240 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_220
timestamp 1586364061
transform 1 0 21344 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_3  PHY_51
timestamp 1586364061
transform -1 0 22816 0 1 15776
box -38 -48 314 592
use scs8hd_fill_1  FILLER_25_232
timestamp 1586364061
transform 1 0 22448 0 1 15776
box -38 -48 130 592
use scs8hd_decap_3  PHY_52
timestamp 1586364061
transform 1 0 1104 0 -1 16864
box -38 -48 314 592
use scs8hd_decap_3  PHY_54
timestamp 1586364061
transform 1 0 1104 0 1 16864
box -38 -48 314 592
use scs8hd_decap_12  FILLER_26_3
timestamp 1586364061
transform 1 0 1380 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_26_15
timestamp 1586364061
transform 1 0 2484 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_3
timestamp 1586364061
transform 1 0 1380 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_15
timestamp 1586364061
transform 1 0 2484 0 1 16864
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_166
timestamp 1586364061
transform 1 0 3956 0 -1 16864
box -38 -48 130 592
use scs8hd_decap_4  FILLER_26_27
timestamp 1586364061
transform 1 0 3588 0 -1 16864
box -38 -48 406 592
use scs8hd_decap_12  FILLER_26_32
timestamp 1586364061
transform 1 0 4048 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_27
timestamp 1586364061
transform 1 0 3588 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_26_44
timestamp 1586364061
transform 1 0 5152 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_39
timestamp 1586364061
transform 1 0 4692 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_27_51
timestamp 1586364061
transform 1 0 5796 0 1 16864
box -38 -48 774 592
use scs8hd_buf_2  _80_
timestamp 1586364061
transform 1 0 6808 0 1 16864
box -38 -48 406 592
use scs8hd_inv_1  mux_bottom_ipin_0.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 7636 0 -1 16864
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_170
timestamp 1586364061
transform 1 0 6716 0 1 16864
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__80__A
timestamp 1586364061
transform 1 0 7360 0 1 16864
box -38 -48 222 592
use scs8hd_decap_12  FILLER_26_56
timestamp 1586364061
transform 1 0 6256 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_26_68
timestamp 1586364061
transform 1 0 7360 0 -1 16864
box -38 -48 314 592
use scs8hd_fill_2  FILLER_27_59
timestamp 1586364061
transform 1 0 6532 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_66
timestamp 1586364061
transform 1 0 7176 0 1 16864
box -38 -48 222 592
use scs8hd_decap_4  FILLER_27_70
timestamp 1586364061
transform 1 0 7544 0 1 16864
box -38 -48 406 592
use scs8hd_inv_1  mux_bottom_ipin_0.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 7912 0 1 16864
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 8372 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 8096 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_74
timestamp 1586364061
transform 1 0 7912 0 -1 16864
box -38 -48 222 592
use scs8hd_decap_12  FILLER_26_78
timestamp 1586364061
transform 1 0 8280 0 -1 16864
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_27_77
timestamp 1586364061
transform 1 0 8188 0 1 16864
box -38 -48 222 592
use scs8hd_decap_12  FILLER_27_81
timestamp 1586364061
transform 1 0 8556 0 1 16864
box -38 -48 1142 592
use scs8hd_inv_1  mux_bottom_ipin_0.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 10672 0 -1 16864
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_167
timestamp 1586364061
transform 1 0 9568 0 -1 16864
box -38 -48 130 592
use scs8hd_fill_2  FILLER_26_90
timestamp 1586364061
transform 1 0 9384 0 -1 16864
box -38 -48 222 592
use scs8hd_decap_8  FILLER_26_93
timestamp 1586364061
transform 1 0 9660 0 -1 16864
box -38 -48 774 592
use scs8hd_decap_3  FILLER_26_101
timestamp 1586364061
transform 1 0 10396 0 -1 16864
box -38 -48 314 592
use scs8hd_decap_12  FILLER_26_107
timestamp 1586364061
transform 1 0 10948 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_93
timestamp 1586364061
transform 1 0 9660 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_105
timestamp 1586364061
transform 1 0 10764 0 1 16864
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_171
timestamp 1586364061
transform 1 0 12328 0 1 16864
box -38 -48 130 592
use scs8hd_decap_12  FILLER_26_119
timestamp 1586364061
transform 1 0 12052 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_27_117
timestamp 1586364061
transform 1 0 11868 0 1 16864
box -38 -48 406 592
use scs8hd_fill_1  FILLER_27_121
timestamp 1586364061
transform 1 0 12236 0 1 16864
box -38 -48 130 592
use scs8hd_decap_12  FILLER_27_123
timestamp 1586364061
transform 1 0 12420 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_26_131
timestamp 1586364061
transform 1 0 13156 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_135
timestamp 1586364061
transform 1 0 13524 0 1 16864
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_168
timestamp 1586364061
transform 1 0 15180 0 -1 16864
box -38 -48 130 592
use scs8hd_decap_8  FILLER_26_143
timestamp 1586364061
transform 1 0 14260 0 -1 16864
box -38 -48 774 592
use scs8hd_fill_2  FILLER_26_151
timestamp 1586364061
transform 1 0 14996 0 -1 16864
box -38 -48 222 592
use scs8hd_decap_12  FILLER_26_154
timestamp 1586364061
transform 1 0 15272 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_147
timestamp 1586364061
transform 1 0 14628 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_159
timestamp 1586364061
transform 1 0 15732 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_26_166
timestamp 1586364061
transform 1 0 16376 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_26_178
timestamp 1586364061
transform 1 0 17480 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_171
timestamp 1586364061
transform 1 0 16836 0 1 16864
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_172
timestamp 1586364061
transform 1 0 17940 0 1 16864
box -38 -48 130 592
use scs8hd_decap_12  FILLER_26_190
timestamp 1586364061
transform 1 0 18584 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_184
timestamp 1586364061
transform 1 0 18032 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_196
timestamp 1586364061
transform 1 0 19136 0 1 16864
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_169
timestamp 1586364061
transform 1 0 20792 0 -1 16864
box -38 -48 130 592
use scs8hd_decap_12  FILLER_26_202
timestamp 1586364061
transform 1 0 19688 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_208
timestamp 1586364061
transform 1 0 20240 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_26_215
timestamp 1586364061
transform 1 0 20884 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_26_227
timestamp 1586364061
transform 1 0 21988 0 -1 16864
box -38 -48 590 592
use scs8hd_decap_12  FILLER_27_220
timestamp 1586364061
transform 1 0 21344 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_3  PHY_53
timestamp 1586364061
transform -1 0 22816 0 -1 16864
box -38 -48 314 592
use scs8hd_decap_3  PHY_55
timestamp 1586364061
transform -1 0 22816 0 1 16864
box -38 -48 314 592
use scs8hd_fill_1  FILLER_27_232
timestamp 1586364061
transform 1 0 22448 0 1 16864
box -38 -48 130 592
use scs8hd_decap_3  PHY_56
timestamp 1586364061
transform 1 0 1104 0 -1 17952
box -38 -48 314 592
use scs8hd_decap_12  FILLER_28_3
timestamp 1586364061
transform 1 0 1380 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_15
timestamp 1586364061
transform 1 0 2484 0 -1 17952
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_173
timestamp 1586364061
transform 1 0 3956 0 -1 17952
box -38 -48 130 592
use scs8hd_decap_4  FILLER_28_27
timestamp 1586364061
transform 1 0 3588 0 -1 17952
box -38 -48 406 592
use scs8hd_decap_12  FILLER_28_32
timestamp 1586364061
transform 1 0 4048 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_44
timestamp 1586364061
transform 1 0 5152 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_56
timestamp 1586364061
transform 1 0 6256 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_68
timestamp 1586364061
transform 1 0 7360 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_80
timestamp 1586364061
transform 1 0 8464 0 -1 17952
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_174
timestamp 1586364061
transform 1 0 9568 0 -1 17952
box -38 -48 130 592
use scs8hd_decap_12  FILLER_28_93
timestamp 1586364061
transform 1 0 9660 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_105
timestamp 1586364061
transform 1 0 10764 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_117
timestamp 1586364061
transform 1 0 11868 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_129
timestamp 1586364061
transform 1 0 12972 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_141
timestamp 1586364061
transform 1 0 14076 0 -1 17952
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_175
timestamp 1586364061
transform 1 0 15180 0 -1 17952
box -38 -48 130 592
use scs8hd_decap_12  FILLER_28_154
timestamp 1586364061
transform 1 0 15272 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_166
timestamp 1586364061
transform 1 0 16376 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_178
timestamp 1586364061
transform 1 0 17480 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_190
timestamp 1586364061
transform 1 0 18584 0 -1 17952
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_176
timestamp 1586364061
transform 1 0 20792 0 -1 17952
box -38 -48 130 592
use scs8hd_decap_12  FILLER_28_202
timestamp 1586364061
transform 1 0 19688 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_215
timestamp 1586364061
transform 1 0 20884 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_28_227
timestamp 1586364061
transform 1 0 21988 0 -1 17952
box -38 -48 590 592
use scs8hd_decap_3  PHY_57
timestamp 1586364061
transform -1 0 22816 0 -1 17952
box -38 -48 314 592
use scs8hd_decap_3  PHY_58
timestamp 1586364061
transform 1 0 1104 0 1 17952
box -38 -48 314 592
use scs8hd_decap_12  FILLER_29_3
timestamp 1586364061
transform 1 0 1380 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_15
timestamp 1586364061
transform 1 0 2484 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_27
timestamp 1586364061
transform 1 0 3588 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_39
timestamp 1586364061
transform 1 0 4692 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_29_51
timestamp 1586364061
transform 1 0 5796 0 1 17952
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_177
timestamp 1586364061
transform 1 0 6716 0 1 17952
box -38 -48 130 592
use scs8hd_fill_2  FILLER_29_59
timestamp 1586364061
transform 1 0 6532 0 1 17952
box -38 -48 222 592
use scs8hd_decap_12  FILLER_29_62
timestamp 1586364061
transform 1 0 6808 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_74
timestamp 1586364061
transform 1 0 7912 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_86
timestamp 1586364061
transform 1 0 9016 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_98
timestamp 1586364061
transform 1 0 10120 0 1 17952
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_178
timestamp 1586364061
transform 1 0 12328 0 1 17952
box -38 -48 130 592
use scs8hd_decap_12  FILLER_29_110
timestamp 1586364061
transform 1 0 11224 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_123
timestamp 1586364061
transform 1 0 12420 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_135
timestamp 1586364061
transform 1 0 13524 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_147
timestamp 1586364061
transform 1 0 14628 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_159
timestamp 1586364061
transform 1 0 15732 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_171
timestamp 1586364061
transform 1 0 16836 0 1 17952
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_179
timestamp 1586364061
transform 1 0 17940 0 1 17952
box -38 -48 130 592
use scs8hd_decap_12  FILLER_29_184
timestamp 1586364061
transform 1 0 18032 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_196
timestamp 1586364061
transform 1 0 19136 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_208
timestamp 1586364061
transform 1 0 20240 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_220
timestamp 1586364061
transform 1 0 21344 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_3  PHY_59
timestamp 1586364061
transform -1 0 22816 0 1 17952
box -38 -48 314 592
use scs8hd_fill_1  FILLER_29_232
timestamp 1586364061
transform 1 0 22448 0 1 17952
box -38 -48 130 592
use scs8hd_decap_3  PHY_60
timestamp 1586364061
transform 1 0 1104 0 -1 19040
box -38 -48 314 592
use scs8hd_decap_12  FILLER_30_3
timestamp 1586364061
transform 1 0 1380 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_15
timestamp 1586364061
transform 1 0 2484 0 -1 19040
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_180
timestamp 1586364061
transform 1 0 3956 0 -1 19040
box -38 -48 130 592
use scs8hd_decap_4  FILLER_30_27
timestamp 1586364061
transform 1 0 3588 0 -1 19040
box -38 -48 406 592
use scs8hd_decap_12  FILLER_30_32
timestamp 1586364061
transform 1 0 4048 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_44
timestamp 1586364061
transform 1 0 5152 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_56
timestamp 1586364061
transform 1 0 6256 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_68
timestamp 1586364061
transform 1 0 7360 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_80
timestamp 1586364061
transform 1 0 8464 0 -1 19040
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_181
timestamp 1586364061
transform 1 0 9568 0 -1 19040
box -38 -48 130 592
use scs8hd_decap_12  FILLER_30_93
timestamp 1586364061
transform 1 0 9660 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_105
timestamp 1586364061
transform 1 0 10764 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_117
timestamp 1586364061
transform 1 0 11868 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_129
timestamp 1586364061
transform 1 0 12972 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_141
timestamp 1586364061
transform 1 0 14076 0 -1 19040
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_182
timestamp 1586364061
transform 1 0 15180 0 -1 19040
box -38 -48 130 592
use scs8hd_decap_12  FILLER_30_154
timestamp 1586364061
transform 1 0 15272 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_166
timestamp 1586364061
transform 1 0 16376 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_178
timestamp 1586364061
transform 1 0 17480 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_190
timestamp 1586364061
transform 1 0 18584 0 -1 19040
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_183
timestamp 1586364061
transform 1 0 20792 0 -1 19040
box -38 -48 130 592
use scs8hd_decap_12  FILLER_30_202
timestamp 1586364061
transform 1 0 19688 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_215
timestamp 1586364061
transform 1 0 20884 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_30_227
timestamp 1586364061
transform 1 0 21988 0 -1 19040
box -38 -48 590 592
use scs8hd_decap_3  PHY_61
timestamp 1586364061
transform -1 0 22816 0 -1 19040
box -38 -48 314 592
use scs8hd_decap_3  PHY_62
timestamp 1586364061
transform 1 0 1104 0 1 19040
box -38 -48 314 592
use scs8hd_decap_12  FILLER_31_3
timestamp 1586364061
transform 1 0 1380 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_15
timestamp 1586364061
transform 1 0 2484 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_27
timestamp 1586364061
transform 1 0 3588 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_39
timestamp 1586364061
transform 1 0 4692 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_31_51
timestamp 1586364061
transform 1 0 5796 0 1 19040
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_184
timestamp 1586364061
transform 1 0 6716 0 1 19040
box -38 -48 130 592
use scs8hd_fill_2  FILLER_31_59
timestamp 1586364061
transform 1 0 6532 0 1 19040
box -38 -48 222 592
use scs8hd_decap_12  FILLER_31_62
timestamp 1586364061
transform 1 0 6808 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_74
timestamp 1586364061
transform 1 0 7912 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_86
timestamp 1586364061
transform 1 0 9016 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_98
timestamp 1586364061
transform 1 0 10120 0 1 19040
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_185
timestamp 1586364061
transform 1 0 12328 0 1 19040
box -38 -48 130 592
use scs8hd_decap_12  FILLER_31_110
timestamp 1586364061
transform 1 0 11224 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_123
timestamp 1586364061
transform 1 0 12420 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_135
timestamp 1586364061
transform 1 0 13524 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_147
timestamp 1586364061
transform 1 0 14628 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_159
timestamp 1586364061
transform 1 0 15732 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_171
timestamp 1586364061
transform 1 0 16836 0 1 19040
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_186
timestamp 1586364061
transform 1 0 17940 0 1 19040
box -38 -48 130 592
use scs8hd_decap_12  FILLER_31_184
timestamp 1586364061
transform 1 0 18032 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_196
timestamp 1586364061
transform 1 0 19136 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_208
timestamp 1586364061
transform 1 0 20240 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_220
timestamp 1586364061
transform 1 0 21344 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_3  PHY_63
timestamp 1586364061
transform -1 0 22816 0 1 19040
box -38 -48 314 592
use scs8hd_fill_1  FILLER_31_232
timestamp 1586364061
transform 1 0 22448 0 1 19040
box -38 -48 130 592
use scs8hd_decap_3  PHY_64
timestamp 1586364061
transform 1 0 1104 0 -1 20128
box -38 -48 314 592
use scs8hd_decap_12  FILLER_32_3
timestamp 1586364061
transform 1 0 1380 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_15
timestamp 1586364061
transform 1 0 2484 0 -1 20128
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_187
timestamp 1586364061
transform 1 0 3956 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_4  FILLER_32_27
timestamp 1586364061
transform 1 0 3588 0 -1 20128
box -38 -48 406 592
use scs8hd_decap_12  FILLER_32_32
timestamp 1586364061
transform 1 0 4048 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_44
timestamp 1586364061
transform 1 0 5152 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_56
timestamp 1586364061
transform 1 0 6256 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_68
timestamp 1586364061
transform 1 0 7360 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_80
timestamp 1586364061
transform 1 0 8464 0 -1 20128
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_188
timestamp 1586364061
transform 1 0 9568 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_12  FILLER_32_93
timestamp 1586364061
transform 1 0 9660 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_105
timestamp 1586364061
transform 1 0 10764 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_117
timestamp 1586364061
transform 1 0 11868 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_129
timestamp 1586364061
transform 1 0 12972 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_141
timestamp 1586364061
transform 1 0 14076 0 -1 20128
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_189
timestamp 1586364061
transform 1 0 15180 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_12  FILLER_32_154
timestamp 1586364061
transform 1 0 15272 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_166
timestamp 1586364061
transform 1 0 16376 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_178
timestamp 1586364061
transform 1 0 17480 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_190
timestamp 1586364061
transform 1 0 18584 0 -1 20128
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_190
timestamp 1586364061
transform 1 0 20792 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_12  FILLER_32_202
timestamp 1586364061
transform 1 0 19688 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_215
timestamp 1586364061
transform 1 0 20884 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_32_227
timestamp 1586364061
transform 1 0 21988 0 -1 20128
box -38 -48 590 592
use scs8hd_decap_3  PHY_65
timestamp 1586364061
transform -1 0 22816 0 -1 20128
box -38 -48 314 592
use scs8hd_decap_3  PHY_66
timestamp 1586364061
transform 1 0 1104 0 1 20128
box -38 -48 314 592
use scs8hd_decap_3  PHY_68
timestamp 1586364061
transform 1 0 1104 0 -1 21216
box -38 -48 314 592
use scs8hd_decap_12  FILLER_33_3
timestamp 1586364061
transform 1 0 1380 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_15
timestamp 1586364061
transform 1 0 2484 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_3
timestamp 1586364061
transform 1 0 1380 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_15
timestamp 1586364061
transform 1 0 2484 0 -1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_194
timestamp 1586364061
transform 1 0 3956 0 -1 21216
box -38 -48 130 592
use scs8hd_decap_12  FILLER_33_27
timestamp 1586364061
transform 1 0 3588 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_34_27
timestamp 1586364061
transform 1 0 3588 0 -1 21216
box -38 -48 406 592
use scs8hd_decap_12  FILLER_34_32
timestamp 1586364061
transform 1 0 4048 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_39
timestamp 1586364061
transform 1 0 4692 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_33_51
timestamp 1586364061
transform 1 0 5796 0 1 20128
box -38 -48 774 592
use scs8hd_decap_12  FILLER_34_44
timestamp 1586364061
transform 1 0 5152 0 -1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_191
timestamp 1586364061
transform 1 0 6716 0 1 20128
box -38 -48 130 592
use scs8hd_fill_2  FILLER_33_59
timestamp 1586364061
transform 1 0 6532 0 1 20128
box -38 -48 222 592
use scs8hd_decap_12  FILLER_33_62
timestamp 1586364061
transform 1 0 6808 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_56
timestamp 1586364061
transform 1 0 6256 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_68
timestamp 1586364061
transform 1 0 7360 0 -1 21216
box -38 -48 1142 592
use scs8hd_buf_2  _76_
timestamp 1586364061
transform 1 0 8648 0 1 20128
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__76__A
timestamp 1586364061
transform 1 0 9200 0 1 20128
box -38 -48 222 592
use scs8hd_decap_8  FILLER_33_74
timestamp 1586364061
transform 1 0 7912 0 1 20128
box -38 -48 774 592
use scs8hd_fill_2  FILLER_33_86
timestamp 1586364061
transform 1 0 9016 0 1 20128
box -38 -48 222 592
use scs8hd_decap_12  FILLER_34_80
timestamp 1586364061
transform 1 0 8464 0 -1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_195
timestamp 1586364061
transform 1 0 9568 0 -1 21216
box -38 -48 130 592
use scs8hd_decap_12  FILLER_33_90
timestamp 1586364061
transform 1 0 9384 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_102
timestamp 1586364061
transform 1 0 10488 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_93
timestamp 1586364061
transform 1 0 9660 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_105
timestamp 1586364061
transform 1 0 10764 0 -1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_192
timestamp 1586364061
transform 1 0 12328 0 1 20128
box -38 -48 130 592
use scs8hd_decap_8  FILLER_33_114
timestamp 1586364061
transform 1 0 11592 0 1 20128
box -38 -48 774 592
use scs8hd_decap_12  FILLER_33_123
timestamp 1586364061
transform 1 0 12420 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_117
timestamp 1586364061
transform 1 0 11868 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_135
timestamp 1586364061
transform 1 0 13524 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_129
timestamp 1586364061
transform 1 0 12972 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_141
timestamp 1586364061
transform 1 0 14076 0 -1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_196
timestamp 1586364061
transform 1 0 15180 0 -1 21216
box -38 -48 130 592
use scs8hd_decap_12  FILLER_33_147
timestamp 1586364061
transform 1 0 14628 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_159
timestamp 1586364061
transform 1 0 15732 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_154
timestamp 1586364061
transform 1 0 15272 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_171
timestamp 1586364061
transform 1 0 16836 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_166
timestamp 1586364061
transform 1 0 16376 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_178
timestamp 1586364061
transform 1 0 17480 0 -1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_193
timestamp 1586364061
transform 1 0 17940 0 1 20128
box -38 -48 130 592
use scs8hd_decap_12  FILLER_33_184
timestamp 1586364061
transform 1 0 18032 0 1 20128
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_33_196
timestamp 1586364061
transform 1 0 19136 0 1 20128
box -38 -48 130 592
use scs8hd_decap_12  FILLER_34_190
timestamp 1586364061
transform 1 0 18584 0 -1 21216
box -38 -48 1142 592
use scs8hd_buf_2  _85_
timestamp 1586364061
transform 1 0 19228 0 1 20128
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_197
timestamp 1586364061
transform 1 0 20792 0 -1 21216
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__85__A
timestamp 1586364061
transform 1 0 19780 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_201
timestamp 1586364061
transform 1 0 19596 0 1 20128
box -38 -48 222 592
use scs8hd_decap_8  FILLER_33_205
timestamp 1586364061
transform 1 0 19964 0 1 20128
box -38 -48 774 592
use scs8hd_fill_2  FILLER_33_213
timestamp 1586364061
transform 1 0 20700 0 1 20128
box -38 -48 222 592
use scs8hd_decap_12  FILLER_34_202
timestamp 1586364061
transform 1 0 19688 0 -1 21216
box -38 -48 1142 592
use scs8hd_buf_2  _81_
timestamp 1586364061
transform 1 0 20884 0 1 20128
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__81__A
timestamp 1586364061
transform 1 0 21436 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_219
timestamp 1586364061
transform 1 0 21252 0 1 20128
box -38 -48 222 592
use scs8hd_decap_8  FILLER_33_223
timestamp 1586364061
transform 1 0 21620 0 1 20128
box -38 -48 774 592
use scs8hd_fill_2  FILLER_33_231
timestamp 1586364061
transform 1 0 22356 0 1 20128
box -38 -48 222 592
use scs8hd_decap_12  FILLER_34_215
timestamp 1586364061
transform 1 0 20884 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_34_227
timestamp 1586364061
transform 1 0 21988 0 -1 21216
box -38 -48 590 592
use scs8hd_decap_3  PHY_67
timestamp 1586364061
transform -1 0 22816 0 1 20128
box -38 -48 314 592
use scs8hd_decap_3  PHY_69
timestamp 1586364061
transform -1 0 22816 0 -1 21216
box -38 -48 314 592
use scs8hd_decap_3  PHY_70
timestamp 1586364061
transform 1 0 1104 0 1 21216
box -38 -48 314 592
use scs8hd_decap_12  FILLER_35_3
timestamp 1586364061
transform 1 0 1380 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_15
timestamp 1586364061
transform 1 0 2484 0 1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_198
timestamp 1586364061
transform 1 0 3956 0 1 21216
box -38 -48 130 592
use scs8hd_decap_4  FILLER_35_27
timestamp 1586364061
transform 1 0 3588 0 1 21216
box -38 -48 406 592
use scs8hd_decap_12  FILLER_35_32
timestamp 1586364061
transform 1 0 4048 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_44
timestamp 1586364061
transform 1 0 5152 0 1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_199
timestamp 1586364061
transform 1 0 6808 0 1 21216
box -38 -48 130 592
use scs8hd_decap_6  FILLER_35_56
timestamp 1586364061
transform 1 0 6256 0 1 21216
box -38 -48 590 592
use scs8hd_decap_12  FILLER_35_63
timestamp 1586364061
transform 1 0 6900 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_75
timestamp 1586364061
transform 1 0 8004 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_35_87
timestamp 1586364061
transform 1 0 9108 0 1 21216
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_200
timestamp 1586364061
transform 1 0 9660 0 1 21216
box -38 -48 130 592
use scs8hd_decap_12  FILLER_35_94
timestamp 1586364061
transform 1 0 9752 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_106
timestamp 1586364061
transform 1 0 10856 0 1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_201
timestamp 1586364061
transform 1 0 12512 0 1 21216
box -38 -48 130 592
use scs8hd_decap_6  FILLER_35_118
timestamp 1586364061
transform 1 0 11960 0 1 21216
box -38 -48 590 592
use scs8hd_decap_12  FILLER_35_125
timestamp 1586364061
transform 1 0 12604 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_137
timestamp 1586364061
transform 1 0 13708 0 1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_202
timestamp 1586364061
transform 1 0 15364 0 1 21216
box -38 -48 130 592
use scs8hd_decap_6  FILLER_35_149
timestamp 1586364061
transform 1 0 14812 0 1 21216
box -38 -48 590 592
use scs8hd_decap_12  FILLER_35_156
timestamp 1586364061
transform 1 0 15456 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_168
timestamp 1586364061
transform 1 0 16560 0 1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_203
timestamp 1586364061
transform 1 0 18216 0 1 21216
box -38 -48 130 592
use scs8hd_decap_6  FILLER_35_180
timestamp 1586364061
transform 1 0 17664 0 1 21216
box -38 -48 590 592
use scs8hd_decap_12  FILLER_35_187
timestamp 1586364061
transform 1 0 18308 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_199
timestamp 1586364061
transform 1 0 19412 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_35_211
timestamp 1586364061
transform 1 0 20516 0 1 21216
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_204
timestamp 1586364061
transform 1 0 21068 0 1 21216
box -38 -48 130 592
use scs8hd_decap_12  FILLER_35_218
timestamp 1586364061
transform 1 0 21160 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_35_230
timestamp 1586364061
transform 1 0 22264 0 1 21216
box -38 -48 314 592
use scs8hd_decap_3  PHY_71
timestamp 1586364061
transform -1 0 22816 0 1 21216
box -38 -48 314 592
<< labels >>
rlabel metal3 s 0 1232 480 1352 6 address[0]
port 0 nsew default input
rlabel metal3 s 23520 688 24000 808 6 address[1]
port 1 nsew default input
rlabel metal2 s 4618 0 4674 480 6 address[2]
port 2 nsew default input
rlabel metal3 s 23520 2184 24000 2304 6 address[3]
port 3 nsew default input
rlabel metal3 s 0 3816 480 3936 6 address[4]
port 4 nsew default input
rlabel metal3 s 0 6536 480 6656 6 address[5]
port 5 nsew default input
rlabel metal3 s 0 9120 480 9240 6 bottom_grid_pin_0_
port 6 nsew default tristate
rlabel metal3 s 23520 3680 24000 3800 6 bottom_grid_pin_4_
port 7 nsew default tristate
rlabel metal2 s 6458 0 6514 480 6 bottom_grid_pin_8_
port 8 nsew default tristate
rlabel metal3 s 23520 5176 24000 5296 6 chanx_left_in[0]
port 9 nsew default input
rlabel metal3 s 23520 6672 24000 6792 6 chanx_left_in[1]
port 10 nsew default input
rlabel metal2 s 8298 0 8354 480 6 chanx_left_in[2]
port 11 nsew default input
rlabel metal3 s 0 11840 480 11960 6 chanx_left_in[3]
port 12 nsew default input
rlabel metal2 s 938 23520 994 24000 6 chanx_left_in[4]
port 13 nsew default input
rlabel metal3 s 23520 8168 24000 8288 6 chanx_left_in[5]
port 14 nsew default input
rlabel metal3 s 23520 9664 24000 9784 6 chanx_left_in[6]
port 15 nsew default input
rlabel metal2 s 2870 23520 2926 24000 6 chanx_left_in[7]
port 16 nsew default input
rlabel metal2 s 4894 23520 4950 24000 6 chanx_left_in[8]
port 17 nsew default input
rlabel metal2 s 6918 23520 6974 24000 6 chanx_left_out[0]
port 18 nsew default tristate
rlabel metal3 s 23520 11160 24000 11280 6 chanx_left_out[1]
port 19 nsew default tristate
rlabel metal2 s 10138 0 10194 480 6 chanx_left_out[2]
port 20 nsew default tristate
rlabel metal3 s 23520 12656 24000 12776 6 chanx_left_out[3]
port 21 nsew default tristate
rlabel metal2 s 8942 23520 8998 24000 6 chanx_left_out[4]
port 22 nsew default tristate
rlabel metal3 s 23520 14152 24000 14272 6 chanx_left_out[5]
port 23 nsew default tristate
rlabel metal3 s 23520 15648 24000 15768 6 chanx_left_out[6]
port 24 nsew default tristate
rlabel metal2 s 11978 0 12034 480 6 chanx_left_out[7]
port 25 nsew default tristate
rlabel metal2 s 13818 0 13874 480 6 chanx_left_out[8]
port 26 nsew default tristate
rlabel metal3 s 23520 17144 24000 17264 6 chanx_right_in[0]
port 27 nsew default input
rlabel metal2 s 10874 23520 10930 24000 6 chanx_right_in[1]
port 28 nsew default input
rlabel metal2 s 12898 23520 12954 24000 6 chanx_right_in[2]
port 29 nsew default input
rlabel metal2 s 14922 23520 14978 24000 6 chanx_right_in[3]
port 30 nsew default input
rlabel metal3 s 23520 18640 24000 18760 6 chanx_right_in[4]
port 31 nsew default input
rlabel metal2 s 15658 0 15714 480 6 chanx_right_in[5]
port 32 nsew default input
rlabel metal3 s 23520 20136 24000 20256 6 chanx_right_in[6]
port 33 nsew default input
rlabel metal2 s 16946 23520 17002 24000 6 chanx_right_in[7]
port 34 nsew default input
rlabel metal2 s 18878 23520 18934 24000 6 chanx_right_in[8]
port 35 nsew default input
rlabel metal3 s 0 14424 480 14544 6 chanx_right_out[0]
port 36 nsew default tristate
rlabel metal2 s 17498 0 17554 480 6 chanx_right_out[1]
port 37 nsew default tristate
rlabel metal2 s 19338 0 19394 480 6 chanx_right_out[2]
port 38 nsew default tristate
rlabel metal3 s 0 17144 480 17264 6 chanx_right_out[3]
port 39 nsew default tristate
rlabel metal2 s 20902 23520 20958 24000 6 chanx_right_out[4]
port 40 nsew default tristate
rlabel metal3 s 0 19728 480 19848 6 chanx_right_out[5]
port 41 nsew default tristate
rlabel metal2 s 21178 0 21234 480 6 chanx_right_out[6]
port 42 nsew default tristate
rlabel metal2 s 23018 0 23074 480 6 chanx_right_out[7]
port 43 nsew default tristate
rlabel metal2 s 22926 23520 22982 24000 6 chanx_right_out[8]
port 44 nsew default tristate
rlabel metal2 s 2778 0 2834 480 6 data_in
port 45 nsew default input
rlabel metal2 s 938 0 994 480 6 enable
port 46 nsew default input
rlabel metal3 s 23520 23128 24000 23248 6 top_grid_pin_14_
port 47 nsew default tristate
rlabel metal3 s 0 22448 480 22568 6 top_grid_pin_2_
port 48 nsew default tristate
rlabel metal3 s 23520 21632 24000 21752 6 top_grid_pin_6_
port 49 nsew default tristate
rlabel metal4 s 4944 2128 5264 21808 6 vpwr
port 50 nsew default input
rlabel metal4 s 8944 2128 9264 21808 6 vgnd
port 51 nsew default input
<< end >>
