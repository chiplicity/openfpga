* NGSPICE file created from sb_0__0_.ext - technology: EFS8A

* Black-box entry subcircuit for scs8hd_lpflow_inputisolatch_1 abstract view
.subckt scs8hd_lpflow_inputisolatch_1 D Q SLEEPB vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_decap_8 abstract view
.subckt scs8hd_decap_8 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_diode_2 abstract view
.subckt scs8hd_diode_2 DIODE vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_decap_6 abstract view
.subckt scs8hd_decap_6 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_fill_1 abstract view
.subckt scs8hd_fill_1 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_fill_2 abstract view
.subckt scs8hd_fill_2 vpwr vgnd
.ends

* Black-box entry subcircuit for scs8hd_inv_1 abstract view
.subckt scs8hd_inv_1 A Y vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_decap_12 abstract view
.subckt scs8hd_decap_12 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_ebufn_2 abstract view
.subckt scs8hd_ebufn_2 A TEB Z vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_inv_8 abstract view
.subckt scs8hd_inv_8 A Y vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_nor2_4 abstract view
.subckt scs8hd_nor2_4 A B Y vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_decap_4 abstract view
.subckt scs8hd_decap_4 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_buf_1 abstract view
.subckt scs8hd_buf_1 A X vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_decap_3 abstract view
.subckt scs8hd_decap_3 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_tapvpwrvgnd_1 abstract view
.subckt scs8hd_tapvpwrvgnd_1 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_or4_4 abstract view
.subckt scs8hd_or4_4 A B C D X vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_buf_2 abstract view
.subckt scs8hd_buf_2 A X vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_nor3_4 abstract view
.subckt scs8hd_nor3_4 A B C Y vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_or2_4 abstract view
.subckt scs8hd_or2_4 A B X vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_conb_1 abstract view
.subckt scs8hd_conb_1 HI LO vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_nand2_4 abstract view
.subckt scs8hd_nand2_4 A B Y vgnd vpwr
.ends

.subckt sb_0__0_ address[0] address[1] address[2] address[3] address[4] address[5]
+ chanx_right_in[0] chanx_right_in[1] chanx_right_in[2] chanx_right_in[3] chanx_right_in[4]
+ chanx_right_in[5] chanx_right_in[6] chanx_right_in[7] chanx_right_in[8] chanx_right_out[0]
+ chanx_right_out[1] chanx_right_out[2] chanx_right_out[3] chanx_right_out[4] chanx_right_out[5]
+ chanx_right_out[6] chanx_right_out[7] chanx_right_out[8] chany_top_in[0] chany_top_in[1]
+ chany_top_in[2] chany_top_in[3] chany_top_in[4] chany_top_in[5] chany_top_in[6]
+ chany_top_in[7] chany_top_in[8] chany_top_out[0] chany_top_out[1] chany_top_out[2]
+ chany_top_out[3] chany_top_out[4] chany_top_out[5] chany_top_out[6] chany_top_out[7]
+ chany_top_out[8] data_in enable right_bottom_grid_pin_11_ right_bottom_grid_pin_13_
+ right_bottom_grid_pin_15_ right_bottom_grid_pin_1_ right_bottom_grid_pin_3_ right_bottom_grid_pin_5_
+ right_bottom_grid_pin_7_ right_bottom_grid_pin_9_ right_top_grid_pin_10_ top_left_grid_pin_11_
+ top_left_grid_pin_13_ top_left_grid_pin_15_ top_left_grid_pin_1_ top_left_grid_pin_3_
+ top_left_grid_pin_5_ top_left_grid_pin_7_ top_left_grid_pin_9_ top_right_grid_pin_11_
+ vpwr vgnd
Xmem_right_track_12.LATCH_1_.latch data_in _202_/A _164_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_22_144 vgnd vpwr scs8hd_decap_8
XANTENNA_mem_top_track_2.LATCH_1_.latch_SLEEPB _111_/Y vgnd vpwr scs8hd_diode_2
XFILLER_26_41 vgnd vpwr scs8hd_decap_6
XFILLER_26_30 vgnd vpwr scs8hd_fill_1
XFILLER_13_100 vpwr vgnd scs8hd_fill_2
XFILLER_9_148 vpwr vgnd scs8hd_fill_2
XFILLER_13_144 vgnd vpwr scs8hd_fill_1
Xmux_top_track_8.INVTX1_0_.scs8hd_inv_1 top_left_grid_pin_9_ mux_top_track_8.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_27_269 vgnd vpwr scs8hd_decap_8
XFILLER_10_125 vpwr vgnd scs8hd_fill_2
XFILLER_10_158 vpwr vgnd scs8hd_fill_2
XFILLER_12_32 vgnd vpwr scs8hd_decap_12
Xmux_right_track_12.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_12.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ _202_/A mux_right_track_12.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XANTENNA_mem_top_track_16.LATCH_0_.latch_SLEEPB _142_/Y vgnd vpwr scs8hd_diode_2
XFILLER_37_95 vpwr vgnd scs8hd_fill_2
XANTENNA__108__B enable vgnd vpwr scs8hd_diode_2
XFILLER_5_162 vpwr vgnd scs8hd_fill_2
XANTENNA__124__A _127_/A vgnd vpwr scs8hd_diode_2
XFILLER_5_184 vgnd vpwr scs8hd_fill_1
XFILLER_24_239 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_right_track_4.tap_buf4_0_.scs8hd_inv_1_A mux_right_track_4.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
X_200_ _200_/A _200_/Y vgnd vpwr scs8hd_inv_8
X_131_ _150_/A _133_/B _131_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_23_86 vpwr vgnd scs8hd_fill_2
XFILLER_2_110 vpwr vgnd scs8hd_fill_2
XANTENNA__110__C _123_/C vgnd vpwr scs8hd_diode_2
XFILLER_17_9 vpwr vgnd scs8hd_fill_2
XANTENNA__119__A _127_/A vgnd vpwr scs8hd_diode_2
XFILLER_9_22 vgnd vpwr scs8hd_decap_12
XFILLER_9_66 vpwr vgnd scs8hd_fill_2
XFILLER_14_261 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_top_track_16.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_18_64 vpwr vgnd scs8hd_fill_2
XFILLER_18_75 vgnd vpwr scs8hd_decap_4
X_114_ _114_/A _115_/B vgnd vpwr scs8hd_buf_1
Xmux_right_track_16.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 _212_/HI _206_/Y mux_right_track_16.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_22_7 vgnd vpwr scs8hd_decap_12
Xmux_top_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 _217_/HI _172_/Y mux_top_track_0.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mem_top_track_6.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_39_19 vgnd vpwr scs8hd_decap_12
XFILLER_4_227 vgnd vpwr scs8hd_decap_12
XFILLER_35_109 vpwr vgnd scs8hd_fill_2
XANTENNA__116__B _116_/B vgnd vpwr scs8hd_diode_2
XFILLER_6_56 vgnd vpwr scs8hd_decap_3
XANTENNA__132__A address[0] vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_track_14.LATCH_1_.latch_SLEEPB _135_/Y vgnd vpwr scs8hd_diode_2
XFILLER_13_3 vgnd vpwr scs8hd_decap_12
XFILLER_19_172 vgnd vpwr scs8hd_decap_8
Xmem_right_track_8.LATCH_1_.latch data_in _198_/A _158_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_40_101 vgnd vpwr scs8hd_decap_12
XFILLER_25_164 vgnd vpwr scs8hd_decap_8
XFILLER_25_131 vgnd vpwr scs8hd_fill_1
XFILLER_17_109 vpwr vgnd scs8hd_fill_2
XFILLER_40_178 vgnd vpwr scs8hd_decap_12
XFILLER_31_53 vpwr vgnd scs8hd_fill_2
XFILLER_25_197 vgnd vpwr scs8hd_decap_12
XFILLER_15_87 vpwr vgnd scs8hd_fill_2
Xmux_right_track_6.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_6.INVTX1_0_.scs8hd_inv_1/Y
+ _197_/A mux_right_track_6.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XFILLER_31_134 vgnd vpwr scs8hd_decap_6
XFILLER_31_112 vgnd vpwr scs8hd_decap_8
XANTENNA__127__A _127_/A vgnd vpwr scs8hd_diode_2
XPHY_170 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_right_track_10.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _201_/Y vgnd
+ vpwr scs8hd_diode_2
XPHY_181 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_192 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_39_223 vpwr vgnd scs8hd_fill_2
XFILLER_39_245 vgnd vpwr scs8hd_decap_8
Xmem_top_track_4.LATCH_0_.latch data_in _177_/A _117_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_13_156 vpwr vgnd scs8hd_fill_2
XFILLER_42_63 vgnd vpwr scs8hd_decap_12
XFILLER_36_215 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_12.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_12.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_42_218 vgnd vpwr scs8hd_decap_12
XFILLER_12_44 vgnd vpwr scs8hd_decap_8
XFILLER_12_88 vpwr vgnd scs8hd_fill_2
XANTENNA__230__A _230_/A vgnd vpwr scs8hd_diode_2
XFILLER_18_215 vgnd vpwr scs8hd_decap_12
XANTENNA__124__B _124_/B vgnd vpwr scs8hd_diode_2
XANTENNA__140__A _115_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_0.INVTX1_0_.scs8hd_inv_1_A top_left_grid_pin_1_ vgnd vpwr scs8hd_diode_2
XFILLER_32_251 vgnd vpwr scs8hd_decap_12
Xmux_top_track_6.INVTX1_0_.scs8hd_inv_1 top_left_grid_pin_7_ mux_top_track_6.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_23_262 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_4.INVTX1_1_.scs8hd_inv_1_A chanx_right_in[3] vgnd vpwr scs8hd_diode_2
X_130_ _123_/A _115_/B _134_/C _123_/D _133_/B vgnd vpwr scs8hd_or4_4
XFILLER_23_21 vgnd vpwr scs8hd_fill_1
XFILLER_23_54 vgnd vpwr scs8hd_decap_3
XFILLER_2_144 vgnd vpwr scs8hd_fill_1
XANTENNA__110__D _110_/D vgnd vpwr scs8hd_diode_2
XANTENNA__119__B _119_/B vgnd vpwr scs8hd_diode_2
XFILLER_9_34 vgnd vpwr scs8hd_decap_12
XFILLER_14_273 vpwr vgnd scs8hd_fill_2
XANTENNA__135__A _150_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_track_2.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_20_276 vgnd vpwr scs8hd_fill_1
XFILLER_18_32 vpwr vgnd scs8hd_fill_2
XFILLER_34_64 vgnd vpwr scs8hd_decap_3
XFILLER_7_203 vgnd vpwr scs8hd_decap_4
XFILLER_7_236 vpwr vgnd scs8hd_fill_2
X_113_ address[2] _114_/A vgnd vpwr scs8hd_inv_8
XFILLER_11_254 vpwr vgnd scs8hd_fill_2
XFILLER_7_258 vgnd vpwr scs8hd_decap_4
XFILLER_15_7 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_12.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _203_/A vgnd
+ vpwr scs8hd_diode_2
Xmux_right_track_14.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_14.INVTX1_0_.scs8hd_inv_1/Y
+ _205_/A mux_right_track_14.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
Xmux_top_track_6.tap_buf4_0_.scs8hd_inv_1 mux_top_track_6.tap_buf4_0_.scs8hd_inv_1/A
+ _240_/A vgnd vpwr scs8hd_inv_1
XFILLER_29_118 vpwr vgnd scs8hd_fill_2
XFILLER_37_184 vgnd vpwr scs8hd_decap_12
XFILLER_1_90 vgnd vpwr scs8hd_decap_4
XFILLER_4_239 vgnd vpwr scs8hd_decap_12
XFILLER_4_206 vgnd vpwr scs8hd_decap_8
XFILLER_29_86 vgnd vpwr scs8hd_decap_12
XFILLER_29_53 vpwr vgnd scs8hd_fill_2
XFILLER_29_31 vpwr vgnd scs8hd_fill_2
XFILLER_28_184 vgnd vpwr scs8hd_fill_1
XANTENNA_mem_right_track_16.LATCH_0_.latch_SLEEPB _171_/Y vgnd vpwr scs8hd_diode_2
XFILLER_19_184 vgnd vpwr scs8hd_decap_12
XFILLER_34_154 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _189_/Y vgnd vpwr
+ scs8hd_diode_2
XFILLER_40_113 vgnd vpwr scs8hd_decap_12
XFILLER_25_176 vpwr vgnd scs8hd_fill_2
XFILLER_31_98 vpwr vgnd scs8hd_fill_2
XANTENNA__233__A _233_/A vgnd vpwr scs8hd_diode_2
XFILLER_31_102 vgnd vpwr scs8hd_decap_8
XANTENNA__127__B _128_/B vgnd vpwr scs8hd_diode_2
Xmux_right_track_16.INVTX1_0_.scs8hd_inv_1 chany_top_in[7] mux_right_track_16.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XPHY_160 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_16_154 vpwr vgnd scs8hd_fill_2
XFILLER_16_187 vgnd vpwr scs8hd_decap_12
XPHY_171 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_182 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_193 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__143__A _115_/A vgnd vpwr scs8hd_diode_2
XFILLER_39_202 vpwr vgnd scs8hd_fill_2
XFILLER_30_190 vgnd vpwr scs8hd_decap_12
XFILLER_22_179 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_right_track_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _192_/Y vgnd vpwr
+ scs8hd_diode_2
XFILLER_26_32 vgnd vpwr scs8hd_decap_6
XFILLER_26_21 vgnd vpwr scs8hd_fill_1
Xmux_top_track_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_top_track_2.INVTX1_1_.scs8hd_inv_1/Y
+ _175_/Y mux_top_track_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XANTENNA__228__A _228_/A vgnd vpwr scs8hd_diode_2
XFILLER_13_179 vpwr vgnd scs8hd_fill_2
XFILLER_42_75 vgnd vpwr scs8hd_decap_12
XFILLER_3_58 vgnd vpwr scs8hd_decap_3
XFILLER_36_227 vgnd vpwr scs8hd_decap_12
XANTENNA__138__A address[4] vgnd vpwr scs8hd_diode_2
XFILLER_27_205 vgnd vpwr scs8hd_decap_12
XFILLER_10_105 vpwr vgnd scs8hd_fill_2
XFILLER_12_56 vpwr vgnd scs8hd_fill_2
XFILLER_12_67 vgnd vpwr scs8hd_decap_4
XFILLER_37_53 vpwr vgnd scs8hd_fill_2
XFILLER_37_31 vgnd vpwr scs8hd_decap_8
XFILLER_33_208 vgnd vpwr scs8hd_decap_12
XFILLER_18_227 vgnd vpwr scs8hd_decap_12
XFILLER_5_120 vpwr vgnd scs8hd_fill_2
XFILLER_38_6 vgnd vpwr scs8hd_decap_12
XANTENNA__140__B _123_/B vgnd vpwr scs8hd_diode_2
XFILLER_32_263 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_right_track_14.LATCH_1_.latch_SLEEPB _168_/Y vgnd vpwr scs8hd_diode_2
XFILLER_15_208 vgnd vpwr scs8hd_decap_12
XFILLER_23_274 vgnd vpwr scs8hd_decap_3
XFILLER_23_241 vgnd vpwr scs8hd_fill_1
XFILLER_23_33 vgnd vpwr scs8hd_decap_4
XFILLER_23_66 vgnd vpwr scs8hd_decap_3
XANTENNA__241__A _241_/A vgnd vpwr scs8hd_diode_2
XFILLER_3_3 vpwr vgnd scs8hd_fill_2
XFILLER_2_123 vpwr vgnd scs8hd_fill_2
XFILLER_0_15 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_12.INVTX1_1_.scs8hd_inv_1_A right_bottom_grid_pin_11_ vgnd
+ vpwr scs8hd_diode_2
XFILLER_9_46 vgnd vpwr scs8hd_decap_4
XFILLER_9_57 vpwr vgnd scs8hd_fill_2
X_189_ _189_/A _189_/Y vgnd vpwr scs8hd_inv_8
XANTENNA__135__B _135_/B vgnd vpwr scs8hd_diode_2
XFILLER_36_3 vgnd vpwr scs8hd_decap_12
XANTENNA__151__A _151_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _175_/Y vgnd vpwr
+ scs8hd_diode_2
XFILLER_20_211 vgnd vpwr scs8hd_decap_3
XFILLER_18_44 vgnd vpwr scs8hd_decap_3
XFILLER_34_32 vgnd vpwr scs8hd_decap_12
XANTENNA__236__A _236_/A vgnd vpwr scs8hd_diode_2
XFILLER_11_233 vgnd vpwr scs8hd_decap_3
XFILLER_11_266 vgnd vpwr scs8hd_decap_8
X_112_ _128_/A _111_/B _112_/Y vgnd vpwr scs8hd_nor2_4
Xmux_top_track_4.INVTX1_0_.scs8hd_inv_1 top_left_grid_pin_5_ mux_top_track_4.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA__146__A address[3] vgnd vpwr scs8hd_diode_2
XFILLER_37_196 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_4.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _194_/A vgnd vpwr
+ scs8hd_diode_2
Xmux_right_track_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ _192_/A mux_right_track_2.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XFILLER_20_23 vgnd vpwr scs8hd_decap_8
XFILLER_20_67 vpwr vgnd scs8hd_fill_2
XFILLER_29_98 vgnd vpwr scs8hd_decap_4
XFILLER_3_262 vgnd vpwr scs8hd_decap_12
XFILLER_3_240 vgnd vpwr scs8hd_decap_4
XFILLER_34_166 vgnd vpwr scs8hd_decap_12
XFILLER_19_196 vgnd vpwr scs8hd_decap_12
XFILLER_40_125 vgnd vpwr scs8hd_decap_12
XFILLER_15_45 vpwr vgnd scs8hd_fill_2
XFILLER_31_77 vgnd vpwr scs8hd_decap_4
XFILLER_0_221 vpwr vgnd scs8hd_fill_2
XPHY_150 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_161 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_16_199 vgnd vpwr scs8hd_decap_12
XPHY_172 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_183 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_194 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__143__B _123_/B vgnd vpwr scs8hd_diode_2
XFILLER_39_258 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_4.INVTX1_0_.scs8hd_inv_1_A chany_top_in[1] vgnd vpwr scs8hd_diode_2
XFILLER_22_125 vgnd vpwr scs8hd_decap_6
XFILLER_22_158 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_top_track_12.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_top_track_12.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
Xmem_right_track_4.LATCH_1_.latch data_in _194_/A _150_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mem_right_track_2.LATCH_0_.latch_SLEEPB _148_/Y vgnd vpwr scs8hd_diode_2
XFILLER_42_87 vgnd vpwr scs8hd_decap_6
XFILLER_42_32 vgnd vpwr scs8hd_decap_12
XFILLER_9_118 vpwr vgnd scs8hd_fill_2
XFILLER_13_114 vpwr vgnd scs8hd_fill_2
XFILLER_13_136 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_8.INVTX1_1_.scs8hd_inv_1_A right_bottom_grid_pin_7_ vgnd
+ vpwr scs8hd_diode_2
Xmux_right_track_6.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 _215_/HI _196_/Y mux_right_track_6.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_36_239 vgnd vpwr scs8hd_decap_12
XANTENNA__138__B _166_/D vgnd vpwr scs8hd_diode_2
XANTENNA__154__A _170_/C vgnd vpwr scs8hd_diode_2
XFILLER_8_151 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_4.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _177_/A vgnd vpwr
+ scs8hd_diode_2
Xmux_right_track_14.INVTX1_0_.scs8hd_inv_1 chany_top_in[6] mux_right_track_14.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_27_217 vgnd vpwr scs8hd_decap_12
XFILLER_41_220 vgnd vpwr scs8hd_decap_12
XANTENNA__239__A _239_/A vgnd vpwr scs8hd_diode_2
XFILLER_18_239 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A _225_/HI vgnd vpwr
+ scs8hd_diode_2
Xmem_top_track_0.LATCH_0_.latch data_in _173_/A _107_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_5_132 vpwr vgnd scs8hd_fill_2
XANTENNA__140__C _149_/C vgnd vpwr scs8hd_diode_2
XANTENNA__149__A address[3] vgnd vpwr scs8hd_diode_2
XFILLER_4_91 vgnd vpwr scs8hd_fill_1
XFILLER_23_78 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_4.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_top_track_4.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_2_157 vpwr vgnd scs8hd_fill_2
XFILLER_0_27 vgnd vpwr scs8hd_decap_4
X_188_ _188_/A _188_/Y vgnd vpwr scs8hd_inv_8
XANTENNA__151__B _151_/B vgnd vpwr scs8hd_diode_2
Xmux_right_track_10.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_10.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ _200_/A mux_right_track_10.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XFILLER_34_44 vgnd vpwr scs8hd_decap_12
XFILLER_11_201 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_right_track_0.LATCH_1_.latch_SLEEPB _144_/Y vgnd vpwr scs8hd_diode_2
X_111_ _127_/A _111_/B _111_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA__146__B _115_/B vgnd vpwr scs8hd_diode_2
XFILLER_6_271 vgnd vpwr scs8hd_decap_4
XANTENNA__162__A _171_/C vgnd vpwr scs8hd_diode_2
XFILLER_37_131 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_right_track_14.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_29_11 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_right_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A _216_/HI vgnd vpwr
+ scs8hd_diode_2
XFILLER_6_15 vgnd vpwr scs8hd_decap_12
XFILLER_3_274 vgnd vpwr scs8hd_decap_3
XFILLER_19_120 vpwr vgnd scs8hd_fill_2
XFILLER_34_178 vgnd vpwr scs8hd_decap_12
XANTENNA__157__A _123_/A vgnd vpwr scs8hd_diode_2
XFILLER_19_153 vgnd vpwr scs8hd_fill_1
Xmux_top_track_2.INVTX1_0_.scs8hd_inv_1 top_left_grid_pin_3_ mux_top_track_2.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
Xmux_right_track_14.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 _211_/HI _204_/Y mux_right_track_14.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_25_123 vgnd vpwr scs8hd_decap_8
XFILLER_25_112 vpwr vgnd scs8hd_fill_2
XFILLER_40_137 vgnd vpwr scs8hd_decap_12
XFILLER_15_57 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_4.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_right_track_4.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_16_101 vpwr vgnd scs8hd_fill_2
XFILLER_16_134 vpwr vgnd scs8hd_fill_2
XFILLER_16_145 vgnd vpwr scs8hd_decap_8
XFILLER_31_148 vgnd vpwr scs8hd_decap_12
XFILLER_31_126 vpwr vgnd scs8hd_fill_2
XPHY_140 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_151 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_162 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_173 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_184 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_195 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__143__C _149_/C vgnd vpwr scs8hd_diode_2
XFILLER_11_3 vpwr vgnd scs8hd_fill_2
XFILLER_22_104 vgnd vpwr scs8hd_decap_8
XFILLER_38_270 vgnd vpwr scs8hd_decap_4
XFILLER_13_104 vpwr vgnd scs8hd_fill_2
XFILLER_42_44 vgnd vpwr scs8hd_decap_12
XFILLER_21_170 vpwr vgnd scs8hd_fill_2
Xmux_right_track_4.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_4.INVTX1_0_.scs8hd_inv_1/Y
+ _195_/A mux_right_track_4.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XANTENNA__154__B _153_/X vgnd vpwr scs8hd_diode_2
XANTENNA__170__A _110_/D vgnd vpwr scs8hd_diode_2
XFILLER_27_229 vgnd vpwr scs8hd_decap_12
XFILLER_10_129 vgnd vpwr scs8hd_decap_4
XFILLER_41_232 vgnd vpwr scs8hd_decap_12
XFILLER_37_99 vgnd vpwr scs8hd_decap_12
XFILLER_37_77 vgnd vpwr scs8hd_decap_3
XFILLER_26_251 vgnd vpwr scs8hd_decap_12
XFILLER_5_111 vgnd vpwr scs8hd_decap_3
XFILLER_5_166 vpwr vgnd scs8hd_fill_2
XANTENNA__140__D _140_/D vgnd vpwr scs8hd_diode_2
XANTENNA__149__B _115_/B vgnd vpwr scs8hd_diode_2
XFILLER_32_276 vgnd vpwr scs8hd_fill_1
XANTENNA__165__A _171_/C vgnd vpwr scs8hd_diode_2
XFILLER_4_81 vpwr vgnd scs8hd_fill_2
XFILLER_23_254 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_top_track_8.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_2_147 vgnd vpwr scs8hd_decap_6
Xmux_right_track_12.INVTX1_0_.scs8hd_inv_1 chany_top_in[5] mux_right_track_12.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_14_276 vgnd vpwr scs8hd_fill_1
X_187_ _187_/A _187_/Y vgnd vpwr scs8hd_inv_8
XFILLER_1_191 vpwr vgnd scs8hd_fill_2
Xmux_right_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_right_track_8.INVTX1_1_.scs8hd_inv_1/Y
+ _199_/Y mux_right_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XFILLER_34_78 vpwr vgnd scs8hd_fill_2
XFILLER_34_56 vgnd vpwr scs8hd_decap_8
XFILLER_11_213 vgnd vpwr scs8hd_decap_12
X_110_ _115_/A _123_/B _123_/C _110_/D _111_/B vgnd vpwr scs8hd_or4_4
XANTENNA_mux_right_track_10.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _200_/Y vgnd
+ vpwr scs8hd_diode_2
X_239_ _239_/A chany_top_out[4] vgnd vpwr scs8hd_buf_2
XANTENNA__146__C _149_/C vgnd vpwr scs8hd_diode_2
XFILLER_41_3 vgnd vpwr scs8hd_decap_12
XANTENNA__162__B _162_/B vgnd vpwr scs8hd_diode_2
XFILLER_37_143 vgnd vpwr scs8hd_decap_12
XFILLER_1_60 vgnd vpwr scs8hd_fill_1
XFILLER_1_71 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_16.tap_buf4_0_.scs8hd_inv_1_A mux_top_track_16.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_29_67 vpwr vgnd scs8hd_fill_2
XFILLER_28_154 vgnd vpwr scs8hd_decap_12
XFILLER_3_253 vpwr vgnd scs8hd_fill_2
XFILLER_6_27 vgnd vpwr scs8hd_decap_4
XFILLER_19_132 vpwr vgnd scs8hd_fill_2
XFILLER_34_102 vgnd vpwr scs8hd_decap_12
XANTENNA__157__B address[2] vgnd vpwr scs8hd_diode_2
XANTENNA__173__A _173_/A vgnd vpwr scs8hd_diode_2
XFILLER_25_135 vpwr vgnd scs8hd_fill_2
XFILLER_40_149 vgnd vpwr scs8hd_decap_4
Xmux_right_track_12.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_12.INVTX1_0_.scs8hd_inv_1/Y
+ _203_/A mux_right_track_12.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XFILLER_31_57 vpwr vgnd scs8hd_fill_2
XFILLER_0_245 vgnd vpwr scs8hd_decap_3
XPHY_130 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_141 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_152 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_196 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__143__D _149_/D vgnd vpwr scs8hd_diode_2
XPHY_163 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_174 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_185 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_39_227 vgnd vpwr scs8hd_decap_12
XANTENNA__168__A _123_/D vgnd vpwr scs8hd_diode_2
Xmux_top_track_0.INVTX1_0_.scs8hd_inv_1 top_left_grid_pin_1_ mux_top_track_0.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_26_57 vgnd vpwr scs8hd_decap_12
XFILLER_26_24 vgnd vpwr scs8hd_decap_4
XFILLER_42_56 vgnd vpwr scs8hd_decap_6
XFILLER_21_182 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_top_track_12.INVTX1_1_.scs8hd_inv_1_A chanx_right_in[7] vgnd vpwr scs8hd_diode_2
XFILLER_16_90 vpwr vgnd scs8hd_fill_2
XFILLER_8_186 vpwr vgnd scs8hd_fill_2
XFILLER_8_197 vgnd vpwr scs8hd_decap_12
XANTENNA__170__B _171_/B vgnd vpwr scs8hd_diode_2
XFILLER_12_182 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_14.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_14.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_37_89 vgnd vpwr scs8hd_decap_4
Xmux_right_track_8.INVTX1_1_.scs8hd_inv_1 right_bottom_grid_pin_7_ mux_right_track_8.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_26_263 vgnd vpwr scs8hd_decap_12
Xmem_right_track_0.LATCH_1_.latch data_in _190_/A _144_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
Xmem_top_track_8.LATCH_1_.latch data_in _180_/A _124_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_5_178 vgnd vpwr scs8hd_decap_3
XFILLER_5_145 vpwr vgnd scs8hd_fill_2
XFILLER_5_123 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_right_track_12.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _202_/A vgnd
+ vpwr scs8hd_diode_2
Xmux_right_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_right_track_16.INVTX1_1_.scs8hd_inv_1/Y
+ _207_/Y mux_right_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
Xmux_top_track_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_top_track_0.INVTX1_1_.scs8hd_inv_1/Y
+ _173_/Y mux_top_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_right_track_10.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_10.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__149__C _149_/C vgnd vpwr scs8hd_diode_2
XFILLER_17_241 vgnd vpwr scs8hd_decap_3
XANTENNA__165__B _165_/B vgnd vpwr scs8hd_diode_2
XANTENNA__181__A _181_/A vgnd vpwr scs8hd_diode_2
XFILLER_4_93 vgnd vpwr scs8hd_decap_4
XFILLER_2_104 vgnd vpwr scs8hd_decap_4
X_186_ _186_/A _186_/Y vgnd vpwr scs8hd_inv_8
XANTENNA_mux_right_track_4.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _195_/Y vgnd vpwr
+ scs8hd_diode_2
XFILLER_1_181 vpwr vgnd scs8hd_fill_2
XANTENNA__176__A _176_/A vgnd vpwr scs8hd_diode_2
XFILLER_9_270 vgnd vpwr scs8hd_decap_6
XANTENNA_mux_top_track_16.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _188_/Y vgnd vpwr
+ scs8hd_diode_2
XFILLER_18_36 vgnd vpwr scs8hd_decap_8
XFILLER_18_58 vgnd vpwr scs8hd_decap_4
XFILLER_11_225 vgnd vpwr scs8hd_decap_8
XFILLER_11_258 vpwr vgnd scs8hd_fill_2
XFILLER_1_3 vgnd vpwr scs8hd_decap_12
X_238_ _238_/A chany_top_out[5] vgnd vpwr scs8hd_buf_2
XANTENNA__146__D _140_/D vgnd vpwr scs8hd_diode_2
Xmux_right_track_10.INVTX1_0_.scs8hd_inv_1 chany_top_in[4] mux_right_track_10.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
X_169_ _123_/D _171_/B _171_/C _169_/Y vgnd vpwr scs8hd_nor3_4
XFILLER_34_3 vgnd vpwr scs8hd_decap_12
XFILLER_37_155 vgnd vpwr scs8hd_decap_12
XFILLER_37_111 vgnd vpwr scs8hd_decap_8
XANTENNA_mem_right_track_8.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_20_15 vgnd vpwr scs8hd_decap_4
XFILLER_29_57 vgnd vpwr scs8hd_decap_4
XFILLER_29_35 vgnd vpwr scs8hd_decap_3
XFILLER_28_188 vgnd vpwr scs8hd_decap_12
XFILLER_28_166 vgnd vpwr scs8hd_decap_12
XFILLER_10_81 vpwr vgnd scs8hd_fill_2
XFILLER_34_114 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_top_track_10.LATCH_0_.latch_SLEEPB _128_/Y vgnd vpwr scs8hd_diode_2
XFILLER_42_180 vgnd vpwr scs8hd_decap_6
XFILLER_34_125 vgnd vpwr scs8hd_decap_12
XANTENNA__157__C _149_/C vgnd vpwr scs8hd_diode_2
XFILLER_25_103 vgnd vpwr scs8hd_decap_6
XFILLER_33_180 vgnd vpwr scs8hd_decap_3
XFILLER_0_202 vpwr vgnd scs8hd_fill_2
XFILLER_16_114 vgnd vpwr scs8hd_decap_8
XPHY_120 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_131 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_142 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_153 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_16_125 vgnd vpwr scs8hd_decap_3
XFILLER_16_158 vgnd vpwr scs8hd_fill_1
XPHY_164 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_175 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_197 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmux_right_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ _190_/A mux_right_track_0.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XPHY_186 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_39_239 vgnd vpwr scs8hd_decap_4
XFILLER_39_206 vgnd vpwr scs8hd_decap_12
XPHY_0 vgnd vpwr scs8hd_decap_3
XANTENNA__168__B _171_/B vgnd vpwr scs8hd_diode_2
XANTENNA__184__A _184_/A vgnd vpwr scs8hd_diode_2
XFILLER_15_180 vgnd vpwr scs8hd_decap_3
XFILLER_7_60 vgnd vpwr scs8hd_fill_1
XFILLER_26_69 vpwr vgnd scs8hd_fill_2
XFILLER_26_47 vgnd vpwr scs8hd_fill_1
XFILLER_21_161 vgnd vpwr scs8hd_decap_6
Xmem_top_track_14.LATCH_0_.latch data_in _187_/A _136_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_right_track_6.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _197_/A vgnd vpwr
+ scs8hd_diode_2
XFILLER_8_132 vgnd vpwr scs8hd_decap_3
XFILLER_8_143 vgnd vpwr scs8hd_decap_8
XFILLER_8_154 vgnd vpwr scs8hd_decap_3
XANTENNA__170__C _170_/C vgnd vpwr scs8hd_diode_2
XANTENNA__179__A _179_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _174_/Y vgnd vpwr
+ scs8hd_diode_2
XFILLER_35_220 vgnd vpwr scs8hd_decap_12
XFILLER_10_109 vpwr vgnd scs8hd_fill_2
Xmux_right_track_12.tap_buf4_0_.scs8hd_inv_1 mux_right_track_12.tap_buf4_0_.scs8hd_inv_1/A
+ _228_/A vgnd vpwr scs8hd_inv_1
XFILLER_37_57 vpwr vgnd scs8hd_fill_2
XFILLER_41_245 vgnd vpwr scs8hd_decap_12
Xmux_top_track_14.tap_buf4_0_.scs8hd_inv_1 mux_top_track_14.tap_buf4_0_.scs8hd_inv_1/A
+ _236_/A vgnd vpwr scs8hd_inv_1
XFILLER_27_90 vgnd vpwr scs8hd_decap_6
XANTENNA__149__D _149_/D vgnd vpwr scs8hd_diode_2
Xmux_right_track_4.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 _214_/HI _194_/Y mux_right_track_4.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_23_15 vgnd vpwr scs8hd_decap_6
XFILLER_23_37 vgnd vpwr scs8hd_fill_1
XFILLER_23_59 vpwr vgnd scs8hd_fill_2
XFILLER_23_201 vgnd vpwr scs8hd_decap_12
XFILLER_3_7 vgnd vpwr scs8hd_decap_12
XFILLER_2_127 vgnd vpwr scs8hd_decap_4
X_185_ _185_/A _185_/Y vgnd vpwr scs8hd_inv_8
XFILLER_13_70 vpwr vgnd scs8hd_fill_2
Xmux_right_track_6.INVTX1_1_.scs8hd_inv_1 right_bottom_grid_pin_5_ mux_right_track_6.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_20_215 vgnd vpwr scs8hd_decap_12
XANTENNA__192__A _192_/A vgnd vpwr scs8hd_diode_2
XFILLER_18_15 vgnd vpwr scs8hd_decap_12
XFILLER_40_90 vpwr vgnd scs8hd_fill_2
XFILLER_24_91 vgnd vpwr scs8hd_fill_1
X_237_ _237_/A chany_top_out[6] vgnd vpwr scs8hd_buf_2
X_168_ _123_/D _171_/B _170_/C _168_/Y vgnd vpwr scs8hd_nor3_4
XFILLER_27_3 vgnd vpwr scs8hd_decap_8
X_099_ address[4] address[5] _134_/C vgnd vpwr scs8hd_or2_4
XFILLER_37_167 vgnd vpwr scs8hd_decap_12
XFILLER_1_51 vgnd vpwr scs8hd_fill_1
XFILLER_1_62 vpwr vgnd scs8hd_fill_2
XANTENNA__187__A _187_/A vgnd vpwr scs8hd_diode_2
XFILLER_28_145 vgnd vpwr scs8hd_decap_8
XFILLER_28_134 vgnd vpwr scs8hd_decap_8
XFILLER_28_101 vpwr vgnd scs8hd_fill_2
XFILLER_28_178 vgnd vpwr scs8hd_decap_6
XANTENNA__097__A address[3] vgnd vpwr scs8hd_diode_2
XFILLER_34_137 vgnd vpwr scs8hd_decap_12
XFILLER_19_156 vpwr vgnd scs8hd_fill_2
XANTENNA__157__D _149_/D vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_4.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _176_/A vgnd vpwr
+ scs8hd_diode_2
XFILLER_15_49 vgnd vpwr scs8hd_decap_8
XFILLER_31_15 vgnd vpwr scs8hd_decap_12
XFILLER_0_225 vgnd vpwr scs8hd_decap_12
XFILLER_0_214 vgnd vpwr scs8hd_decap_3
XFILLER_24_192 vgnd vpwr scs8hd_decap_12
XPHY_198 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_110 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_121 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_132 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_143 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_154 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_165 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_176 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_187 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_39_218 vpwr vgnd scs8hd_fill_2
XPHY_1 vgnd vpwr scs8hd_decap_3
XANTENNA__168__C _170_/C vgnd vpwr scs8hd_diode_2
XFILLER_38_251 vgnd vpwr scs8hd_decap_4
XFILLER_26_15 vgnd vpwr scs8hd_decap_6
XANTENNA_mux_top_track_14.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_top_track_14.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
Xmux_right_track_6.tap_buf4_0_.scs8hd_inv_1 mux_right_track_6.tap_buf4_0_.scs8hd_inv_1/A
+ _231_/A vgnd vpwr scs8hd_inv_1
XFILLER_13_118 vpwr vgnd scs8hd_fill_2
Xmux_right_track_12.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 _210_/HI _202_/Y mux_right_track_12.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_21_184 vgnd vpwr scs8hd_decap_3
XFILLER_3_19 vgnd vpwr scs8hd_decap_12
XFILLER_29_240 vgnd vpwr scs8hd_decap_4
XFILLER_8_111 vgnd vpwr scs8hd_decap_8
XANTENNA__195__A _195_/A vgnd vpwr scs8hd_diode_2
XFILLER_35_232 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_10.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_top_track_10.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_26_276 vgnd vpwr scs8hd_fill_1
XFILLER_26_210 vgnd vpwr scs8hd_decap_4
XFILLER_41_257 vgnd vpwr scs8hd_decap_12
XFILLER_32_202 vgnd vpwr scs8hd_decap_12
XFILLER_4_191 vgnd vpwr scs8hd_decap_8
XFILLER_4_73 vpwr vgnd scs8hd_fill_2
XFILLER_23_213 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_right_track_10.LATCH_0_.latch_SLEEPB _162_/Y vgnd vpwr scs8hd_diode_2
Xmux_right_track_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_2.INVTX1_0_.scs8hd_inv_1/Y
+ _193_/A mux_right_track_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_top_track_6.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_top_track_6.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_14_213 vgnd vpwr scs8hd_fill_1
X_184_ _184_/A _184_/Y vgnd vpwr scs8hd_inv_8
XFILLER_29_7 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_right_track_16.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
Xmem_top_track_4.LATCH_1_.latch data_in _176_/A _116_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_20_227 vgnd vpwr scs8hd_decap_12
XFILLER_18_27 vgnd vpwr scs8hd_decap_4
XFILLER_34_15 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_top_track_14.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_11_238 vgnd vpwr scs8hd_decap_4
XFILLER_24_70 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_top_track_4.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
X_236_ _236_/A chany_top_out[7] vgnd vpwr scs8hd_buf_2
XFILLER_6_231 vgnd vpwr scs8hd_decap_4
X_167_ _167_/A _171_/B vgnd vpwr scs8hd_buf_1
X_098_ address[2] _123_/B vgnd vpwr scs8hd_buf_1
XFILLER_37_179 vgnd vpwr scs8hd_decap_4
Xmux_right_track_4.INVTX1_1_.scs8hd_inv_1 right_bottom_grid_pin_3_ mux_right_track_4.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_36_190 vgnd vpwr scs8hd_decap_12
Xmux_right_track_6.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_right_track_6.INVTX1_1_.scs8hd_inv_1/Y
+ _197_/Y mux_right_track_6.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XANTENNA_mem_top_track_8.LATCH_0_.latch_SLEEPB _125_/Y vgnd vpwr scs8hd_diode_2
XFILLER_3_245 vgnd vpwr scs8hd_decap_8
XFILLER_34_149 vgnd vpwr scs8hd_decap_4
XFILLER_19_92 vgnd vpwr scs8hd_decap_4
X_219_ _219_/HI _219_/LO vgnd vpwr scs8hd_conb_1
XANTENNA__198__A _198_/A vgnd vpwr scs8hd_diode_2
XFILLER_25_116 vgnd vpwr scs8hd_decap_6
XFILLER_31_27 vgnd vpwr scs8hd_decap_12
XFILLER_0_237 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_right_track_6.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_right_track_6.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XPHY_100 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_16_138 vgnd vpwr scs8hd_decap_4
XPHY_199 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_111 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_122 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_133 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_144 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_155 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_166 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_177 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_188 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_21_82 vpwr vgnd scs8hd_fill_2
XFILLER_11_7 vgnd vpwr scs8hd_decap_8
XPHY_2 vgnd vpwr scs8hd_decap_3
XFILLER_15_171 vgnd vpwr scs8hd_decap_6
XFILLER_30_152 vgnd vpwr scs8hd_fill_1
XFILLER_7_51 vgnd vpwr scs8hd_decap_3
XFILLER_7_62 vgnd vpwr scs8hd_decap_3
XFILLER_7_73 vgnd vpwr scs8hd_decap_3
XFILLER_7_95 vpwr vgnd scs8hd_fill_2
XFILLER_38_274 vgnd vpwr scs8hd_fill_1
XFILLER_26_38 vgnd vpwr scs8hd_fill_1
XFILLER_42_15 vgnd vpwr scs8hd_decap_12
XFILLER_13_108 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_right_track_12.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _203_/Y vgnd
+ vpwr scs8hd_diode_2
XFILLER_21_174 vgnd vpwr scs8hd_decap_8
XFILLER_29_252 vgnd vpwr scs8hd_decap_12
XFILLER_16_60 vpwr vgnd scs8hd_fill_2
XFILLER_16_82 vpwr vgnd scs8hd_fill_2
XFILLER_16_93 vgnd vpwr scs8hd_fill_1
XFILLER_8_167 vpwr vgnd scs8hd_fill_2
Xmux_right_track_10.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_10.INVTX1_0_.scs8hd_inv_1/Y
+ _201_/A mux_right_track_10.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XFILLER_12_163 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_0.INVTX1_1_.scs8hd_inv_1_A chanx_right_in[1] vgnd vpwr scs8hd_diode_2
XFILLER_12_18 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_16.tap_buf4_0_.scs8hd_inv_1_A mux_right_track_16.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_41_269 vgnd vpwr scs8hd_decap_8
Xmem_top_track_10.LATCH_0_.latch data_in _183_/A _128_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mem_top_track_6.LATCH_1_.latch_SLEEPB _119_/Y vgnd vpwr scs8hd_diode_2
XFILLER_4_85 vgnd vpwr scs8hd_decap_6
XFILLER_4_30 vgnd vpwr scs8hd_fill_1
XFILLER_23_225 vgnd vpwr scs8hd_decap_12
XFILLER_23_258 vpwr vgnd scs8hd_fill_2
Xmux_top_track_2.tap_buf4_0_.scs8hd_inv_1 mux_top_track_2.tap_buf4_0_.scs8hd_inv_1/A
+ _242_/A vgnd vpwr scs8hd_inv_1
X_183_ _183_/A _183_/Y vgnd vpwr scs8hd_inv_8
XFILLER_13_83 vpwr vgnd scs8hd_fill_2
XFILLER_1_173 vgnd vpwr scs8hd_decap_8
XANTENNA_mem_right_track_0.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
Xmux_right_track_14.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_right_track_14.INVTX1_1_.scs8hd_inv_1/Y
+ _205_/Y mux_right_track_14.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XFILLER_20_239 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_8.tap_buf4_0_.scs8hd_inv_1_A mux_top_track_8.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_34_27 vgnd vpwr scs8hd_decap_4
Xmux_top_track_16.INVTX1_1_.scs8hd_inv_1 chanx_right_in[0] mux_top_track_16.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_24_93 vpwr vgnd scs8hd_fill_2
X_235_ _235_/A chany_top_out[8] vgnd vpwr scs8hd_buf_2
XFILLER_6_276 vgnd vpwr scs8hd_fill_1
X_166_ address[3] address[2] address[4] _166_/D _167_/A vgnd vpwr scs8hd_or4_4
X_097_ address[3] _115_/A vgnd vpwr scs8hd_buf_1
XFILLER_1_86 vpwr vgnd scs8hd_fill_2
XFILLER_1_97 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_14.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _205_/A vgnd
+ vpwr scs8hd_diode_2
XFILLER_29_16 vgnd vpwr scs8hd_decap_4
XFILLER_19_71 vpwr vgnd scs8hd_fill_2
XFILLER_19_114 vgnd vpwr scs8hd_decap_4
XFILLER_19_136 vpwr vgnd scs8hd_fill_2
X_218_ _218_/HI _218_/LO vgnd vpwr scs8hd_conb_1
X_149_ address[3] _115_/B _149_/C _149_/D _151_/B vgnd vpwr scs8hd_or4_4
XFILLER_32_3 vgnd vpwr scs8hd_decap_12
XFILLER_25_139 vpwr vgnd scs8hd_fill_2
XFILLER_31_39 vgnd vpwr scs8hd_decap_3
XFILLER_0_249 vgnd vpwr scs8hd_decap_12
Xmux_right_track_2.INVTX1_1_.scs8hd_inv_1 right_bottom_grid_pin_1_ mux_right_track_2.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XPHY_112 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_101 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_123 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_134 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_145 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_156 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_167 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_178 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_189 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_3 vgnd vpwr scs8hd_decap_3
XFILLER_15_150 vpwr vgnd scs8hd_fill_2
XFILLER_7_85 vpwr vgnd scs8hd_fill_2
XFILLER_42_27 vgnd vpwr scs8hd_decap_4
XFILLER_21_120 vpwr vgnd scs8hd_fill_2
XFILLER_29_264 vgnd vpwr scs8hd_decap_12
XFILLER_8_102 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_right_track_4.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _194_/Y vgnd vpwr
+ scs8hd_diode_2
XFILLER_32_60 vgnd vpwr scs8hd_decap_12
XFILLER_12_186 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_top_track_6.INVTX1_0_.scs8hd_inv_1_A top_left_grid_pin_7_ vgnd vpwr scs8hd_diode_2
XFILLER_35_245 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_16.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_5_149 vpwr vgnd scs8hd_fill_2
XFILLER_5_116 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_8.tap_buf4_0_.scs8hd_inv_1_A mux_right_track_8.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_27_71 vpwr vgnd scs8hd_fill_2
XFILLER_17_245 vgnd vpwr scs8hd_decap_12
XFILLER_32_215 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_10.tap_buf4_0_.scs8hd_inv_1_A mux_top_track_10.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_4_182 vgnd vpwr scs8hd_decap_3
XFILLER_4_97 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_right_track_12.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_12.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_23_237 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_top_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_top_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
X_182_ _182_/A _182_/Y vgnd vpwr scs8hd_inv_8
XFILLER_14_215 vgnd vpwr scs8hd_decap_12
XFILLER_22_270 vgnd vpwr scs8hd_decap_4
XFILLER_13_62 vgnd vpwr scs8hd_fill_1
XFILLER_1_152 vpwr vgnd scs8hd_fill_2
XANTENNA__100__A _134_/C vgnd vpwr scs8hd_diode_2
XFILLER_9_241 vgnd vpwr scs8hd_fill_1
Xmux_right_track_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 _213_/HI _192_/Y mux_right_track_2.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_top_track_4.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _177_/Y vgnd vpwr
+ scs8hd_diode_2
XFILLER_24_83 vgnd vpwr scs8hd_decap_8
X_234_ _234_/A chanx_right_out[0] vgnd vpwr scs8hd_buf_2
XFILLER_6_211 vgnd vpwr scs8hd_decap_3
XFILLER_10_273 vpwr vgnd scs8hd_fill_2
X_165_ _171_/C _165_/B _165_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_40_93 vgnd vpwr scs8hd_decap_4
XFILLER_40_82 vgnd vpwr scs8hd_decap_8
XFILLER_40_71 vgnd vpwr scs8hd_decap_8
XFILLER_40_60 vgnd vpwr scs8hd_decap_8
X_096_ _096_/A _127_/A vgnd vpwr scs8hd_buf_1
XFILLER_1_54 vgnd vpwr scs8hd_decap_6
Xmem_top_track_0.LATCH_1_.latch data_in _172_/A _105_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_20_19 vgnd vpwr scs8hd_fill_1
XFILLER_3_258 vpwr vgnd scs8hd_fill_2
XFILLER_10_52 vgnd vpwr scs8hd_decap_3
XFILLER_10_85 vpwr vgnd scs8hd_fill_2
XFILLER_10_96 vgnd vpwr scs8hd_decap_6
XANTENNA_mux_right_track_6.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _196_/A vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_right_track_0.INVTX1_0_.scs8hd_inv_1_A chany_top_in[8] vgnd vpwr scs8hd_diode_2
Xmux_top_track_14.INVTX1_1_.scs8hd_inv_1 chanx_right_in[8] mux_top_track_14.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
X_217_ _217_/HI _217_/LO vgnd vpwr scs8hd_conb_1
X_148_ _151_/A _147_/B _148_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_25_3 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_4.INVTX1_1_.scs8hd_inv_1_A right_bottom_grid_pin_3_ vgnd
+ vpwr scs8hd_diode_2
XFILLER_15_19 vgnd vpwr scs8hd_decap_12
XFILLER_33_184 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_0_206 vgnd vpwr scs8hd_decap_8
XFILLER_24_162 vpwr vgnd scs8hd_fill_2
XPHY_113 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_102 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_124 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_135 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_146 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_157 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_168 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_179 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_21_51 vgnd vpwr scs8hd_fill_1
XFILLER_21_62 vgnd vpwr scs8hd_decap_4
XFILLER_21_95 vpwr vgnd scs8hd_fill_2
XFILLER_30_154 vgnd vpwr scs8hd_decap_12
XFILLER_30_132 vgnd vpwr scs8hd_decap_12
XFILLER_30_121 vgnd vpwr scs8hd_decap_8
XPHY_4 vgnd vpwr scs8hd_decap_3
XFILLER_15_184 vgnd vpwr scs8hd_decap_12
XFILLER_38_276 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_top_track_10.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _183_/A vgnd vpwr
+ scs8hd_diode_2
XFILLER_29_276 vgnd vpwr scs8hd_fill_1
XFILLER_16_40 vgnd vpwr scs8hd_decap_3
XFILLER_32_72 vgnd vpwr scs8hd_fill_1
Xmux_right_track_0.INVTX1_1_.scs8hd_inv_1 right_top_grid_pin_10_ mux_right_track_0.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA__103__A _140_/D vgnd vpwr scs8hd_diode_2
XFILLER_35_257 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_14.INVTX1_0_.scs8hd_inv_1_A chany_top_in[6] vgnd vpwr scs8hd_diode_2
XFILLER_7_180 vgnd vpwr scs8hd_fill_1
XFILLER_37_39 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_top_track_6.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _179_/A vgnd vpwr
+ scs8hd_diode_2
XFILLER_5_128 vpwr vgnd scs8hd_fill_2
XFILLER_32_227 vgnd vpwr scs8hd_decap_12
XFILLER_17_257 vgnd vpwr scs8hd_decap_12
Xmux_right_track_10.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 _209_/HI _200_/Y mux_right_track_10.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_4_65 vpwr vgnd scs8hd_fill_2
XFILLER_4_32 vgnd vpwr scs8hd_decap_12
XFILLER_14_227 vgnd vpwr scs8hd_decap_12
X_181_ _181_/A _181_/Y vgnd vpwr scs8hd_inv_8
XFILLER_14_249 vgnd vpwr scs8hd_decap_12
Xmem_right_track_14.LATCH_0_.latch data_in _205_/A _169_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_38_71 vgnd vpwr scs8hd_decap_4
XANTENNA__201__A _201_/A vgnd vpwr scs8hd_diode_2
Xmux_right_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_0.INVTX1_0_.scs8hd_inv_1/Y
+ _191_/A mux_right_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
X_233_ _233_/A chanx_right_out[1] vgnd vpwr scs8hd_buf_2
X_164_ _170_/C _165_/B _164_/Y vgnd vpwr scs8hd_nor2_4
X_095_ address[0] _096_/A vgnd vpwr scs8hd_inv_8
XFILLER_37_127 vpwr vgnd scs8hd_fill_2
XANTENNA__111__A _127_/A vgnd vpwr scs8hd_diode_2
XFILLER_28_105 vgnd vpwr scs8hd_fill_1
XANTENNA_mem_right_track_12.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_3_204 vgnd vpwr scs8hd_decap_12
XFILLER_10_64 vpwr vgnd scs8hd_fill_2
XFILLER_19_149 vgnd vpwr scs8hd_decap_4
XFILLER_27_193 vgnd vpwr scs8hd_decap_12
X_216_ _216_/HI _216_/LO vgnd vpwr scs8hd_conb_1
XANTENNA__106__A address[0] vgnd vpwr scs8hd_diode_2
X_147_ _150_/A _147_/B _147_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA_mux_right_track_10.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A _209_/HI vgnd vpwr
+ scs8hd_diode_2
XFILLER_18_3 vgnd vpwr scs8hd_decap_12
XFILLER_33_196 vgnd vpwr scs8hd_decap_12
XPHY_114 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_103 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_125 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_136 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_147 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_158 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_169 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_21_30 vpwr vgnd scs8hd_fill_2
Xmux_top_track_16.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_top_track_16.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ _188_/A mux_top_track_16.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XPHY_5 vgnd vpwr scs8hd_decap_3
Xmux_right_track_4.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_right_track_4.INVTX1_1_.scs8hd_inv_1/Y
+ _195_/Y mux_right_track_4.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XFILLER_30_166 vgnd vpwr scs8hd_decap_12
XFILLER_30_144 vgnd vpwr scs8hd_decap_8
XFILLER_15_163 vpwr vgnd scs8hd_fill_2
XFILLER_15_196 vgnd vpwr scs8hd_decap_12
Xmux_top_track_12.INVTX1_1_.scs8hd_inv_1 chanx_right_in[7] mux_top_track_12.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_21_133 vpwr vgnd scs8hd_fill_2
XFILLER_21_144 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_16.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_top_track_16.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_16_52 vpwr vgnd scs8hd_fill_2
XFILLER_8_137 vgnd vpwr scs8hd_decap_3
XFILLER_8_159 vgnd vpwr scs8hd_decap_8
XFILLER_12_199 vgnd vpwr scs8hd_decap_12
XFILLER_32_84 vgnd vpwr scs8hd_decap_8
XFILLER_35_269 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_top_track_12.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_top_track_12.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_5_107 vpwr vgnd scs8hd_fill_2
XANTENNA__204__A _204_/A vgnd vpwr scs8hd_diode_2
XFILLER_32_239 vgnd vpwr scs8hd_decap_12
XFILLER_27_62 vgnd vpwr scs8hd_decap_3
XFILLER_27_51 vpwr vgnd scs8hd_fill_2
XFILLER_17_269 vgnd vpwr scs8hd_decap_8
XANTENNA_mem_right_track_6.LATCH_0_.latch_SLEEPB _156_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_track_16.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_4_140 vgnd vpwr scs8hd_decap_12
XFILLER_4_77 vpwr vgnd scs8hd_fill_2
XFILLER_4_44 vgnd vpwr scs8hd_decap_12
XANTENNA__114__A _114_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_track_6.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_14_239 vgnd vpwr scs8hd_decap_8
XFILLER_13_53 vpwr vgnd scs8hd_fill_2
X_180_ _180_/A _180_/Y vgnd vpwr scs8hd_inv_8
XANTENNA_mux_top_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_top_track_8.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_1_132 vpwr vgnd scs8hd_fill_2
XFILLER_1_165 vpwr vgnd scs8hd_fill_2
XFILLER_38_61 vgnd vpwr scs8hd_fill_1
XFILLER_1_198 vpwr vgnd scs8hd_fill_2
XFILLER_1_187 vpwr vgnd scs8hd_fill_2
XANTENNA__109__A _149_/D vgnd vpwr scs8hd_diode_2
XFILLER_9_254 vpwr vgnd scs8hd_fill_2
XFILLER_9_276 vgnd vpwr scs8hd_fill_1
XFILLER_39_191 vgnd vpwr scs8hd_decap_8
X_232_ _232_/A chanx_right_out[2] vgnd vpwr scs8hd_buf_2
XFILLER_6_235 vgnd vpwr scs8hd_fill_1
X_163_ _121_/Y _114_/A _163_/C _149_/D _165_/B vgnd vpwr scs8hd_or4_4
XFILLER_10_253 vgnd vpwr scs8hd_decap_12
XANTENNA__111__B _111_/B vgnd vpwr scs8hd_diode_2
XFILLER_1_67 vpwr vgnd scs8hd_fill_2
XFILLER_28_117 vgnd vpwr scs8hd_decap_6
XANTENNA_mux_right_track_12.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _202_/Y vgnd
+ vpwr scs8hd_diode_2
Xmux_right_track_12.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_right_track_12.INVTX1_1_.scs8hd_inv_1/Y
+ _203_/Y mux_right_track_12.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XFILLER_3_216 vgnd vpwr scs8hd_decap_12
XFILLER_10_32 vgnd vpwr scs8hd_decap_12
XFILLER_35_51 vgnd vpwr scs8hd_decap_8
XFILLER_19_96 vgnd vpwr scs8hd_fill_1
XFILLER_35_62 vgnd vpwr scs8hd_decap_12
X_215_ _215_/HI _215_/LO vgnd vpwr scs8hd_conb_1
XANTENNA__122__A _121_/Y vgnd vpwr scs8hd_diode_2
X_146_ address[3] _115_/B _149_/C _140_/D _147_/B vgnd vpwr scs8hd_or4_4
XFILLER_25_109 vgnd vpwr scs8hd_fill_1
XFILLER_18_183 vgnd vpwr scs8hd_fill_1
XANTENNA_mem_right_track_4.LATCH_1_.latch_SLEEPB _150_/Y vgnd vpwr scs8hd_diode_2
XFILLER_24_175 vgnd vpwr scs8hd_decap_8
XPHY_115 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_104 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_126 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_137 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_148 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__207__A _207_/A vgnd vpwr scs8hd_diode_2
XPHY_159 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_right_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_right_track_8.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XPHY_6 vgnd vpwr scs8hd_decap_3
XFILLER_30_178 vgnd vpwr scs8hd_decap_12
XANTENNA__117__A _128_/A vgnd vpwr scs8hd_diode_2
XFILLER_7_99 vpwr vgnd scs8hd_fill_2
X_129_ _096_/A _150_/A vgnd vpwr scs8hd_buf_1
XFILLER_21_112 vpwr vgnd scs8hd_fill_2
XFILLER_21_167 vgnd vpwr scs8hd_fill_1
XFILLER_21_189 vgnd vpwr scs8hd_decap_12
XFILLER_12_101 vpwr vgnd scs8hd_fill_2
XFILLER_16_64 vgnd vpwr scs8hd_decap_3
XFILLER_16_86 vpwr vgnd scs8hd_fill_2
XFILLER_12_167 vgnd vpwr scs8hd_decap_4
XFILLER_16_97 vpwr vgnd scs8hd_fill_2
XFILLER_37_19 vgnd vpwr scs8hd_decap_12
XFILLER_26_215 vgnd vpwr scs8hd_decap_12
Xmux_top_track_10.INVTX1_1_.scs8hd_inv_1 chanx_right_in[6] mux_top_track_10.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_40_251 vgnd vpwr scs8hd_decap_12
XFILLER_27_96 vgnd vpwr scs8hd_fill_1
XFILLER_4_152 vgnd vpwr scs8hd_fill_1
XANTENNA__130__A _123_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_14.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _204_/A vgnd
+ vpwr scs8hd_diode_2
XFILLER_16_270 vgnd vpwr scs8hd_decap_4
XFILLER_14_207 vgnd vpwr scs8hd_decap_6
XFILLER_13_87 vpwr vgnd scs8hd_fill_2
XFILLER_1_144 vpwr vgnd scs8hd_fill_2
XFILLER_8_3 vgnd vpwr scs8hd_decap_12
XFILLER_38_84 vpwr vgnd scs8hd_fill_2
Xmem_top_track_14.LATCH_1_.latch data_in _186_/A _135_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA__125__A _128_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_6.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _197_/Y vgnd vpwr
+ scs8hd_diode_2
XFILLER_39_170 vgnd vpwr scs8hd_decap_12
XFILLER_24_97 vpwr vgnd scs8hd_fill_2
X_231_ _231_/A chanx_right_out[3] vgnd vpwr scs8hd_buf_2
X_162_ _171_/C _162_/B _162_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_10_265 vgnd vpwr scs8hd_decap_8
XFILLER_10_276 vgnd vpwr scs8hd_fill_1
Xmem_right_track_10.LATCH_0_.latch data_in _201_/A _162_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mem_right_track_6.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_10.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A _218_/HI vgnd vpwr
+ scs8hd_diode_2
XFILLER_3_228 vgnd vpwr scs8hd_decap_12
XFILLER_10_44 vgnd vpwr scs8hd_decap_8
XFILLER_19_53 vpwr vgnd scs8hd_fill_2
XFILLER_35_74 vgnd vpwr scs8hd_fill_1
XFILLER_19_75 vpwr vgnd scs8hd_fill_2
XFILLER_42_187 vgnd vpwr scs8hd_decap_12
X_214_ _214_/HI _214_/LO vgnd vpwr scs8hd_conb_1
XFILLER_35_96 vgnd vpwr scs8hd_decap_8
Xmux_right_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 _208_/HI _190_/Y mux_right_track_0.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
X_145_ _151_/A _144_/B _145_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA_mux_top_track_14.INVTX1_0_.scs8hd_inv_1_A top_left_grid_pin_15_ vgnd vpwr
+ scs8hd_diode_2
XFILLER_33_132 vgnd vpwr scs8hd_decap_12
XFILLER_33_110 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_10.tap_buf4_0_.scs8hd_inv_1_A mux_right_track_10.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XPHY_105 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_116 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_154 vgnd vpwr scs8hd_decap_8
XPHY_127 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_138 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_149 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_21_21 vgnd vpwr scs8hd_decap_3
XFILLER_21_43 vgnd vpwr scs8hd_decap_8
XFILLER_21_54 vgnd vpwr scs8hd_decap_4
XPHY_7 vgnd vpwr scs8hd_decap_3
X_128_ _128_/A _128_/B _128_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_7_56 vgnd vpwr scs8hd_decap_4
XFILLER_7_89 vgnd vpwr scs8hd_decap_4
XANTENNA__133__A _151_/A vgnd vpwr scs8hd_diode_2
XANTENNA__117__B _116_/B vgnd vpwr scs8hd_diode_2
XFILLER_38_202 vgnd vpwr scs8hd_decap_12
XFILLER_23_3 vgnd vpwr scs8hd_decap_12
Xmux_top_track_10.tap_buf4_0_.scs8hd_inv_1 mux_top_track_10.tap_buf4_0_.scs8hd_inv_1/A
+ _238_/A vgnd vpwr scs8hd_inv_1
XFILLER_12_135 vpwr vgnd scs8hd_fill_2
XFILLER_16_32 vgnd vpwr scs8hd_decap_6
XANTENNA_mux_top_track_2.tap_buf4_0_.scs8hd_inv_1_A mux_top_track_2.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XANTENNA__128__A _128_/A vgnd vpwr scs8hd_diode_2
XFILLER_7_172 vpwr vgnd scs8hd_fill_2
XFILLER_41_208 vgnd vpwr scs8hd_decap_12
XFILLER_26_227 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _199_/A vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_top_track_4.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _176_/Y vgnd vpwr
+ scs8hd_diode_2
XFILLER_27_86 vpwr vgnd scs8hd_fill_2
XFILLER_27_20 vgnd vpwr scs8hd_decap_6
XFILLER_17_205 vgnd vpwr scs8hd_decap_12
XFILLER_40_263 vgnd vpwr scs8hd_decap_12
XFILLER_4_131 vgnd vpwr scs8hd_fill_1
XANTENNA__130__B _115_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_track_2.LATCH_0_.latch_SLEEPB _112_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_14.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_14.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_top_track_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_22_274 vgnd vpwr scs8hd_fill_1
XFILLER_13_66 vpwr vgnd scs8hd_fill_2
XFILLER_38_30 vgnd vpwr scs8hd_fill_1
XFILLER_1_101 vpwr vgnd scs8hd_fill_2
XANTENNA__231__A _231_/A vgnd vpwr scs8hd_diode_2
XANTENNA__125__B _124_/B vgnd vpwr scs8hd_diode_2
Xmem_right_track_6.LATCH_0_.latch data_in _197_/A _156_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_13_241 vgnd vpwr scs8hd_fill_1
XANTENNA__141__A _150_/A vgnd vpwr scs8hd_diode_2
XFILLER_39_182 vgnd vpwr scs8hd_fill_1
XFILLER_24_32 vgnd vpwr scs8hd_decap_6
X_230_ _230_/A chanx_right_out[4] vgnd vpwr scs8hd_buf_2
X_161_ _170_/C _162_/B _161_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_6_215 vgnd vpwr scs8hd_decap_12
XANTENNA__226__A _226_/A vgnd vpwr scs8hd_diode_2
XFILLER_40_97 vgnd vpwr scs8hd_fill_1
XFILLER_6_248 vgnd vpwr scs8hd_decap_8
XFILLER_6_259 vgnd vpwr scs8hd_decap_12
XFILLER_37_119 vgnd vpwr scs8hd_decap_3
XANTENNA__136__A _151_/A vgnd vpwr scs8hd_diode_2
XFILLER_36_141 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_10.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _182_/A vgnd vpwr
+ scs8hd_diode_2
XFILLER_10_89 vgnd vpwr scs8hd_decap_3
XFILLER_19_10 vgnd vpwr scs8hd_decap_12
XFILLER_19_43 vgnd vpwr scs8hd_decap_4
XFILLER_42_199 vgnd vpwr scs8hd_decap_12
X_213_ _213_/HI _213_/LO vgnd vpwr scs8hd_conb_1
X_144_ _150_/A _144_/B _144_/Y vgnd vpwr scs8hd_nor2_4
Xmux_right_track_2.tap_buf4_0_.scs8hd_inv_1 mux_right_track_2.tap_buf4_0_.scs8hd_inv_1/A
+ _233_/A vgnd vpwr scs8hd_inv_1
XFILLER_2_251 vgnd vpwr scs8hd_decap_12
XFILLER_18_141 vgnd vpwr scs8hd_fill_1
XFILLER_18_152 vgnd vpwr scs8hd_fill_1
XFILLER_18_163 vgnd vpwr scs8hd_decap_12
XFILLER_33_144 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_2.tap_buf4_0_.scs8hd_inv_1_A mux_right_track_2.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_track_0.LATCH_1_.latch_SLEEPB _105_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_6.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _178_/A vgnd vpwr
+ scs8hd_diode_2
XPHY_106 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_117 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_128 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_139 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_21_66 vgnd vpwr scs8hd_fill_1
XFILLER_21_99 vpwr vgnd scs8hd_fill_2
XPHY_8 vgnd vpwr scs8hd_decap_3
XFILLER_15_177 vgnd vpwr scs8hd_fill_1
X_127_ _127_/A _128_/B _127_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_7_68 vgnd vpwr scs8hd_decap_3
XANTENNA__133__B _133_/B vgnd vpwr scs8hd_diode_2
XFILLER_38_258 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_top_track_14.LATCH_0_.latch_SLEEPB _136_/Y vgnd vpwr scs8hd_diode_2
XFILLER_8_107 vpwr vgnd scs8hd_fill_2
XFILLER_32_43 vgnd vpwr scs8hd_decap_6
XFILLER_32_32 vgnd vpwr scs8hd_decap_8
XANTENNA__234__A _234_/A vgnd vpwr scs8hd_diode_2
XANTENNA__128__B _128_/B vgnd vpwr scs8hd_diode_2
XANTENNA__144__A _150_/A vgnd vpwr scs8hd_diode_2
XFILLER_7_184 vgnd vpwr scs8hd_decap_4
Xmux_top_track_14.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_top_track_14.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ _186_/A mux_top_track_14.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XFILLER_26_239 vgnd vpwr scs8hd_decap_12
Xmux_right_track_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_right_track_2.INVTX1_1_.scs8hd_inv_1/Y
+ _193_/Y mux_right_track_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XFILLER_27_43 vgnd vpwr scs8hd_decap_6
XANTENNA__229__A _229_/A vgnd vpwr scs8hd_diode_2
XFILLER_17_217 vgnd vpwr scs8hd_decap_12
XFILLER_4_187 vpwr vgnd scs8hd_fill_2
XFILLER_4_165 vgnd vpwr scs8hd_decap_8
XFILLER_4_69 vpwr vgnd scs8hd_fill_2
XANTENNA__130__C _134_/C vgnd vpwr scs8hd_diode_2
XFILLER_31_220 vgnd vpwr scs8hd_decap_12
XANTENNA__139__A _163_/C vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_track_14.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA__141__B _141_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_track_12.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_40_32 vgnd vpwr scs8hd_decap_12
XFILLER_24_66 vpwr vgnd scs8hd_fill_2
X_160_ _121_/Y _114_/A _163_/C _140_/D _162_/B vgnd vpwr scs8hd_or4_4
XFILLER_6_227 vgnd vpwr scs8hd_fill_1
XFILLER_6_238 vgnd vpwr scs8hd_fill_1
XANTENNA_mem_top_track_12.LATCH_1_.latch_SLEEPB _131_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_track_2.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA__242__A _242_/A vgnd vpwr scs8hd_diode_2
XFILLER_1_15 vgnd vpwr scs8hd_decap_12
XANTENNA__136__B _135_/B vgnd vpwr scs8hd_diode_2
XANTENNA__152__A _096_/A vgnd vpwr scs8hd_diode_2
Xmem_top_track_10.LATCH_1_.latch data_in _182_/A _127_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_10_68 vpwr vgnd scs8hd_fill_2
XFILLER_27_153 vgnd vpwr scs8hd_decap_12
XFILLER_19_88 vpwr vgnd scs8hd_fill_2
XFILLER_19_99 vpwr vgnd scs8hd_fill_2
XFILLER_42_156 vgnd vpwr scs8hd_decap_12
XANTENNA__237__A _237_/A vgnd vpwr scs8hd_diode_2
X_212_ _212_/HI _212_/LO vgnd vpwr scs8hd_conb_1
X_143_ _115_/A _123_/B _149_/C _149_/D _144_/B vgnd vpwr scs8hd_or4_4
XFILLER_2_263 vgnd vpwr scs8hd_decap_12
XFILLER_18_175 vgnd vpwr scs8hd_decap_8
XFILLER_18_186 vgnd vpwr scs8hd_decap_12
XFILLER_33_156 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_12.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A _210_/HI vgnd vpwr
+ scs8hd_diode_2
XANTENNA__147__A _150_/A vgnd vpwr scs8hd_diode_2
XFILLER_24_145 vpwr vgnd scs8hd_fill_2
XFILLER_24_101 vgnd vpwr scs8hd_fill_1
XPHY_107 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_118 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_129 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_21_78 vpwr vgnd scs8hd_fill_2
XPHY_9 vgnd vpwr scs8hd_decap_3
Xmux_right_track_10.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_right_track_10.INVTX1_1_.scs8hd_inv_1/Y
+ _201_/Y mux_right_track_10.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XFILLER_15_123 vpwr vgnd scs8hd_fill_2
XFILLER_15_145 vgnd vpwr scs8hd_decap_3
XFILLER_15_167 vpwr vgnd scs8hd_fill_2
X_126_ _123_/A _123_/B _123_/C _110_/D _128_/B vgnd vpwr scs8hd_or4_4
XFILLER_38_215 vgnd vpwr scs8hd_decap_12
XFILLER_30_6 vgnd vpwr scs8hd_decap_8
XFILLER_21_148 vpwr vgnd scs8hd_fill_2
XFILLER_29_248 vpwr vgnd scs8hd_fill_2
XFILLER_29_204 vgnd vpwr scs8hd_decap_12
XFILLER_8_119 vpwr vgnd scs8hd_fill_2
XFILLER_16_56 vpwr vgnd scs8hd_fill_2
XFILLER_16_78 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_14.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _205_/Y vgnd
+ vpwr scs8hd_diode_2
XFILLER_28_270 vgnd vpwr scs8hd_decap_4
XFILLER_7_130 vpwr vgnd scs8hd_fill_2
XANTENNA__144__B _144_/B vgnd vpwr scs8hd_diode_2
XANTENNA__160__A _121_/Y vgnd vpwr scs8hd_diode_2
X_109_ _149_/D _110_/D vgnd vpwr scs8hd_buf_1
XFILLER_34_251 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_14.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_top_track_14.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_27_11 vgnd vpwr scs8hd_decap_3
XFILLER_27_99 vpwr vgnd scs8hd_fill_2
XFILLER_27_55 vgnd vpwr scs8hd_decap_6
XFILLER_25_262 vgnd vpwr scs8hd_decap_12
XFILLER_17_229 vgnd vpwr scs8hd_decap_12
XFILLER_40_276 vgnd vpwr scs8hd_fill_1
XFILLER_4_199 vgnd vpwr scs8hd_decap_3
XFILLER_4_100 vgnd vpwr scs8hd_decap_4
XANTENNA__130__D _123_/D vgnd vpwr scs8hd_diode_2
XFILLER_31_232 vgnd vpwr scs8hd_decap_12
XANTENNA__155__A address[0] vgnd vpwr scs8hd_diode_2
XFILLER_16_251 vgnd vpwr scs8hd_decap_4
XFILLER_13_57 vpwr vgnd scs8hd_fill_2
XFILLER_22_276 vgnd vpwr scs8hd_fill_1
XFILLER_1_114 vpwr vgnd scs8hd_fill_2
XFILLER_1_136 vpwr vgnd scs8hd_fill_2
XFILLER_38_32 vgnd vpwr scs8hd_decap_12
XFILLER_1_169 vpwr vgnd scs8hd_fill_2
XFILLER_13_276 vgnd vpwr scs8hd_fill_1
XFILLER_9_258 vgnd vpwr scs8hd_decap_12
XFILLER_0_191 vpwr vgnd scs8hd_fill_2
XFILLER_24_23 vgnd vpwr scs8hd_decap_8
XFILLER_40_44 vgnd vpwr scs8hd_decap_12
XFILLER_10_213 vgnd vpwr scs8hd_fill_1
XFILLER_6_3 vgnd vpwr scs8hd_decap_12
Xmux_top_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_top_track_16.INVTX1_0_.scs8hd_inv_1/Y
+ _189_/A mux_top_track_16.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A vgnd vpwr scs8hd_ebufn_2
XFILLER_1_27 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_right_track_14.LATCH_0_.latch_SLEEPB _169_/Y vgnd vpwr scs8hd_diode_2
XFILLER_39_3 vgnd vpwr scs8hd_decap_8
XFILLER_36_154 vgnd vpwr scs8hd_decap_12
XFILLER_36_121 vpwr vgnd scs8hd_fill_2
Xmem_right_track_2.LATCH_0_.latch data_in _193_/A _148_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_27_165 vgnd vpwr scs8hd_decap_12
XFILLER_27_132 vpwr vgnd scs8hd_fill_2
XFILLER_42_168 vgnd vpwr scs8hd_decap_12
XFILLER_35_77 vgnd vpwr scs8hd_decap_12
X_211_ _211_/HI _211_/LO vgnd vpwr scs8hd_conb_1
X_142_ _151_/A _141_/B _142_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA_mux_right_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _207_/A vgnd
+ vpwr scs8hd_diode_2
XFILLER_33_168 vgnd vpwr scs8hd_decap_12
XFILLER_18_110 vgnd vpwr scs8hd_decap_6
XFILLER_18_198 vgnd vpwr scs8hd_decap_12
XANTENNA__147__B _147_/B vgnd vpwr scs8hd_diode_2
XANTENNA__163__A _121_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_2.INVTX1_0_.scs8hd_inv_1_A top_left_grid_pin_3_ vgnd vpwr scs8hd_diode_2
XFILLER_32_190 vgnd vpwr scs8hd_decap_12
XPHY_108 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_119 vgnd vpwr scs8hd_tapvpwrvgnd_1
X_125_ _128_/A _124_/B _125_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_7_15 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_6.INVTX1_1_.scs8hd_inv_1_A chanx_right_in[4] vgnd vpwr scs8hd_diode_2
XFILLER_11_90 vpwr vgnd scs8hd_fill_2
XFILLER_38_227 vgnd vpwr scs8hd_decap_12
XANTENNA__158__A _170_/C vgnd vpwr scs8hd_diode_2
XFILLER_21_116 vpwr vgnd scs8hd_fill_2
XFILLER_21_127 vgnd vpwr scs8hd_decap_4
XFILLER_29_216 vgnd vpwr scs8hd_decap_12
XFILLER_12_116 vgnd vpwr scs8hd_decap_8
XFILLER_12_149 vpwr vgnd scs8hd_fill_2
XFILLER_35_208 vgnd vpwr scs8hd_decap_12
X_108_ address[1] enable _149_/D vgnd vpwr scs8hd_nand2_4
XFILLER_11_193 vpwr vgnd scs8hd_fill_2
XANTENNA__160__B _114_/A vgnd vpwr scs8hd_diode_2
XFILLER_21_3 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_right_track_12.LATCH_1_.latch_SLEEPB _164_/Y vgnd vpwr scs8hd_diode_2
XFILLER_34_263 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_6.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _196_/Y vgnd vpwr
+ scs8hd_diode_2
Xmux_top_track_8.tap_buf4_0_.scs8hd_inv_1 mux_top_track_8.tap_buf4_0_.scs8hd_inv_1/A
+ _239_/A vgnd vpwr scs8hd_inv_1
XFILLER_8_80 vpwr vgnd scs8hd_fill_2
XFILLER_27_67 vpwr vgnd scs8hd_fill_2
XFILLER_25_274 vgnd vpwr scs8hd_decap_3
XFILLER_25_241 vgnd vpwr scs8hd_decap_3
XPHY_280 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_16_274 vgnd vpwr scs8hd_fill_1
XANTENNA__171__A _110_/D vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_track_8.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_1_148 vpwr vgnd scs8hd_fill_2
XFILLER_38_88 vgnd vpwr scs8hd_decap_4
XFILLER_38_55 vgnd vpwr scs8hd_decap_6
XFILLER_38_44 vpwr vgnd scs8hd_fill_2
XANTENNA__166__A address[3] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_10.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _183_/Y vgnd vpwr
+ scs8hd_diode_2
XFILLER_5_92 vgnd vpwr scs8hd_decap_3
XFILLER_40_56 vgnd vpwr scs8hd_fill_1
XFILLER_10_247 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_right_track_0.INVTX1_1_.scs8hd_inv_1_A right_top_grid_pin_10_ vgnd vpwr
+ scs8hd_diode_2
XFILLER_1_39 vgnd vpwr scs8hd_decap_12
XFILLER_5_262 vpwr vgnd scs8hd_fill_2
XFILLER_5_240 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_6.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _179_/Y vgnd vpwr
+ scs8hd_diode_2
XFILLER_36_166 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_12.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A _219_/HI vgnd vpwr
+ scs8hd_diode_2
XFILLER_10_15 vgnd vpwr scs8hd_decap_12
XFILLER_19_24 vpwr vgnd scs8hd_fill_2
XFILLER_42_125 vgnd vpwr scs8hd_decap_12
XFILLER_19_57 vpwr vgnd scs8hd_fill_2
XFILLER_35_89 vgnd vpwr scs8hd_decap_4
X_210_ _210_/HI _210_/LO vgnd vpwr scs8hd_conb_1
X_141_ _150_/A _141_/B _141_/Y vgnd vpwr scs8hd_nor2_4
Xmux_top_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_top_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ _180_/A mux_top_track_8.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XFILLER_2_276 vgnd vpwr scs8hd_fill_1
XFILLER_33_114 vpwr vgnd scs8hd_fill_2
XFILLER_18_144 vpwr vgnd scs8hd_fill_2
XANTENNA__163__B _114_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _198_/A vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mem_right_track_0.LATCH_0_.latch_SLEEPB _145_/Y vgnd vpwr scs8hd_diode_2
Xmem_right_track_14.LATCH_1_.latch data_in _204_/A _168_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_2_93 vgnd vpwr scs8hd_decap_8
XPHY_109 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_21_58 vgnd vpwr scs8hd_fill_1
XFILLER_15_114 vpwr vgnd scs8hd_fill_2
X_124_ _127_/A _124_/B _124_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_7_27 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_10.INVTX1_0_.scs8hd_inv_1_A chany_top_in[4] vgnd vpwr scs8hd_diode_2
XFILLER_38_239 vgnd vpwr scs8hd_decap_12
XANTENNA__158__B _159_/B vgnd vpwr scs8hd_diode_2
XANTENNA__174__A _174_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_14.INVTX1_1_.scs8hd_inv_1_A right_bottom_grid_pin_13_ vgnd
+ vpwr scs8hd_diode_2
XFILLER_29_228 vgnd vpwr scs8hd_decap_12
XFILLER_12_139 vgnd vpwr scs8hd_decap_8
X_107_ _128_/A _105_/B _107_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_7_143 vgnd vpwr scs8hd_decap_12
XFILLER_7_176 vgnd vpwr scs8hd_decap_4
XANTENNA__160__C _163_/C vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_12.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _185_/A vgnd vpwr
+ scs8hd_diode_2
XFILLER_14_3 vgnd vpwr scs8hd_decap_12
XANTENNA__169__A _123_/D vgnd vpwr scs8hd_diode_2
XFILLER_25_253 vpwr vgnd scs8hd_fill_2
XPHY_281 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_270 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_31_245 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _181_/A vgnd vpwr
+ scs8hd_diode_2
XANTENNA__171__B _171_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_16.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_13_15 vgnd vpwr scs8hd_decap_12
Xmux_top_track_12.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_top_track_12.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ _184_/A mux_top_track_12.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_top_track_4.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_top_track_4.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_38_67 vpwr vgnd scs8hd_fill_2
Xmux_right_track_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_right_track_0.INVTX1_1_.scs8hd_inv_1/Y
+ _191_/Y mux_right_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XFILLER_9_205 vgnd vpwr scs8hd_decap_12
XFILLER_13_245 vpwr vgnd scs8hd_fill_2
XFILLER_13_256 vgnd vpwr scs8hd_decap_12
XFILLER_0_182 vgnd vpwr scs8hd_decap_4
XANTENNA__166__B address[2] vgnd vpwr scs8hd_diode_2
XANTENNA__182__A _182_/A vgnd vpwr scs8hd_diode_2
XFILLER_39_142 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_top_track_0.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_10_215 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_6.INVTX1_0_.scs8hd_inv_1_A chany_top_in[2] vgnd vpwr scs8hd_diode_2
XFILLER_5_274 vgnd vpwr scs8hd_decap_3
XFILLER_36_178 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_right_track_10.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA__177__A _177_/A vgnd vpwr scs8hd_diode_2
XFILLER_10_27 vgnd vpwr scs8hd_decap_4
XFILLER_42_137 vgnd vpwr scs8hd_decap_12
X_140_ _115_/A _123_/B _149_/C _140_/D _141_/B vgnd vpwr scs8hd_or4_4
XFILLER_2_211 vgnd vpwr scs8hd_decap_3
Xmux_top_track_16.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 _221_/HI _188_/Y mux_top_track_16.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_18_123 vpwr vgnd scs8hd_fill_2
XFILLER_25_90 vpwr vgnd scs8hd_fill_2
XPHY_90 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__163__C _163_/C vgnd vpwr scs8hd_diode_2
XFILLER_2_61 vgnd vpwr scs8hd_fill_1
XFILLER_21_15 vgnd vpwr scs8hd_fill_1
XFILLER_21_26 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_4.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_4.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
Xmem_top_track_6.LATCH_0_.latch data_in _179_/A _120_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_30_107 vgnd vpwr scs8hd_decap_3
XFILLER_7_39 vgnd vpwr scs8hd_decap_12
X_123_ _123_/A _123_/B _123_/C _123_/D _124_/B vgnd vpwr scs8hd_or4_4
XFILLER_16_7 vgnd vpwr scs8hd_decap_12
XANTENNA__190__A _190_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_0.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_28_251 vgnd vpwr scs8hd_decap_4
XANTENNA__160__D _140_/D vgnd vpwr scs8hd_diode_2
XFILLER_7_199 vpwr vgnd scs8hd_fill_2
X_106_ address[0] _128_/A vgnd vpwr scs8hd_buf_1
XFILLER_22_80 vgnd vpwr scs8hd_decap_6
XANTENNA__169__B _171_/B vgnd vpwr scs8hd_diode_2
XFILLER_34_276 vgnd vpwr scs8hd_fill_1
XANTENNA__185__A _185_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_14.tap_buf4_0_.scs8hd_inv_1_A mux_top_track_14.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_25_221 vgnd vpwr scs8hd_decap_12
XFILLER_40_202 vgnd vpwr scs8hd_decap_12
XANTENNA__095__A address[0] vgnd vpwr scs8hd_diode_2
XFILLER_4_136 vpwr vgnd scs8hd_fill_2
XFILLER_4_18 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_top_track_14.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_16_276 vgnd vpwr scs8hd_fill_1
XPHY_282 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_271 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_260 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_31_257 vgnd vpwr scs8hd_decap_12
XFILLER_3_191 vgnd vpwr scs8hd_decap_8
XANTENNA__171__C _171_/C vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_track_4.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_13_27 vgnd vpwr scs8hd_decap_12
XFILLER_13_49 vpwr vgnd scs8hd_fill_2
XFILLER_9_217 vgnd vpwr scs8hd_decap_12
XFILLER_13_268 vgnd vpwr scs8hd_decap_8
Xmux_right_track_8.INVTX1_0_.scs8hd_inv_1 chany_top_in[3] mux_right_track_8.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA__166__C address[4] vgnd vpwr scs8hd_diode_2
XFILLER_39_121 vgnd vpwr scs8hd_fill_1
XFILLER_39_187 vpwr vgnd scs8hd_fill_2
XFILLER_24_15 vgnd vpwr scs8hd_decap_4
XFILLER_10_205 vgnd vpwr scs8hd_decap_8
XFILLER_10_227 vgnd vpwr scs8hd_decap_12
XFILLER_14_81 vpwr vgnd scs8hd_fill_2
XFILLER_30_91 vgnd vpwr scs8hd_fill_1
XFILLER_36_113 vgnd vpwr scs8hd_decap_8
XANTENNA__193__A _193_/A vgnd vpwr scs8hd_diode_2
XFILLER_42_149 vgnd vpwr scs8hd_decap_6
XFILLER_27_179 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_14.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _204_/Y vgnd
+ vpwr scs8hd_diode_2
XFILLER_18_102 vpwr vgnd scs8hd_fill_2
XFILLER_41_171 vgnd vpwr scs8hd_decap_12
XPHY_80 vgnd vpwr scs8hd_decap_3
XPHY_91 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmux_top_track_14.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_top_track_14.INVTX1_0_.scs8hd_inv_1/Y
+ _187_/A mux_top_track_14.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
X_199_ _199_/A _199_/Y vgnd vpwr scs8hd_inv_8
XANTENNA__163__D _149_/D vgnd vpwr scs8hd_diode_2
XFILLER_37_3 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_14.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A _211_/HI vgnd vpwr
+ scs8hd_diode_2
XANTENNA__188__A _188_/A vgnd vpwr scs8hd_diode_2
XFILLER_24_149 vgnd vpwr scs8hd_decap_4
XFILLER_24_116 vgnd vpwr scs8hd_decap_12
XFILLER_24_105 vgnd vpwr scs8hd_decap_8
XANTENNA__098__A address[2] vgnd vpwr scs8hd_diode_2
XFILLER_15_127 vgnd vpwr scs8hd_decap_3
XFILLER_23_193 vpwr vgnd scs8hd_fill_2
X_122_ _121_/Y _123_/A vgnd vpwr scs8hd_buf_1
XANTENNA_mux_right_track_10.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_right_track_10.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_32_15 vgnd vpwr scs8hd_decap_12
Xmem_right_track_10.LATCH_1_.latch data_in _200_/A _161_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_20_152 vgnd vpwr scs8hd_fill_1
XFILLER_20_163 vgnd vpwr scs8hd_decap_12
XFILLER_28_274 vgnd vpwr scs8hd_fill_1
X_105_ _127_/A _105_/B _105_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_11_163 vpwr vgnd scs8hd_fill_2
XANTENNA__169__C _171_/C vgnd vpwr scs8hd_diode_2
XFILLER_25_233 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_top_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_top_track_16.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_4_104 vgnd vpwr scs8hd_fill_1
XPHY_261 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_250 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_16_211 vgnd vpwr scs8hd_decap_3
XFILLER_17_92 vgnd vpwr scs8hd_fill_1
XPHY_283 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_272 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_31_269 vgnd vpwr scs8hd_decap_8
XANTENNA__196__A _196_/A vgnd vpwr scs8hd_diode_2
XFILLER_13_39 vgnd vpwr scs8hd_decap_8
XFILLER_22_247 vpwr vgnd scs8hd_fill_2
XFILLER_22_258 vgnd vpwr scs8hd_decap_12
XFILLER_1_118 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_16.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _206_/A vgnd
+ vpwr scs8hd_diode_2
XFILLER_9_229 vgnd vpwr scs8hd_decap_12
XFILLER_0_151 vpwr vgnd scs8hd_fill_2
XFILLER_0_195 vgnd vpwr scs8hd_decap_4
XFILLER_0_173 vpwr vgnd scs8hd_fill_2
XANTENNA__166__D _166_/D vgnd vpwr scs8hd_diode_2
XFILLER_5_73 vgnd vpwr scs8hd_decap_4
XFILLER_5_51 vgnd vpwr scs8hd_decap_4
XFILLER_8_262 vgnd vpwr scs8hd_decap_12
XFILLER_24_49 vgnd vpwr scs8hd_decap_8
XFILLER_40_15 vgnd vpwr scs8hd_decap_12
XFILLER_10_239 vgnd vpwr scs8hd_decap_6
XANTENNA_mux_top_track_10.INVTX1_0_.scs8hd_inv_1_A top_left_grid_pin_11_ vgnd vpwr
+ scs8hd_diode_2
XFILLER_14_71 vgnd vpwr scs8hd_fill_1
XFILLER_30_81 vpwr vgnd scs8hd_fill_2
XFILLER_5_221 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _199_/Y vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mem_right_track_4.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_36_125 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_top_track_14.INVTX1_1_.scs8hd_inv_1_A chanx_right_in[8] vgnd vpwr scs8hd_diode_2
XFILLER_35_15 vgnd vpwr scs8hd_decap_12
XFILLER_27_136 vpwr vgnd scs8hd_fill_2
XFILLER_27_114 vgnd vpwr scs8hd_decap_6
Xmux_right_track_6.INVTX1_0_.scs8hd_inv_1 chany_top_in[2] mux_right_track_6.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_19_49 vpwr vgnd scs8hd_fill_2
XFILLER_42_106 vgnd vpwr scs8hd_decap_12
XFILLER_35_180 vgnd vpwr scs8hd_decap_3
XFILLER_35_59 vpwr vgnd scs8hd_fill_2
XFILLER_33_106 vpwr vgnd scs8hd_fill_2
XFILLER_26_191 vgnd vpwr scs8hd_decap_4
XPHY_81 vgnd vpwr scs8hd_decap_3
XPHY_70 vgnd vpwr scs8hd_decap_3
XPHY_92 vgnd vpwr scs8hd_tapvpwrvgnd_1
X_198_ _198_/A _198_/Y vgnd vpwr scs8hd_inv_8
XFILLER_24_128 vgnd vpwr scs8hd_decap_8
Xmem_right_track_6.LATCH_1_.latch data_in _196_/A _154_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
X_121_ address[3] _121_/Y vgnd vpwr scs8hd_inv_8
XFILLER_14_183 vgnd vpwr scs8hd_decap_12
Xmux_top_track_6.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_top_track_6.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ _178_/A mux_top_track_6.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XANTENNA__199__A _199_/A vgnd vpwr scs8hd_diode_2
XFILLER_37_253 vpwr vgnd scs8hd_fill_2
XFILLER_37_220 vgnd vpwr scs8hd_decap_12
XFILLER_32_27 vgnd vpwr scs8hd_decap_4
XFILLER_20_175 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_right_track_8.LATCH_1_.latch_SLEEPB _158_/Y vgnd vpwr scs8hd_diode_2
XFILLER_7_168 vpwr vgnd scs8hd_fill_2
XFILLER_11_175 vpwr vgnd scs8hd_fill_2
XFILLER_11_197 vpwr vgnd scs8hd_fill_2
X_104_ _115_/A _123_/B _123_/C _123_/D _105_/B vgnd vpwr scs8hd_or4_4
Xmem_top_track_2.LATCH_0_.latch data_in _175_/A _112_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_top_track_10.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _182_/Y vgnd vpwr
+ scs8hd_diode_2
XFILLER_19_220 vgnd vpwr scs8hd_decap_12
XFILLER_21_7 vgnd vpwr scs8hd_decap_8
XFILLER_8_84 vgnd vpwr scs8hd_decap_8
XFILLER_27_16 vpwr vgnd scs8hd_fill_2
XFILLER_40_215 vgnd vpwr scs8hd_decap_12
XFILLER_25_245 vgnd vpwr scs8hd_decap_8
XPHY_284 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_273 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_262 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_251 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_240 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_17_71 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_6.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _178_/Y vgnd vpwr
+ scs8hd_diode_2
XFILLER_3_182 vgnd vpwr scs8hd_fill_1
XFILLER_3_160 vgnd vpwr scs8hd_decap_3
XFILLER_22_215 vgnd vpwr scs8hd_decap_12
XFILLER_8_274 vgnd vpwr scs8hd_fill_1
XFILLER_39_123 vgnd vpwr scs8hd_decap_12
XFILLER_40_27 vgnd vpwr scs8hd_decap_4
Xmux_top_track_10.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_top_track_10.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ _182_/A mux_top_track_10.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XFILLER_30_93 vgnd vpwr scs8hd_decap_12
XFILLER_30_71 vgnd vpwr scs8hd_fill_1
XFILLER_5_266 vgnd vpwr scs8hd_decap_8
XFILLER_19_28 vpwr vgnd scs8hd_fill_2
XFILLER_42_118 vgnd vpwr scs8hd_decap_6
XFILLER_35_27 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_14.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A _220_/HI vgnd vpwr
+ scs8hd_diode_2
XFILLER_2_203 vgnd vpwr scs8hd_decap_8
Xmux_right_track_14.tap_buf4_0_.scs8hd_inv_1 mux_right_track_14.tap_buf4_0_.scs8hd_inv_1/A
+ _227_/A vgnd vpwr scs8hd_inv_1
XANTENNA_mux_right_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _191_/A vgnd vpwr
+ scs8hd_diode_2
XPHY_82 vgnd vpwr scs8hd_decap_3
XPHY_71 vgnd vpwr scs8hd_decap_3
XFILLER_33_118 vpwr vgnd scs8hd_fill_2
XPHY_60 vgnd vpwr scs8hd_decap_3
XFILLER_25_60 vgnd vpwr scs8hd_fill_1
XFILLER_18_137 vgnd vpwr scs8hd_decap_4
XFILLER_18_148 vgnd vpwr scs8hd_decap_4
XFILLER_41_184 vgnd vpwr scs8hd_decap_12
XFILLER_25_82 vpwr vgnd scs8hd_fill_2
X_197_ _197_/A _197_/Y vgnd vpwr scs8hd_inv_8
XPHY_93 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_top_track_12.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _184_/A vgnd vpwr
+ scs8hd_diode_2
Xmux_top_track_16.tap_buf4_0_.scs8hd_inv_1 mux_top_track_16.tap_buf4_0_.scs8hd_inv_1/A
+ _235_/A vgnd vpwr scs8hd_inv_1
XFILLER_2_64 vgnd vpwr scs8hd_decap_12
XFILLER_17_170 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_top_track_10.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_top_track_10.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_15_118 vpwr vgnd scs8hd_fill_2
X_120_ _128_/A _119_/B _120_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_23_151 vgnd vpwr scs8hd_decap_6
Xmux_right_track_4.INVTX1_0_.scs8hd_inv_1 chany_top_in[1] mux_right_track_4.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_11_62 vpwr vgnd scs8hd_fill_2
XFILLER_11_73 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _180_/A vgnd vpwr
+ scs8hd_diode_2
XFILLER_14_195 vgnd vpwr scs8hd_decap_12
Xmux_top_track_14.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 _220_/HI _186_/Y mux_top_track_14.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_42_3 vgnd vpwr scs8hd_decap_12
XFILLER_37_232 vgnd vpwr scs8hd_decap_12
XFILLER_20_110 vgnd vpwr scs8hd_decap_6
XFILLER_20_187 vgnd vpwr scs8hd_decap_12
XFILLER_28_276 vgnd vpwr scs8hd_fill_1
XFILLER_11_132 vpwr vgnd scs8hd_fill_2
XFILLER_7_103 vpwr vgnd scs8hd_fill_2
XFILLER_7_114 vpwr vgnd scs8hd_fill_2
X_103_ _140_/D _123_/D vgnd vpwr scs8hd_buf_1
XFILLER_22_61 vgnd vpwr scs8hd_decap_6
XFILLER_34_202 vgnd vpwr scs8hd_decap_12
XFILLER_19_232 vgnd vpwr scs8hd_decap_12
XFILLER_8_52 vpwr vgnd scs8hd_fill_2
XFILLER_8_63 vpwr vgnd scs8hd_fill_2
XFILLER_27_39 vpwr vgnd scs8hd_fill_2
XFILLER_40_227 vgnd vpwr scs8hd_decap_12
XPHY_285 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_274 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_263 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_252 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_241 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_33_93 vpwr vgnd scs8hd_fill_2
XPHY_230 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_22_227 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_6.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_top_track_6.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_13_205 vgnd vpwr scs8hd_decap_12
Xmux_top_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_top_track_8.INVTX1_0_.scs8hd_inv_1/Y
+ _181_/A mux_top_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XANTENNA_mem_right_track_12.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_0_120 vpwr vgnd scs8hd_fill_2
XFILLER_28_93 vgnd vpwr scs8hd_decap_8
XFILLER_28_60 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_top_track_10.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_5_97 vgnd vpwr scs8hd_fill_1
XFILLER_39_146 vgnd vpwr scs8hd_decap_12
XFILLER_39_135 vgnd vpwr scs8hd_decap_3
XANTENNA_mem_top_track_6.LATCH_0_.latch_SLEEPB _120_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_track_0.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_top_track_2.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_38_190 vgnd vpwr scs8hd_decap_12
Xmux_right_track_8.tap_buf4_0_.scs8hd_inv_1 mux_right_track_8.tap_buf4_0_.scs8hd_inv_1/A
+ _230_/A vgnd vpwr scs8hd_inv_1
XFILLER_5_245 vpwr vgnd scs8hd_fill_2
XFILLER_36_105 vgnd vpwr scs8hd_decap_4
XANTENNA__101__A enable vgnd vpwr scs8hd_diode_2
XFILLER_35_160 vgnd vpwr scs8hd_decap_12
XFILLER_35_39 vgnd vpwr scs8hd_decap_12
XFILLER_27_149 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_14.tap_buf4_0_.scs8hd_inv_1_A mux_right_track_14.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_4_6 vgnd vpwr scs8hd_decap_12
XFILLER_2_215 vgnd vpwr scs8hd_decap_12
XFILLER_18_127 vgnd vpwr scs8hd_fill_1
XPHY_83 vgnd vpwr scs8hd_decap_3
XPHY_72 vgnd vpwr scs8hd_decap_3
XPHY_61 vgnd vpwr scs8hd_decap_3
XPHY_50 vgnd vpwr scs8hd_decap_3
XPHY_94 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_41_196 vgnd vpwr scs8hd_decap_12
X_196_ _196_/A _196_/Y vgnd vpwr scs8hd_inv_8
Xmux_top_track_16.INVTX1_0_.scs8hd_inv_1 top_right_grid_pin_11_ mux_top_track_16.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_2_32 vgnd vpwr scs8hd_decap_12
XFILLER_2_76 vgnd vpwr scs8hd_decap_12
XFILLER_32_152 vgnd vpwr scs8hd_fill_1
XFILLER_17_193 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_6.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_6.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_23_174 vpwr vgnd scs8hd_fill_2
XFILLER_11_41 vgnd vpwr scs8hd_decap_12
XFILLER_2_3 vgnd vpwr scs8hd_decap_12
XFILLER_36_60 vpwr vgnd scs8hd_fill_2
XFILLER_36_93 vgnd vpwr scs8hd_decap_12
XFILLER_14_152 vgnd vpwr scs8hd_fill_1
X_179_ _179_/A _179_/Y vgnd vpwr scs8hd_inv_8
XFILLER_35_3 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_6.tap_buf4_0_.scs8hd_inv_1_A mux_top_track_6.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_16_19 vgnd vpwr scs8hd_decap_12
Xmux_top_track_12.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_top_track_12.INVTX1_0_.scs8hd_inv_1/Y
+ _185_/A mux_top_track_12.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XFILLER_20_133 vpwr vgnd scs8hd_fill_2
XFILLER_20_144 vgnd vpwr scs8hd_decap_8
XFILLER_20_199 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_2.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_28_200 vgnd vpwr scs8hd_decap_12
Xmem_right_track_2.LATCH_1_.latch data_in _192_/A _147_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
X_102_ address[1] _102_/B _140_/D vgnd vpwr scs8hd_or2_4
XFILLER_7_126 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_top_track_4.LATCH_1_.latch_SLEEPB _116_/Y vgnd vpwr scs8hd_diode_2
Xmux_right_track_2.INVTX1_0_.scs8hd_inv_1 chany_top_in[0] mux_right_track_2.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_6_181 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_right_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _207_/Y vgnd
+ vpwr scs8hd_diode_2
XFILLER_40_239 vgnd vpwr scs8hd_decap_12
XFILLER_25_258 vpwr vgnd scs8hd_fill_2
XFILLER_4_107 vgnd vpwr scs8hd_fill_1
XFILLER_16_258 vgnd vpwr scs8hd_decap_12
XFILLER_17_51 vgnd vpwr scs8hd_decap_4
XFILLER_17_95 vgnd vpwr scs8hd_fill_1
XPHY_275 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_264 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_253 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_242 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_231 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_220 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__104__A _115_/A vgnd vpwr scs8hd_diode_2
XFILLER_22_239 vgnd vpwr scs8hd_decap_8
XFILLER_13_217 vgnd vpwr scs8hd_decap_12
Xmux_top_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_top_track_16.INVTX1_1_.scs8hd_inv_1/Y
+ _189_/Y mux_top_track_16.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A vgnd vpwr scs8hd_ebufn_2
XFILLER_0_165 vgnd vpwr scs8hd_decap_8
XFILLER_8_276 vgnd vpwr scs8hd_fill_1
XFILLER_39_158 vgnd vpwr scs8hd_decap_12
XFILLER_24_19 vgnd vpwr scs8hd_fill_1
XFILLER_14_52 vgnd vpwr scs8hd_decap_3
XFILLER_14_85 vpwr vgnd scs8hd_fill_2
XFILLER_39_71 vpwr vgnd scs8hd_fill_2
XFILLER_29_180 vgnd vpwr scs8hd_decap_3
XFILLER_35_172 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_top_track_2.INVTX1_1_.scs8hd_inv_1_A chanx_right_in[2] vgnd vpwr scs8hd_diode_2
XFILLER_2_227 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_6.tap_buf4_0_.scs8hd_inv_1_A mux_right_track_6.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XANTENNA__202__A _202_/A vgnd vpwr scs8hd_diode_2
Xmux_top_track_8.INVTX1_1_.scs8hd_inv_1 chanx_right_in[5] mux_top_track_8.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_18_106 vpwr vgnd scs8hd_fill_2
XPHY_84 vgnd vpwr scs8hd_decap_3
XPHY_73 vgnd vpwr scs8hd_decap_3
XPHY_62 vgnd vpwr scs8hd_decap_3
XPHY_51 vgnd vpwr scs8hd_decap_3
XFILLER_25_62 vgnd vpwr scs8hd_decap_4
XPHY_95 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_40 vgnd vpwr scs8hd_decap_3
X_195_ _195_/A _195_/Y vgnd vpwr scs8hd_inv_8
XFILLER_37_7 vgnd vpwr scs8hd_decap_12
XFILLER_2_55 vgnd vpwr scs8hd_decap_6
XFILLER_2_44 vgnd vpwr scs8hd_decap_8
XANTENNA__112__A _128_/A vgnd vpwr scs8hd_diode_2
XFILLER_2_88 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_right_track_16.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A _212_/HI vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mem_top_track_16.LATCH_1_.latch_SLEEPB _141_/Y vgnd vpwr scs8hd_diode_2
Xmem_top_track_16.LATCH_0_.latch data_in _189_/A _142_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_23_197 vpwr vgnd scs8hd_fill_2
XFILLER_11_86 vpwr vgnd scs8hd_fill_2
XFILLER_11_97 vpwr vgnd scs8hd_fill_2
XFILLER_36_72 vgnd vpwr scs8hd_fill_1
XANTENNA__107__A _128_/A vgnd vpwr scs8hd_diode_2
XFILLER_14_164 vgnd vpwr scs8hd_decap_8
Xmux_top_track_4.tap_buf4_0_.scs8hd_inv_1 mux_top_track_4.tap_buf4_0_.scs8hd_inv_1/A
+ _241_/A vgnd vpwr scs8hd_inv_1
X_178_ _178_/A _178_/Y vgnd vpwr scs8hd_inv_8
XFILLER_37_245 vgnd vpwr scs8hd_decap_8
XFILLER_28_3 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_12.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_right_track_12.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xmux_top_track_14.INVTX1_0_.scs8hd_inv_1 top_left_grid_pin_15_ mux_top_track_14.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_top_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A _217_/HI vgnd vpwr
+ scs8hd_diode_2
XFILLER_28_212 vpwr vgnd scs8hd_fill_2
X_101_ enable _102_/B vgnd vpwr scs8hd_inv_8
XFILLER_11_101 vpwr vgnd scs8hd_fill_2
XFILLER_11_145 vpwr vgnd scs8hd_fill_2
XFILLER_11_167 vgnd vpwr scs8hd_decap_3
XFILLER_22_41 vpwr vgnd scs8hd_fill_2
XFILLER_19_245 vgnd vpwr scs8hd_decap_12
XFILLER_34_215 vgnd vpwr scs8hd_decap_12
XFILLER_8_32 vgnd vpwr scs8hd_decap_12
XFILLER_4_119 vgnd vpwr scs8hd_decap_12
Xmux_top_track_4.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_top_track_4.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ _176_/A mux_top_track_4.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XPHY_243 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_232 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_221 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_210 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_right_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _198_/Y vgnd vpwr
+ scs8hd_diode_2
XFILLER_16_215 vgnd vpwr scs8hd_decap_12
XPHY_276 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_265 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_254 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_33_62 vgnd vpwr scs8hd_decap_4
XFILLER_33_51 vgnd vpwr scs8hd_decap_8
XFILLER_3_174 vpwr vgnd scs8hd_fill_2
XANTENNA__104__B _123_/B vgnd vpwr scs8hd_diode_2
XANTENNA__120__A _128_/A vgnd vpwr scs8hd_diode_2
XFILLER_30_251 vgnd vpwr scs8hd_decap_12
XFILLER_38_18 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_right_track_6.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_13_229 vgnd vpwr scs8hd_decap_12
Xmux_right_track_0.INVTX1_0_.scs8hd_inv_1 chany_top_in[8] mux_right_track_0.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_21_251 vpwr vgnd scs8hd_fill_2
XANTENNA__205__A _205_/A vgnd vpwr scs8hd_diode_2
XFILLER_28_84 vgnd vpwr scs8hd_decap_8
XANTENNA__115__A _115_/A vgnd vpwr scs8hd_diode_2
XFILLER_5_88 vpwr vgnd scs8hd_fill_2
XFILLER_10_3 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A _208_/HI vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_top_track_12.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _185_/Y vgnd vpwr
+ scs8hd_diode_2
XFILLER_30_30 vgnd vpwr scs8hd_fill_1
XFILLER_5_258 vpwr vgnd scs8hd_fill_2
XFILLER_5_236 vpwr vgnd scs8hd_fill_2
XFILLER_14_64 vgnd vpwr scs8hd_decap_4
Xmux_top_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 _225_/HI _180_/Y mux_top_track_8.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_30_85 vgnd vpwr scs8hd_decap_6
XFILLER_36_129 vgnd vpwr scs8hd_decap_12
XFILLER_29_192 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_8.INVTX1_0_.scs8hd_inv_1_A top_left_grid_pin_9_ vgnd vpwr scs8hd_diode_2
XFILLER_35_184 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _181_/Y vgnd vpwr
+ scs8hd_diode_2
XFILLER_2_239 vgnd vpwr scs8hd_decap_12
XPHY_30 vgnd vpwr scs8hd_decap_3
XPHY_85 vgnd vpwr scs8hd_decap_3
XFILLER_41_110 vgnd vpwr scs8hd_decap_12
XPHY_74 vgnd vpwr scs8hd_decap_3
XPHY_63 vgnd vpwr scs8hd_decap_3
XPHY_52 vgnd vpwr scs8hd_decap_3
XFILLER_25_52 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_10.INVTX1_1_.scs8hd_inv_1_A right_bottom_grid_pin_9_ vgnd
+ vpwr scs8hd_diode_2
XPHY_96 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_41 vgnd vpwr scs8hd_decap_3
XFILLER_41_62 vgnd vpwr scs8hd_decap_12
XFILLER_41_51 vgnd vpwr scs8hd_decap_8
X_194_ _194_/A _194_/Y vgnd vpwr scs8hd_inv_8
XANTENNA__112__B _111_/B vgnd vpwr scs8hd_diode_2
XFILLER_32_154 vgnd vpwr scs8hd_decap_12
XFILLER_32_132 vgnd vpwr scs8hd_decap_12
XFILLER_23_132 vpwr vgnd scs8hd_fill_2
XFILLER_36_84 vpwr vgnd scs8hd_fill_2
XFILLER_14_121 vpwr vgnd scs8hd_fill_2
XFILLER_14_154 vgnd vpwr scs8hd_fill_1
XANTENNA__107__B _105_/B vgnd vpwr scs8hd_diode_2
X_177_ _177_/A _177_/Y vgnd vpwr scs8hd_inv_8
Xmux_top_track_6.INVTX1_1_.scs8hd_inv_1 chanx_right_in[4] mux_top_track_6.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA__123__A _123_/A vgnd vpwr scs8hd_diode_2
XFILLER_37_257 vgnd vpwr scs8hd_decap_12
XFILLER_11_179 vpwr vgnd scs8hd_fill_2
X_100_ _134_/C _123_/C vgnd vpwr scs8hd_buf_1
XFILLER_19_257 vgnd vpwr scs8hd_decap_12
XFILLER_34_227 vgnd vpwr scs8hd_decap_12
XANTENNA__118__A _115_/A vgnd vpwr scs8hd_diode_2
X_229_ _229_/A chanx_right_out[5] vgnd vpwr scs8hd_buf_2
XFILLER_8_44 vgnd vpwr scs8hd_decap_8
XFILLER_40_3 vgnd vpwr scs8hd_decap_12
Xmux_top_track_12.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 _219_/HI _184_/Y mux_top_track_12.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_top_track_14.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _187_/A vgnd vpwr
+ scs8hd_diode_2
XPHY_277 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_266 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmux_top_track_12.INVTX1_0_.scs8hd_inv_1 top_left_grid_pin_13_ mux_top_track_12.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XPHY_255 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_244 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_233 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_31_208 vgnd vpwr scs8hd_decap_12
XPHY_222 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_211 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_271 vgnd vpwr scs8hd_decap_4
XPHY_200 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_16_227 vgnd vpwr scs8hd_decap_12
XFILLER_17_75 vpwr vgnd scs8hd_fill_2
Xmem_top_track_6.LATCH_1_.latch data_in _178_/A _119_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_3_142 vgnd vpwr scs8hd_fill_1
XANTENNA__104__C _123_/C vgnd vpwr scs8hd_diode_2
XANTENNA__120__B _119_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_2.INVTX1_0_.scs8hd_inv_1_A chany_top_in[0] vgnd vpwr scs8hd_diode_2
XFILLER_12_7 vgnd vpwr scs8hd_decap_8
XFILLER_30_263 vgnd vpwr scs8hd_decap_12
XFILLER_22_208 vgnd vpwr scs8hd_decap_6
XANTENNA_mux_right_track_6.INVTX1_1_.scs8hd_inv_1_A right_bottom_grid_pin_5_ vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mux_right_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _190_/A vgnd vpwr
+ scs8hd_diode_2
XFILLER_0_134 vpwr vgnd scs8hd_fill_2
XFILLER_0_178 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_right_track_16.LATCH_1_.latch_SLEEPB _170_/Y vgnd vpwr scs8hd_diode_2
XFILLER_28_74 vgnd vpwr scs8hd_fill_1
XFILLER_28_41 vgnd vpwr scs8hd_decap_3
XFILLER_8_245 vpwr vgnd scs8hd_fill_2
XANTENNA__115__B _115_/B vgnd vpwr scs8hd_diode_2
XFILLER_39_105 vpwr vgnd scs8hd_fill_2
XANTENNA__131__A _150_/A vgnd vpwr scs8hd_diode_2
Xmux_right_track_16.INVTX1_1_.scs8hd_inv_1 right_bottom_grid_pin_15_ mux_right_track_16.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_14_32 vgnd vpwr scs8hd_decap_12
XFILLER_39_40 vgnd vpwr scs8hd_decap_12
Xmux_top_track_6.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_top_track_6.INVTX1_0_.scs8hd_inv_1/Y
+ _179_/A mux_top_track_6.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XANTENNA__126__A _123_/A vgnd vpwr scs8hd_diode_2
XFILLER_35_196 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_16.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A _221_/HI vgnd vpwr
+ scs8hd_diode_2
XPHY_64 vgnd vpwr scs8hd_decap_3
XPHY_53 vgnd vpwr scs8hd_decap_3
XFILLER_25_31 vgnd vpwr scs8hd_decap_6
XANTENNA_mux_right_track_16.INVTX1_0_.scs8hd_inv_1_A chany_top_in[7] vgnd vpwr scs8hd_diode_2
XPHY_20 vgnd vpwr scs8hd_decap_3
XPHY_31 vgnd vpwr scs8hd_decap_3
XFILLER_18_119 vpwr vgnd scs8hd_fill_2
XPHY_42 vgnd vpwr scs8hd_decap_3
XFILLER_41_74 vgnd vpwr scs8hd_decap_12
XPHY_75 vgnd vpwr scs8hd_decap_3
XFILLER_25_86 vpwr vgnd scs8hd_fill_2
X_193_ _193_/A _193_/Y vgnd vpwr scs8hd_inv_8
XPHY_97 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_86 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_32_166 vgnd vpwr scs8hd_decap_12
XFILLER_32_144 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_top_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _173_/A vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_top_track_12.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_top_track_12.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_11_55 vgnd vpwr scs8hd_decap_4
XFILLER_14_144 vgnd vpwr scs8hd_decap_8
X_176_ _176_/A _176_/Y vgnd vpwr scs8hd_inv_8
XANTENNA__123__B _123_/B vgnd vpwr scs8hd_diode_2
XFILLER_37_269 vgnd vpwr scs8hd_decap_8
XFILLER_28_258 vgnd vpwr scs8hd_decap_12
XFILLER_11_114 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_right_track_4.LATCH_0_.latch_SLEEPB _151_/Y vgnd vpwr scs8hd_diode_2
XFILLER_7_118 vpwr vgnd scs8hd_fill_2
XFILLER_11_136 vgnd vpwr scs8hd_decap_6
XFILLER_0_3 vgnd vpwr scs8hd_decap_12
Xmem_top_track_12.LATCH_0_.latch data_in _185_/A _133_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_34_239 vgnd vpwr scs8hd_decap_12
XFILLER_19_269 vgnd vpwr scs8hd_decap_8
XFILLER_42_261 vgnd vpwr scs8hd_decap_12
XFILLER_8_67 vpwr vgnd scs8hd_fill_2
XANTENNA__118__B _115_/B vgnd vpwr scs8hd_diode_2
X_228_ _228_/A chanx_right_out[6] vgnd vpwr scs8hd_buf_2
X_159_ _171_/C _159_/B _159_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_6_195 vpwr vgnd scs8hd_fill_2
XANTENNA__134__A _123_/A vgnd vpwr scs8hd_diode_2
XFILLER_33_3 vgnd vpwr scs8hd_decap_12
Xmux_top_track_4.INVTX1_1_.scs8hd_inv_1 chanx_right_in[3] mux_top_track_4.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mem_top_track_12.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_16_239 vgnd vpwr scs8hd_decap_12
XPHY_278 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_267 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_256 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_245 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmux_top_track_10.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_top_track_10.INVTX1_0_.scs8hd_inv_1/Y
+ _183_/A mux_top_track_10.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XPHY_234 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_223 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_212 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_201 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_3_132 vpwr vgnd scs8hd_fill_2
XANTENNA__104__D _123_/D vgnd vpwr scs8hd_diode_2
XFILLER_3_187 vpwr vgnd scs8hd_fill_2
XANTENNA__129__A _096_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_track_2.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_21_275 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_top_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_8_213 vgnd vpwr scs8hd_fill_1
XFILLER_8_235 vgnd vpwr scs8hd_fill_1
XFILLER_5_57 vpwr vgnd scs8hd_fill_2
XANTENNA__131__B _133_/B vgnd vpwr scs8hd_diode_2
XANTENNA__115__C _123_/C vgnd vpwr scs8hd_diode_2
Xmux_top_track_10.INVTX1_0_.scs8hd_inv_1 top_left_grid_pin_11_ mux_top_track_10.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_38_150 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_top_track_4.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_top_track_4.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_14_44 vgnd vpwr scs8hd_decap_8
XANTENNA__232__A _232_/A vgnd vpwr scs8hd_diode_2
XFILLER_30_21 vgnd vpwr scs8hd_fill_1
XFILLER_5_249 vgnd vpwr scs8hd_decap_6
XFILLER_5_205 vpwr vgnd scs8hd_fill_2
XFILLER_39_52 vgnd vpwr scs8hd_decap_4
XFILLER_36_109 vgnd vpwr scs8hd_fill_1
XANTENNA__126__B _123_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_track_2.LATCH_1_.latch_SLEEPB _147_/Y vgnd vpwr scs8hd_diode_2
Xmux_top_track_14.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_top_track_14.INVTX1_1_.scs8hd_inv_1/Y
+ _187_/Y mux_top_track_14.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XANTENNA__142__A _151_/A vgnd vpwr scs8hd_diode_2
XFILLER_41_123 vgnd vpwr scs8hd_decap_12
XPHY_76 vgnd vpwr scs8hd_decap_3
XPHY_65 vgnd vpwr scs8hd_decap_3
XPHY_54 vgnd vpwr scs8hd_decap_3
XPHY_10 vgnd vpwr scs8hd_decap_3
XPHY_98 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_87 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_21 vgnd vpwr scs8hd_decap_3
XANTENNA__227__A _227_/A vgnd vpwr scs8hd_diode_2
XPHY_32 vgnd vpwr scs8hd_decap_3
XPHY_43 vgnd vpwr scs8hd_decap_3
XFILLER_41_86 vgnd vpwr scs8hd_decap_12
X_192_ _192_/A _192_/Y vgnd vpwr scs8hd_inv_8
Xmux_right_track_14.INVTX1_1_.scs8hd_inv_1 right_bottom_grid_pin_13_ mux_right_track_14.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_17_153 vpwr vgnd scs8hd_fill_2
XFILLER_32_178 vgnd vpwr scs8hd_decap_12
XANTENNA__137__A address[5] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_16.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _206_/Y vgnd
+ vpwr scs8hd_diode_2
XFILLER_23_112 vgnd vpwr scs8hd_fill_1
XFILLER_23_123 vpwr vgnd scs8hd_fill_2
XFILLER_23_178 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_right_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_36_64 vgnd vpwr scs8hd_decap_8
X_175_ _175_/A _175_/Y vgnd vpwr scs8hd_inv_8
XANTENNA__123__C _123_/C vgnd vpwr scs8hd_diode_2
XFILLER_9_171 vgnd vpwr scs8hd_decap_6
XFILLER_9_193 vgnd vpwr scs8hd_decap_12
XFILLER_28_215 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_4.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_4.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_22_88 vgnd vpwr scs8hd_decap_4
XANTENNA__240__A _240_/A vgnd vpwr scs8hd_diode_2
XFILLER_42_273 vgnd vpwr scs8hd_decap_4
X_227_ _227_/A chanx_right_out[7] vgnd vpwr scs8hd_buf_2
XANTENNA__118__C _123_/C vgnd vpwr scs8hd_diode_2
X_158_ _170_/C _159_/B _158_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_6_185 vgnd vpwr scs8hd_fill_1
XANTENNA__134__B _115_/B vgnd vpwr scs8hd_diode_2
XFILLER_26_3 vgnd vpwr scs8hd_decap_12
XANTENNA__150__A _150_/A vgnd vpwr scs8hd_diode_2
XFILLER_17_33 vgnd vpwr scs8hd_decap_3
XFILLER_17_88 vgnd vpwr scs8hd_decap_4
XPHY_279 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_268 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_257 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_246 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_235 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_224 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_213 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_202 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__235__A _235_/A vgnd vpwr scs8hd_diode_2
XFILLER_3_199 vgnd vpwr scs8hd_decap_3
XFILLER_30_276 vgnd vpwr scs8hd_fill_1
XANTENNA__145__A _151_/A vgnd vpwr scs8hd_diode_2
XFILLER_21_243 vgnd vpwr scs8hd_fill_1
XFILLER_0_103 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_10.INVTX1_1_.scs8hd_inv_1_A chanx_right_in[6] vgnd vpwr scs8hd_diode_2
XFILLER_0_147 vpwr vgnd scs8hd_fill_2
Xmux_top_track_2.INVTX1_1_.scs8hd_inv_1 chanx_right_in[2] mux_top_track_2.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_12_276 vgnd vpwr scs8hd_fill_1
XANTENNA__115__D _123_/D vgnd vpwr scs8hd_diode_2
Xmux_top_track_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_top_track_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ _174_/A mux_top_track_2.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XFILLER_5_69 vpwr vgnd scs8hd_fill_2
Xmem_top_track_2.LATCH_1_.latch data_in _174_/A _111_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_14_89 vgnd vpwr scs8hd_decap_3
XFILLER_39_31 vpwr vgnd scs8hd_fill_2
XFILLER_39_75 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_0.tap_buf4_0_.scs8hd_inv_1_A mux_top_track_0.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_track_2.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA__126__C _123_/C vgnd vpwr scs8hd_diode_2
XANTENNA__142__B _141_/B vgnd vpwr scs8hd_diode_2
XFILLER_35_132 vpwr vgnd scs8hd_fill_2
XFILLER_41_135 vgnd vpwr scs8hd_decap_12
XPHY_77 vgnd vpwr scs8hd_decap_3
XPHY_66 vgnd vpwr scs8hd_decap_3
XPHY_55 vgnd vpwr scs8hd_decap_3
XFILLER_26_198 vgnd vpwr scs8hd_decap_12
XFILLER_26_187 vpwr vgnd scs8hd_fill_2
XFILLER_26_154 vgnd vpwr scs8hd_decap_12
XFILLER_25_66 vgnd vpwr scs8hd_fill_1
XPHY_99 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_88 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_11 vgnd vpwr scs8hd_decap_3
XPHY_22 vgnd vpwr scs8hd_decap_3
XPHY_33 vgnd vpwr scs8hd_decap_3
XPHY_44 vgnd vpwr scs8hd_decap_3
XFILLER_41_98 vgnd vpwr scs8hd_decap_12
XANTENNA__243__A _243_/A vgnd vpwr scs8hd_diode_2
X_191_ _191_/A _191_/Y vgnd vpwr scs8hd_inv_8
XFILLER_2_15 vgnd vpwr scs8hd_decap_12
XFILLER_32_102 vgnd vpwr scs8hd_decap_8
XFILLER_40_190 vgnd vpwr scs8hd_decap_12
Xmux_top_track_6.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 _224_/HI _178_/Y mux_top_track_6.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA__153__A _123_/A vgnd vpwr scs8hd_diode_2
XANTENNA__238__A _238_/A vgnd vpwr scs8hd_diode_2
XFILLER_36_32 vgnd vpwr scs8hd_decap_12
XFILLER_14_102 vgnd vpwr scs8hd_decap_3
XFILLER_14_113 vgnd vpwr scs8hd_decap_8
X_243_ _243_/A chany_top_out[0] vgnd vpwr scs8hd_buf_2
XANTENNA__123__D _123_/D vgnd vpwr scs8hd_diode_2
X_174_ _174_/A _174_/Y vgnd vpwr scs8hd_inv_8
XFILLER_28_7 vgnd vpwr scs8hd_decap_6
XANTENNA__148__A _151_/A vgnd vpwr scs8hd_diode_2
Xmux_right_track_12.INVTX1_1_.scs8hd_inv_1 right_bottom_grid_pin_11_ mux_right_track_12.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_9_161 vgnd vpwr scs8hd_decap_4
XFILLER_20_127 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_right_track_14.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_right_track_14.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_28_227 vgnd vpwr scs8hd_decap_12
XFILLER_11_149 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_top_track_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A _222_/HI vgnd vpwr
+ scs8hd_diode_2
XFILLER_22_45 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_top_track_0.LATCH_0_.latch_SLEEPB _107_/Y vgnd vpwr scs8hd_diode_2
XFILLER_42_230 vgnd vpwr scs8hd_decap_12
X_157_ _123_/A address[2] _149_/C _149_/D _159_/B vgnd vpwr scs8hd_or4_4
XFILLER_6_131 vgnd vpwr scs8hd_decap_3
XFILLER_10_193 vgnd vpwr scs8hd_decap_12
X_226_ _226_/A chanx_right_out[8] vgnd vpwr scs8hd_buf_2
XANTENNA__134__C _134_/C vgnd vpwr scs8hd_diode_2
XANTENNA__118__D _110_/D vgnd vpwr scs8hd_diode_2
XANTENNA__150__B _151_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _191_/Y vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_top_track_12.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _184_/Y vgnd vpwr
+ scs8hd_diode_2
XPHY_225 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_214 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_203 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_269 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_258 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_247 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_33_77 vgnd vpwr scs8hd_fill_1
XFILLER_33_66 vgnd vpwr scs8hd_fill_1
XPHY_236 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmem_right_track_16.LATCH_0_.latch data_in _207_/A _171_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_3_178 vpwr vgnd scs8hd_fill_2
XFILLER_3_156 vpwr vgnd scs8hd_fill_2
XFILLER_3_101 vpwr vgnd scs8hd_fill_2
XANTENNA__161__A _170_/C vgnd vpwr scs8hd_diode_2
X_209_ _209_/HI _209_/LO vgnd vpwr scs8hd_conb_1
XANTENNA__145__B _144_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_0.tap_buf4_0_.scs8hd_inv_1_A mux_right_track_0.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_0_70 vgnd vpwr scs8hd_decap_12
XFILLER_21_255 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _180_/Y vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_top_track_16.INVTX1_0_.scs8hd_inv_1_A top_right_grid_pin_11_ vgnd vpwr
+ scs8hd_diode_2
XFILLER_12_211 vgnd vpwr scs8hd_decap_3
Xmux_top_track_10.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 _218_/HI _182_/Y mux_top_track_10.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_5_15 vgnd vpwr scs8hd_decap_12
XFILLER_8_215 vgnd vpwr scs8hd_decap_12
XANTENNA__156__A _171_/C vgnd vpwr scs8hd_diode_2
Xmux_right_track_10.tap_buf4_0_.scs8hd_inv_1 mux_right_track_10.tap_buf4_0_.scs8hd_inv_1/A
+ _229_/A vgnd vpwr scs8hd_inv_1
XFILLER_7_270 vgnd vpwr scs8hd_decap_6
XANTENNA_mux_right_track_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A _213_/HI vgnd vpwr
+ scs8hd_diode_2
XFILLER_14_68 vgnd vpwr scs8hd_fill_1
Xmux_top_track_12.tap_buf4_0_.scs8hd_inv_1 mux_top_track_12.tap_buf4_0_.scs8hd_inv_1/A
+ _237_/A vgnd vpwr scs8hd_inv_1
XANTENNA__126__D _110_/D vgnd vpwr scs8hd_diode_2
XFILLER_4_251 vgnd vpwr scs8hd_decap_12
Xmux_top_track_0.INVTX1_1_.scs8hd_inv_1 chanx_right_in[1] mux_top_track_0.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XPHY_12 vgnd vpwr scs8hd_decap_3
XFILLER_41_147 vgnd vpwr scs8hd_decap_12
XPHY_78 vgnd vpwr scs8hd_decap_3
XPHY_67 vgnd vpwr scs8hd_decap_3
XPHY_56 vgnd vpwr scs8hd_decap_3
XFILLER_26_166 vgnd vpwr scs8hd_decap_12
XFILLER_25_56 vgnd vpwr scs8hd_decap_4
XPHY_89 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_23 vgnd vpwr scs8hd_decap_3
X_190_ _190_/A _190_/Y vgnd vpwr scs8hd_inv_8
XPHY_34 vgnd vpwr scs8hd_decap_3
XPHY_45 vgnd vpwr scs8hd_decap_3
XFILLER_2_27 vgnd vpwr scs8hd_decap_4
XANTENNA__153__B address[2] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _193_/A vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mem_top_track_12.LATCH_0_.latch_SLEEPB _133_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_14.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _186_/A vgnd vpwr
+ scs8hd_diode_2
Xmux_top_track_4.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_top_track_4.INVTX1_0_.scs8hd_inv_1/Y
+ _177_/A mux_top_track_4.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A vgnd vpwr scs8hd_ebufn_2
XFILLER_23_147 vpwr vgnd scs8hd_fill_2
XFILLER_31_180 vgnd vpwr scs8hd_decap_3
XFILLER_11_69 vpwr vgnd scs8hd_fill_2
XFILLER_36_88 vgnd vpwr scs8hd_decap_4
XFILLER_36_44 vpwr vgnd scs8hd_fill_2
XFILLER_14_125 vgnd vpwr scs8hd_decap_6
X_173_ _173_/A _173_/Y vgnd vpwr scs8hd_inv_8
X_242_ _242_/A chany_top_out[1] vgnd vpwr scs8hd_buf_2
XANTENNA__148__B _147_/B vgnd vpwr scs8hd_diode_2
XANTENNA__164__A _170_/C vgnd vpwr scs8hd_diode_2
XFILLER_28_239 vgnd vpwr scs8hd_decap_12
XFILLER_42_242 vgnd vpwr scs8hd_decap_6
XFILLER_8_15 vgnd vpwr scs8hd_decap_12
X_225_ _225_/HI _225_/LO vgnd vpwr scs8hd_conb_1
X_156_ _171_/C _153_/X _156_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_6_110 vgnd vpwr scs8hd_decap_4
XFILLER_6_154 vgnd vpwr scs8hd_decap_4
XFILLER_10_150 vgnd vpwr scs8hd_decap_3
XANTENNA__134__D _110_/D vgnd vpwr scs8hd_diode_2
XFILLER_33_220 vgnd vpwr scs8hd_decap_12
XFILLER_25_209 vgnd vpwr scs8hd_decap_12
XANTENNA__159__A _171_/C vgnd vpwr scs8hd_diode_2
XFILLER_17_13 vgnd vpwr scs8hd_decap_12
XPHY_259 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_248 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_237 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_226 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_215 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_204 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmux_right_track_10.INVTX1_1_.scs8hd_inv_1 right_bottom_grid_pin_9_ mux_right_track_10.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_17_57 vpwr vgnd scs8hd_fill_2
XFILLER_33_89 vpwr vgnd scs8hd_fill_2
Xmux_top_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_top_track_8.INVTX1_1_.scs8hd_inv_1/Y
+ _181_/Y mux_top_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XFILLER_15_220 vgnd vpwr scs8hd_decap_12
XFILLER_15_253 vpwr vgnd scs8hd_fill_2
XANTENNA__161__B _162_/B vgnd vpwr scs8hd_diode_2
X_139_ _163_/C _149_/C vgnd vpwr scs8hd_buf_1
X_208_ _208_/HI _208_/LO vgnd vpwr scs8hd_conb_1
Xmux_right_track_4.tap_buf4_0_.scs8hd_inv_1 mux_right_track_4.tap_buf4_0_.scs8hd_inv_1/A
+ _232_/A vgnd vpwr scs8hd_inv_1
XFILLER_31_3 vgnd vpwr scs8hd_decap_12
XFILLER_21_201 vgnd vpwr scs8hd_decap_12
XFILLER_21_245 vgnd vpwr scs8hd_decap_4
XFILLER_21_267 vgnd vpwr scs8hd_decap_8
XFILLER_0_116 vpwr vgnd scs8hd_fill_2
XFILLER_0_138 vgnd vpwr scs8hd_decap_3
XANTENNA_mem_right_track_10.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_track_10.LATCH_1_.latch_SLEEPB _127_/Y vgnd vpwr scs8hd_diode_2
XFILLER_28_23 vgnd vpwr scs8hd_decap_8
XFILLER_8_227 vgnd vpwr scs8hd_decap_8
XFILLER_12_256 vgnd vpwr scs8hd_decap_8
XFILLER_12_267 vgnd vpwr scs8hd_decap_8
XFILLER_5_27 vgnd vpwr scs8hd_decap_12
XFILLER_8_249 vgnd vpwr scs8hd_decap_4
XFILLER_39_109 vgnd vpwr scs8hd_decap_12
XANTENNA__172__A _172_/A vgnd vpwr scs8hd_diode_2
XANTENNA__156__B _153_/X vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _172_/A vgnd vpwr
+ scs8hd_diode_2
XFILLER_30_46 vpwr vgnd scs8hd_fill_2
XFILLER_30_24 vgnd vpwr scs8hd_decap_6
XFILLER_39_88 vgnd vpwr scs8hd_decap_6
XFILLER_39_66 vgnd vpwr scs8hd_decap_3
XFILLER_39_11 vgnd vpwr scs8hd_fill_1
XFILLER_4_263 vgnd vpwr scs8hd_decap_12
XANTENNA__167__A _167_/A vgnd vpwr scs8hd_diode_2
XFILLER_26_145 vpwr vgnd scs8hd_fill_2
XPHY_13 vgnd vpwr scs8hd_decap_3
XPHY_24 vgnd vpwr scs8hd_decap_3
XPHY_35 vgnd vpwr scs8hd_decap_3
XPHY_46 vgnd vpwr scs8hd_decap_3
XFILLER_41_159 vgnd vpwr scs8hd_decap_12
XPHY_79 vgnd vpwr scs8hd_decap_3
XPHY_68 vgnd vpwr scs8hd_decap_3
XPHY_57 vgnd vpwr scs8hd_decap_3
XFILLER_17_134 vpwr vgnd scs8hd_fill_2
XFILLER_17_178 vgnd vpwr scs8hd_decap_3
XANTENNA__153__C _149_/C vgnd vpwr scs8hd_diode_2
Xmux_top_track_12.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_top_track_12.INVTX1_1_.scs8hd_inv_1/Y
+ _185_/Y mux_top_track_12.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XFILLER_23_115 vgnd vpwr scs8hd_decap_4
XFILLER_23_159 vpwr vgnd scs8hd_fill_2
Xmux_right_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ _198_/A mux_right_track_8.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_top_track_14.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_top_track_14.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
X_241_ _241_/A chany_top_out[2] vgnd vpwr scs8hd_buf_2
X_172_ _172_/A _172_/Y vgnd vpwr scs8hd_inv_8
XANTENNA__164__B _165_/B vgnd vpwr scs8hd_diode_2
XANTENNA__180__A _180_/A vgnd vpwr scs8hd_diode_2
XFILLER_3_71 vgnd vpwr scs8hd_decap_4
XFILLER_36_251 vgnd vpwr scs8hd_decap_12
XFILLER_11_118 vpwr vgnd scs8hd_fill_2
X_224_ _224_/HI _224_/LO vgnd vpwr scs8hd_conb_1
XFILLER_8_27 vgnd vpwr scs8hd_decap_4
X_155_ address[0] _171_/C vgnd vpwr scs8hd_buf_1
XFILLER_6_199 vgnd vpwr scs8hd_decap_12
XFILLER_10_162 vgnd vpwr scs8hd_decap_3
XFILLER_33_232 vgnd vpwr scs8hd_decap_12
XANTENNA__159__B _159_/B vgnd vpwr scs8hd_diode_2
XFILLER_18_251 vgnd vpwr scs8hd_decap_12
XANTENNA__175__A _175_/A vgnd vpwr scs8hd_diode_2
XFILLER_17_25 vgnd vpwr scs8hd_decap_8
XFILLER_17_47 vpwr vgnd scs8hd_fill_2
XPHY_249 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_238 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_227 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_216 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_205 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_276 vgnd vpwr scs8hd_fill_1
XFILLER_3_114 vpwr vgnd scs8hd_fill_2
XFILLER_3_136 vgnd vpwr scs8hd_decap_6
XFILLER_15_232 vgnd vpwr scs8hd_decap_12
Xmem_top_track_16.LATCH_1_.latch data_in _188_/A _141_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_30_202 vgnd vpwr scs8hd_decap_12
X_207_ _207_/A _207_/Y vgnd vpwr scs8hd_inv_8
X_138_ address[4] _166_/D _163_/C vgnd vpwr scs8hd_nand2_4
XFILLER_24_3 vgnd vpwr scs8hd_decap_12
XFILLER_2_191 vgnd vpwr scs8hd_decap_12
XFILLER_0_94 vgnd vpwr scs8hd_fill_1
XFILLER_21_213 vgnd vpwr scs8hd_decap_12
XFILLER_9_70 vpwr vgnd scs8hd_fill_2
XFILLER_28_13 vgnd vpwr scs8hd_fill_1
XFILLER_28_46 vgnd vpwr scs8hd_decap_3
XFILLER_12_235 vgnd vpwr scs8hd_fill_1
XANTENNA_mem_right_track_12.LATCH_0_.latch_SLEEPB _165_/Y vgnd vpwr scs8hd_diode_2
XFILLER_5_39 vgnd vpwr scs8hd_decap_12
Xmem_right_track_12.LATCH_0_.latch data_in _203_/A _165_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mem_top_track_8.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_38_154 vgnd vpwr scs8hd_decap_12
XFILLER_14_15 vgnd vpwr scs8hd_decap_12
XFILLER_30_36 vgnd vpwr scs8hd_decap_8
XFILLER_5_209 vgnd vpwr scs8hd_decap_12
XFILLER_39_56 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_top_track_6.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_top_track_6.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_29_132 vgnd vpwr scs8hd_decap_12
XFILLER_20_91 vgnd vpwr scs8hd_fill_1
XFILLER_35_113 vpwr vgnd scs8hd_fill_2
Xmux_right_track_16.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ _206_/A mux_right_track_16.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XANTENNA__183__A _183_/A vgnd vpwr scs8hd_diode_2
Xmux_top_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_top_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ _172_/A mux_top_track_0.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XFILLER_6_71 vpwr vgnd scs8hd_fill_2
XFILLER_6_93 vpwr vgnd scs8hd_fill_2
Xmux_top_track_0.tap_buf4_0_.scs8hd_inv_1 mux_top_track_0.tap_buf4_0_.scs8hd_inv_1/A
+ _243_/A vgnd vpwr scs8hd_inv_1
XPHY_69 vgnd vpwr scs8hd_decap_3
XPHY_58 vgnd vpwr scs8hd_decap_3
XFILLER_26_135 vgnd vpwr scs8hd_fill_1
XFILLER_26_102 vgnd vpwr scs8hd_decap_4
XFILLER_25_69 vpwr vgnd scs8hd_fill_2
XPHY_47 vgnd vpwr scs8hd_decap_3
XPHY_14 vgnd vpwr scs8hd_decap_3
XPHY_25 vgnd vpwr scs8hd_decap_3
XPHY_36 vgnd vpwr scs8hd_decap_3
XFILLER_34_190 vgnd vpwr scs8hd_decap_12
XFILLER_1_245 vgnd vpwr scs8hd_decap_12
XFILLER_17_113 vgnd vpwr scs8hd_decap_3
XFILLER_32_127 vgnd vpwr scs8hd_fill_1
XFILLER_15_91 vgnd vpwr scs8hd_decap_3
XFILLER_17_157 vpwr vgnd scs8hd_fill_2
XANTENNA__153__D _140_/D vgnd vpwr scs8hd_diode_2
XANTENNA__178__A _178_/A vgnd vpwr scs8hd_diode_2
XFILLER_31_160 vgnd vpwr scs8hd_decap_12
X_240_ _240_/A chany_top_out[3] vgnd vpwr scs8hd_buf_2
X_171_ _110_/D _171_/B _171_/C _171_/Y vgnd vpwr scs8hd_nor3_4
XFILLER_37_208 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_right_track_10.LATCH_1_.latch_SLEEPB _161_/Y vgnd vpwr scs8hd_diode_2
XFILLER_9_131 vpwr vgnd scs8hd_fill_2
XFILLER_13_160 vpwr vgnd scs8hd_fill_2
XFILLER_13_193 vgnd vpwr scs8hd_decap_12
XFILLER_36_263 vgnd vpwr scs8hd_decap_12
Xmux_top_track_4.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 _223_/HI _176_/Y mux_top_track_4.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_right_track_6.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_6.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_42_211 vgnd vpwr scs8hd_decap_6
XFILLER_27_241 vgnd vpwr scs8hd_decap_3
XFILLER_19_208 vgnd vpwr scs8hd_decap_12
X_223_ _223_/HI _223_/LO vgnd vpwr scs8hd_conb_1
X_154_ _170_/C _153_/X _154_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_6_123 vgnd vpwr scs8hd_decap_8
XFILLER_6_145 vgnd vpwr scs8hd_decap_8
XFILLER_19_6 vpwr vgnd scs8hd_fill_2
XFILLER_18_263 vgnd vpwr scs8hd_decap_12
XANTENNA__191__A _191_/A vgnd vpwr scs8hd_diode_2
XPHY_239 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_33_69 vgnd vpwr scs8hd_decap_8
XPHY_228 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_217 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_206 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmem_right_track_8.LATCH_0_.latch data_in _199_/A _159_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
X_137_ address[5] _166_/D vgnd vpwr scs8hd_inv_8
X_206_ _206_/A _206_/Y vgnd vpwr scs8hd_inv_8
XFILLER_23_91 vpwr vgnd scs8hd_fill_2
XFILLER_17_3 vgnd vpwr scs8hd_decap_3
XANTENNA__186__A _186_/A vgnd vpwr scs8hd_diode_2
XFILLER_21_225 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_top_track_8.LATCH_1_.latch_SLEEPB _124_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_track_4.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_10.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _201_/A vgnd
+ vpwr scs8hd_diode_2
XANTENNA__096__A _096_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_4.INVTX1_0_.scs8hd_inv_1_A top_left_grid_pin_5_ vgnd vpwr scs8hd_diode_2
XFILLER_34_90 vpwr vgnd scs8hd_fill_2
XFILLER_18_91 vgnd vpwr scs8hd_fill_1
XFILLER_7_240 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_8.INVTX1_1_.scs8hd_inv_1_A chanx_right_in[5] vgnd vpwr scs8hd_diode_2
XFILLER_38_166 vgnd vpwr scs8hd_decap_12
XFILLER_14_27 vgnd vpwr scs8hd_decap_4
XFILLER_30_59 vgnd vpwr scs8hd_decap_12
XFILLER_29_188 vpwr vgnd scs8hd_fill_2
XFILLER_29_144 vgnd vpwr scs8hd_decap_12
XFILLER_4_276 vgnd vpwr scs8hd_fill_1
XFILLER_20_81 vpwr vgnd scs8hd_fill_2
XFILLER_35_136 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_14.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _187_/Y vgnd vpwr
+ scs8hd_diode_2
XPHY_59 vgnd vpwr scs8hd_decap_3
XFILLER_26_125 vpwr vgnd scs8hd_fill_2
XFILLER_25_48 vpwr vgnd scs8hd_fill_2
XFILLER_25_15 vgnd vpwr scs8hd_decap_4
XPHY_48 vgnd vpwr scs8hd_decap_3
XPHY_15 vgnd vpwr scs8hd_decap_3
XPHY_26 vgnd vpwr scs8hd_decap_3
XPHY_37 vgnd vpwr scs8hd_decap_3
XFILLER_1_257 vgnd vpwr scs8hd_decap_12
XFILLER_1_202 vgnd vpwr scs8hd_decap_12
XFILLER_25_180 vgnd vpwr scs8hd_decap_3
XFILLER_15_70 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _190_/Y vgnd vpwr
+ scs8hd_diode_2
XANTENNA__194__A _194_/A vgnd vpwr scs8hd_diode_2
XFILLER_23_128 vpwr vgnd scs8hd_fill_2
XFILLER_31_172 vgnd vpwr scs8hd_decap_8
XFILLER_11_17 vgnd vpwr scs8hd_decap_12
X_170_ _110_/D _171_/B _170_/C _170_/Y vgnd vpwr scs8hd_nor3_4
XFILLER_3_51 vgnd vpwr scs8hd_fill_1
XANTENNA__189__A _189_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_right_track_16.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_22_49 vgnd vpwr scs8hd_decap_3
XANTENNA__099__A address[4] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_4.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A _223_/HI vgnd vpwr
+ scs8hd_diode_2
XFILLER_27_253 vpwr vgnd scs8hd_fill_2
X_153_ _123_/A address[2] _149_/C _140_/D _153_/X vgnd vpwr scs8hd_or4_4
XFILLER_10_142 vgnd vpwr scs8hd_decap_8
X_222_ _222_/HI _222_/LO vgnd vpwr scs8hd_conb_1
Xmux_top_track_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_top_track_2.INVTX1_0_.scs8hd_inv_1/Y
+ _175_/A mux_top_track_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XFILLER_12_60 vpwr vgnd scs8hd_fill_2
XFILLER_12_71 vgnd vpwr scs8hd_fill_1
XFILLER_12_93 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_2.INVTX1_1_.scs8hd_inv_1_A right_bottom_grid_pin_1_ vgnd
+ vpwr scs8hd_diode_2
XFILLER_33_245 vgnd vpwr scs8hd_decap_12
XPHY_207 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_212 vpwr vgnd scs8hd_fill_2
XFILLER_33_59 vpwr vgnd scs8hd_fill_2
XFILLER_33_15 vgnd vpwr scs8hd_decap_12
XPHY_229 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_218 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_top_track_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_top_track_0.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_30_215 vgnd vpwr scs8hd_decap_12
XFILLER_15_245 vgnd vpwr scs8hd_decap_8
X_205_ _205_/A _205_/Y vgnd vpwr scs8hd_inv_8
XANTENNA_mux_top_track_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _173_/Y vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_top_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _189_/A vgnd vpwr
+ scs8hd_diode_2
X_136_ _151_/A _135_/B _136_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_0_85 vpwr vgnd scs8hd_fill_2
XFILLER_9_50 vgnd vpwr scs8hd_fill_1
XFILLER_9_83 vgnd vpwr scs8hd_decap_6
XFILLER_9_94 vpwr vgnd scs8hd_fill_2
XFILLER_21_237 vgnd vpwr scs8hd_decap_6
XFILLER_12_215 vgnd vpwr scs8hd_decap_12
XFILLER_18_81 vpwr vgnd scs8hd_fill_2
Xmux_top_track_6.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_top_track_6.INVTX1_1_.scs8hd_inv_1/Y
+ _179_/Y mux_top_track_6.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_right_track_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _192_/A vgnd vpwr
+ scs8hd_diode_2
X_119_ _127_/A _119_/B _119_/Y vgnd vpwr scs8hd_nor2_4
Xmem_top_track_12.LATCH_1_.latch data_in _184_/A _131_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_right_track_12.INVTX1_0_.scs8hd_inv_1_A chany_top_in[5] vgnd vpwr scs8hd_diode_2
XFILLER_38_178 vgnd vpwr scs8hd_decap_12
XANTENNA__197__A _197_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_16.INVTX1_1_.scs8hd_inv_1_A right_bottom_grid_pin_15_ vgnd
+ vpwr scs8hd_diode_2
XFILLER_39_36 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_4.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A _214_/HI vgnd vpwr
+ scs8hd_diode_2
XFILLER_29_156 vgnd vpwr scs8hd_decap_12
XFILLER_20_71 vgnd vpwr scs8hd_fill_1
XFILLER_20_93 vpwr vgnd scs8hd_fill_2
XFILLER_35_148 vgnd vpwr scs8hd_decap_12
XFILLER_35_104 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_12.tap_buf4_0_.scs8hd_inv_1_A mux_top_track_12.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_6_84 vpwr vgnd scs8hd_fill_2
XPHY_49 vgnd vpwr scs8hd_decap_3
XPHY_16 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_right_track_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_right_track_0.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XPHY_27 vgnd vpwr scs8hd_decap_3
XPHY_38 vgnd vpwr scs8hd_decap_3
XFILLER_41_59 vpwr vgnd scs8hd_fill_2
XFILLER_41_15 vgnd vpwr scs8hd_decap_12
XFILLER_1_269 vgnd vpwr scs8hd_decap_8
XFILLER_1_214 vgnd vpwr scs8hd_decap_12
XFILLER_9_6 vpwr vgnd scs8hd_fill_2
XFILLER_31_140 vgnd vpwr scs8hd_fill_1
XFILLER_16_170 vgnd vpwr scs8hd_decap_8
XFILLER_31_184 vgnd vpwr scs8hd_decap_12
XFILLER_11_29 vgnd vpwr scs8hd_decap_12
XFILLER_39_262 vgnd vpwr scs8hd_decap_12
XFILLER_36_48 vgnd vpwr scs8hd_decap_12
XFILLER_36_15 vgnd vpwr scs8hd_decap_12
XFILLER_14_107 vgnd vpwr scs8hd_decap_3
XFILLER_22_140 vpwr vgnd scs8hd_fill_2
XFILLER_22_162 vgnd vpwr scs8hd_fill_1
XFILLER_7_3 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _175_/A vgnd vpwr
+ scs8hd_diode_2
XFILLER_13_140 vgnd vpwr scs8hd_decap_4
XFILLER_9_144 vpwr vgnd scs8hd_fill_2
XFILLER_36_276 vgnd vpwr scs8hd_fill_1
XFILLER_3_85 vgnd vpwr scs8hd_fill_1
XANTENNA__099__B address[5] vgnd vpwr scs8hd_diode_2
Xmux_top_track_10.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_top_track_10.INVTX1_1_.scs8hd_inv_1/Y
+ _183_/Y mux_top_track_10.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
X_221_ _221_/HI _221_/LO vgnd vpwr scs8hd_conb_1
XFILLER_10_154 vpwr vgnd scs8hd_fill_2
XFILLER_10_176 vgnd vpwr scs8hd_decap_8
X_152_ _096_/A _170_/C vgnd vpwr scs8hd_buf_1
XANTENNA_mux_right_track_8.INVTX1_0_.scs8hd_inv_1_A chany_top_in[3] vgnd vpwr scs8hd_diode_2
XFILLER_6_169 vgnd vpwr scs8hd_decap_12
Xmux_right_track_6.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_6.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ _196_/A mux_right_track_6.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XFILLER_18_210 vgnd vpwr scs8hd_decap_4
XFILLER_18_276 vgnd vpwr scs8hd_fill_1
XFILLER_33_257 vgnd vpwr scs8hd_decap_12
XPHY_219 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_208 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_33_27 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_top_track_10.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_30_227 vgnd vpwr scs8hd_decap_12
X_204_ _204_/A _204_/Y vgnd vpwr scs8hd_inv_8
XFILLER_15_257 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_top_track_0.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
X_135_ _150_/A _135_/B _135_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_23_82 vpwr vgnd scs8hd_fill_2
XFILLER_2_161 vgnd vpwr scs8hd_decap_4
XFILLER_9_62 vpwr vgnd scs8hd_fill_2
XFILLER_8_209 vgnd vpwr scs8hd_decap_4
XFILLER_12_227 vgnd vpwr scs8hd_decap_8
XFILLER_34_70 vgnd vpwr scs8hd_decap_8
X_118_ _115_/A _115_/B _123_/C _110_/D _119_/B vgnd vpwr scs8hd_or4_4
XFILLER_38_102 vgnd vpwr scs8hd_decap_12
Xmem_right_track_4.LATCH_0_.latch data_in _195_/A _151_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_30_17 vgnd vpwr scs8hd_decap_4
XFILLER_39_59 vpwr vgnd scs8hd_fill_2
XFILLER_39_15 vpwr vgnd scs8hd_fill_2
XFILLER_29_102 vgnd vpwr scs8hd_fill_1
XFILLER_29_168 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_right_track_16.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_26_149 vgnd vpwr scs8hd_decap_4
XPHY_17 vgnd vpwr scs8hd_decap_3
XPHY_28 vgnd vpwr scs8hd_decap_3
XFILLER_41_27 vgnd vpwr scs8hd_decap_12
XPHY_39 vgnd vpwr scs8hd_decap_3
XFILLER_1_226 vgnd vpwr scs8hd_decap_12
XFILLER_32_119 vgnd vpwr scs8hd_decap_8
XFILLER_25_193 vpwr vgnd scs8hd_fill_2
XFILLER_17_105 vpwr vgnd scs8hd_fill_2
XFILLER_17_138 vpwr vgnd scs8hd_fill_2
XFILLER_31_71 vgnd vpwr scs8hd_decap_4
XFILLER_31_130 vpwr vgnd scs8hd_fill_2
XFILLER_23_108 vgnd vpwr scs8hd_decap_4
XFILLER_23_119 vgnd vpwr scs8hd_fill_1
XFILLER_31_196 vgnd vpwr scs8hd_decap_12
Xmux_right_track_14.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_14.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ _204_/A mux_right_track_14.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XFILLER_39_274 vgnd vpwr scs8hd_decap_3
XFILLER_36_27 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_top_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_top_track_16.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_22_152 vgnd vpwr scs8hd_fill_1
XFILLER_22_185 vpwr vgnd scs8hd_fill_2
XFILLER_22_196 vgnd vpwr scs8hd_decap_12
XFILLER_9_123 vgnd vpwr scs8hd_decap_6
XANTENNA_mux_right_track_10.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_10.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_9_167 vpwr vgnd scs8hd_fill_2
XFILLER_3_97 vpwr vgnd scs8hd_fill_2
XFILLER_3_31 vgnd vpwr scs8hd_decap_12
X_220_ _220_/HI _220_/LO vgnd vpwr scs8hd_conb_1
X_151_ _151_/A _151_/B _151_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_12_84 vpwr vgnd scs8hd_fill_2
XFILLER_33_269 vgnd vpwr scs8hd_decap_8
XFILLER_5_170 vgnd vpwr scs8hd_decap_8
XFILLER_33_39 vgnd vpwr scs8hd_decap_12
XPHY_209 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_247 vgnd vpwr scs8hd_decap_3
XFILLER_3_118 vpwr vgnd scs8hd_fill_2
XFILLER_30_239 vgnd vpwr scs8hd_decap_12
XFILLER_15_269 vgnd vpwr scs8hd_decap_8
Xmux_top_track_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 _222_/HI _174_/Y mux_top_track_2.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
X_203_ _203_/A _203_/Y vgnd vpwr scs8hd_inv_8
XFILLER_23_50 vpwr vgnd scs8hd_fill_2
XFILLER_2_140 vgnd vpwr scs8hd_decap_4
X_134_ _123_/A _115_/B _134_/C _110_/D _135_/B vgnd vpwr scs8hd_or4_4
XFILLER_0_32 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_right_track_8.LATCH_0_.latch_SLEEPB _159_/Y vgnd vpwr scs8hd_diode_2
XFILLER_12_239 vgnd vpwr scs8hd_decap_8
XFILLER_34_82 vgnd vpwr scs8hd_decap_8
XFILLER_7_210 vgnd vpwr scs8hd_decap_12
XFILLER_7_254 vpwr vgnd scs8hd_fill_2
X_117_ _128_/A _116_/B _117_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_7_276 vgnd vpwr scs8hd_fill_1
XFILLER_38_114 vgnd vpwr scs8hd_decap_12
XFILLER_15_3 vpwr vgnd scs8hd_fill_2
Xmux_right_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_8.INVTX1_0_.scs8hd_inv_1/Y
+ _199_/A mux_right_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XFILLER_29_114 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_top_track_8.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_track_0.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_20_62 vgnd vpwr scs8hd_decap_3
XFILLER_35_117 vgnd vpwr scs8hd_decap_3
XFILLER_29_71 vpwr vgnd scs8hd_fill_2
Xmem_right_track_16.LATCH_1_.latch data_in _206_/A _170_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XPHY_18 vgnd vpwr scs8hd_decap_3
XPHY_29 vgnd vpwr scs8hd_decap_3
XFILLER_19_180 vgnd vpwr scs8hd_decap_3
XFILLER_41_39 vgnd vpwr scs8hd_decap_12
XFILLER_1_238 vgnd vpwr scs8hd_decap_6
XFILLER_25_172 vpwr vgnd scs8hd_fill_2
XFILLER_15_62 vgnd vpwr scs8hd_decap_3
XFILLER_31_94 vpwr vgnd scs8hd_fill_2
XANTENNA__102__A address[1] vgnd vpwr scs8hd_diode_2
XFILLER_31_120 vpwr vgnd scs8hd_fill_2
XFILLER_39_253 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_right_track_6.LATCH_1_.latch_SLEEPB _154_/Y vgnd vpwr scs8hd_diode_2
XFILLER_9_102 vgnd vpwr scs8hd_fill_1
XFILLER_13_175 vpwr vgnd scs8hd_fill_2
XFILLER_9_179 vpwr vgnd scs8hd_fill_2
XFILLER_3_54 vpwr vgnd scs8hd_fill_2
XFILLER_3_43 vgnd vpwr scs8hd_decap_8
XFILLER_22_19 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_10.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _200_/A vgnd
+ vpwr scs8hd_diode_2
XFILLER_27_245 vgnd vpwr scs8hd_decap_8
X_150_ _150_/A _151_/B _150_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA_mux_right_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_8.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_12_30 vgnd vpwr scs8hd_fill_1
XFILLER_12_52 vgnd vpwr scs8hd_fill_1
XFILLER_12_74 vgnd vpwr scs8hd_fill_1
XFILLER_37_71 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_top_track_12.INVTX1_0_.scs8hd_inv_1_A top_left_grid_pin_13_ vgnd vpwr
+ scs8hd_diode_2
XFILLER_24_259 vgnd vpwr scs8hd_decap_12
XFILLER_24_215 vgnd vpwr scs8hd_decap_12
XFILLER_24_204 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_top_track_16.INVTX1_1_.scs8hd_inv_1_A chanx_right_in[0] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _193_/Y vgnd vpwr
+ scs8hd_diode_2
XANTENNA__200__A _200_/A vgnd vpwr scs8hd_diode_2
X_202_ _202_/A _202_/Y vgnd vpwr scs8hd_inv_8
X_133_ _151_/A _133_/B _133_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_23_40 vgnd vpwr scs8hd_fill_1
XFILLER_23_62 vpwr vgnd scs8hd_fill_2
XFILLER_23_95 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_14.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _186_/Y vgnd vpwr
+ scs8hd_diode_2
XFILLER_2_174 vgnd vpwr scs8hd_decap_8
Xmux_right_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_16.INVTX1_0_.scs8hd_inv_1/Y
+ _207_/A mux_right_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XFILLER_0_44 vgnd vpwr scs8hd_decap_12
XANTENNA__110__A _115_/A vgnd vpwr scs8hd_diode_2
Xmux_top_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_top_track_0.INVTX1_0_.scs8hd_inv_1/Y
+ _173_/A mux_top_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A vgnd vpwr scs8hd_ebufn_2
XFILLER_0_66 vpwr vgnd scs8hd_fill_2
XFILLER_0_99 vpwr vgnd scs8hd_fill_2
XFILLER_9_53 vpwr vgnd scs8hd_fill_2
XFILLER_20_251 vgnd vpwr scs8hd_decap_12
XANTENNA__105__A _127_/A vgnd vpwr scs8hd_diode_2
XFILLER_7_222 vgnd vpwr scs8hd_decap_3
XFILLER_7_266 vpwr vgnd scs8hd_fill_2
XFILLER_11_262 vpwr vgnd scs8hd_fill_2
X_116_ _127_/A _116_/B _116_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_38_126 vgnd vpwr scs8hd_decap_12
XFILLER_20_41 vgnd vpwr scs8hd_decap_12
XFILLER_20_85 vgnd vpwr scs8hd_decap_6
XFILLER_6_32 vgnd vpwr scs8hd_decap_12
XFILLER_26_129 vgnd vpwr scs8hd_decap_6
XFILLER_25_19 vgnd vpwr scs8hd_fill_1
Xmux_top_track_4.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_top_track_4.INVTX1_1_.scs8hd_inv_1/Y
+ _177_/Y mux_top_track_4.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A vgnd vpwr scs8hd_ebufn_2
XPHY_19 vgnd vpwr scs8hd_decap_3
Xmem_top_track_8.LATCH_0_.latch data_in _181_/A _125_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
Xmem_right_track_0.LATCH_0_.latch data_in _191_/A _145_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_17_118 vpwr vgnd scs8hd_fill_2
XFILLER_40_154 vgnd vpwr scs8hd_decap_12
XFILLER_15_74 vpwr vgnd scs8hd_fill_2
XFILLER_15_96 vgnd vpwr scs8hd_decap_3
XANTENNA__102__B _102_/B vgnd vpwr scs8hd_diode_2
XFILLER_0_261 vgnd vpwr scs8hd_decap_12
XPHY_190 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_top_track_10.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_top_track_10.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_39_243 vgnd vpwr scs8hd_fill_1
XFILLER_22_121 vpwr vgnd scs8hd_fill_2
XFILLER_22_154 vpwr vgnd scs8hd_fill_2
XFILLER_22_165 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_right_track_4.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _195_/A vgnd vpwr
+ scs8hd_diode_2
XANTENNA__203__A _203_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _172_/Y vgnd vpwr
+ scs8hd_diode_2
XFILLER_26_84 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_top_track_16.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _188_/A vgnd vpwr
+ scs8hd_diode_2
XFILLER_42_94 vgnd vpwr scs8hd_decap_12
XFILLER_9_114 vpwr vgnd scs8hd_fill_2
XFILLER_13_132 vpwr vgnd scs8hd_fill_2
XANTENNA__113__A address[2] vgnd vpwr scs8hd_diode_2
XFILLER_36_202 vgnd vpwr scs8hd_decap_12
XFILLER_3_77 vgnd vpwr scs8hd_decap_8
XFILLER_8_180 vgnd vpwr scs8hd_decap_4
XFILLER_27_257 vgnd vpwr scs8hd_decap_12
XFILLER_42_249 vgnd vpwr scs8hd_decap_12
XFILLER_6_106 vpwr vgnd scs8hd_fill_2
XFILLER_10_102 vgnd vpwr scs8hd_fill_1
XFILLER_10_113 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_top_track_6.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A _224_/HI vgnd vpwr
+ scs8hd_diode_2
XFILLER_5_3 vgnd vpwr scs8hd_decap_12
Xmux_right_track_0.tap_buf4_0_.scs8hd_inv_1 mux_right_track_0.tap_buf4_0_.scs8hd_inv_1/A
+ _234_/A vgnd vpwr scs8hd_inv_1
XFILLER_12_97 vpwr vgnd scs8hd_fill_2
XANTENNA__108__A address[1] vgnd vpwr scs8hd_diode_2
XFILLER_5_194 vgnd vpwr scs8hd_decap_8
XFILLER_24_227 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_12.tap_buf4_0_.scs8hd_inv_1_A mux_right_track_12.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_top_track_2.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
X_201_ _201_/A _201_/Y vgnd vpwr scs8hd_inv_8
X_132_ address[0] _151_/A vgnd vpwr scs8hd_buf_1
XFILLER_0_56 vgnd vpwr scs8hd_decap_6
XANTENNA__110__B _123_/B vgnd vpwr scs8hd_diode_2
Xmux_right_track_16.tap_buf4_0_.scs8hd_inv_1 mux_right_track_16.tap_buf4_0_.scs8hd_inv_1/A
+ _226_/A vgnd vpwr scs8hd_inv_1
XFILLER_0_89 vpwr vgnd scs8hd_fill_2
XFILLER_9_10 vgnd vpwr scs8hd_decap_12
XFILLER_9_98 vgnd vpwr scs8hd_decap_4
Xmux_right_track_4.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_4.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ _194_/A mux_right_track_4.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XANTENNA_mem_top_track_4.LATCH_0_.latch_SLEEPB _117_/Y vgnd vpwr scs8hd_diode_2
XFILLER_20_263 vgnd vpwr scs8hd_decap_12
XFILLER_18_85 vgnd vpwr scs8hd_decap_6
XANTENNA__105__B _105_/B vgnd vpwr scs8hd_diode_2
XFILLER_11_274 vgnd vpwr scs8hd_decap_3
X_115_ _115_/A _115_/B _123_/C _123_/D _116_/B vgnd vpwr scs8hd_or4_4
XANTENNA__121__A address[3] vgnd vpwr scs8hd_diode_2
XFILLER_38_138 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_4.tap_buf4_0_.scs8hd_inv_1_A mux_top_track_4.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_4_215 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_6.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A _215_/HI vgnd vpwr
+ scs8hd_diode_2
XANTENNA__206__A _206_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _174_/A vgnd vpwr
+ scs8hd_diode_2
XFILLER_29_62 vgnd vpwr scs8hd_decap_3
XFILLER_29_40 vpwr vgnd scs8hd_fill_2
XFILLER_20_97 vgnd vpwr scs8hd_decap_4
XANTENNA__116__A _127_/A vgnd vpwr scs8hd_diode_2
XFILLER_6_44 vgnd vpwr scs8hd_decap_12
XFILLER_6_66 vgnd vpwr scs8hd_decap_3
XFILLER_6_88 vpwr vgnd scs8hd_fill_2
XFILLER_26_119 vgnd vpwr scs8hd_decap_4
XFILLER_26_108 vpwr vgnd scs8hd_fill_2
XFILLER_20_3 vgnd vpwr scs8hd_decap_12
XFILLER_19_160 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_right_track_2.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xmux_right_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 _216_/HI _198_/Y mux_right_track_8.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_40_166 vgnd vpwr scs8hd_decap_12
XFILLER_25_152 vgnd vpwr scs8hd_decap_12
XFILLER_15_31 vgnd vpwr scs8hd_decap_12
XFILLER_0_273 vgnd vpwr scs8hd_decap_4
XFILLER_16_130 vpwr vgnd scs8hd_fill_2
XFILLER_31_144 vpwr vgnd scs8hd_fill_2
XPHY_180 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_191 vgnd vpwr scs8hd_tapvpwrvgnd_1
.ends

